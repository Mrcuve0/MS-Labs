
module register_file ( CLK, RESET, ENABLE, RD1, RD2, WR, ADD_WR, ADD_RD1, 
        ADD_RD2, DATAIN, OUT1, OUT2 );
  input [4:0] ADD_WR;
  input [4:0] ADD_RD1;
  input [4:0] ADD_RD2;
  input [63:0] DATAIN;
  output [63:0] OUT1;
  output [63:0] OUT2;
  input CLK, RESET, ENABLE, RD1, RD2, WR;
  wire   n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107,
         n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117,
         n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127,
         n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137,
         n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147,
         n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157,
         n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167,
         n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177,
         n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187,
         n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197,
         n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207,
         n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217,
         n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227,
         n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237,
         n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247,
         n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257,
         n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267,
         n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277,
         n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287,
         n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297,
         n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307,
         n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
         n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
         n4348, n4349, n4350, n4351, n4352, n4353, n5763, n5765, n5767, n5769,
         n5771, n5773, n5775, n5777, n5779, n5781, n5783, n5785, n5787, n5789,
         n5791, n5793, n5795, n5797, n5799, n5801, n5803, n5805, n5807, n5809,
         n5811, n5813, n5815, n5817, n5819, n5821, n5823, n5825, n5827, n5829,
         n5831, n5833, n5835, n5837, n5839, n5841, n5843, n5845, n5847, n5849,
         n5851, n5853, n5855, n5857, n5859, n5861, n5863, n5865, n5867, n5869,
         n5871, n5873, n5875, n5877, n5879, n5881, n5883, n5885, n5887, n5889,
         n5891, n5893, n5895, n5897, n5899, n5901, n5903, n5905, n5907, n5909,
         n5911, n5913, n5915, n5917, n5919, n5921, n5923, n5925, n5927, n5929,
         n5931, n5933, n5935, n5937, n5939, n5941, n5943, n5945, n5947, n5949,
         n5951, n5953, n5955, n5957, n5959, n5961, n5963, n5965, n5967, n5969,
         n5971, n5973, n5975, n5977, n5979, n5981, n5983, n5985, n5987, n5989,
         n5991, n5993, n5995, n5997, n5999, n6001, n6003, n6005, n6007, n6009,
         n6011, n6013, n6015, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
         n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
         n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
         n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
         n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
         n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
         n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
         n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
         n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
         n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
         n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
         n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
         n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
         n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
         n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8450, n8453, n8456, n8459, n8462, n8465, n8468, n8471,
         n8474, n8477, n8480, n8483, n8486, n8489, n8492, n8495, n8498, n8501,
         n8504, n8507, n8510, n8513, n8516, n8519, n8522, n8525, n8528, n8531,
         n8534, n8537, n8540, n8543, n8546, n8549, n8552, n8555, n8558, n8561,
         n8564, n8567, n8570, n8573, n8576, n8579, n8582, n8585, n8588, n8591,
         n8594, n8597, n8600, n8603, n8606, n8609, n8612, n8615, n8618, n8621,
         n8624, n8627, n8630, n8633, n8636, n8639, n9249, n9252, n9255, n9258,
         n9261, n9264, n9267, n9270, n9273, n9276, n9279, n9282, n9285, n9288,
         n9291, n9294, n9297, n9300, n9303, n9306, n9309, n9312, n9315, n9318,
         n9321, n9324, n9327, n9330, n9333, n9336, n9339, n9342, n9345, n9348,
         n9351, n9354, n9357, n9360, n9363, n9366, n9369, n9372, n9375, n9378,
         n9381, n9384, n9387, n9390, n9393, n9396, n9399, n9402, n9405, n9408,
         n9411, n9414, n9417, n9420, n9423, n9426, n9429, n9432, n9435, n9438,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18382, n18383,
         n18384, n18399, n18400, n18401, n18416, n18417, n18418, n18433,
         n18434, n18435, n18450, n18451, n18452, n18467, n18468, n18469,
         n18484, n18485, n18486, n18501, n18502, n18503, n18518, n18519,
         n18520, n18535, n18536, n18537, n18552, n18553, n18554, n18569,
         n18570, n18571, n18586, n18587, n18588, n18603, n18604, n18605,
         n18620, n18621, n18622, n18637, n18638, n18639, n18654, n18655,
         n18656, n18671, n18672, n18673, n18688, n18689, n18690, n18705,
         n18706, n18707, n18722, n18723, n18724, n18739, n18740, n18741,
         n18756, n18757, n18758, n18773, n18774, n18775, n18790, n18791,
         n18792, n18807, n18808, n18809, n18824, n18825, n18826, n18841,
         n18842, n18843, n18858, n18859, n18860, n18875, n18876, n18877,
         n18892, n18893, n18894, n18909, n18910, n18911, n18926, n18927,
         n18928, n18943, n18944, n18945, n18960, n18961, n18962, n18977,
         n18978, n18979, n18994, n18995, n18996, n19011, n19012, n19013,
         n19028, n19029, n19030, n19045, n19046, n19047, n19062, n19063,
         n19064, n19079, n19080, n19081, n19096, n19097, n19098, n19113,
         n19114, n19115, n19130, n19131, n19132, n19147, n19148, n19149,
         n19164, n19165, n19166, n19181, n19182, n19183, n19198, n19199,
         n19200, n19215, n19216, n19217, n19232, n19233, n19234, n19249,
         n19250, n19251, n19266, n19267, n19268, n19283, n19284, n19285,
         n19300, n19301, n19302, n19317, n19318, n19319, n19334, n19335,
         n19336, n19351, n19352, n19353, n19368, n19369, n19370, n19385,
         n19386, n19387, n19402, n19403, n19404, n19419, n19420, n19421,
         n19436, n19437, n19438, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n20626, n20630, n20631,
         n20632, n20633, n20634, n20635, n20636, n20637, n20638, n20639,
         n20640, n20641, n20642, n20643, n20644, n20645, n20646, n20647,
         n20648, n20649, n20650, n20651, n20652, n20653, n20654, n20655,
         n20656, n20657, n20658, n20659, n20660, n20661, n20662, n20663,
         n20664, n20665, n20666, n20667, n20668, n20669, n20670, n20671,
         n20672, n20673, n20674, n20675, n20676, n20677, n20678, n20679,
         n20680, n20681, n20682, n20683, n20684, n20685, n20686, n20687,
         n20688, n20689, n20690, n20691, n20692, n20693, n20694, n20695,
         n20696, n20697, n20698, n20699, n20700, n20701, n20702, n20703,
         n20704, n20705, n20706, n20707, n20708, n20709, n20710, n20711,
         n20712, n20713, n20714, n20715, n20716, n20717, n20718, n20719,
         n20720, n20721, n20722, n20723, n20724, n20725, n20726, n20727,
         n20728, n20729, n20730, n20731, n20732, n20733, n20734, n20735,
         n20736, n20737, n20738, n20739, n20740, n20741, n20742, n20743,
         n20744, n20745, n20746, n20747, n20748, n20749, n20750, n20751,
         n20752, n20753, n20754, n20755, n20756, n20757, n20758, n20759,
         n20760, n20761, n20762, n20763, n20764, n20765, n20766, n20767,
         n20768, n20769, n20770, n20771, n20772, n20773, n20774, n20775,
         n20776, n20777, n20778, n20779, n20780, n20781, n20782, n20783,
         n20784, n20785, n20786, n20787, n20788, n20789, n20790, n20791,
         n20792, n20793, n20794, n20795, n20796, n20797, n20798, n20799,
         n20800, n20801, n20802, n20803, n20804, n20805, n20806, n20807,
         n20808, n20809, n20810, n20811, n20812, n20813, n20814, n20815,
         n20816, n20817, n20818, n20819, n20820, n20821, n20822, n20823,
         n20824, n20825, n20826, n20827, n20828, n20829, n20830, n20831,
         n20832, n20833, n20834, n20835, n20836, n20837, n20838, n20839,
         n20840, n20841, n20842, n20843, n20844, n20845, n20846, n20847,
         n20848, n20849, n20850, n20851, n20852, n20853, n20854, n20855,
         n20856, n20857, n20858, n20859, n20860, n20861, n20862, n20863,
         n20864, n20865, n20866, n20867, n20868, n20869, n20870, n20871,
         n20872, n20873, n20874, n20875, n20876, n20877, n20878, n20879,
         n20880, n20881, n20882, n20883, n20884, n20885, n20886, n20887,
         n20888, n20889, n20890, n20891, n20892, n20893, n20894, n20895,
         n20896, n20897, n20898, n20899, n20900, n20901, n20902, n20903,
         n20904, n20905, n20906, n20907, n20908, n20909, n20910, n20911,
         n20912, n20913, n20914, n20915, n20916, n20917, n20918, n20919,
         n20920, n20921, n20922, n20923, n20924, n20925, n20926, n20927,
         n20928, n20929, n20930, n20931, n20932, n20933, n20934, n20935,
         n20936, n20937, n20938, n20939, n20940, n20941, n20942, n20943,
         n20944, n20945, n20946, n20947, n20948, n20949, n20950, n20951,
         n20952, n20953, n20954, n20955, n20956, n20957, n20958, n20959,
         n20960, n20961, n20962, n20963, n20964, n20965, n20966, n20967,
         n20968, n20969, n20970, n20971, n20972, n20973, n20974, n20975,
         n20976, n20977, n20978, n20979, n20980, n20981, n20982, n20983,
         n20984, n20985, n20986, n20987, n20988, n20989, n20990, n20991,
         n20992, n20993, n20994, n20995, n20996, n20997, n20998, n20999,
         n21000, n21001, n21002, n21003, n21004, n21005, n21006, n21007,
         n21008, n21009, n21010, n21011, n21012, n21013, n21014, n21015,
         n21016, n21017, n21018, n21019, n21020, n21021, n21022, n21023,
         n21024, n21025, n21026, n21027, n21028, n21029, n21030, n21031,
         n21032, n21033, n21034, n21035, n21036, n21037, n21038, n21039,
         n21040, n21041, n21042, n21043, n21044, n21045, n21046, n21047,
         n21048, n21049, n21050, n21051, n21052, n21053, n21054, n21055,
         n21056, n21057, n21058, n21059, n21060, n21061, n21062, n21063,
         n21064, n21065, n21066, n21067, n21068, n21069, n21070, n21071,
         n21072, n21073, n21074, n21075, n21076, n21077, n21078, n21079,
         n21080, n21081, n21082, n21083, n21084, n21085, n21086, n21087,
         n21088, n21089, n21090, n21091, n21092, n21093, n21094, n21095,
         n21096, n21097, n21098, n21099, n21100, n21101, n21102, n21103,
         n21104, n21105, n21106, n21107, n21108, n21109, n21110, n21111,
         n21112, n21113, n21114, n21115, n21116, n21117, n21118, n21119,
         n21120, n21121, n21122, n21123, n21124, n21125, n21126, n21127,
         n21128, n21129, n21130, n21131, n21132, n21133, n21134, n21135,
         n21136, n21137, n21138, n21139, n21140, n21141, n21142, n21143,
         n21144, n21145, n21146, n21147, n21148, n21149, n21150, n21151,
         n21152, n21153, n21154, n21155, n21156, n21157, n21158, n21159,
         n21160, n21161, n21162, n21163, n21164, n21165, n21166, n21167,
         n21168, n21169, n21170, n21171, n21172, n21173, n21174, n21175,
         n21176, n21177, n21178, n21179, n21180, n21181, n21182, n21183,
         n21184, n21185, n21186, n21187, n21188, n21189, n21190, n21191,
         n21192, n21193, n21194, n21195, n21196, n21197, n21198, n21199,
         n21200, n21201, n21202, n21203, n21204, n21205, n21206, n21207,
         n21208, n21209, n21210, n21211, n21212, n21213, n21214, n21215,
         n21216, n21217, n21218, n21219, n21220, n21221, n21222, n21223,
         n21224, n21225, n21226, n21227, n21228, n21229, n21230, n21231,
         n21232, n21233, n21234, n21235, n21236, n21237, n21238, n21239,
         n21240, n21241, n21242, n21243, n21244, n21245, n21246, n21247,
         n21248, n21249, n21250, n21251, n21252, n21253, n21254, n21255,
         n21256, n21257, n21258, n21259, n21260, n21261, n21262, n21263,
         n21264, n21265, n21266, n21267, n21268, n21269, n21270, n21271,
         n21272, n21273, n21274, n21275, n21276, n21277, n21278, n21279,
         n21280, n21281, n21282, n21283, n21284, n21285, n21286, n21287,
         n21288, n21289, n21290, n21291, n21292, n21293, n21294, n21295,
         n21296, n21297, n21298, n21299, n21300, n21301, n21302, n21303,
         n21304, n21305, n21306, n21307, n21308, n21309, n21310, n21311,
         n21312, n21313, n21314, n21315, n21316, n21317, n21318, n21319,
         n21320, n21321, n21322, n21323, n21324, n21325, n21326, n21327,
         n21328, n21329, n21330, n21331, n21332, n21333, n21334, n21335,
         n21336, n21337, n21338, n21339, n21340, n21341, n21342, n21343,
         n21344, n21345, n21346, n21347, n21348, n21349, n21350, n21351,
         n21352, n21353, n21354, n21355, n21356, n21357, n21358, n21359,
         n21360, n21361, n21362, n21363, n21364, n21365, n21366, n21367,
         n21368, n21369, n21370, n21371, n21372, n21373, n21374, n21375,
         n21376, n21377, n21378, n21379, n21380, n21381, n21382, n21383,
         n21384, n21385, n21386, n21387, n21388, n21389, n21390, n21391,
         n21392, n21393, n21394, n21395, n21396, n21397, n21398, n21399,
         n21400, n21401, n21402, n21403, n21404, n21405, n21406, n21407,
         n21408, n21409, n21410, n21411, n21412, n21413, n21414, n21415,
         n21416, n21417, n21418, n21419, n21420, n21421, n21422, n21423,
         n21424, n21425, n21426, n21427, n21428, n21429, n21430, n21431,
         n21432, n21433, n21434, n21435, n21436, n21437, n21438, n21439,
         n21440, n21441, n21442, n21443, n21444, n21445, n21446, n21447,
         n21448, n21449, n21450, n21451, n21452, n21453, n21454, n21455,
         n21456, n21457, n21458, n21459, n21460, n21461, n21462, n21463,
         n21464, n21465, n21466, n21467, n21468, n21469, n21470, n21471,
         n21472, n21473, n21474, n21475, n21476, n21477, n21478, n21479,
         n21480, n21481, n21482, n21483, n21484, n21485, n21486, n21487,
         n21488, n21489, n21490, n21491, n21492, n21493, n21494, n21495,
         n21496, n21497, n21498, n21499, n21500, n21501, n21502, n21503,
         n21504, n21505, n21506, n21507, n21508, n21509, n21510, n21511,
         n21512, n21513, n21514, n21515, n21516, n21517, n21518, n21519,
         n21520, n21521, n21522, n21523, n21524, n21525, n21526, n21527,
         n21528, n21529, n21530, n21531, n21532, n21533, n21534, n21535,
         n21536, n21537, n21538, n21539, n21540, n21541, n21542, n21543,
         n21544, n21545, n21546, n21547, n21548, n21549, n21550, n21551,
         n21552, n21553, n21554, n21555, n21556, n21557, n21558, n21559,
         n21560, n21561, n21562, n21563, n21564, n21565, n21566, n21567,
         n21568, n21569, n21570, n21571, n21572, n21573, n21574, n21575,
         n21576, n21577, n21578, n21579, n21580, n21581, n21582, n21583,
         n21584, n21585, n21586, n21587, n21588, n21589, n21590, n21591,
         n21592, n21593, n21594, n21595, n21596, n21597, n21598, n21599,
         n21600, n21601, n21602, n21603, n21604, n21605, n21606, n21607,
         n21608, n21609, n21610, n21611, n21612, n21613, n21614, n21615,
         n21616, n21617, n21618, n21619, n21620, n21621, n21622, n21623,
         n21624, n21625, n21626, n21627, n21628, n21629, n21630, n21631,
         n21632, n21633, n21634, n21635, n21636, n21637, n21638, n21639,
         n21640, n21641, n21642, n21643, n21644, n21645, n21646, n21647,
         n21648, n21649, n21650, n21651, n21652, n21653, n21654, n21655,
         n21656, n21657, n21658, n21659, n21660, n21661, n21662, n21663,
         n21664, n21665, n21666, n21667, n21668, n21669, n21670, n21671,
         n21672, n21673, n21674, n21675, n21676, n21677, n21678, n21679,
         n21680, n21681, n21682, n21683, n21684, n21685, n21686, n21687,
         n21688, n21689, n21690, n21691, n21692, n21693, n21694, n21695,
         n21696, n21697, n21698, n21699, n21700, n21701, n21702, n21703,
         n21704, n21705, n21706, n21707, n21708, n21709, n21710, n21711,
         n21712, n21713, n21714, n21715, n21716, n21717, n21718, n21719,
         n21720, n21721, n21722, n21723, n21724, n21725, n21726, n21727,
         n21728, n21729, n21730, n21731, n21732, n21733, n21734, n21735,
         n21736, n21737, n21738, n21739, n21740, n21741, n21742, n21743,
         n21744, n21745, n21746, n21747, n21748, n21749, n21750, n21751,
         n21752, n21753, n21754, n21755, n21756, n21757, n21758, n21759,
         n21760, n21761, n21762, n21763, n21764, n21765, n21766, n21767,
         n21768, n21769, n21770, n21771, n21772, n21773, n21774, n21775,
         n21776, n21777, n21778, n21779, n21780, n21781, n21782, n21783,
         n21784, n21785, n21786, n21787, n21788, n21789, n21790, n21791,
         n21792, n21793, n21794, n21795, n21796, n21797, n21798, n21799,
         n21800, n21801, n21802, n21803, n21804, n21805, n21806, n21807,
         n21808, n21809, n21810, n21811, n21812, n21813, n21814, n21815,
         n21816, n21817, n21818, n21819, n21820, n21821, n21822, n21823,
         n21824, n21825, n21826, n21827, n21828, n21829, n21830, n21831,
         n21832, n21833, n21834, n21835, n21836, n21837, n21838, n21839,
         n21840, n21841, n21842, n21843, n21844, n21845, n21846, n21847,
         n21848, n21849, n21850, n21851, n21852, n21853, n21854, n21855,
         n21856, n21857, n21858, n21859, n21860, n21861, n21862, n21863,
         n21864, n21865, n21866, n21867, n21868, n21869, n21870, n21871,
         n21872, n21873, n21874, n21875, n21876, n21877, n21878, n21879,
         n21880, n21881, n21882, n21883, n21884, n21885, n21886, n21887,
         n21888, n21889, n21890, n21891, n21892, n21893, n21894, n21895,
         n21896, n21897, n21898, n21899, n21900, n21901, n21902, n21903,
         n21904, n21905, n21906, n21907, n21908, n21909, n21910, n21911,
         n21912, n21913, n21914, n21915, n21916, n21917, n21918, n21919,
         n21920, n21921, n21922, n21923, n21924, n21925, n21926, n21927,
         n21928, n21929, n21930, n21931, n21932, n21933, n21934, n21935,
         n21936, n21937, n21938, n21939, n21940, n21941, n21942, n21943,
         n21944, n21945, n21946, n21947, n21948, n21949, n21950, n21951,
         n21952, n21953, n21954, n21955, n21956, n21957, n21958, n21959,
         n21960, n21961, n21962, n21963, n21964, n21965, n21966, n21967,
         n21968, n21969, n21970, n21971, n21972, n21973, n21974, n21975,
         n21976, n21977, n21978, n21979, n21980, n21981, n21982, n21983,
         n21984, n21985, n21986, n21987, n21988, n21989, n21990, n21991,
         n21992, n21993, n21994, n21995, n21996, n21997, n21998, n21999,
         n22000, n22001, n22002, n22003, n22004, n22005, n22006, n22007,
         n22008, n22009, n22010, n22011, n22012, n22013, n22014, n22015,
         n22016, n22017, n22018, n22019, n22020, n22021, n22022, n22023,
         n22024, n22025, n22026, n22027, n22028, n22029, n22030, n22031,
         n22032, n22033, n22034, n22035, n22036, n22037, n22038, n22039,
         n22040, n22041, n22042, n22043, n22044, n22045, n22046, n22047,
         n22048, n22049, n22050, n22051, n22052, n22053, n22054, n22055,
         n22056, n22057, n22058, n22059, n22060, n22061, n22062, n22063,
         n22064, n22065, n22066, n22067, n22068, n22069, n22070, n22071,
         n22072, n22073, n22074, n22075, n22076, n22077, n22078, n22079,
         n22080, n22081, n22082, n22083, n22084, n22085, n22086, n22087,
         n22088, n22089, n22090, n22091, n22092, n22093, n22094, n22095,
         n22096, n22097, n22098, n22099, n22100, n22101, n22102, n22103,
         n22104, n22105, n22106, n22107, n22108, n22109, n22110, n22111,
         n22112, n22113, n22114, n22115, n22116, n22117, n22118, n22119,
         n22120, n22121, n22122, n22123, n22124, n22125, n22126, n22127,
         n22128, n22129, n22130, n22131, n22132, n22133, n22134, n22135,
         n22136, n22137, n22138, n22139, n22140, n22141, n22142, n22143,
         n22144, n22145, n22146, n22147, n22148, n22149, n22150, n22151,
         n22152, n22153, n22154, n22155, n22156, n22157, n22158, n22159,
         n22160, n22161, n22162, n22163, n22164, n22165, n22166, n22167,
         n22168, n22169, n22170, n22171, n22172, n22173, n22174, n22175,
         n22176, n22177, n22178, n22179, n22180, n22181, n22182, n22183,
         n22184, n22185, n22186, n22187, n22188, n22189, n22190, n22191,
         n22192, n22193, n22194, n22195, n22196, n22197, n22198, n22199,
         n22200, n22201, n22202, n22203, n22204, n22205, n22206, n22207,
         n22208, n22209, n22210, n22211, n22212, n22213, n22214, n22215,
         n22216, n22217, n22218, n22219, n22220, n22221, n22222, n22223,
         n22224, n22225, n22226, n22227, n22228, n22229, n22230, n22231,
         n22232, n22233, n22234, n22235, n22236, n22237, n22238, n22239,
         n22240, n22241, n22242, n22243, n22244, n22245, n22246, n22247,
         n22248, n22249, n22250, n22251, n22252, n22253, n22254, n22255,
         n22256, n22257, n22258, n22259, n22260, n22261, n22262, n22263,
         n22264, n22265, n22266, n22267, n22268, n22269, n22270, n22271,
         n22272, n22273, n22274, n22275, n22276, n22277, n22278, n22279,
         n22280, n22281, n22282, n22283, n22284, n22285, n22286, n22287,
         n22288, n22289, n22290, n22291, n22292, n22293, n22294, n22295,
         n22296, n22297, n22298, n22299, n22300, n22301, n22302, n22303,
         n22304, n22305, n22306, n22307, n22308, n22309, n22310, n22311,
         n22312, n22313, n22314, n22315, n22316, n22317, n22318, n22319,
         n22320, n22321, n22322, n22323, n22324, n22325, n22326, n22327,
         n22328, n22329, n22330, n22331, n22332, n22333, n22334, n22335,
         n22336, n22337, n22338, n22339, n22340, n22341, n22342, n22343,
         n22344, n22345, n22346, n22347, n22348, n22349, n22350, n22351,
         n22352, n22353, n22354, n22355, n22356, n22357, n22358, n22359,
         n22360, n22361, n22362, n22363, n22364, n22365, n22366, n22367,
         n22368, n22369, n22370, n22371, n22372, n22373, n22374, n22375,
         n22376, n22377, n22378, n22379, n22380, n22381, n22382, n22383,
         n22384, n22385, n22386, n22387, n22388, n22389, n22390, n22391,
         n22392, n22393, n22394, n22395, n22396, n22397, n22398, n22399,
         n22400, n22401, n22402, n22403, n22404, n22405, n22406, n22407,
         n22408, n22409, n22410, n22411, n22412, n22413, n22414, n22415,
         n22416, n22417, n22418, n22419, n22420, n22421, n22422, n22423,
         n22424, n22425, n22426, n22427, n22428, n22429, n22430, n22431,
         n22432, n22433, n22434, n22435, n22436, n22437, n22438, n22439,
         n22440, n22441, n22442, n22443, n22444, n22445, n22446, n22447,
         n22448, n22449, n22450, n22451, n22452, n22453, n22454, n22455,
         n22456, n22457, n22458, n22459, n22460, n22461, n22462, n22463,
         n22464, n22465, n22466, n22467, n22468, n22469, n22470, n22471,
         n22472, n22473, n22474, n22475, n22476, n22477, n22478, n22479,
         n22480, n22481, n22482, n22483, n22484, n22485, n22486, n22487,
         n22488, n22489, n22490, n22491, n22492, n22493, n22494, n22495,
         n22496, n22497, n22498, n22499, n22500, n22501, n22502, n22503,
         n22504, n22505, n22506, n22507, n22508, n22509, n22510, n22511,
         n22512, n22513, n22514, n22515, n22516, n22517, n22518, n22519,
         n22520, n22521, n22522, n22523, n22524, n22525, n22526, n22527,
         n22528, n22529, n22530, n22531, n22532, n22533, n22534, n22535,
         n22536, n22537, n22538, n22539, n22540, n22541, n22542, n22543,
         n22544, n22545, n22546, n22547, n22548, n22549, n22550, n22551,
         n22552, n22553, n22554, n22555, n22556, n22557, n22558, n22559,
         n22560, n22561, n22562, n22563, n22564, n22565, n22566, n22567,
         n22568, n22569, n22570, n22571, n22572, n22573, n22574, n22575,
         n22576, n22577, n22578, n22579, n22580, n22581, n22582, n22583,
         n22584, n22585, n22586, n22587, n22588, n22589, n22590, n22591,
         n22592, n22593, n22594, n22595, n22596, n22597, n22598, n22599,
         n22600, n22601, n22602, n22603, n22604, n22605, n22606, n22607,
         n22608, n22609, n22610, n22611, n22612, n22613, n22614, n22615,
         n22616, n22617, n22618, n22619, n22620, n22621, n22622, n22623,
         n22624, n22625, n22626, n22627, n22628, n22629, n22630, n22631,
         n22632, n22633, n22634, n22635, n22636, n22637, n22638, n22639,
         n22640, n22641, n22642, n22643, n22644, n22645, n22646, n22647,
         n22648, n22649, n22650, n22651, n22652, n22653, n22654, n22655,
         n22656, n22657, n22658, n22659, n22660, n22661, n22662, n22663,
         n22664, n22665, n22666, n22667, n22668, n22669, n22670, n22671,
         n22672, n22673, n22674, n22675, n22676, n22677, n22678, n22679,
         n22680, n22681, n22682, n22683, n22684, n22685, n22686, n22687,
         n22688, n22689, n22690, n22691, n22692, n22693, n22694, n22695,
         n22696, n22697, n22698, n22699, n22700, n22701, n22702, n22703,
         n22704, n22705, n22706, n22707, n22708, n22709, n22710, n22711,
         n22712, n22713, n22714, n22715, n22716, n22717, n22718, n22719,
         n22720, n22721, n22722, n22723, n22724, n22725, n22726, n22727,
         n22728, n22729, n22730, n22731, n22732, n22733, n22734, n22735,
         n22736, n22737, n22738, n22739, n22740, n22741, n22742, n22743,
         n22744, n22745, n22746, n22747, n22748, n22749, n22750, n22751,
         n22752, n22753, n22754, n22755, n22756, n22757, n22758, n22759,
         n22760, n22761, n22762, n22763, n22764, n22765, n22766, n22767,
         n22768, n22769, n22770, n22771, n22772, n22773, n22774, n22775,
         n22776, n22777, n22778, n22779, n22780, n22781, n22782, n22783,
         n22784, n22785, n22786, n22787, n22788, n22789, n22790, n22791,
         n22792, n22793, n22794, n22795, n22796, n22797, n22798, n22799,
         n22800, n22801, n22802, n22803, n22804, n22805, n22806, n22807,
         n22808, n22809, n22810, n22811, n22812, n22813, n22814, n22815,
         n22816, n22817, n22818, n22819, n22820, n22821, n22822, n22823,
         n22824, n22825, n22826, n22827, n22828, n22829, n22830, n22831,
         n22832, n22833, n22834, n22835, n22836, n22837, n22838, n22839,
         n22840, n22841, n22842, n22843, n22844, n22845, n22846, n22847,
         n22848, n22849, n22850, n22851, n22852, n22853, n22854, n22855,
         n22856, n22857, n22858, n22859, n22860, n22861, n22862, n22863,
         n22864, n22865, n22866, n22867, n22868, n22869, n22870, n22871,
         n22872, n22873, n22874, n22875, n22876, n22877, n22878, n22879,
         n22880, n22881, n22882, n22883, n22884, n22885, n22886, n22887,
         n22888, n22889, n22890, n22891, n22892, n22893, n22894, n22895,
         n22896, n22897, n22898, n22899, n22900, n22901, n22902, n22903,
         n22904, n22905, n22906, n22907, n22908, n22909, n22910, n22911,
         n22912, n22913, n22914, n22915, n22916, n22917, n22918, n22919,
         n22920, n22921, n22922, n22923, n22924, n22925, n22926, n22927,
         n22928, n22929, n22930, n22931, n22932, n22933, n22934, n22935,
         n22936, n22937, n22938, n22939, n22940, n22941, n22942, n22943,
         n22944, n22945, n22946, n22947, n22948, n22949, n22950, n22951,
         n22952, n22953, n22954, n22955, n22956, n22957, n22958, n22959,
         n22960, n22961, n22962, n22963, n22964, n22965, n22966, n22967,
         n22968, n22969, n22970, n22971, n22972, n22973, n22974, n22975,
         n22976, n22977, n22978, n22979, n22980, n22981, n22982, n22983,
         n22984, n22985, n22986, n22987, n22988, n22989, n22990, n22991,
         n22992, n22993, n22994, n22995, n22996, n22997, n22998, n22999,
         n23000, n23001, n23002, n23003, n23004, n23005, n23006, n23007,
         n23008, n23009, n23010, n23011, n23012, n23013, n23014, n23015,
         n23016, n23017, n23018, n23019, n23020, n23021, n23022, n23023,
         n23024, n23025, n23026, n23027, n23028, n23029, n23030, n23031,
         n23032, n23033, n23034, n23035, n23036, n23037, n23038, n23039,
         n23040, n23041, n23042, n23043, n23044, n23045, n23046, n23047,
         n23048, n23049, n23050, n23051, n23052, n23053, n23054, n23055,
         n23056, n23057, n23058, n23059, n23060, n23061, n23062, n23063,
         n23064, n23065, n23066, n23067, n23068, n23069, n23070, n23071,
         n23072, n23073, n23074, n23075, n23076, n23077, n23078, n23079,
         n23080, n23081, n23082, n23083, n23084, n23085, n23086, n23087,
         n23088, n23089, n23090, n23091, n23092, n23093, n23094, n23095,
         n23096, n23097, n23098, n23099, n23100, n23101, n23102, n23103,
         n23104, n23105, n23106, n23107, n23108, n23109, n23110, n23111,
         n23112, n23113, n23114, n23115, n23116, n23117, n23118, n23119,
         n23120, n23121, n23122, n23123, n23124, n23125, n23126, n23127,
         n23128, n23129, n23130, n23131, n23132, n23133, n23134, n23135,
         n23136, n23137, n23138, n23139, n23140, n23141, n23142, n23143,
         n23144, n23145, n23146, n23147, n23148, n23149, n23150, n23151,
         n23152, n23153, n23154, n23155, n23156, n23157, n23158, n23159,
         n23160, n23161, n23162, n23163, n23164, n23165, n23166, n23167,
         n23168, n23169, n23170, n23171, n23172, n23173, n23174, n23175,
         n23176, n23177, n23178, n23179, n23180, n23181, n23182, n23183,
         n23184, n23185, n23186, n23187, n23188, n23189, n23190, n23191,
         n23192, n23193, n23194, n23195, n23196, n23197, n23198, n23199,
         n23200, n23201, n23202, n23203, n23204, n23205, n23206, n23207,
         n23208, n23209, n23210, n23211, n23212, n23213, n23214, n23215,
         n23216, n23217, n23218, n23219, n23220, n23221, n23222, n23223,
         n23224, n23225, n23226, n23227, n23228, n23229, n23230, n23231,
         n23232, n23233, n23234, n23235, n23236, n23237, n23238, n23239,
         n23240, n23241, n23242, n23243, n23244, n23245, n23246, n23247,
         n23248, n23249, n23250, n23251, n23252, n23253, n23254, n23255,
         n23256, n23257, n23258, n23259, n23260, n23261, n23262, n23263,
         n23264, n23265, n23266, n23267, n23268, n23269, n23270, n23271,
         n23272, n23273, n23274, n23275, n23276, n23277, n23278, n23279,
         n23280, n23281, n23282, n23283, n23284, n23285, n23286, n23287,
         n23288, n23289, n23290, n23291, n23292, n23293, n23294, n23295,
         n23296, n23297, n23298, n23299, n23300, n23301, n23302, n23303,
         n23304, n23305, n23306, n23307, n23308, n23309, n23310, n23311,
         n23312, n23313, n23314, n23315, n23316, n23317, n23318, n23319,
         n23320, n23321, n23322, n23323, n23324, n23325, n23326, n23327,
         n23328, n23329, n23330, n23331, n23332, n23333, n23334, n23335,
         n23336, n23337, n23338, n23339, n23340, n23341, n23342, n23343,
         n23344, n23345, n23346, n23347, n23348, n23349, n23350, n23351,
         n23352, n23353, n23354, n23355, n23356, n23357, n23358, n23359,
         n23360, n23361, n23362, n23363, n23364, n23365, n23366, n23367,
         n23368, n23369, n23370, n23371, n23372, n23373, n23374, n23375,
         n23376, n23377, n23378, n23379, n23380, n23381, n23382, n23383,
         n23384, n23385, n23386, n23387, n23388, n23389, n23390, n23391,
         n23392, n23393, n23394, n23395, n23396, n23397, n23398, n23399,
         n23400, n23401, n23402, n23403, n23404, n23405, n23406, n23407,
         n23408, n23409, n23410, n23411, n23412, n23413, n23414, n23415,
         n23416, n23417, n23418, n23419, n23420, n23421, n23422, n23423,
         n23424, n23425, n23426, n23427, n23428, n23429, n23430, n23431,
         n23432, n23433, n23434, n23435, n23436, n23437, n23438, n23439,
         n23440, n23441, n23442, n23443, n23444, n23445, n23446, n23447,
         n23448, n23449, n23450, n23451, n23452, n23453, n23454, n23455,
         n23456, n23457, n23458, n23459, n23460, n23461, n23462, n23463,
         n23464, n23465, n23466, n23467, n23468, n23469, n23470, n23471,
         n23472, n23473, n23474, n23475, n23476, n23477, n23478, n23479,
         n23480, n23481, n23482, n23483, n23484, n23485, n23486, n23487,
         n23488, n23489, n23490, n23491, n23492, n23493, n23494, n23495,
         n23496, n23497, n23498, n23499, n23500, n23501, n23502, n23503,
         n23504, n23505, n23506, n23507, n23508, n23509, n23510, n23511,
         n23512, n23513, n23514, n23515, n23516, n23517, n23518, n23519,
         n23520, n23521, n23522, n23523, n23524, n23525, n23526, n23527,
         n23528, n23529, n23530, n23531, n23532, n23533, n23534, n23535,
         n23536, n23537, n23538, n23539, n23540, n23541, n23542, n23543,
         n23544, n23545, n23546, n23547, n23548, n23549, n23550, n23551,
         n23552, n23553, n23554, n23555, n23556, n23557, n23558, n23559,
         n23560, n23561, n23562, n23563, n23564, n23565, n23566, n23567,
         n23568, n23569, n23570, n23571, n23572, n23573, n23574, n23575,
         n23576, n23577, n23578, n23579, n23580, n23581, n23582, n23583,
         n23584, n23585, n23586, n23587, n23588, n23589, n23590, n23591,
         n23592, n23593, n23594, n23595, n23596, n23597, n23598, n23599,
         n23600, n23601, n23602, n23603, n23604, n23605, n23606, n23607,
         n23608, n23609, n23610, n23611, n23612, n23613, n23614, n23615,
         n23616, n23617, n23618, n23619, n23620, n23621, n23622, n23623,
         n23624, n23625, n23626, n23627, n23628, n23629, n23630, n23631,
         n23632, n23633, n23634, n23635, n23636, n23637, n23638, n23639,
         n23640, n23641, n23642, n23643, n23644, n23645, n23646, n23647,
         n23648, n23649, n23650, n23651, n23652, n23653, n23654, n23655,
         n23656, n23657, n23658, n23659, n23660, n23661, n23662, n23663,
         n23664, n23665, n23666, n23667, n23668, n23669, n23670, n23671,
         n23672, n23673, n23674, n23675, n23676, n23677, n23678, n23679,
         n23680, n23681, n23682, n23683, n23684, n23685, n23686, n23687,
         n23688, n23689, n23690, n23691, n23692, n23693, n23694, n23695,
         n23696, n23697, n23698, n23699, n23700, n23701, n23702, n23703,
         n23704, n23705, n23706, n23707, n23708, n23709, n23710, n23711,
         n23712, n23713, n23714, n23715, n23716, n23717, n23718, n23719,
         n23720, n23721, n23722, n23723, n23724, n23725, n23726, n23727,
         n23728, n23729, n23730, n23731, n23732, n23733, n23734, n23735,
         n23736, n23737, n23738, n23739, n23740, n23741, n23742, n23743,
         n23744, n23745, n23746, n23747, n23748, n23749, n23750, n23751,
         n23752, n23753, n23754, n23755, n23756, n23757, n23758, n23759,
         n23760, n23761, n23762, n23763, n23764, n23765, n23766, n23767,
         n23768, n23769, n23770, n23771, n23772, n23773, n23774, n23775,
         n23776, n23777, n23778, n23779, n23780, n23781, n23782, n23783,
         n23784, n23785, n23786, n23787, n23788, n23789, n23790, n23791,
         n23792, n23793, n23794, n23795, n23796, n23797, n23798, n23799,
         n23800, n23801, n23802, n23803, n23804, n23805, n23806, n23807,
         n23808, n23809, n23810, n23811, n23812, n23813, n23814, n23815,
         n23816, n23817, n23818, n23819, n23820, n23821, n23822, n23823,
         n23824, n23825, n23826, n23827, n23828, n23829, n23830, n23831,
         n23832, n23833, n23834, n23835, n23836, n23837, n23838, n23839,
         n23840, n23841, n23842, n23843, n23844, n23845, n23846, n23847,
         n23848, n23849, n23850, n23851, n23852, n23853, n23854, n23855,
         n23856, n23857, n23858, n23859, n23860, n23861, n23862, n23863,
         n23864, n23865, n23866, n23867, n23868, n23869, n23870, n23871,
         n23872, n23873, n23874, n23875, n23876, n23877, n23878, n23879,
         n23880, n23881, n23882, n23883, n23884, n23885, n23886, n23887,
         n23888, n23889, n23890, n23891, n23892, n23893, n23894, n23895,
         n23896, n23897, n23898, n23899, n23900, n23901, n23902, n23903,
         n23904, n23905, n23906, n23907, n23908, n23909, n23910, n23911,
         n23912, n23913, n23914, n23915, n23916, n23917, n23918, n23919,
         n23920, n23921, n23922, n23923, n23924, n23925, n23926, n23927,
         n23928, n23929, n23930, n23931, n23932, n23933, n23934, n23935,
         n23936, n23937, n23938, n23939, n23940, n23941, n23942, n23943,
         n23944, n23945, n23946, n23947, n23948, n23949, n23950, n23951,
         n23952, n23953, n23954, n23955, n23956, n23957, n23958, n23959,
         n23960, n23961, n23962, n23963, n23964, n23965, n23966, n23967,
         n23968, n23969, n23970, n23971, n23972, n23973, n23974, n23975,
         n23976, n23977, n23978, n23979, n23980, n23981, n23982, n23983,
         n23984, n23985, n23986, n23987, n23988, n23989, n23990, n23991,
         n23992, n23993, n23994, n23995, n23996, n23997, n23998, n23999,
         n24000, n24001, n24002, n24003, n24004, n24005, n24006, n24007,
         n24008, n24009, n24010, n24011, n24012, n24013, n24014, n24015,
         n24016, n24017, n24018, n24019, n24020, n24021, n24022, n24023,
         n24024, n24025, n24026, n24027, n24028, n24029, n24030, n24031,
         n24032, n24033, n24034, n24035, n24036, n24037, n24038, n24039,
         n24040, n24041, n24042, n24043, n24044, n24045, n24046, n24047,
         n24048, n24049, n24050, n24051, n24052, n24053, n24054, n24055,
         n24056, n24057, n24058, n24059, n24060, n24061, n24062, n24063,
         n24064, n24065, n24066, n24067, n24068, n24069, n24070, n24071,
         n24072, n24073, n24074, n24075, n24076, n24077, n24078, n24079,
         n24080, n24081, n24082, n24083, n24084, n24085, n24086, n24087,
         n24088, n24089, n24090, n24091, n24092, n24093, n24094, n24095,
         n24096, n24097, n24098, n24099, n24100, n24101, n24102, n24103,
         n24104, n24105, n24106, n24107, n24108, n24109, n24110, n24111,
         n24112, n24113, n24114, n24115, n24116, n24117, n24118, n24119,
         n24120, n24121, n24122, n24123, n24124, n24125, n24126, n24127,
         n24128, n24129, n24130, n24131, n24132, n24133, n24134, n24135,
         n24136, n24137, n24138, n24139, n24140, n24141, n24142, n24143,
         n24144, n24145, n24146, n24147, n24148, n24149, n24150, n24151,
         n24152, n24153, n24154, n24155, n24156, n24157, n24158, n24159,
         n24160, n24161, n24162, n24163, n24164, n24165, n24166, n24167,
         n24168, n24169, n24170, n24171, n24172, n24173, n24174, n24175,
         n24176, n24177, n24178, n24179, n24180, n24181, n24182, n24183,
         n24184, n24185, n24186, n24187, n24188, n24189, n24190, n24191,
         n24192, n24193, n24194, n24195, n24196, n24197, n24198, n24199,
         n24200, n24201, n24202, n24203, n24204, n24205, n24206, n24207,
         n24208, n24209, n24210, n24211, n24212, n24213, n24214, n24215,
         n24216, n24217, n24218, n24219, n24220, n24221, n24222, n24223,
         n24224, n24225, n24226, n24227, n24228, n24229, n24230, n24231,
         n24232, n24233, n24234, n24235, n24236, n24237, n24238, n24239,
         n24240, n24241, n24242, n24243, n24244, n24245, n24246, n24247,
         n24248, n24249, n24250, n24251, n24252, n24253, n24254, n24255,
         n24256, n24257, n24258, n24259, n24260, n24261, n24262, n24263,
         n24264, n24265, n24266, n24267, n24268, n24269, n24270, n24271,
         n24272, n24273, n24274, n24275, n24276, n24277, n24278, n24279,
         n24280, n24281, n24282, n24283, n24284, n24285, n24286, n24287,
         n24288, n24289, n24290, n24291, n24292, n24293, n24294, n24295,
         n24296, n24297, n24298, n24299, n24300, n24301, n24302, n24303,
         n24304, n24305, n24306, n24307, n24308, n24309, n24310, n24311,
         n24312, n24313, n24314, n24315, n24316, n24317, n24318, n24319,
         n24320, n24321, n24322, n24323, n24324, n24325, n24326, n24327,
         n24328, n24329, n24330, n24331, n24332, n24333, n24334, n24335,
         n24336, n24337, n24338, n24339, n24340, n24341, n24342, n24343,
         n24344, n24345, n24346, n24347, n24348, n24349, n24350, n24351,
         n24352, n24353, n24354, n24355, n24356, n24357, n24358, n24359,
         n24360, n24361, n24362, n24363, n24364, n24365, n24366, n24367,
         n24368, n24369, n24370, n24371, n24372, n24373, n24374, n24375,
         n24376, n24377, n24378, n24379, n24380, n24381, n24382, n24383,
         n24384, n24385, n24386, n24387, n24388, n24389, n24390, n24391,
         n24392, n24393, n24394, n24395, n24396, n24397, n24398, n24399,
         n24400, n24401, n24402, n24403, n24404, n24405, n24406, n24407,
         n24408, n24409, n24410, n24411, n24412, n24413, n24414, n24415,
         n24416, n24417, n24418, n24419, n24420, n24421, n24422, n24423,
         n24424, n24425, n24426, n24427, n24428, n24429, n24430, n24431,
         n24432, n24433, n24434, n24435, n24436, n24437, n24438, n24439,
         n24440, n24441, n24442, n24443, n24444, n24445, n24446, n24447,
         n24448, n24449, n24450, n24451, n24452, n24453, n24454, n24455,
         n24456, n24457, n24458, n24459, n24460, n24461, n24462, n24463,
         n24464, n24465, n24466, n24467, n24468, n24469, n24470, n24471,
         n24472, n24473, n24474, n24475, n24476, n24477, n24478, n24479,
         n24480, n24481, n24482, n24483, n24484, n24485, n24486, n24487,
         n24488, n24489, n24490, n24491, n24492, n24493, n24494, n24495,
         n24496, n24497, n24498, n24499, n24500, n24501, n24502, n24503,
         n24504, n24505, n24506, n24507, n24508, n24509, n24510, n24511,
         n24512, n24513, n24514, n24515, n24516, n24517, n24518, n24519,
         n24520, n24521, n24522, n24523, n24524, n24525, n24526, n24527,
         n24528, n24529, n24530, n24531, n24532, n24533, n24534, n24535,
         n24536, n24537, n24538, n24539, n24540, n24541, n24542, n24543,
         n24544, n24545, n24546, n24547, n24548, n24549, n24550, n24551,
         n24552, n24553, n24554, n24555, n24556, n24557, n24558, n24559,
         n24560, n24561, n24562, n24563, n24564, n24565, n24566, n24567,
         n24568, n24569, n24570, n24571, n24572, n24573, n24574, n24575,
         n24576, n24577, n24578, n24579, n24580, n24581, n24582, n24583,
         n24584, n24585, n24586, n24587, n24588, n24589, n24590, n24591,
         n24592, n24593, n24594, n24595, n24596, n24597, n24598, n24599,
         n24600, n24601, n24602, n24603, n24604, n24605, n24606, n24607,
         n24608, n24609, n24610, n24611, n24612, n24613, n24614, n24615,
         n24616, n24617, n24618, n24619, n24620, n24621, n24622, n24623,
         n24624, n24625, n24626, n24627, n24628, n24629, n24630, n24631,
         n24632, n24633, n24634, n24635, n24636, n24637, n24638, n24639,
         n24640, n24641, n24642, n24643, n24644, n24645, n24646, n24647,
         n24648, n24649, n24650, n24651, n24652, n24653, n24654, n24655,
         n24656, n24657, n24658, n24659, n24660, n24661, n24662, n24663,
         n24664, n24665, n24666, n24667, n24668, n24669, n24670, n24671,
         n24672, n24673, n24674, n24675, n24676, n24677, n24678, n24679,
         n24680, n24681, n24682, n24683, n24684, n24685, n24686, n24687,
         n24688, n24689, n24690, n24691, n24692, n24693, n24694, n24695,
         n24696, n24697, n24698, n24699, n24700, n24701, n24702, n24703,
         n24704, n24705, n24706, n24707, n24708, n24709, n24710, n24711,
         n24712, n24713, n24714, n24715, n24716, n24717, n24718, n24719,
         n24720, n24721, n24722, n24723, n24724, n24725, n24726, n24727,
         n24728, n24729, n24730, n24731, n24732, n24733, n24734, n24735,
         n24736, n24737, n24738, n24739, n24740, n24741, n24742, n24743,
         n24744, n24745, n24746, n24747, n24748, n24749, n24750, n24751,
         n24752, n24753, n24754, n24755, n24756, n24757, n24758, n24759,
         n24760, n24761, n24762, n24763, n24764, n24765, n24766, n24767,
         n24768, n24769, n24770, n24771, n24772, n24773, n24774, n24775,
         n24776, n24777, n24778, n24779, n24780, n24781, n24782, n24783,
         n24784, n24785, n24786, n24787, n24788, n24789, n24790, n24791,
         n24792, n24793, n24794, n24795, n24796, n24797, n24798, n24799,
         n24800, n24801, n24802, n24803, n24804, n24805, n24806, n24807,
         n24808, n24809, n24810, n24811, n24812, n24813, n24814, n24815,
         n24816, n24817, n24818, n24819, n24820, n24821, n24822, n24823,
         n24824, n24825, n24826, n24827, n24828, n24829, n24830, n24831,
         n24832, n24833, n24834, n24835, n24836, n24837, n24838, n24839,
         n24840, n24841, n24842, n24843, n24844, n24845, n24846, n24847,
         n24848, n24849, n24850, n24851, n24852, n24853, n24854, n24855,
         n24856, n24857, n24858, n24859, n24860, n24861, n24862, n24863,
         n24864, n24865, n24866, n24867, n24868, n24869, n24870, n24871,
         n24872, n24873, n24874, n24875, n24876, n24877, n24878, n24879,
         n24880, n24881, n24882, n24883, n24884, n24885, n24886, n24887,
         n24888, n24889, n24890, n24891, n24892, n24893, n24894, n24895,
         n24896, n24897, n24898, n24899, n24900, n24901, n24902, n24903,
         n24904, n24905, n24906, n24907, n24908, n24909, n24910, n24911,
         n24912, n24913, n24914, n24915, n24916, n24917, n24918, n24919,
         n24920, n24921, n24922, n24923, n24924, n24925, n24926, n24927,
         n24928, n24929, n24930, n24931, n24932, n24933, n24934, n24935,
         n24936, n24937, n24938, n24939, n24940, n24941, n24942, n24943,
         n24944, n24945, n24946, n24947, n24948, n24949, n24950, n24951,
         n24952, n24953, n24954, n24955, n24956, n24957, n24958, n24959,
         n24960, n24961, n24962, n24963, n24964, n24965, n24966, n24967,
         n24968, n24969, n24970, n24971, n24972, n24973, n24974, n24975,
         n24976, n24977, n24978, n24979, n24980, n24981, n24982, n24983,
         n24984, n24985, n24986, n24987, n24988, n24989, n24990, n24991,
         n24992, n24993, n24994, n24995, n24996, n24997, n24998, n24999,
         n25000, n25001, n25002, n25003, n25004, n25005, n25006, n25007,
         n25008, n25009, n25010, n25011, n25012, n25013, n25014, n25015,
         n25016, n25017, n25018, n25019, n25020, n25021, n25022, n25023,
         n25024, n25025, n25026, n25027, n25028, n25029, n25030, n25031,
         n25032, n25033, n25034, n25035, n25036, n25037, n25038, n25039,
         n25040, n25041, n25042, n25043, n25044, n25045, n25046, n25047,
         n25048, n25049, n25050, n25051, n25052, n25053, n25054, n25055,
         n25056, n25057, n25058, n25059, n25060, n25061, n25062, n25063,
         n25064, n25065, n25066, n25067, n25068, n25069, n25070, n25071,
         n25072, n25073, n25074, n25075, n25076, n25077, n25078, n25079,
         n25080, n25081, n25082, n25083, n25084, n25085, n25086, n25087,
         n25088, n25089, n25090, n25091, n25092, n25093, n25094, n25095,
         n25096, n25097, n25098, n25099, n25100, n25101, n25102, n25103,
         n25104, n25105, n25106, n25107, n25108, n25109, n25110, n25111,
         n25112, n25113, n25114, n25115, n25116, n25117, n25118, n25119,
         n25120, n25121, n25122, n25123, n25124, n25125, n25126, n25127,
         n25128, n25129, n25130, n25131, n25132, n25133, n25134, n25135,
         n25136, n25137, n25138, n25139, n25140, n25141, n25142, n25143,
         n25144, n25145, n25146, n25147, n25148, n25149, n25150, n25151,
         n25152, n25153, n25154, n25155, n25156, n25157, n25158, n25159,
         n25160, n25161, n25162, n25163, n25164, n25165, n25166, n25215,
         n25216, n25217, n25218, n25219, n25220, n25221, n25222, n25223,
         n25224, n25225, n25226, n25227, n25228, n25229, n25230, n25231,
         n25232, n25233, n25234, n25235, n25236, n25237, n25238, n25239,
         n25240, n25241, n25242, n25243, n25244, n25245, n25246, n25247,
         n25248, n25249, n25250, n25251, n25252, n25253, n25254, n25255,
         n25256, n25257, n25258, n25259, n25260, n25261, n25262, n25311,
         n25312, n25313, n25314, n25315, n25316, n25317, n25318, n25319,
         n25320, n25321, n25322, n25323, n25324, n25325, n25326, n25327,
         n25328, n25329, n25330, n25331, n25332, n25333, n25334, n25335,
         n25336, n25337, n25338, n25339, n25340, n25341, n25342, n25343,
         n25344, n25345, n25346, n25347, n25348, n25349, n25350, n25351,
         n25352, n25353, n25354, n25355, n25356, n25357, n25358, n25407,
         n25408, n25409, n25410, n25411, n25412, n25413, n25414, n25415,
         n25416, n25417, n25418, n25419, n25420, n25421, n25422, n25423,
         n25424, n25425, n25426, n25427, n25428, n25429, n25430, n25431,
         n25432, n25433, n25434, n25435, n25436, n25437, n25438, n25439,
         n25440, n25441, n25442, n25443, n25444, n25445, n25446, n25447,
         n25448, n25449, n25450, n25451, n25452, n25453, n25454, n25455,
         n25456, n25457, n25458, n25459, n25460, n25461, n25462, n25463,
         n25464, n25465, n25466, n25467, n25468, n25469, n25470, n25471,
         n25472, n25473, n25474, n25475, n25476, n25477, n25478, n25479,
         n25480, n25481, n25482, n25483, n25484, n25485, n25486, n25487,
         n25488, n25489, n25490, n25491, n25492, n25493, n25494, n25495,
         n25496, n25497, n25498, n25499, n25500, n25501, n25502, n25503,
         n25504, n25505, n25506, n25507, n25508, n25509, n25510, n25511,
         n25512, n25513, n25514, n25515, n25516, n25517, n25518, n25519,
         n25520, n25521, n25522, n25523, n25524, n25525, n25526, n25527,
         n25528, n25529, n25530, n25531, n25532, n25533, n25534, n25535,
         n25536, n25537, n25538, n25539, n25540, n25541, n25542, n25543,
         n25544, n25545, n25546, n25547, n25548, n25549, n25550, n25555,
         n25556, n25557, n25558, n25563, n25564, n25565, n25566, n25571,
         n25572, n25573, n25574, n25575, n25576, n25577, n25578, n25579,
         n25580, n25581, n25582, n25595, n25596, n25597, n25598, n25599,
         n25600, n25601, n25602, n25603, n25604, n25605, n25606, n25619,
         n25620, n25621, n25622, n25623, n25624, n25625, n25626, n25627,
         n25628, n25629, n25630, n25643, n25644, n25645, n25646, n25647,
         n25648, n25649, n25650, n25651, n25652, n25653, n25654, n25655,
         n25656, n25657, n25658, n25659, n25660, n25661, n25662, n25663,
         n25664, n25665, n25666, n25667, n25668, n25669, n25670, n25671,
         n25672, n25673, n25674, n25675, n25676, n25677, n25678, n25680,
         n25681, n25682, n25685, n25686, n25687, n25690, n25691, n25692,
         n25695, n25696, n25697, n25700, n25701, n25702, n25705, n25706,
         n25707, n25710, n25711, n25712, n25715, n25716, n25717, n25720,
         n25721, n25722, n25725, n25726, n25727, n25730, n25731, n25732,
         n25735, n25736, n25737, n25740, n25741, n25742, n25745, n25746,
         n25747, n25750, n25751, n25752, n25755, n25756, n25757, n25760,
         n25761, n25762, n25765, n25766, n25767, n25770, n25771, n25772,
         n25775, n25776, n25777, n25780, n25781, n25782, n25785, n25786,
         n25787, n25790, n25791, n25792, n25795, n25796, n25797, n25800,
         n25801, n25802, n25805, n25806, n25807, n25810, n25811, n25812,
         n25815, n25816, n25817, n25820, n25821, n25822, n25825, n25826,
         n25827, n25830, n25831, n25832, n25835, n25836, n25837, n25840,
         n25841, n25842, n25845, n25846, n25847, n25850, n25851, n25852,
         n25855, n25856, n25857, n25860, n25861, n25862, n25865, n25866,
         n25867, n25870, n25871, n25872, n25875, n25876, n25877, n25880,
         n25881, n25882, n25885, n25886, n25887, n25890, n25891, n25892,
         n25895, n25896, n25897, n25900, n25901, n25902, n25905, n25906,
         n25907, n25910, n25911, n25912, n25915, n25916, n25917, n25920,
         n25921, n25922, n25925, n25926, n25927, n25930, n25931, n25932,
         n25935, n25936, n25937, n25940, n25941, n25942, n25945, n25946,
         n25947, n25950, n25951, n25952, n25955, n25956, n25957, n25960,
         n25961, n25962, n25965, n25966, n25967, n25970, n25971, n25972,
         n25975, n25976, n25977, n25980, n25981, n25982, n25985, n25986,
         n25987, n25990, n25991, n25992, n25995, n25996, n25997, n26191,
         n26192, n26193, n26194, n26195, n26196, n26197, n26198, n26207,
         n26208, n26209, n26210, n26211, n26212, n26213, n26214, n26215,
         n26216, n26217, n26218, n26219, n26220, n26221, n26222, n26223,
         n26224, n26225, n26226, n26227, n26228, n26229, n26230, n26231,
         n26232, n26233, n26234, n26235, n26236, n26237, n26238, n26239,
         n26240, n26241, n26242, n26243, n26244, n26245, n26246, n26247,
         n26248, n26249, n26250, n26251, n26252, n26253, n26254, n26255,
         n26256, n26257, n26258, n26259, n26260, n26261, n26262, n26263,
         n26264, n26265, n26266, n26327, n26328, n26329, n26330, n26331,
         n26332, n26333, n26334, n26335, n26336, n26337, n26338, n26339,
         n26340, n26341, n26342, n26343, n26344, n26345, n26346, n26347,
         n26348, n26349, n26350, n26351, n26352, n26353, n26354, n26355,
         n26356, n26357, n26358, n26359, n26360, n26361, n26362, n26363,
         n26364, n26365, n26366, n26367, n26368, n26369, n26370, n26371,
         n26372, n26373, n26374, n26375, n26376, n26377, n26378, n26379,
         n26380, n26381, n26382, n26383, n26384, n26385, n26386, n26447,
         n26448, n26449, n26450, n26451, n26452, n26453, n26454, n26455,
         n26456, n26457, n26458, n26459, n26460, n26461, n26462, n26463,
         n26464, n26465, n26466, n26467, n26468, n26469, n26470, n26471,
         n26472, n26473, n26474, n26475, n26476, n26477, n26478, n26479,
         n26480, n26481, n26482, n26483, n26484, n26485, n26486, n26487,
         n26488, n26489, n26490, n26491, n26492, n26493, n26494, n26495,
         n26496, n26497, n26498, n26499, n26500, n26501, n26502, n26503,
         n26504, n26505, n26506, n26507, n26508, n26509, n26510, n26511,
         n26512, n26513, n26514, n26515, n26516, n26517, n26518, n26519,
         n26520, n26521, n26522, n26523, n26524, n26525, n26526, n26527,
         n26528, n26529, n26530, n26531, n26532, n26533, n26534, n26535,
         n26536, n26537, n26538, n26539, n26540, n26541, n26542, n26543,
         n26544, n26545, n26546, n26547, n26548, n26549, n26550, n26551,
         n26552, n26553, n26554, n26555, n26556, n26557, n26558, n26559,
         n26560, n26561, n26562, n26563, n26564, n26565, n26566, n26567,
         n26568, n26569, n26570, n26571, n26572, n26573, n26574, n26575,
         n26576, n26577, n26578, n26579, n26580, n26581, n26582, n26583,
         n26584, n26585, n26586, n26587, n26588, n26589, n26590, n26591,
         n26592, n26593, n26594, n26595, n26596, n26597, n26598, n26599,
         n26600, n26601, n26602, n26603, n26604, n26605, n26606, n26607,
         n26608, n26609, n26610, n26611, n26612, n26613, n26614, n26615,
         n26616, n26617, n26618, n26619, n26620, n26621, n26622, n26623,
         n26624, n26625, n26626, n26627, n26628, n26629, n26630, n26631,
         n26632, n26633, n26634, n26635, n26636, n26637, n26638, n26639,
         n26640, n26641, n26642, n26643, n26644, n26645, n26646, n26647,
         n26648, n26649, n26650, n26651, n26652, n26653, n26654, n26655,
         n26656, n26657, n26658, n26659, n26660, n26661, n26662, n26663,
         n26664, n26665, n26666, n26667, n26668, n26669, n26670, n26671,
         n26672, n26673, n26674, n26675, n26676, n26677, n26678, n26679,
         n26680, n26681, n26682, n26683, n26684, n26685, n26686, n26687,
         n26688, n26689, n26690, n26691, n26692, n26693, n26694, n26695,
         n26696, n26697, n26698, n26699, n26700, n26701, n26702, n26703,
         n26704, n26705, n26706, n26707, n26708, n26709, n26710, n26711,
         n26712, n26713, n26714, n26715, n26716, n26717, n26718, n26719,
         n26720, n26721, n26722, n26723, n26724, n26725, n26726, n26727,
         n26728, n26729, n26730, n26731, n26732, n26733, n26734, n26735,
         n26736, n26737, n26738, n26739, n26740, n26741, n26742, n26743,
         n26744, n26745, n26746, n26747, n26748, n26749, n26750, n26751,
         n26752, n26753, n26754, n26755, n26756, n26757, n26758, n26759,
         n26760, n26761, n26762, n26763, n26764, n26765, n26766, n26767,
         n26768, n26769, n26770, n26771, n26772, n26773, n26774, n26775,
         n26776, n26777, n26778, n26779, n26780, n26781, n26782, n26783,
         n26784, n26785, n26786, n26787, n26788, n26789, n26790, n26791,
         n26792, n26793, n26794, n26795, n26796, n26797, n26798, n26799,
         n26800, n26801, n26802, n26803, n26804, n26805, n26806, n26807,
         n26808, n26809, n26810, n26811, n26812, n26813, n26814, n26815,
         n26816, n26817, n26818, n26819, n26820, n26821, n26822, n26823,
         n26824, n26825, n26826, n26827, n26828, n26829, n26830, n26831,
         n26832, n26833, n26834, n26835, n26836, n26837, n26838, n26839,
         n26840, n26841, n26842, n26843, n26844, n26845, n26846, n26847,
         n26848, n26849, n26850, n26851, n26852, n26853, n26854, n26855,
         n26856, n26857, n26858, n26859, n26860, n26861, n26862, n26863,
         n26864, n26865, n26866, n26867, n26868, n26869, n26870, n26871,
         n26872, n26873, n26874, n26875, n26876, n26877, n26878, n26879,
         n26880, n26881, n26882, n26883, n26884, n26885, n26886, n26887,
         n26888, n26889, n26890, n26891, n26892, n26893, n26894, n26895,
         n26896, n26897, n26898, n26899, n26900, n26901, n26902, n26903,
         n26904, n26905, n26906, n26907, n26908, n26909, n26910, n26911,
         n26912, n26913, n26914, n26915, n26916, n26917, n26918, n26919,
         n26920, n26921, n26922, n26923, n26924, n26925, n26926, n26927,
         n26928, n26929, n26930, n26931, n26932, n26933, n26934, n26935,
         n26936, n26937, n26938, n26939, n26940, n26941, n26942, n26943,
         n26944, n26945, n26946, n26947, n26948, n26949, n26950, n26951,
         n26952, n26953, n26954, n26955, n26956, n26957, n26958, n26959,
         n26960, n26961, n26962, n26963, n26964, n26965, n26966, n26967,
         n26968, n26969, n26970, n26971, n26972, n26973, n26974, n26975,
         n26976, n26977, n26978, n26979, n26980, n26981, n26982, n26983,
         n26984, n26985, n26986, n26987, n26988, n26989, n26990, n26991,
         n26992, n26993, n26994, n26995, n26996, n26997, n26998, n26999,
         n27000, n27001, n27002, n27003, n27004, n27005, n27006, n27007,
         n27008, n27009, n27010, n27011, n27012, n27013, n27014, n27015,
         n27016, n27017, n27018, n27019, n27020, n27021, n27022, n27023,
         n27024, n27025, n27026, n27027, n27028, n27029, n27030, n27031,
         n27032, n27033, n27034, n27035, n27036, n27037, n27038, n27039,
         n27040, n27041, n27042, n27043, n27044, n27045, n27046, n27047,
         n27048, n27049, n27050, n27051, n27052, n27053, n27054, n27055,
         n27056, n27057, n27058, n27059, n27060, n27061, n27062, n27063,
         n27064, n27065, n27066, n27067, n27068, n27069, n27070, n27071,
         n27072, n27073, n27074, n27075, n27076, n27077, n27078, n27079,
         n27080, n27081, n27082, n27083, n27084, n27085, n27086, n27087,
         n27088, n27089, n27090, n27091, n27092, n27093, n27094, n27095,
         n27096, n27097, n27098, n27099, n27100, n27101, n27102, n27103,
         n27104, n27105, n27106, n27107, n27108, n27109, n27110, n27111,
         n27112, n27113, n27114, n27115, n27116, n27117, n27118, n27119,
         n27120, n27121, n27122, n27123, n27124, n27125, n27126, n27127,
         n27128, n27129, n27130, n27131, n27132, n27133, n27134, n27135,
         n27136, n27137, n27138, n27139, n27140, n27141, n27142, n27143,
         n27144, n27145, n27146, n27147, n27148, n27149, n27150, n27151,
         n27152, n27153, n27154, n27155, n27156, n27157, n27158, n27159,
         n27160, n27161, n27162, n27163, n27164, n27165, n27166, n27167,
         n27168, n27169, n27170, n27171, n27172, n27173, n27174, n27175,
         n27176, n27177, n27178, n27179, n27180, n27181, n27182, n27183,
         n27184, n27185, n27186, n27187, n27188, n27189, n27190, n27191,
         n27192, n27193, n27194, n27195, n27196, n27197, n27198, n27199,
         n27200, n27201, n27202, n27203, n27204, n27205, n27206, n27207,
         n27208, n27209, n27210, n27211, n27212, n27213, n27214, n27215,
         n27216, n27217, n27218, n27219, n27220, n27221, n27222, n27223,
         n27224, n27225, n27226, n27227, n27228, n27229, n27230, n27231,
         n27232, n27233, n27234, n27235, n27236, n27237, n27238, n27239,
         n27240, n27241, n27242, n27243, n27244, n27245, n27246, n27247,
         n27248, n27249, n27250, n27251, n27252, n27253, n27254, n27255,
         n27256, n27257, n27258, n27259, n27260, n27261, n27262, n27263,
         n27264, n27265, n27266, n27267, n27268, n27269, n27270, n27271,
         n27272, n27273, n27274, n27275, n27276, n27277, n27278, n27279,
         n27280, n27281, n27282, n27283, n27284, n27285, n27286, n27287,
         n27288, n27289, n27290, n27291, n27292, n27293, n27294, n27295,
         n27296, n27297, n27298, n27299, n27300, n27301, n27302, n27303,
         n27304, n27305, n27306, n27307, n27308, n27309, n27310, n27311,
         n27312, n27313, n27314, n27315, n27316, n27317, n27318, n27319,
         n27320, n27321, n27322, n27323, n27324, n27325, n27326, n27327,
         n27328, n27329, n27330, n27331, n27332, n27333, n27334, n27335,
         n27336, n27337, n27338, n27339, n27340, n27341, n27342, n27343,
         n27344, n27345, n27346, n27347, n27348, n27349, n27350, n27351,
         n27352, n27353, n27354, n27355, n27356, n27357, n27358, n27359,
         n27360, n27361, n27362, n27363, n27364, n27365, n27366, n27367,
         n27368, n27369, n27370, n27371, n27372, n27373, n27374, n27375,
         n27376, n27377, n27378, n27379, n27380, n27381, n27382, n27383,
         n27384, n27385, n27386, n27387, n27388, n27389, n27390, n27391,
         n27392, n27393, n27394, n27395, n27396, n27397, n27398, n27399,
         n27400, n27401, n27402, n27403, n27404, n27405, n27406, n27407,
         n27408, n27409, n27410, n27411, n27412, n27413, n27414, n27415,
         n27416, n27417, n27418, n27419, n27420, n27421, n27422, n27423,
         n27424, n27425, n27426, n27427, n27428, n27429, n27430, n27431,
         n27432, n27433, n27434, n27435, n27436, n27437, n27438, n27439,
         n27440, n27441, n27442, n27443, n27444, n27445, n27446, n27447,
         n27448, n27449, n27450, n27451, n27452, n27453, n27454, n27455,
         n27456, n27457, n27458, n27459, n27460, n27461, n27462, n27463,
         n27464, n27465, n27466, n27467, n27468, n27469, n27470, n27471,
         n27472, n27473, n27474, n27475, n27476, n27477, n27478, n27479,
         n27480, n27481, n27482, n27483, n27484, n27485, n27486, n27487;
  tri   [63:0] OUT1;
  tri   [63:0] OUT2;

  DFF_X1 \OUT1_reg[63]  ( .D(n6017), .CK(CLK), .Q(n4098) );
  DFF_X1 \OUT1_tri_enable_reg[63]  ( .D(n19582), .CK(CLK), .Q(n4099), .QN(
        n18303) );
  DFF_X1 \OUT1_reg[62]  ( .D(n6015), .CK(CLK), .Q(n4100) );
  DFF_X1 \OUT1_tri_enable_reg[62]  ( .D(n19578), .CK(CLK), .Q(n4101), .QN(
        n18304) );
  DFF_X1 \OUT1_reg[61]  ( .D(n6013), .CK(CLK), .Q(n4102) );
  DFF_X1 \OUT1_tri_enable_reg[61]  ( .D(n19581), .CK(CLK), .Q(n4103), .QN(
        n18305) );
  DFF_X1 \OUT1_reg[60]  ( .D(n6011), .CK(CLK), .Q(n4104) );
  DFF_X1 \OUT1_tri_enable_reg[60]  ( .D(n19576), .CK(CLK), .Q(n4105), .QN(
        n18306) );
  DFF_X1 \OUT1_reg[59]  ( .D(n6009), .CK(CLK), .Q(n4106) );
  DFF_X1 \OUT1_tri_enable_reg[59]  ( .D(n19579), .CK(CLK), .Q(n4107), .QN(
        n18307) );
  DFF_X1 \OUT1_reg[58]  ( .D(n6007), .CK(CLK), .Q(n4108) );
  DFF_X1 \OUT1_tri_enable_reg[58]  ( .D(n19549), .CK(CLK), .Q(n4109), .QN(
        n18308) );
  DFF_X1 \OUT1_reg[57]  ( .D(n6005), .CK(CLK), .Q(n4110) );
  DFF_X1 \OUT1_tri_enable_reg[57]  ( .D(n19577), .CK(CLK), .Q(n4111), .QN(
        n18309) );
  DFF_X1 \OUT1_reg[56]  ( .D(n6003), .CK(CLK), .Q(n4112) );
  DFF_X1 \OUT1_tri_enable_reg[56]  ( .D(n19574), .CK(CLK), .Q(n4113), .QN(
        n18310) );
  DFF_X1 \OUT1_reg[55]  ( .D(n6001), .CK(CLK), .Q(n4114) );
  DFF_X1 \OUT1_tri_enable_reg[55]  ( .D(n19575), .CK(CLK), .Q(n4115), .QN(
        n18311) );
  DFF_X1 \OUT1_reg[54]  ( .D(n5999), .CK(CLK), .Q(n4116) );
  DFF_X1 \OUT1_tri_enable_reg[54]  ( .D(n19572), .CK(CLK), .Q(n4117), .QN(
        n18312) );
  DFF_X1 \OUT1_reg[53]  ( .D(n5997), .CK(CLK), .Q(n4118) );
  DFF_X1 \OUT1_tri_enable_reg[53]  ( .D(n19573), .CK(CLK), .Q(n4119), .QN(
        n18313) );
  DFF_X1 \OUT1_reg[52]  ( .D(n5995), .CK(CLK), .Q(n4120) );
  DFF_X1 \OUT1_tri_enable_reg[52]  ( .D(n19570), .CK(CLK), .Q(n4121), .QN(
        n18314) );
  DFF_X1 \OUT1_reg[51]  ( .D(n5993), .CK(CLK), .Q(n4122) );
  DFF_X1 \OUT1_tri_enable_reg[51]  ( .D(n19571), .CK(CLK), .Q(n4123), .QN(
        n18315) );
  DFF_X1 \OUT1_reg[50]  ( .D(n5991), .CK(CLK), .Q(n4124) );
  DFF_X1 \OUT1_tri_enable_reg[50]  ( .D(n19568), .CK(CLK), .Q(n4125), .QN(
        n18316) );
  DFF_X1 \OUT1_reg[49]  ( .D(n5989), .CK(CLK), .Q(n4126) );
  DFF_X1 \OUT1_tri_enable_reg[49]  ( .D(n19569), .CK(CLK), .Q(n4127), .QN(
        n18317) );
  DFF_X1 \OUT1_reg[48]  ( .D(n5987), .CK(CLK), .Q(n4128) );
  DFF_X1 \OUT1_tri_enable_reg[48]  ( .D(n19566), .CK(CLK), .Q(n4129), .QN(
        n18318) );
  DFF_X1 \OUT1_reg[47]  ( .D(n5985), .CK(CLK), .Q(n4130) );
  DFF_X1 \OUT1_tri_enable_reg[47]  ( .D(n19567), .CK(CLK), .Q(n4131), .QN(
        n18319) );
  DFF_X1 \OUT1_reg[46]  ( .D(n5983), .CK(CLK), .Q(n4132) );
  DFF_X1 \OUT1_tri_enable_reg[46]  ( .D(n19564), .CK(CLK), .Q(n4133), .QN(
        n18320) );
  DFF_X1 \OUT1_reg[45]  ( .D(n5981), .CK(CLK), .Q(n4134) );
  DFF_X1 \OUT1_tri_enable_reg[45]  ( .D(n19565), .CK(CLK), .Q(n4135), .QN(
        n18321) );
  DFF_X1 \OUT1_reg[44]  ( .D(n5979), .CK(CLK), .Q(n4136) );
  DFF_X1 \OUT1_tri_enable_reg[44]  ( .D(n19562), .CK(CLK), .Q(n4137), .QN(
        n18322) );
  DFF_X1 \OUT1_reg[43]  ( .D(n5977), .CK(CLK), .Q(n4138) );
  DFF_X1 \OUT1_tri_enable_reg[43]  ( .D(n19563), .CK(CLK), .Q(n4139), .QN(
        n18323) );
  DFF_X1 \OUT1_reg[42]  ( .D(n5975), .CK(CLK), .Q(n4140) );
  DFF_X1 \OUT1_tri_enable_reg[42]  ( .D(n19560), .CK(CLK), .Q(n4141), .QN(
        n18324) );
  DFF_X1 \OUT1_reg[41]  ( .D(n5973), .CK(CLK), .Q(n4142) );
  DFF_X1 \OUT1_tri_enable_reg[41]  ( .D(n19561), .CK(CLK), .Q(n4143), .QN(
        n18325) );
  DFF_X1 \OUT1_reg[40]  ( .D(n5971), .CK(CLK), .Q(n4144) );
  DFF_X1 \OUT1_tri_enable_reg[40]  ( .D(n19558), .CK(CLK), .Q(n4145), .QN(
        n18326) );
  DFF_X1 \OUT1_reg[39]  ( .D(n5969), .CK(CLK), .Q(n4146) );
  DFF_X1 \OUT1_tri_enable_reg[39]  ( .D(n19559), .CK(CLK), .Q(n4147), .QN(
        n18327) );
  DFF_X1 \OUT1_reg[38]  ( .D(n5967), .CK(CLK), .Q(n4148) );
  DFF_X1 \OUT1_tri_enable_reg[38]  ( .D(n19556), .CK(CLK), .Q(n4149), .QN(
        n18328) );
  DFF_X1 \OUT1_reg[37]  ( .D(n5965), .CK(CLK), .Q(n4150) );
  DFF_X1 \OUT1_tri_enable_reg[37]  ( .D(n19557), .CK(CLK), .Q(n4151), .QN(
        n18329) );
  DFF_X1 \OUT1_reg[36]  ( .D(n5963), .CK(CLK), .Q(n4152) );
  DFF_X1 \OUT1_tri_enable_reg[36]  ( .D(n19554), .CK(CLK), .Q(n4153), .QN(
        n18330) );
  DFF_X1 \OUT1_reg[35]  ( .D(n5961), .CK(CLK), .Q(n4154) );
  DFF_X1 \OUT1_tri_enable_reg[35]  ( .D(n19555), .CK(CLK), .Q(n4155), .QN(
        n18331) );
  DFF_X1 \OUT1_reg[34]  ( .D(n5959), .CK(CLK), .Q(n4156) );
  DFF_X1 \OUT1_tri_enable_reg[34]  ( .D(n19552), .CK(CLK), .Q(n4157), .QN(
        n18332) );
  DFF_X1 \OUT1_reg[33]  ( .D(n5957), .CK(CLK), .Q(n4158) );
  DFF_X1 \OUT1_tri_enable_reg[33]  ( .D(n19553), .CK(CLK), .Q(n4159), .QN(
        n18333) );
  DFF_X1 \OUT1_reg[32]  ( .D(n5955), .CK(CLK), .Q(n4160) );
  DFF_X1 \OUT1_tri_enable_reg[32]  ( .D(n19519), .CK(CLK), .Q(n4161), .QN(
        n18334) );
  DFF_X1 \OUT1_reg[31]  ( .D(n5953), .CK(CLK), .Q(n4162) );
  DFF_X1 \OUT1_tri_enable_reg[31]  ( .D(n19551), .CK(CLK), .Q(n4163), .QN(
        n18335) );
  DFF_X1 \OUT1_reg[30]  ( .D(n5951), .CK(CLK), .Q(n4164) );
  DFF_X1 \OUT1_tri_enable_reg[30]  ( .D(n19550), .CK(CLK), .Q(n4165), .QN(
        n18336) );
  DFF_X1 \OUT1_reg[29]  ( .D(n5949), .CK(CLK), .Q(n4166) );
  DFF_X1 \OUT1_tri_enable_reg[29]  ( .D(n19520), .CK(CLK), .Q(n4167), .QN(
        n18337) );
  DFF_X1 \OUT1_reg[28]  ( .D(n5947), .CK(CLK), .Q(n4168) );
  DFF_X1 \OUT1_tri_enable_reg[28]  ( .D(n19548), .CK(CLK), .Q(n4169), .QN(
        n18338) );
  DFF_X1 \OUT1_reg[27]  ( .D(n5945), .CK(CLK), .Q(n4170) );
  DFF_X1 \OUT1_tri_enable_reg[27]  ( .D(n19547), .CK(CLK), .Q(n4171), .QN(
        n18339) );
  DFF_X1 \OUT1_reg[26]  ( .D(n5943), .CK(CLK), .Q(n4172) );
  DFF_X1 \OUT1_tri_enable_reg[26]  ( .D(n19546), .CK(CLK), .Q(n4173), .QN(
        n18340) );
  DFF_X1 \OUT1_reg[25]  ( .D(n5941), .CK(CLK), .Q(n4174) );
  DFF_X1 \OUT1_tri_enable_reg[25]  ( .D(n19545), .CK(CLK), .Q(n4175), .QN(
        n18341) );
  DFF_X1 \OUT1_reg[24]  ( .D(n5939), .CK(CLK), .Q(n4176) );
  DFF_X1 \OUT1_tri_enable_reg[24]  ( .D(n19544), .CK(CLK), .Q(n4177), .QN(
        n18342) );
  DFF_X1 \OUT1_reg[23]  ( .D(n5937), .CK(CLK), .Q(n4178) );
  DFF_X1 \OUT1_tri_enable_reg[23]  ( .D(n19543), .CK(CLK), .Q(n4179), .QN(
        n18343) );
  DFF_X1 \OUT1_reg[22]  ( .D(n5935), .CK(CLK), .Q(n4180) );
  DFF_X1 \OUT1_tri_enable_reg[22]  ( .D(n19542), .CK(CLK), .Q(n4181), .QN(
        n18344) );
  DFF_X1 \OUT1_reg[21]  ( .D(n5933), .CK(CLK), .Q(n4182) );
  DFF_X1 \OUT1_tri_enable_reg[21]  ( .D(n19541), .CK(CLK), .Q(n4183), .QN(
        n18345) );
  DFF_X1 \OUT1_reg[20]  ( .D(n5931), .CK(CLK), .Q(n4184) );
  DFF_X1 \OUT1_tri_enable_reg[20]  ( .D(n19540), .CK(CLK), .Q(n4185), .QN(
        n18346) );
  DFF_X1 \OUT1_reg[19]  ( .D(n5929), .CK(CLK), .Q(n4186) );
  DFF_X1 \OUT1_tri_enable_reg[19]  ( .D(n19539), .CK(CLK), .Q(n4187), .QN(
        n18347) );
  DFF_X1 \OUT1_reg[18]  ( .D(n5927), .CK(CLK), .Q(n4188) );
  DFF_X1 \OUT1_tri_enable_reg[18]  ( .D(n19538), .CK(CLK), .Q(n4189), .QN(
        n18348) );
  DFF_X1 \OUT1_reg[17]  ( .D(n5925), .CK(CLK), .Q(n4190) );
  DFF_X1 \OUT1_tri_enable_reg[17]  ( .D(n19537), .CK(CLK), .Q(n4191), .QN(
        n18349) );
  DFF_X1 \OUT1_reg[16]  ( .D(n5923), .CK(CLK), .Q(n4192) );
  DFF_X1 \OUT1_tri_enable_reg[16]  ( .D(n19536), .CK(CLK), .Q(n4193), .QN(
        n18350) );
  DFF_X1 \OUT1_reg[15]  ( .D(n5921), .CK(CLK), .Q(n4194) );
  DFF_X1 \OUT1_tri_enable_reg[15]  ( .D(n19535), .CK(CLK), .Q(n4195), .QN(
        n18351) );
  DFF_X1 \OUT1_reg[14]  ( .D(n5919), .CK(CLK), .Q(n4196) );
  DFF_X1 \OUT1_tri_enable_reg[14]  ( .D(n19534), .CK(CLK), .Q(n4197), .QN(
        n18352) );
  DFF_X1 \OUT1_reg[13]  ( .D(n5917), .CK(CLK), .Q(n4198) );
  DFF_X1 \OUT1_tri_enable_reg[13]  ( .D(n19533), .CK(CLK), .Q(n4199), .QN(
        n18353) );
  DFF_X1 \OUT1_reg[12]  ( .D(n5915), .CK(CLK), .Q(n4200) );
  DFF_X1 \OUT1_tri_enable_reg[12]  ( .D(n19532), .CK(CLK), .Q(n4201), .QN(
        n18354) );
  DFF_X1 \OUT1_reg[11]  ( .D(n5913), .CK(CLK), .Q(n4202) );
  DFF_X1 \OUT1_tri_enable_reg[11]  ( .D(n19531), .CK(CLK), .Q(n4203), .QN(
        n18355) );
  DFF_X1 \OUT1_reg[10]  ( .D(n5911), .CK(CLK), .Q(n4204) );
  DFF_X1 \OUT1_tri_enable_reg[10]  ( .D(n19530), .CK(CLK), .Q(n4205), .QN(
        n18356) );
  DFF_X1 \OUT1_reg[9]  ( .D(n5909), .CK(CLK), .Q(n4206) );
  DFF_X1 \OUT1_tri_enable_reg[9]  ( .D(n19529), .CK(CLK), .Q(n4207), .QN(
        n18357) );
  DFF_X1 \OUT1_reg[8]  ( .D(n5907), .CK(CLK), .Q(n4208) );
  DFF_X1 \OUT1_tri_enable_reg[8]  ( .D(n19528), .CK(CLK), .Q(n4209), .QN(
        n18358) );
  DFF_X1 \OUT1_reg[7]  ( .D(n5905), .CK(CLK), .Q(n4210) );
  DFF_X1 \OUT1_tri_enable_reg[7]  ( .D(n19527), .CK(CLK), .Q(n4211), .QN(
        n18359) );
  DFF_X1 \OUT1_reg[6]  ( .D(n5903), .CK(CLK), .Q(n4212) );
  DFF_X1 \OUT1_tri_enable_reg[6]  ( .D(n19526), .CK(CLK), .Q(n4213), .QN(
        n18360) );
  DFF_X1 \OUT1_reg[5]  ( .D(n5901), .CK(CLK), .Q(n4214) );
  DFF_X1 \OUT1_tri_enable_reg[5]  ( .D(n19525), .CK(CLK), .Q(n4215), .QN(
        n18361) );
  DFF_X1 \OUT1_reg[4]  ( .D(n5899), .CK(CLK), .Q(n4216) );
  DFF_X1 \OUT1_tri_enable_reg[4]  ( .D(n19524), .CK(CLK), .Q(n4217), .QN(
        n18362) );
  DFF_X1 \OUT1_reg[3]  ( .D(n5897), .CK(CLK), .Q(n4218) );
  DFF_X1 \OUT1_tri_enable_reg[3]  ( .D(n19523), .CK(CLK), .Q(n4219), .QN(
        n18363) );
  DFF_X1 \OUT1_reg[2]  ( .D(n5895), .CK(CLK), .Q(n4220) );
  DFF_X1 \OUT1_tri_enable_reg[2]  ( .D(n19522), .CK(CLK), .Q(n4221), .QN(
        n18364) );
  DFF_X1 \OUT1_reg[1]  ( .D(n5893), .CK(CLK), .Q(n4222) );
  DFF_X1 \OUT1_tri_enable_reg[1]  ( .D(n19521), .CK(CLK), .Q(n4223), .QN(
        n18365) );
  DFF_X1 \OUT1_reg[0]  ( .D(n5891), .CK(CLK), .Q(n4224) );
  DFF_X1 \OUT1_tri_enable_reg[0]  ( .D(n19518), .CK(CLK), .Q(n4225), .QN(
        n18366) );
  DFF_X1 \OUT2_tri_enable_reg[63]  ( .D(n19517), .CK(CLK), .Q(n4227), .QN(
        n18383) );
  DFF_X1 \OUT2_reg[62]  ( .D(n5887), .CK(CLK), .Q(n4228) );
  DFF_X1 \OUT2_tri_enable_reg[62]  ( .D(n19516), .CK(CLK), .Q(n4229), .QN(
        n18400) );
  DFF_X1 \OUT2_reg[61]  ( .D(n5885), .CK(CLK), .Q(n4230) );
  DFF_X1 \OUT2_tri_enable_reg[61]  ( .D(n19515), .CK(CLK), .Q(n4231), .QN(
        n18417) );
  DFF_X1 \OUT2_reg[60]  ( .D(n5883), .CK(CLK), .Q(n4232) );
  DFF_X1 \OUT2_tri_enable_reg[60]  ( .D(n19514), .CK(CLK), .Q(n4233), .QN(
        n18434) );
  DFF_X1 \OUT2_reg[59]  ( .D(n5881), .CK(CLK), .Q(n4234) );
  DFF_X1 \OUT2_tri_enable_reg[59]  ( .D(n19513), .CK(CLK), .Q(n4235), .QN(
        n18451) );
  DFF_X1 \OUT2_reg[58]  ( .D(n5879), .CK(CLK), .Q(n4236) );
  DFF_X1 \OUT2_tri_enable_reg[58]  ( .D(n19512), .CK(CLK), .Q(n4237), .QN(
        n18468) );
  DFF_X1 \OUT2_reg[57]  ( .D(n5877), .CK(CLK), .Q(n4238) );
  DFF_X1 \OUT2_tri_enable_reg[57]  ( .D(n19511), .CK(CLK), .Q(n4239), .QN(
        n18485) );
  DFF_X1 \OUT2_reg[56]  ( .D(n5875), .CK(CLK), .Q(n4240) );
  DFF_X1 \OUT2_tri_enable_reg[56]  ( .D(n19510), .CK(CLK), .Q(n4241), .QN(
        n18502) );
  DFF_X1 \OUT2_reg[55]  ( .D(n5873), .CK(CLK), .Q(n4242) );
  DFF_X1 \OUT2_tri_enable_reg[55]  ( .D(n19509), .CK(CLK), .Q(n4243), .QN(
        n18519) );
  DFF_X1 \OUT2_reg[54]  ( .D(n5871), .CK(CLK), .Q(n4244) );
  DFF_X1 \OUT2_tri_enable_reg[54]  ( .D(n19508), .CK(CLK), .Q(n4245), .QN(
        n18536) );
  DFF_X1 \OUT2_reg[53]  ( .D(n5869), .CK(CLK), .Q(n4246) );
  DFF_X1 \OUT2_tri_enable_reg[53]  ( .D(n19507), .CK(CLK), .Q(n4247), .QN(
        n18553) );
  DFF_X1 \OUT2_reg[52]  ( .D(n5867), .CK(CLK), .Q(n4248) );
  DFF_X1 \OUT2_tri_enable_reg[52]  ( .D(n19506), .CK(CLK), .Q(n4249), .QN(
        n18570) );
  DFF_X1 \OUT2_reg[51]  ( .D(n5865), .CK(CLK), .Q(n4250) );
  DFF_X1 \OUT2_tri_enable_reg[51]  ( .D(n19505), .CK(CLK), .Q(n4251), .QN(
        n18587) );
  DFF_X1 \OUT2_reg[50]  ( .D(n5863), .CK(CLK), .Q(n4252) );
  DFF_X1 \OUT2_tri_enable_reg[50]  ( .D(n19504), .CK(CLK), .Q(n4253), .QN(
        n18604) );
  DFF_X1 \OUT2_reg[49]  ( .D(n5861), .CK(CLK), .Q(n4254) );
  DFF_X1 \OUT2_tri_enable_reg[49]  ( .D(n19503), .CK(CLK), .Q(n4255), .QN(
        n18621) );
  DFF_X1 \OUT2_reg[48]  ( .D(n5859), .CK(CLK), .Q(n4256) );
  DFF_X1 \OUT2_tri_enable_reg[48]  ( .D(n19502), .CK(CLK), .Q(n4257), .QN(
        n18638) );
  DFF_X1 \OUT2_reg[47]  ( .D(n5857), .CK(CLK), .Q(n4258) );
  DFF_X1 \OUT2_tri_enable_reg[47]  ( .D(n19501), .CK(CLK), .Q(n4259), .QN(
        n18655) );
  DFF_X1 \OUT2_reg[46]  ( .D(n5855), .CK(CLK), .Q(n4260) );
  DFF_X1 \OUT2_tri_enable_reg[46]  ( .D(n19500), .CK(CLK), .Q(n4261), .QN(
        n18672) );
  DFF_X1 \OUT2_reg[45]  ( .D(n5853), .CK(CLK), .Q(n4262) );
  DFF_X1 \OUT2_tri_enable_reg[45]  ( .D(n19499), .CK(CLK), .Q(n4263), .QN(
        n18689) );
  DFF_X1 \OUT2_reg[44]  ( .D(n5851), .CK(CLK), .Q(n4264) );
  DFF_X1 \OUT2_tri_enable_reg[44]  ( .D(n19498), .CK(CLK), .Q(n4265), .QN(
        n18706) );
  DFF_X1 \OUT2_reg[43]  ( .D(n5849), .CK(CLK), .Q(n4266) );
  DFF_X1 \OUT2_tri_enable_reg[43]  ( .D(n19497), .CK(CLK), .Q(n4267), .QN(
        n18723) );
  DFF_X1 \OUT2_reg[42]  ( .D(n5847), .CK(CLK), .Q(n4268) );
  DFF_X1 \OUT2_tri_enable_reg[42]  ( .D(n19496), .CK(CLK), .Q(n4269), .QN(
        n18740) );
  DFF_X1 \OUT2_reg[41]  ( .D(n5845), .CK(CLK), .Q(n4270) );
  DFF_X1 \OUT2_tri_enable_reg[41]  ( .D(n19495), .CK(CLK), .Q(n4271), .QN(
        n18757) );
  DFF_X1 \OUT2_reg[40]  ( .D(n5843), .CK(CLK), .Q(n4272) );
  DFF_X1 \OUT2_tri_enable_reg[40]  ( .D(n19494), .CK(CLK), .Q(n4273), .QN(
        n18774) );
  DFF_X1 \OUT2_reg[39]  ( .D(n5841), .CK(CLK), .Q(n4274) );
  DFF_X1 \OUT2_tri_enable_reg[39]  ( .D(n19493), .CK(CLK), .Q(n4275), .QN(
        n18791) );
  DFF_X1 \OUT2_reg[38]  ( .D(n5839), .CK(CLK), .Q(n4276) );
  DFF_X1 \OUT2_tri_enable_reg[38]  ( .D(n19492), .CK(CLK), .Q(n4277), .QN(
        n18808) );
  DFF_X1 \OUT2_reg[37]  ( .D(n5837), .CK(CLK), .Q(n4278) );
  DFF_X1 \OUT2_tri_enable_reg[37]  ( .D(n19491), .CK(CLK), .Q(n4279), .QN(
        n18825) );
  DFF_X1 \OUT2_reg[36]  ( .D(n5835), .CK(CLK), .Q(n4280) );
  DFF_X1 \OUT2_tri_enable_reg[36]  ( .D(n19490), .CK(CLK), .Q(n4281), .QN(
        n18842) );
  DFF_X1 \OUT2_reg[35]  ( .D(n5833), .CK(CLK), .Q(n4282) );
  DFF_X1 \OUT2_tri_enable_reg[35]  ( .D(n19489), .CK(CLK), .Q(n4283), .QN(
        n18859) );
  DFF_X1 \OUT2_reg[34]  ( .D(n5831), .CK(CLK), .Q(n4284) );
  DFF_X1 \OUT2_tri_enable_reg[34]  ( .D(n19488), .CK(CLK), .Q(n4285), .QN(
        n18876) );
  DFF_X1 \OUT2_reg[33]  ( .D(n5829), .CK(CLK), .Q(n4286) );
  DFF_X1 \OUT2_tri_enable_reg[33]  ( .D(n19487), .CK(CLK), .Q(n4287), .QN(
        n18893) );
  DFF_X1 \OUT2_reg[32]  ( .D(n5827), .CK(CLK), .Q(n4288) );
  DFF_X1 \OUT2_tri_enable_reg[32]  ( .D(n19486), .CK(CLK), .Q(n4289), .QN(
        n18910) );
  DFF_X1 \OUT2_reg[31]  ( .D(n5825), .CK(CLK), .Q(n4290) );
  DFF_X1 \OUT2_tri_enable_reg[31]  ( .D(n19485), .CK(CLK), .Q(n4291), .QN(
        n18927) );
  DFF_X1 \OUT2_reg[30]  ( .D(n5823), .CK(CLK), .Q(n4292) );
  DFF_X1 \OUT2_tri_enable_reg[30]  ( .D(n19484), .CK(CLK), .Q(n4293), .QN(
        n18944) );
  DFF_X1 \OUT2_reg[29]  ( .D(n5821), .CK(CLK), .Q(n4294) );
  DFF_X1 \OUT2_tri_enable_reg[29]  ( .D(n19483), .CK(CLK), .Q(n4295), .QN(
        n18961) );
  DFF_X1 \OUT2_reg[28]  ( .D(n5819), .CK(CLK), .Q(n4296) );
  DFF_X1 \OUT2_tri_enable_reg[28]  ( .D(n19482), .CK(CLK), .Q(n4297), .QN(
        n18978) );
  DFF_X1 \OUT2_reg[27]  ( .D(n5817), .CK(CLK), .Q(n4298) );
  DFF_X1 \OUT2_tri_enable_reg[27]  ( .D(n19481), .CK(CLK), .Q(n4299), .QN(
        n18995) );
  DFF_X1 \OUT2_reg[26]  ( .D(n5815), .CK(CLK), .Q(n4300) );
  DFF_X1 \OUT2_tri_enable_reg[26]  ( .D(n19480), .CK(CLK), .Q(n4301), .QN(
        n19012) );
  DFF_X1 \OUT2_reg[25]  ( .D(n5813), .CK(CLK), .Q(n4302) );
  DFF_X1 \OUT2_tri_enable_reg[25]  ( .D(n19479), .CK(CLK), .Q(n4303), .QN(
        n19029) );
  DFF_X1 \OUT2_reg[24]  ( .D(n5811), .CK(CLK), .Q(n4304) );
  DFF_X1 \OUT2_tri_enable_reg[24]  ( .D(n19478), .CK(CLK), .Q(n4305), .QN(
        n19046) );
  DFF_X1 \OUT2_reg[23]  ( .D(n5809), .CK(CLK), .Q(n4306) );
  DFF_X1 \OUT2_tri_enable_reg[23]  ( .D(n19477), .CK(CLK), .Q(n4307), .QN(
        n19063) );
  DFF_X1 \OUT2_reg[22]  ( .D(n5807), .CK(CLK), .Q(n4308) );
  DFF_X1 \OUT2_tri_enable_reg[22]  ( .D(n19476), .CK(CLK), .Q(n4309), .QN(
        n19080) );
  DFF_X1 \OUT2_reg[21]  ( .D(n5805), .CK(CLK), .Q(n4310) );
  DFF_X1 \OUT2_tri_enable_reg[21]  ( .D(n19475), .CK(CLK), .Q(n4311), .QN(
        n19097) );
  DFF_X1 \OUT2_reg[20]  ( .D(n5803), .CK(CLK), .Q(n4312) );
  DFF_X1 \OUT2_tri_enable_reg[20]  ( .D(n19474), .CK(CLK), .Q(n4313), .QN(
        n19114) );
  DFF_X1 \OUT2_reg[19]  ( .D(n5801), .CK(CLK), .Q(n4314) );
  DFF_X1 \OUT2_tri_enable_reg[19]  ( .D(n19473), .CK(CLK), .Q(n4315), .QN(
        n19131) );
  DFF_X1 \OUT2_reg[18]  ( .D(n5799), .CK(CLK), .Q(n4316) );
  DFF_X1 \OUT2_tri_enable_reg[18]  ( .D(n19472), .CK(CLK), .Q(n4317), .QN(
        n19148) );
  DFF_X1 \OUT2_reg[17]  ( .D(n5797), .CK(CLK), .Q(n4318) );
  DFF_X1 \OUT2_tri_enable_reg[17]  ( .D(n19471), .CK(CLK), .Q(n4319), .QN(
        n19165) );
  DFF_X1 \OUT2_reg[16]  ( .D(n5795), .CK(CLK), .Q(n4320) );
  DFF_X1 \OUT2_tri_enable_reg[16]  ( .D(n19470), .CK(CLK), .Q(n4321), .QN(
        n19182) );
  DFF_X1 \OUT2_reg[15]  ( .D(n5793), .CK(CLK), .Q(n4322) );
  DFF_X1 \OUT2_tri_enable_reg[15]  ( .D(n19469), .CK(CLK), .Q(n4323), .QN(
        n19199) );
  DFF_X1 \OUT2_reg[14]  ( .D(n5791), .CK(CLK), .Q(n4324) );
  DFF_X1 \OUT2_tri_enable_reg[14]  ( .D(n19468), .CK(CLK), .Q(n4325), .QN(
        n19216) );
  DFF_X1 \OUT2_reg[13]  ( .D(n5789), .CK(CLK), .Q(n4326) );
  DFF_X1 \OUT2_tri_enable_reg[13]  ( .D(n19467), .CK(CLK), .Q(n4327), .QN(
        n19233) );
  DFF_X1 \OUT2_reg[12]  ( .D(n5787), .CK(CLK), .Q(n4328) );
  DFF_X1 \OUT2_tri_enable_reg[12]  ( .D(n19466), .CK(CLK), .Q(n4329), .QN(
        n19250) );
  DFF_X1 \OUT2_reg[11]  ( .D(n5785), .CK(CLK), .Q(n4330) );
  DFF_X1 \OUT2_tri_enable_reg[11]  ( .D(n19465), .CK(CLK), .Q(n4331), .QN(
        n19267) );
  DFF_X1 \OUT2_reg[10]  ( .D(n5783), .CK(CLK), .Q(n4332) );
  DFF_X1 \OUT2_tri_enable_reg[10]  ( .D(n19464), .CK(CLK), .Q(n4333), .QN(
        n19284) );
  DFF_X1 \OUT2_reg[9]  ( .D(n5781), .CK(CLK), .Q(n4334) );
  DFF_X1 \OUT2_tri_enable_reg[9]  ( .D(n19463), .CK(CLK), .Q(n4335), .QN(
        n19301) );
  DFF_X1 \OUT2_reg[8]  ( .D(n5779), .CK(CLK), .Q(n4336) );
  DFF_X1 \OUT2_tri_enable_reg[8]  ( .D(n19462), .CK(CLK), .Q(n4337), .QN(
        n19318) );
  DFF_X1 \OUT2_reg[7]  ( .D(n5777), .CK(CLK), .Q(n4338) );
  DFF_X1 \OUT2_tri_enable_reg[7]  ( .D(n19461), .CK(CLK), .Q(n4339), .QN(
        n19335) );
  DFF_X1 \OUT2_reg[6]  ( .D(n5775), .CK(CLK), .Q(n4340) );
  DFF_X1 \OUT2_tri_enable_reg[6]  ( .D(n19460), .CK(CLK), .Q(n4341), .QN(
        n19352) );
  DFF_X1 \OUT2_reg[5]  ( .D(n5773), .CK(CLK), .Q(n4342) );
  DFF_X1 \OUT2_tri_enable_reg[5]  ( .D(n19459), .CK(CLK), .Q(n4343), .QN(
        n19369) );
  DFF_X1 \OUT2_reg[4]  ( .D(n5771), .CK(CLK), .Q(n4344) );
  DFF_X1 \OUT2_tri_enable_reg[4]  ( .D(n19458), .CK(CLK), .Q(n4345), .QN(
        n19386) );
  DFF_X1 \OUT2_reg[3]  ( .D(n5769), .CK(CLK), .Q(n4346) );
  DFF_X1 \OUT2_tri_enable_reg[3]  ( .D(n19457), .CK(CLK), .Q(n4347), .QN(
        n19403) );
  DFF_X1 \OUT2_reg[2]  ( .D(n5767), .CK(CLK), .Q(n4348) );
  DFF_X1 \OUT2_tri_enable_reg[2]  ( .D(n19456), .CK(CLK), .Q(n4349), .QN(
        n19420) );
  DFF_X1 \OUT2_reg[1]  ( .D(n5765), .CK(CLK), .Q(n4350) );
  DFF_X1 \OUT2_tri_enable_reg[1]  ( .D(n19455), .CK(CLK), .Q(n4351), .QN(
        n19437) );
  DFF_X1 \OUT2_reg[0]  ( .D(n5763), .CK(CLK), .Q(n4352) );
  DFF_X1 \OUT2_tri_enable_reg[0]  ( .D(n19580), .CK(CLK), .Q(n4353), .QN(
        n19454) );
  DFF_X1 \REGISTERS_reg[20][62]  ( .D(n6784), .CK(CLK), .QN(n9570) );
  DFF_X1 \REGISTERS_reg[20][61]  ( .D(n6783), .CK(CLK), .QN(n9571) );
  DFF_X1 \REGISTERS_reg[20][60]  ( .D(n6782), .CK(CLK), .QN(n9572) );
  DFF_X1 \REGISTERS_reg[20][59]  ( .D(n6781), .CK(CLK), .QN(n9573) );
  DFF_X1 \REGISTERS_reg[20][58]  ( .D(n6780), .CK(CLK), .QN(n9574) );
  DFF_X1 \REGISTERS_reg[20][57]  ( .D(n6779), .CK(CLK), .QN(n9575) );
  DFF_X1 \REGISTERS_reg[20][56]  ( .D(n6778), .CK(CLK), .QN(n9576) );
  DFF_X1 \REGISTERS_reg[20][55]  ( .D(n6777), .CK(CLK), .QN(n9577) );
  DFF_X1 \REGISTERS_reg[20][54]  ( .D(n6776), .CK(CLK), .QN(n9578) );
  DFF_X1 \REGISTERS_reg[20][53]  ( .D(n6775), .CK(CLK), .QN(n9579) );
  DFF_X1 \REGISTERS_reg[20][52]  ( .D(n6774), .CK(CLK), .QN(n9580) );
  DFF_X1 \REGISTERS_reg[20][51]  ( .D(n6773), .CK(CLK), .QN(n9581) );
  DFF_X1 \REGISTERS_reg[20][50]  ( .D(n6772), .CK(CLK), .QN(n9582) );
  DFF_X1 \REGISTERS_reg[20][49]  ( .D(n6771), .CK(CLK), .QN(n9583) );
  DFF_X1 \REGISTERS_reg[20][48]  ( .D(n6770), .CK(CLK), .QN(n9584) );
  DFF_X1 \REGISTERS_reg[20][47]  ( .D(n6769), .CK(CLK), .QN(n9585) );
  DFF_X1 \REGISTERS_reg[20][46]  ( .D(n6768), .CK(CLK), .QN(n9586) );
  DFF_X1 \REGISTERS_reg[20][45]  ( .D(n6767), .CK(CLK), .QN(n9587) );
  DFF_X1 \REGISTERS_reg[20][44]  ( .D(n6766), .CK(CLK), .QN(n9588) );
  DFF_X1 \REGISTERS_reg[20][43]  ( .D(n6765), .CK(CLK), .QN(n9589) );
  DFF_X1 \REGISTERS_reg[20][42]  ( .D(n6764), .CK(CLK), .QN(n9590) );
  DFF_X1 \REGISTERS_reg[20][41]  ( .D(n6763), .CK(CLK), .QN(n9591) );
  DFF_X1 \REGISTERS_reg[20][40]  ( .D(n6762), .CK(CLK), .QN(n9592) );
  DFF_X1 \REGISTERS_reg[20][39]  ( .D(n6761), .CK(CLK), .QN(n9593) );
  DFF_X1 \REGISTERS_reg[20][38]  ( .D(n6760), .CK(CLK), .QN(n9594) );
  DFF_X1 \REGISTERS_reg[20][37]  ( .D(n6759), .CK(CLK), .QN(n9595) );
  DFF_X1 \REGISTERS_reg[20][36]  ( .D(n6758), .CK(CLK), .QN(n9596) );
  DFF_X1 \REGISTERS_reg[20][35]  ( .D(n6757), .CK(CLK), .QN(n9597) );
  DFF_X1 \REGISTERS_reg[20][34]  ( .D(n6756), .CK(CLK), .QN(n9598) );
  DFF_X1 \REGISTERS_reg[20][33]  ( .D(n6755), .CK(CLK), .QN(n9599) );
  DFF_X1 \REGISTERS_reg[20][32]  ( .D(n6754), .CK(CLK), .QN(n9600) );
  DFF_X1 \REGISTERS_reg[20][31]  ( .D(n6753), .CK(CLK), .QN(n9601) );
  DFF_X1 \REGISTERS_reg[20][30]  ( .D(n6752), .CK(CLK), .QN(n9602) );
  DFF_X1 \REGISTERS_reg[20][29]  ( .D(n6751), .CK(CLK), .QN(n9603) );
  DFF_X1 \REGISTERS_reg[20][28]  ( .D(n6750), .CK(CLK), .QN(n9604) );
  DFF_X1 \REGISTERS_reg[20][27]  ( .D(n6749), .CK(CLK), .QN(n9605) );
  DFF_X1 \REGISTERS_reg[20][26]  ( .D(n6748), .CK(CLK), .QN(n9606) );
  DFF_X1 \REGISTERS_reg[20][25]  ( .D(n6747), .CK(CLK), .QN(n9607) );
  DFF_X1 \REGISTERS_reg[20][24]  ( .D(n6746), .CK(CLK), .QN(n9608) );
  DFF_X1 \REGISTERS_reg[20][23]  ( .D(n6745), .CK(CLK), .QN(n9609) );
  DFF_X1 \REGISTERS_reg[20][22]  ( .D(n6744), .CK(CLK), .QN(n9610) );
  DFF_X1 \REGISTERS_reg[20][21]  ( .D(n6743), .CK(CLK), .QN(n9611) );
  DFF_X1 \REGISTERS_reg[20][20]  ( .D(n6742), .CK(CLK), .QN(n9612) );
  DFF_X1 \REGISTERS_reg[20][19]  ( .D(n6741), .CK(CLK), .QN(n9613) );
  DFF_X1 \REGISTERS_reg[20][18]  ( .D(n6740), .CK(CLK), .QN(n9614) );
  DFF_X1 \REGISTERS_reg[20][17]  ( .D(n6739), .CK(CLK), .QN(n9615) );
  DFF_X1 \REGISTERS_reg[20][16]  ( .D(n6738), .CK(CLK), .QN(n9616) );
  DFF_X1 \REGISTERS_reg[20][15]  ( .D(n6737), .CK(CLK), .QN(n9617) );
  DFF_X1 \REGISTERS_reg[20][14]  ( .D(n6736), .CK(CLK), .QN(n9618) );
  DFF_X1 \REGISTERS_reg[20][13]  ( .D(n6735), .CK(CLK), .QN(n9619) );
  DFF_X1 \REGISTERS_reg[20][12]  ( .D(n6734), .CK(CLK), .QN(n9620) );
  DFF_X1 \REGISTERS_reg[20][11]  ( .D(n6733), .CK(CLK), .QN(n9621) );
  DFF_X1 \REGISTERS_reg[20][10]  ( .D(n6732), .CK(CLK), .QN(n9622) );
  DFF_X1 \REGISTERS_reg[20][9]  ( .D(n6731), .CK(CLK), .QN(n9623) );
  DFF_X1 \REGISTERS_reg[20][8]  ( .D(n6730), .CK(CLK), .QN(n9624) );
  DFF_X1 \REGISTERS_reg[20][7]  ( .D(n6729), .CK(CLK), .QN(n9625) );
  DFF_X1 \REGISTERS_reg[20][6]  ( .D(n6728), .CK(CLK), .QN(n9626) );
  DFF_X1 \REGISTERS_reg[20][5]  ( .D(n6727), .CK(CLK), .QN(n9627) );
  DFF_X1 \REGISTERS_reg[20][4]  ( .D(n6726), .CK(CLK), .QN(n9628) );
  DFF_X1 \REGISTERS_reg[20][3]  ( .D(n6725), .CK(CLK), .QN(n9629) );
  DFF_X1 \REGISTERS_reg[20][2]  ( .D(n6724), .CK(CLK), .QN(n9630) );
  DFF_X1 \REGISTERS_reg[20][1]  ( .D(n6723), .CK(CLK), .QN(n9631) );
  DFF_X1 \REGISTERS_reg[20][0]  ( .D(n6722), .CK(CLK), .QN(n9632) );
  NAND3_X1 U19260 ( .A1(ADD_RD1[1]), .A2(n20636), .A3(n23966), .ZN(n22811) );
  NAND3_X1 U19261 ( .A1(ADD_RD1[2]), .A2(n20637), .A3(n23966), .ZN(n22810) );
  NAND3_X1 U19262 ( .A1(ADD_RD1[2]), .A2(ADD_RD1[1]), .A3(n23966), .ZN(n22815)
         );
  NAND3_X1 U19263 ( .A1(ADD_RD2[1]), .A2(n20641), .A3(n25165), .ZN(n24010) );
  NAND3_X1 U19264 ( .A1(ADD_RD2[2]), .A2(n20642), .A3(n25165), .ZN(n24009) );
  NAND3_X1 U19265 ( .A1(ADD_RD2[2]), .A2(ADD_RD2[1]), .A3(n25165), .ZN(n24014)
         );
  TBUF_X1 \OUT2_tri[0]  ( .A(n4352), .EN(n4353), .Z(OUT2[0]) );
  TBUF_X1 \OUT2_tri[1]  ( .A(n4350), .EN(n4351), .Z(OUT2[1]) );
  TBUF_X1 \OUT2_tri[2]  ( .A(n4348), .EN(n4349), .Z(OUT2[2]) );
  TBUF_X1 \OUT2_tri[3]  ( .A(n4346), .EN(n4347), .Z(OUT2[3]) );
  TBUF_X1 \OUT2_tri[4]  ( .A(n4344), .EN(n4345), .Z(OUT2[4]) );
  TBUF_X1 \OUT2_tri[5]  ( .A(n4342), .EN(n4343), .Z(OUT2[5]) );
  TBUF_X1 \OUT2_tri[6]  ( .A(n4340), .EN(n4341), .Z(OUT2[6]) );
  TBUF_X1 \OUT2_tri[7]  ( .A(n4338), .EN(n4339), .Z(OUT2[7]) );
  TBUF_X1 \OUT2_tri[8]  ( .A(n4336), .EN(n4337), .Z(OUT2[8]) );
  TBUF_X1 \OUT2_tri[9]  ( .A(n4334), .EN(n4335), .Z(OUT2[9]) );
  TBUF_X1 \OUT2_tri[10]  ( .A(n4332), .EN(n4333), .Z(OUT2[10]) );
  TBUF_X1 \OUT2_tri[11]  ( .A(n4330), .EN(n4331), .Z(OUT2[11]) );
  TBUF_X1 \OUT2_tri[12]  ( .A(n4328), .EN(n4329), .Z(OUT2[12]) );
  TBUF_X1 \OUT2_tri[13]  ( .A(n4326), .EN(n4327), .Z(OUT2[13]) );
  TBUF_X1 \OUT2_tri[14]  ( .A(n4324), .EN(n4325), .Z(OUT2[14]) );
  TBUF_X1 \OUT2_tri[15]  ( .A(n4322), .EN(n4323), .Z(OUT2[15]) );
  TBUF_X1 \OUT2_tri[16]  ( .A(n4320), .EN(n4321), .Z(OUT2[16]) );
  TBUF_X1 \OUT2_tri[17]  ( .A(n4318), .EN(n4319), .Z(OUT2[17]) );
  TBUF_X1 \OUT2_tri[18]  ( .A(n4316), .EN(n4317), .Z(OUT2[18]) );
  TBUF_X1 \OUT2_tri[19]  ( .A(n4314), .EN(n4315), .Z(OUT2[19]) );
  TBUF_X1 \OUT2_tri[20]  ( .A(n4312), .EN(n4313), .Z(OUT2[20]) );
  TBUF_X1 \OUT2_tri[21]  ( .A(n4310), .EN(n4311), .Z(OUT2[21]) );
  TBUF_X1 \OUT2_tri[22]  ( .A(n4308), .EN(n4309), .Z(OUT2[22]) );
  TBUF_X1 \OUT2_tri[23]  ( .A(n4306), .EN(n4307), .Z(OUT2[23]) );
  TBUF_X1 \OUT2_tri[24]  ( .A(n4304), .EN(n4305), .Z(OUT2[24]) );
  TBUF_X1 \OUT2_tri[25]  ( .A(n4302), .EN(n4303), .Z(OUT2[25]) );
  TBUF_X1 \OUT2_tri[26]  ( .A(n4300), .EN(n4301), .Z(OUT2[26]) );
  TBUF_X1 \OUT2_tri[27]  ( .A(n4298), .EN(n4299), .Z(OUT2[27]) );
  TBUF_X1 \OUT2_tri[28]  ( .A(n4296), .EN(n4297), .Z(OUT2[28]) );
  TBUF_X1 \OUT2_tri[29]  ( .A(n4294), .EN(n4295), .Z(OUT2[29]) );
  TBUF_X1 \OUT2_tri[30]  ( .A(n4292), .EN(n4293), .Z(OUT2[30]) );
  TBUF_X1 \OUT2_tri[31]  ( .A(n4290), .EN(n4291), .Z(OUT2[31]) );
  TBUF_X1 \OUT2_tri[32]  ( .A(n4288), .EN(n4289), .Z(OUT2[32]) );
  TBUF_X1 \OUT2_tri[33]  ( .A(n4286), .EN(n4287), .Z(OUT2[33]) );
  TBUF_X1 \OUT2_tri[34]  ( .A(n4284), .EN(n4285), .Z(OUT2[34]) );
  TBUF_X1 \OUT2_tri[35]  ( .A(n4282), .EN(n4283), .Z(OUT2[35]) );
  TBUF_X1 \OUT2_tri[36]  ( .A(n4280), .EN(n4281), .Z(OUT2[36]) );
  TBUF_X1 \OUT2_tri[37]  ( .A(n4278), .EN(n4279), .Z(OUT2[37]) );
  TBUF_X1 \OUT2_tri[38]  ( .A(n4276), .EN(n4277), .Z(OUT2[38]) );
  TBUF_X1 \OUT2_tri[39]  ( .A(n4274), .EN(n4275), .Z(OUT2[39]) );
  TBUF_X1 \OUT2_tri[40]  ( .A(n4272), .EN(n4273), .Z(OUT2[40]) );
  TBUF_X1 \OUT2_tri[41]  ( .A(n4270), .EN(n4271), .Z(OUT2[41]) );
  TBUF_X1 \OUT2_tri[42]  ( .A(n4268), .EN(n4269), .Z(OUT2[42]) );
  TBUF_X1 \OUT2_tri[43]  ( .A(n4266), .EN(n4267), .Z(OUT2[43]) );
  TBUF_X1 \OUT2_tri[44]  ( .A(n4264), .EN(n4265), .Z(OUT2[44]) );
  TBUF_X1 \OUT2_tri[45]  ( .A(n4262), .EN(n4263), .Z(OUT2[45]) );
  TBUF_X1 \OUT2_tri[46]  ( .A(n4260), .EN(n4261), .Z(OUT2[46]) );
  TBUF_X1 \OUT2_tri[47]  ( .A(n4258), .EN(n4259), .Z(OUT2[47]) );
  TBUF_X1 \OUT2_tri[48]  ( .A(n4256), .EN(n4257), .Z(OUT2[48]) );
  TBUF_X1 \OUT2_tri[49]  ( .A(n4254), .EN(n4255), .Z(OUT2[49]) );
  TBUF_X1 \OUT2_tri[50]  ( .A(n4252), .EN(n4253), .Z(OUT2[50]) );
  TBUF_X1 \OUT2_tri[51]  ( .A(n4250), .EN(n4251), .Z(OUT2[51]) );
  TBUF_X1 \OUT2_tri[52]  ( .A(n4248), .EN(n4249), .Z(OUT2[52]) );
  TBUF_X1 \OUT2_tri[53]  ( .A(n4246), .EN(n4247), .Z(OUT2[53]) );
  TBUF_X1 \OUT2_tri[54]  ( .A(n4244), .EN(n4245), .Z(OUT2[54]) );
  TBUF_X1 \OUT2_tri[55]  ( .A(n4242), .EN(n4243), .Z(OUT2[55]) );
  TBUF_X1 \OUT2_tri[56]  ( .A(n4240), .EN(n4241), .Z(OUT2[56]) );
  TBUF_X1 \OUT2_tri[57]  ( .A(n4238), .EN(n4239), .Z(OUT2[57]) );
  TBUF_X1 \OUT2_tri[58]  ( .A(n4236), .EN(n4237), .Z(OUT2[58]) );
  TBUF_X1 \OUT2_tri[59]  ( .A(n4234), .EN(n4235), .Z(OUT2[59]) );
  TBUF_X1 \OUT2_tri[60]  ( .A(n4232), .EN(n4233), .Z(OUT2[60]) );
  TBUF_X1 \OUT2_tri[61]  ( .A(n4230), .EN(n4231), .Z(OUT2[61]) );
  TBUF_X1 \OUT2_tri[62]  ( .A(n4228), .EN(n4229), .Z(OUT2[62]) );
  TBUF_X1 \OUT2_tri[63]  ( .A(n4226), .EN(n4227), .Z(OUT2[63]) );
  TBUF_X1 \OUT1_tri[0]  ( .A(n4224), .EN(n4225), .Z(OUT1[0]) );
  TBUF_X1 \OUT1_tri[1]  ( .A(n4222), .EN(n4223), .Z(OUT1[1]) );
  TBUF_X1 \OUT1_tri[2]  ( .A(n4220), .EN(n4221), .Z(OUT1[2]) );
  TBUF_X1 \OUT1_tri[3]  ( .A(n4218), .EN(n4219), .Z(OUT1[3]) );
  TBUF_X1 \OUT1_tri[4]  ( .A(n4216), .EN(n4217), .Z(OUT1[4]) );
  TBUF_X1 \OUT1_tri[5]  ( .A(n4214), .EN(n4215), .Z(OUT1[5]) );
  TBUF_X1 \OUT1_tri[6]  ( .A(n4212), .EN(n4213), .Z(OUT1[6]) );
  TBUF_X1 \OUT1_tri[7]  ( .A(n4210), .EN(n4211), .Z(OUT1[7]) );
  TBUF_X1 \OUT1_tri[8]  ( .A(n4208), .EN(n4209), .Z(OUT1[8]) );
  TBUF_X1 \OUT1_tri[9]  ( .A(n4206), .EN(n4207), .Z(OUT1[9]) );
  TBUF_X1 \OUT1_tri[10]  ( .A(n4204), .EN(n4205), .Z(OUT1[10]) );
  TBUF_X1 \OUT1_tri[11]  ( .A(n4202), .EN(n4203), .Z(OUT1[11]) );
  TBUF_X1 \OUT1_tri[12]  ( .A(n4200), .EN(n4201), .Z(OUT1[12]) );
  TBUF_X1 \OUT1_tri[13]  ( .A(n4198), .EN(n4199), .Z(OUT1[13]) );
  TBUF_X1 \OUT1_tri[14]  ( .A(n4196), .EN(n4197), .Z(OUT1[14]) );
  TBUF_X1 \OUT1_tri[15]  ( .A(n4194), .EN(n4195), .Z(OUT1[15]) );
  TBUF_X1 \OUT1_tri[16]  ( .A(n4192), .EN(n4193), .Z(OUT1[16]) );
  TBUF_X1 \OUT1_tri[17]  ( .A(n4190), .EN(n4191), .Z(OUT1[17]) );
  TBUF_X1 \OUT1_tri[18]  ( .A(n4188), .EN(n4189), .Z(OUT1[18]) );
  TBUF_X1 \OUT1_tri[19]  ( .A(n4186), .EN(n4187), .Z(OUT1[19]) );
  TBUF_X1 \OUT1_tri[20]  ( .A(n4184), .EN(n4185), .Z(OUT1[20]) );
  TBUF_X1 \OUT1_tri[21]  ( .A(n4182), .EN(n4183), .Z(OUT1[21]) );
  TBUF_X1 \OUT1_tri[22]  ( .A(n4180), .EN(n4181), .Z(OUT1[22]) );
  TBUF_X1 \OUT1_tri[23]  ( .A(n4178), .EN(n4179), .Z(OUT1[23]) );
  TBUF_X1 \OUT1_tri[24]  ( .A(n4176), .EN(n4177), .Z(OUT1[24]) );
  TBUF_X1 \OUT1_tri[25]  ( .A(n4174), .EN(n4175), .Z(OUT1[25]) );
  TBUF_X1 \OUT1_tri[26]  ( .A(n4172), .EN(n4173), .Z(OUT1[26]) );
  TBUF_X1 \OUT1_tri[27]  ( .A(n4170), .EN(n4171), .Z(OUT1[27]) );
  TBUF_X1 \OUT1_tri[28]  ( .A(n4168), .EN(n4169), .Z(OUT1[28]) );
  TBUF_X1 \OUT1_tri[29]  ( .A(n4166), .EN(n4167), .Z(OUT1[29]) );
  TBUF_X1 \OUT1_tri[30]  ( .A(n4164), .EN(n4165), .Z(OUT1[30]) );
  TBUF_X1 \OUT1_tri[31]  ( .A(n4162), .EN(n4163), .Z(OUT1[31]) );
  TBUF_X1 \OUT1_tri[32]  ( .A(n4160), .EN(n4161), .Z(OUT1[32]) );
  TBUF_X1 \OUT1_tri[33]  ( .A(n4158), .EN(n4159), .Z(OUT1[33]) );
  TBUF_X1 \OUT1_tri[34]  ( .A(n4156), .EN(n4157), .Z(OUT1[34]) );
  TBUF_X1 \OUT1_tri[35]  ( .A(n4154), .EN(n4155), .Z(OUT1[35]) );
  TBUF_X1 \OUT1_tri[36]  ( .A(n4152), .EN(n4153), .Z(OUT1[36]) );
  TBUF_X1 \OUT1_tri[37]  ( .A(n4150), .EN(n4151), .Z(OUT1[37]) );
  TBUF_X1 \OUT1_tri[38]  ( .A(n4148), .EN(n4149), .Z(OUT1[38]) );
  TBUF_X1 \OUT1_tri[39]  ( .A(n4146), .EN(n4147), .Z(OUT1[39]) );
  TBUF_X1 \OUT1_tri[40]  ( .A(n4144), .EN(n4145), .Z(OUT1[40]) );
  TBUF_X1 \OUT1_tri[41]  ( .A(n4142), .EN(n4143), .Z(OUT1[41]) );
  TBUF_X1 \OUT1_tri[42]  ( .A(n4140), .EN(n4141), .Z(OUT1[42]) );
  TBUF_X1 \OUT1_tri[43]  ( .A(n4138), .EN(n4139), .Z(OUT1[43]) );
  TBUF_X1 \OUT1_tri[44]  ( .A(n4136), .EN(n4137), .Z(OUT1[44]) );
  TBUF_X1 \OUT1_tri[45]  ( .A(n4134), .EN(n4135), .Z(OUT1[45]) );
  TBUF_X1 \OUT1_tri[46]  ( .A(n4132), .EN(n4133), .Z(OUT1[46]) );
  TBUF_X1 \OUT1_tri[47]  ( .A(n4130), .EN(n4131), .Z(OUT1[47]) );
  TBUF_X1 \OUT1_tri[48]  ( .A(n4128), .EN(n4129), .Z(OUT1[48]) );
  TBUF_X1 \OUT1_tri[49]  ( .A(n4126), .EN(n4127), .Z(OUT1[49]) );
  TBUF_X1 \OUT1_tri[50]  ( .A(n4124), .EN(n4125), .Z(OUT1[50]) );
  TBUF_X1 \OUT1_tri[51]  ( .A(n4122), .EN(n4123), .Z(OUT1[51]) );
  TBUF_X1 \OUT1_tri[52]  ( .A(n4120), .EN(n4121), .Z(OUT1[52]) );
  TBUF_X1 \OUT1_tri[53]  ( .A(n4118), .EN(n4119), .Z(OUT1[53]) );
  TBUF_X1 \OUT1_tri[54]  ( .A(n4116), .EN(n4117), .Z(OUT1[54]) );
  TBUF_X1 \OUT1_tri[55]  ( .A(n4114), .EN(n4115), .Z(OUT1[55]) );
  TBUF_X1 \OUT1_tri[56]  ( .A(n4112), .EN(n4113), .Z(OUT1[56]) );
  TBUF_X1 \OUT1_tri[57]  ( .A(n4110), .EN(n4111), .Z(OUT1[57]) );
  TBUF_X1 \OUT1_tri[58]  ( .A(n4108), .EN(n4109), .Z(OUT1[58]) );
  TBUF_X1 \OUT1_tri[59]  ( .A(n4106), .EN(n4107), .Z(OUT1[59]) );
  TBUF_X1 \OUT1_tri[60]  ( .A(n4104), .EN(n4105), .Z(OUT1[60]) );
  TBUF_X1 \OUT1_tri[61]  ( .A(n4102), .EN(n4103), .Z(OUT1[61]) );
  TBUF_X1 \OUT1_tri[62]  ( .A(n4100), .EN(n4101), .Z(OUT1[62]) );
  TBUF_X1 \OUT1_tri[63]  ( .A(n4098), .EN(n4099), .Z(OUT1[63]) );
  DFF_X1 \REGISTERS_reg[21][63]  ( .D(n6721), .CK(CLK), .Q(n20963), .QN(n9633)
         );
  DFF_X1 \REGISTERS_reg[21][62]  ( .D(n6720), .CK(CLK), .Q(n20964), .QN(n9634)
         );
  DFF_X1 \REGISTERS_reg[21][61]  ( .D(n6719), .CK(CLK), .Q(n20965), .QN(n9635)
         );
  DFF_X1 \REGISTERS_reg[21][60]  ( .D(n6718), .CK(CLK), .Q(n20966), .QN(n9636)
         );
  DFF_X1 \REGISTERS_reg[15][63]  ( .D(n7105), .CK(CLK), .Q(n20967), .QN(n9505)
         );
  DFF_X1 \REGISTERS_reg[15][62]  ( .D(n7104), .CK(CLK), .Q(n20968), .QN(n9506)
         );
  DFF_X1 \REGISTERS_reg[15][61]  ( .D(n7103), .CK(CLK), .Q(n20969), .QN(n9507)
         );
  DFF_X1 \REGISTERS_reg[15][60]  ( .D(n7102), .CK(CLK), .Q(n20970), .QN(n9508)
         );
  DFF_X1 \REGISTERS_reg[13][63]  ( .D(n7233), .CK(CLK), .Q(n20971), .QN(n9697)
         );
  DFF_X1 \REGISTERS_reg[13][62]  ( .D(n7232), .CK(CLK), .Q(n20972), .QN(n9698)
         );
  DFF_X1 \REGISTERS_reg[13][61]  ( .D(n7231), .CK(CLK), .Q(n20973), .QN(n9699)
         );
  DFF_X1 \REGISTERS_reg[13][60]  ( .D(n7230), .CK(CLK), .Q(n20974), .QN(n9700)
         );
  DFF_X1 \REGISTERS_reg[21][59]  ( .D(n6717), .CK(CLK), .Q(n20975), .QN(n9637)
         );
  DFF_X1 \REGISTERS_reg[21][58]  ( .D(n6716), .CK(CLK), .Q(n20976), .QN(n9638)
         );
  DFF_X1 \REGISTERS_reg[21][57]  ( .D(n6715), .CK(CLK), .Q(n20977), .QN(n9639)
         );
  DFF_X1 \REGISTERS_reg[21][56]  ( .D(n6714), .CK(CLK), .Q(n20978), .QN(n9640)
         );
  DFF_X1 \REGISTERS_reg[21][55]  ( .D(n6713), .CK(CLK), .Q(n20979), .QN(n9641)
         );
  DFF_X1 \REGISTERS_reg[21][54]  ( .D(n6712), .CK(CLK), .Q(n20980), .QN(n9642)
         );
  DFF_X1 \REGISTERS_reg[21][53]  ( .D(n6711), .CK(CLK), .Q(n20981), .QN(n9643)
         );
  DFF_X1 \REGISTERS_reg[21][52]  ( .D(n6710), .CK(CLK), .Q(n20982), .QN(n9644)
         );
  DFF_X1 \REGISTERS_reg[21][51]  ( .D(n6709), .CK(CLK), .Q(n20983), .QN(n9645)
         );
  DFF_X1 \REGISTERS_reg[21][50]  ( .D(n6708), .CK(CLK), .Q(n20984), .QN(n9646)
         );
  DFF_X1 \REGISTERS_reg[21][49]  ( .D(n6707), .CK(CLK), .Q(n20985), .QN(n9647)
         );
  DFF_X1 \REGISTERS_reg[21][48]  ( .D(n6706), .CK(CLK), .Q(n20986), .QN(n9648)
         );
  DFF_X1 \REGISTERS_reg[21][47]  ( .D(n6705), .CK(CLK), .Q(n20987), .QN(n9649)
         );
  DFF_X1 \REGISTERS_reg[21][46]  ( .D(n6704), .CK(CLK), .Q(n20988), .QN(n9650)
         );
  DFF_X1 \REGISTERS_reg[21][45]  ( .D(n6703), .CK(CLK), .Q(n20989), .QN(n9651)
         );
  DFF_X1 \REGISTERS_reg[21][44]  ( .D(n6702), .CK(CLK), .Q(n20990), .QN(n9652)
         );
  DFF_X1 \REGISTERS_reg[21][43]  ( .D(n6701), .CK(CLK), .Q(n20991), .QN(n9653)
         );
  DFF_X1 \REGISTERS_reg[21][42]  ( .D(n6700), .CK(CLK), .Q(n20992), .QN(n9654)
         );
  DFF_X1 \REGISTERS_reg[21][41]  ( .D(n6699), .CK(CLK), .Q(n20993), .QN(n9655)
         );
  DFF_X1 \REGISTERS_reg[21][40]  ( .D(n6698), .CK(CLK), .Q(n20994), .QN(n9656)
         );
  DFF_X1 \REGISTERS_reg[21][39]  ( .D(n6697), .CK(CLK), .Q(n20995), .QN(n9657)
         );
  DFF_X1 \REGISTERS_reg[21][38]  ( .D(n6696), .CK(CLK), .Q(n20996), .QN(n9658)
         );
  DFF_X1 \REGISTERS_reg[21][37]  ( .D(n6695), .CK(CLK), .Q(n20997), .QN(n9659)
         );
  DFF_X1 \REGISTERS_reg[21][36]  ( .D(n6694), .CK(CLK), .Q(n20998), .QN(n9660)
         );
  DFF_X1 \REGISTERS_reg[21][35]  ( .D(n6693), .CK(CLK), .Q(n20999), .QN(n9661)
         );
  DFF_X1 \REGISTERS_reg[21][34]  ( .D(n6692), .CK(CLK), .Q(n21000), .QN(n9662)
         );
  DFF_X1 \REGISTERS_reg[21][33]  ( .D(n6691), .CK(CLK), .Q(n21001), .QN(n9663)
         );
  DFF_X1 \REGISTERS_reg[21][32]  ( .D(n6690), .CK(CLK), .Q(n21002), .QN(n9664)
         );
  DFF_X1 \REGISTERS_reg[21][31]  ( .D(n6689), .CK(CLK), .Q(n21003), .QN(n9665)
         );
  DFF_X1 \REGISTERS_reg[21][30]  ( .D(n6688), .CK(CLK), .Q(n21004), .QN(n9666)
         );
  DFF_X1 \REGISTERS_reg[21][29]  ( .D(n6687), .CK(CLK), .Q(n21005), .QN(n9667)
         );
  DFF_X1 \REGISTERS_reg[21][28]  ( .D(n6686), .CK(CLK), .Q(n21006), .QN(n9668)
         );
  DFF_X1 \REGISTERS_reg[21][27]  ( .D(n6685), .CK(CLK), .Q(n21007), .QN(n9669)
         );
  DFF_X1 \REGISTERS_reg[21][26]  ( .D(n6684), .CK(CLK), .Q(n21008), .QN(n9670)
         );
  DFF_X1 \REGISTERS_reg[21][25]  ( .D(n6683), .CK(CLK), .Q(n21009), .QN(n9671)
         );
  DFF_X1 \REGISTERS_reg[21][24]  ( .D(n6682), .CK(CLK), .Q(n21010), .QN(n9672)
         );
  DFF_X1 \REGISTERS_reg[21][23]  ( .D(n6681), .CK(CLK), .Q(n21011), .QN(n9673)
         );
  DFF_X1 \REGISTERS_reg[21][22]  ( .D(n6680), .CK(CLK), .Q(n21012), .QN(n9674)
         );
  DFF_X1 \REGISTERS_reg[21][21]  ( .D(n6679), .CK(CLK), .Q(n21013), .QN(n9675)
         );
  DFF_X1 \REGISTERS_reg[21][20]  ( .D(n6678), .CK(CLK), .Q(n21014), .QN(n9676)
         );
  DFF_X1 \REGISTERS_reg[21][19]  ( .D(n6677), .CK(CLK), .Q(n21015), .QN(n9677)
         );
  DFF_X1 \REGISTERS_reg[21][18]  ( .D(n6676), .CK(CLK), .Q(n21016), .QN(n9678)
         );
  DFF_X1 \REGISTERS_reg[21][17]  ( .D(n6675), .CK(CLK), .Q(n21017), .QN(n9679)
         );
  DFF_X1 \REGISTERS_reg[21][16]  ( .D(n6674), .CK(CLK), .Q(n21018), .QN(n9680)
         );
  DFF_X1 \REGISTERS_reg[21][15]  ( .D(n6673), .CK(CLK), .Q(n21019), .QN(n9681)
         );
  DFF_X1 \REGISTERS_reg[21][14]  ( .D(n6672), .CK(CLK), .Q(n21020), .QN(n9682)
         );
  DFF_X1 \REGISTERS_reg[21][13]  ( .D(n6671), .CK(CLK), .Q(n21021), .QN(n9683)
         );
  DFF_X1 \REGISTERS_reg[21][12]  ( .D(n6670), .CK(CLK), .Q(n21022), .QN(n9684)
         );
  DFF_X1 \REGISTERS_reg[21][11]  ( .D(n6669), .CK(CLK), .Q(n21023), .QN(n9685)
         );
  DFF_X1 \REGISTERS_reg[21][10]  ( .D(n6668), .CK(CLK), .Q(n21024), .QN(n9686)
         );
  DFF_X1 \REGISTERS_reg[21][9]  ( .D(n6667), .CK(CLK), .Q(n21025), .QN(n9687)
         );
  DFF_X1 \REGISTERS_reg[21][8]  ( .D(n6666), .CK(CLK), .Q(n21026), .QN(n9688)
         );
  DFF_X1 \REGISTERS_reg[21][7]  ( .D(n6665), .CK(CLK), .Q(n21027), .QN(n9689)
         );
  DFF_X1 \REGISTERS_reg[21][6]  ( .D(n6664), .CK(CLK), .Q(n21028), .QN(n9690)
         );
  DFF_X1 \REGISTERS_reg[21][5]  ( .D(n6663), .CK(CLK), .Q(n21029), .QN(n9691)
         );
  DFF_X1 \REGISTERS_reg[21][4]  ( .D(n6662), .CK(CLK), .Q(n21030), .QN(n9692)
         );
  DFF_X1 \REGISTERS_reg[21][3]  ( .D(n6661), .CK(CLK), .Q(n21031), .QN(n9693)
         );
  DFF_X1 \REGISTERS_reg[21][2]  ( .D(n6660), .CK(CLK), .Q(n21032), .QN(n9694)
         );
  DFF_X1 \REGISTERS_reg[21][1]  ( .D(n6659), .CK(CLK), .Q(n21033), .QN(n9695)
         );
  DFF_X1 \REGISTERS_reg[21][0]  ( .D(n6658), .CK(CLK), .Q(n21034), .QN(n9696)
         );
  DFF_X1 \REGISTERS_reg[15][59]  ( .D(n7101), .CK(CLK), .Q(n21035), .QN(n9509)
         );
  DFF_X1 \REGISTERS_reg[15][58]  ( .D(n7100), .CK(CLK), .Q(n21036), .QN(n9510)
         );
  DFF_X1 \REGISTERS_reg[15][57]  ( .D(n7099), .CK(CLK), .Q(n21037), .QN(n9511)
         );
  DFF_X1 \REGISTERS_reg[15][56]  ( .D(n7098), .CK(CLK), .Q(n21038), .QN(n9512)
         );
  DFF_X1 \REGISTERS_reg[15][55]  ( .D(n7097), .CK(CLK), .Q(n21039), .QN(n9513)
         );
  DFF_X1 \REGISTERS_reg[15][54]  ( .D(n7096), .CK(CLK), .Q(n21040), .QN(n9514)
         );
  DFF_X1 \REGISTERS_reg[15][53]  ( .D(n7095), .CK(CLK), .Q(n21041), .QN(n9515)
         );
  DFF_X1 \REGISTERS_reg[15][52]  ( .D(n7094), .CK(CLK), .Q(n21042), .QN(n9516)
         );
  DFF_X1 \REGISTERS_reg[15][51]  ( .D(n7093), .CK(CLK), .Q(n21043), .QN(n9517)
         );
  DFF_X1 \REGISTERS_reg[15][50]  ( .D(n7092), .CK(CLK), .Q(n21044), .QN(n9518)
         );
  DFF_X1 \REGISTERS_reg[15][49]  ( .D(n7091), .CK(CLK), .Q(n21045), .QN(n9519)
         );
  DFF_X1 \REGISTERS_reg[15][48]  ( .D(n7090), .CK(CLK), .Q(n21046), .QN(n9520)
         );
  DFF_X1 \REGISTERS_reg[15][47]  ( .D(n7089), .CK(CLK), .Q(n21047), .QN(n9521)
         );
  DFF_X1 \REGISTERS_reg[15][46]  ( .D(n7088), .CK(CLK), .Q(n21048), .QN(n9522)
         );
  DFF_X1 \REGISTERS_reg[15][45]  ( .D(n7087), .CK(CLK), .Q(n21049), .QN(n9523)
         );
  DFF_X1 \REGISTERS_reg[15][44]  ( .D(n7086), .CK(CLK), .Q(n21050), .QN(n9524)
         );
  DFF_X1 \REGISTERS_reg[15][43]  ( .D(n7085), .CK(CLK), .Q(n21051), .QN(n9525)
         );
  DFF_X1 \REGISTERS_reg[15][42]  ( .D(n7084), .CK(CLK), .Q(n21052), .QN(n9526)
         );
  DFF_X1 \REGISTERS_reg[15][41]  ( .D(n7083), .CK(CLK), .Q(n21053), .QN(n9527)
         );
  DFF_X1 \REGISTERS_reg[15][40]  ( .D(n7082), .CK(CLK), .Q(n21054), .QN(n9528)
         );
  DFF_X1 \REGISTERS_reg[15][39]  ( .D(n7081), .CK(CLK), .Q(n21055), .QN(n9529)
         );
  DFF_X1 \REGISTERS_reg[15][38]  ( .D(n7080), .CK(CLK), .Q(n21056), .QN(n9530)
         );
  DFF_X1 \REGISTERS_reg[15][37]  ( .D(n7079), .CK(CLK), .Q(n21057), .QN(n9531)
         );
  DFF_X1 \REGISTERS_reg[15][36]  ( .D(n7078), .CK(CLK), .Q(n21058), .QN(n9532)
         );
  DFF_X1 \REGISTERS_reg[15][35]  ( .D(n7077), .CK(CLK), .Q(n21059), .QN(n9533)
         );
  DFF_X1 \REGISTERS_reg[15][34]  ( .D(n7076), .CK(CLK), .Q(n21060), .QN(n9534)
         );
  DFF_X1 \REGISTERS_reg[15][33]  ( .D(n7075), .CK(CLK), .Q(n21061), .QN(n9535)
         );
  DFF_X1 \REGISTERS_reg[15][32]  ( .D(n7074), .CK(CLK), .Q(n21062), .QN(n9536)
         );
  DFF_X1 \REGISTERS_reg[15][31]  ( .D(n7073), .CK(CLK), .Q(n21063), .QN(n9537)
         );
  DFF_X1 \REGISTERS_reg[15][30]  ( .D(n7072), .CK(CLK), .Q(n21064), .QN(n9538)
         );
  DFF_X1 \REGISTERS_reg[15][29]  ( .D(n7071), .CK(CLK), .Q(n21065), .QN(n9539)
         );
  DFF_X1 \REGISTERS_reg[15][28]  ( .D(n7070), .CK(CLK), .Q(n21066), .QN(n9540)
         );
  DFF_X1 \REGISTERS_reg[15][27]  ( .D(n7069), .CK(CLK), .Q(n21067), .QN(n9541)
         );
  DFF_X1 \REGISTERS_reg[15][26]  ( .D(n7068), .CK(CLK), .Q(n21068), .QN(n9542)
         );
  DFF_X1 \REGISTERS_reg[15][25]  ( .D(n7067), .CK(CLK), .Q(n21069), .QN(n9543)
         );
  DFF_X1 \REGISTERS_reg[15][24]  ( .D(n7066), .CK(CLK), .Q(n21070), .QN(n9544)
         );
  DFF_X1 \REGISTERS_reg[15][23]  ( .D(n7065), .CK(CLK), .Q(n21071), .QN(n9545)
         );
  DFF_X1 \REGISTERS_reg[15][22]  ( .D(n7064), .CK(CLK), .Q(n21072), .QN(n9546)
         );
  DFF_X1 \REGISTERS_reg[15][21]  ( .D(n7063), .CK(CLK), .Q(n21073), .QN(n9547)
         );
  DFF_X1 \REGISTERS_reg[15][20]  ( .D(n7062), .CK(CLK), .Q(n21074), .QN(n9548)
         );
  DFF_X1 \REGISTERS_reg[15][19]  ( .D(n7061), .CK(CLK), .Q(n21075), .QN(n9549)
         );
  DFF_X1 \REGISTERS_reg[15][18]  ( .D(n7060), .CK(CLK), .Q(n21076), .QN(n9550)
         );
  DFF_X1 \REGISTERS_reg[15][17]  ( .D(n7059), .CK(CLK), .Q(n21077), .QN(n9551)
         );
  DFF_X1 \REGISTERS_reg[15][16]  ( .D(n7058), .CK(CLK), .Q(n21078), .QN(n9552)
         );
  DFF_X1 \REGISTERS_reg[15][15]  ( .D(n7057), .CK(CLK), .Q(n21079), .QN(n9553)
         );
  DFF_X1 \REGISTERS_reg[15][14]  ( .D(n7056), .CK(CLK), .Q(n21080), .QN(n9554)
         );
  DFF_X1 \REGISTERS_reg[15][13]  ( .D(n7055), .CK(CLK), .Q(n21081), .QN(n9555)
         );
  DFF_X1 \REGISTERS_reg[15][12]  ( .D(n7054), .CK(CLK), .Q(n21082), .QN(n9556)
         );
  DFF_X1 \REGISTERS_reg[15][11]  ( .D(n7053), .CK(CLK), .Q(n21083), .QN(n9557)
         );
  DFF_X1 \REGISTERS_reg[15][10]  ( .D(n7052), .CK(CLK), .Q(n21084), .QN(n9558)
         );
  DFF_X1 \REGISTERS_reg[15][9]  ( .D(n7051), .CK(CLK), .Q(n21085), .QN(n9559)
         );
  DFF_X1 \REGISTERS_reg[15][8]  ( .D(n7050), .CK(CLK), .Q(n21086), .QN(n9560)
         );
  DFF_X1 \REGISTERS_reg[15][7]  ( .D(n7049), .CK(CLK), .Q(n21087), .QN(n9561)
         );
  DFF_X1 \REGISTERS_reg[15][6]  ( .D(n7048), .CK(CLK), .Q(n21088), .QN(n9562)
         );
  DFF_X1 \REGISTERS_reg[15][5]  ( .D(n7047), .CK(CLK), .Q(n21089), .QN(n9563)
         );
  DFF_X1 \REGISTERS_reg[15][4]  ( .D(n7046), .CK(CLK), .Q(n21090), .QN(n9564)
         );
  DFF_X1 \REGISTERS_reg[15][3]  ( .D(n7045), .CK(CLK), .Q(n21091), .QN(n9565)
         );
  DFF_X1 \REGISTERS_reg[15][2]  ( .D(n7044), .CK(CLK), .Q(n21092), .QN(n9566)
         );
  DFF_X1 \REGISTERS_reg[15][1]  ( .D(n7043), .CK(CLK), .Q(n21093), .QN(n9567)
         );
  DFF_X1 \REGISTERS_reg[15][0]  ( .D(n7042), .CK(CLK), .Q(n21094), .QN(n9568)
         );
  DFF_X1 \REGISTERS_reg[13][59]  ( .D(n7229), .CK(CLK), .Q(n21095), .QN(n9701)
         );
  DFF_X1 \REGISTERS_reg[13][58]  ( .D(n7228), .CK(CLK), .Q(n21096), .QN(n9702)
         );
  DFF_X1 \REGISTERS_reg[13][57]  ( .D(n7227), .CK(CLK), .Q(n21097), .QN(n9703)
         );
  DFF_X1 \REGISTERS_reg[13][56]  ( .D(n7226), .CK(CLK), .Q(n21098), .QN(n9704)
         );
  DFF_X1 \REGISTERS_reg[13][55]  ( .D(n7225), .CK(CLK), .Q(n21099), .QN(n9705)
         );
  DFF_X1 \REGISTERS_reg[13][54]  ( .D(n7224), .CK(CLK), .Q(n21100), .QN(n9706)
         );
  DFF_X1 \REGISTERS_reg[13][53]  ( .D(n7223), .CK(CLK), .Q(n21101), .QN(n9707)
         );
  DFF_X1 \REGISTERS_reg[13][52]  ( .D(n7222), .CK(CLK), .Q(n21102), .QN(n9708)
         );
  DFF_X1 \REGISTERS_reg[13][51]  ( .D(n7221), .CK(CLK), .Q(n21103), .QN(n9709)
         );
  DFF_X1 \REGISTERS_reg[13][50]  ( .D(n7220), .CK(CLK), .Q(n21104), .QN(n9710)
         );
  DFF_X1 \REGISTERS_reg[13][49]  ( .D(n7219), .CK(CLK), .Q(n21105), .QN(n9711)
         );
  DFF_X1 \REGISTERS_reg[13][48]  ( .D(n7218), .CK(CLK), .Q(n21106), .QN(n9712)
         );
  DFF_X1 \REGISTERS_reg[13][47]  ( .D(n7217), .CK(CLK), .Q(n21107), .QN(n9713)
         );
  DFF_X1 \REGISTERS_reg[13][46]  ( .D(n7216), .CK(CLK), .Q(n21108), .QN(n9714)
         );
  DFF_X1 \REGISTERS_reg[13][45]  ( .D(n7215), .CK(CLK), .Q(n21109), .QN(n9715)
         );
  DFF_X1 \REGISTERS_reg[13][44]  ( .D(n7214), .CK(CLK), .Q(n21110), .QN(n9716)
         );
  DFF_X1 \REGISTERS_reg[13][43]  ( .D(n7213), .CK(CLK), .Q(n21111), .QN(n9717)
         );
  DFF_X1 \REGISTERS_reg[13][42]  ( .D(n7212), .CK(CLK), .Q(n21112), .QN(n9718)
         );
  DFF_X1 \REGISTERS_reg[13][41]  ( .D(n7211), .CK(CLK), .Q(n21113), .QN(n9719)
         );
  DFF_X1 \REGISTERS_reg[13][40]  ( .D(n7210), .CK(CLK), .Q(n21114), .QN(n9720)
         );
  DFF_X1 \REGISTERS_reg[13][39]  ( .D(n7209), .CK(CLK), .Q(n21115), .QN(n9721)
         );
  DFF_X1 \REGISTERS_reg[13][38]  ( .D(n7208), .CK(CLK), .Q(n21116), .QN(n9722)
         );
  DFF_X1 \REGISTERS_reg[13][37]  ( .D(n7207), .CK(CLK), .Q(n21117), .QN(n9723)
         );
  DFF_X1 \REGISTERS_reg[13][36]  ( .D(n7206), .CK(CLK), .Q(n21118), .QN(n9724)
         );
  DFF_X1 \REGISTERS_reg[13][35]  ( .D(n7205), .CK(CLK), .Q(n21119), .QN(n9725)
         );
  DFF_X1 \REGISTERS_reg[13][34]  ( .D(n7204), .CK(CLK), .Q(n21120), .QN(n9726)
         );
  DFF_X1 \REGISTERS_reg[13][33]  ( .D(n7203), .CK(CLK), .Q(n21121), .QN(n9727)
         );
  DFF_X1 \REGISTERS_reg[13][32]  ( .D(n7202), .CK(CLK), .Q(n21122), .QN(n9728)
         );
  DFF_X1 \REGISTERS_reg[13][31]  ( .D(n7201), .CK(CLK), .Q(n21123), .QN(n9729)
         );
  DFF_X1 \REGISTERS_reg[13][30]  ( .D(n7200), .CK(CLK), .Q(n21124), .QN(n9730)
         );
  DFF_X1 \REGISTERS_reg[13][29]  ( .D(n7199), .CK(CLK), .Q(n21125), .QN(n9731)
         );
  DFF_X1 \REGISTERS_reg[13][28]  ( .D(n7198), .CK(CLK), .Q(n21126), .QN(n9732)
         );
  DFF_X1 \REGISTERS_reg[13][27]  ( .D(n7197), .CK(CLK), .Q(n21127), .QN(n9733)
         );
  DFF_X1 \REGISTERS_reg[13][26]  ( .D(n7196), .CK(CLK), .Q(n21128), .QN(n9734)
         );
  DFF_X1 \REGISTERS_reg[13][25]  ( .D(n7195), .CK(CLK), .Q(n21129), .QN(n9735)
         );
  DFF_X1 \REGISTERS_reg[13][24]  ( .D(n7194), .CK(CLK), .Q(n21130), .QN(n9736)
         );
  DFF_X1 \REGISTERS_reg[13][23]  ( .D(n7193), .CK(CLK), .Q(n21131), .QN(n9737)
         );
  DFF_X1 \REGISTERS_reg[13][22]  ( .D(n7192), .CK(CLK), .Q(n21132), .QN(n9738)
         );
  DFF_X1 \REGISTERS_reg[13][21]  ( .D(n7191), .CK(CLK), .Q(n21133), .QN(n9739)
         );
  DFF_X1 \REGISTERS_reg[13][20]  ( .D(n7190), .CK(CLK), .Q(n21134), .QN(n9740)
         );
  DFF_X1 \REGISTERS_reg[13][19]  ( .D(n7189), .CK(CLK), .Q(n21135), .QN(n9741)
         );
  DFF_X1 \REGISTERS_reg[13][18]  ( .D(n7188), .CK(CLK), .Q(n21136), .QN(n9742)
         );
  DFF_X1 \REGISTERS_reg[13][17]  ( .D(n7187), .CK(CLK), .Q(n21137), .QN(n9743)
         );
  DFF_X1 \REGISTERS_reg[13][16]  ( .D(n7186), .CK(CLK), .Q(n21138), .QN(n9744)
         );
  DFF_X1 \REGISTERS_reg[13][15]  ( .D(n7185), .CK(CLK), .Q(n21139), .QN(n9745)
         );
  DFF_X1 \REGISTERS_reg[13][14]  ( .D(n7184), .CK(CLK), .Q(n21140), .QN(n9746)
         );
  DFF_X1 \REGISTERS_reg[13][13]  ( .D(n7183), .CK(CLK), .Q(n21141), .QN(n9747)
         );
  DFF_X1 \REGISTERS_reg[13][12]  ( .D(n7182), .CK(CLK), .Q(n21142), .QN(n9748)
         );
  DFF_X1 \REGISTERS_reg[13][11]  ( .D(n7181), .CK(CLK), .Q(n21143), .QN(n9749)
         );
  DFF_X1 \REGISTERS_reg[13][10]  ( .D(n7180), .CK(CLK), .Q(n21144), .QN(n9750)
         );
  DFF_X1 \REGISTERS_reg[13][9]  ( .D(n7179), .CK(CLK), .Q(n21145), .QN(n9751)
         );
  DFF_X1 \REGISTERS_reg[13][8]  ( .D(n7178), .CK(CLK), .Q(n21146), .QN(n9752)
         );
  DFF_X1 \REGISTERS_reg[13][7]  ( .D(n7177), .CK(CLK), .Q(n21147), .QN(n9753)
         );
  DFF_X1 \REGISTERS_reg[13][6]  ( .D(n7176), .CK(CLK), .Q(n21148), .QN(n9754)
         );
  DFF_X1 \REGISTERS_reg[13][5]  ( .D(n7175), .CK(CLK), .Q(n21149), .QN(n9755)
         );
  DFF_X1 \REGISTERS_reg[13][4]  ( .D(n7174), .CK(CLK), .Q(n21150), .QN(n9756)
         );
  DFF_X1 \REGISTERS_reg[13][3]  ( .D(n7173), .CK(CLK), .Q(n21151), .QN(n9757)
         );
  DFF_X1 \REGISTERS_reg[13][2]  ( .D(n7172), .CK(CLK), .Q(n21152), .QN(n9758)
         );
  DFF_X1 \REGISTERS_reg[13][1]  ( .D(n7171), .CK(CLK), .Q(n21153), .QN(n9759)
         );
  DFF_X1 \REGISTERS_reg[13][0]  ( .D(n7170), .CK(CLK), .Q(n21154), .QN(n9760)
         );
  DFF_X1 \REGISTERS_reg[20][63]  ( .D(n6785), .CK(CLK), .QN(n9569) );
  DFF_X1 \REGISTERS_reg[26][63]  ( .D(n6401), .CK(CLK), .QN(n21480) );
  DFF_X1 \REGISTERS_reg[26][62]  ( .D(n6400), .CK(CLK), .QN(n21481) );
  DFF_X1 \REGISTERS_reg[26][61]  ( .D(n6399), .CK(CLK), .QN(n21482) );
  DFF_X1 \REGISTERS_reg[26][60]  ( .D(n6398), .CK(CLK), .QN(n21483) );
  DFF_X1 \REGISTERS_reg[25][63]  ( .D(n6465), .CK(CLK), .QN(n21156) );
  DFF_X1 \REGISTERS_reg[25][62]  ( .D(n6464), .CK(CLK), .QN(n21157) );
  DFF_X1 \REGISTERS_reg[25][61]  ( .D(n6463), .CK(CLK), .QN(n21158) );
  DFF_X1 \REGISTERS_reg[25][60]  ( .D(n6462), .CK(CLK), .QN(n21159) );
  DFF_X1 \REGISTERS_reg[19][63]  ( .D(n6849), .CK(CLK), .QN(n22248) );
  DFF_X1 \REGISTERS_reg[19][62]  ( .D(n6848), .CK(CLK), .QN(n22249) );
  DFF_X1 \REGISTERS_reg[19][61]  ( .D(n6847), .CK(CLK), .QN(n22250) );
  DFF_X1 \REGISTERS_reg[19][60]  ( .D(n6846), .CK(CLK), .QN(n22251) );
  DFF_X1 \REGISTERS_reg[14][63]  ( .D(n7169), .CK(CLK), .QN(n21155) );
  DFF_X1 \REGISTERS_reg[14][62]  ( .D(n7168), .CK(CLK), .QN(n20772) );
  DFF_X1 \REGISTERS_reg[14][61]  ( .D(n7167), .CK(CLK), .QN(n20773) );
  DFF_X1 \REGISTERS_reg[14][60]  ( .D(n7166), .CK(CLK), .QN(n20774) );
  DFF_X1 \REGISTERS_reg[11][63]  ( .D(n7361), .CK(CLK), .QN(n21504) );
  DFF_X1 \REGISTERS_reg[11][62]  ( .D(n7360), .CK(CLK), .QN(n21505) );
  DFF_X1 \REGISTERS_reg[11][61]  ( .D(n7359), .CK(CLK), .QN(n21506) );
  DFF_X1 \REGISTERS_reg[11][60]  ( .D(n7358), .CK(CLK), .QN(n21507) );
  DFF_X1 \REGISTERS_reg[8][63]  ( .D(n7553), .CK(CLK), .QN(n22256) );
  DFF_X1 \REGISTERS_reg[8][62]  ( .D(n7552), .CK(CLK), .QN(n22257) );
  DFF_X1 \REGISTERS_reg[8][61]  ( .D(n7551), .CK(CLK), .QN(n22258) );
  DFF_X1 \REGISTERS_reg[8][60]  ( .D(n7550), .CK(CLK), .QN(n22259) );
  DFF_X1 \REGISTERS_reg[3][63]  ( .D(n7873), .CK(CLK), .QN(n21168) );
  DFF_X1 \REGISTERS_reg[3][62]  ( .D(n7872), .CK(CLK), .QN(n21169) );
  DFF_X1 \REGISTERS_reg[3][61]  ( .D(n7871), .CK(CLK), .QN(n21170) );
  DFF_X1 \REGISTERS_reg[3][60]  ( .D(n7870), .CK(CLK), .QN(n21171) );
  DFF_X1 \REGISTERS_reg[26][59]  ( .D(n6397), .CK(CLK), .QN(n21580) );
  DFF_X1 \REGISTERS_reg[26][58]  ( .D(n6396), .CK(CLK), .QN(n21581) );
  DFF_X1 \REGISTERS_reg[26][57]  ( .D(n6395), .CK(CLK), .QN(n21582) );
  DFF_X1 \REGISTERS_reg[26][56]  ( .D(n6394), .CK(CLK), .QN(n21583) );
  DFF_X1 \REGISTERS_reg[26][55]  ( .D(n6393), .CK(CLK), .QN(n21584) );
  DFF_X1 \REGISTERS_reg[26][54]  ( .D(n6392), .CK(CLK), .QN(n21585) );
  DFF_X1 \REGISTERS_reg[26][53]  ( .D(n6391), .CK(CLK), .QN(n21586) );
  DFF_X1 \REGISTERS_reg[26][52]  ( .D(n6390), .CK(CLK), .QN(n21587) );
  DFF_X1 \REGISTERS_reg[26][51]  ( .D(n6389), .CK(CLK), .QN(n21588) );
  DFF_X1 \REGISTERS_reg[26][50]  ( .D(n6388), .CK(CLK), .QN(n21589) );
  DFF_X1 \REGISTERS_reg[26][49]  ( .D(n6387), .CK(CLK), .QN(n21590) );
  DFF_X1 \REGISTERS_reg[26][48]  ( .D(n6386), .CK(CLK), .QN(n21591) );
  DFF_X1 \REGISTERS_reg[26][47]  ( .D(n6385), .CK(CLK), .QN(n21592) );
  DFF_X1 \REGISTERS_reg[26][46]  ( .D(n6384), .CK(CLK), .QN(n21593) );
  DFF_X1 \REGISTERS_reg[26][45]  ( .D(n6383), .CK(CLK), .QN(n21594) );
  DFF_X1 \REGISTERS_reg[26][44]  ( .D(n6382), .CK(CLK), .QN(n21595) );
  DFF_X1 \REGISTERS_reg[26][43]  ( .D(n6381), .CK(CLK), .QN(n21596) );
  DFF_X1 \REGISTERS_reg[26][42]  ( .D(n6380), .CK(CLK), .QN(n21597) );
  DFF_X1 \REGISTERS_reg[26][41]  ( .D(n6379), .CK(CLK), .QN(n21598) );
  DFF_X1 \REGISTERS_reg[26][40]  ( .D(n6378), .CK(CLK), .QN(n21599) );
  DFF_X1 \REGISTERS_reg[26][39]  ( .D(n6377), .CK(CLK), .QN(n21600) );
  DFF_X1 \REGISTERS_reg[26][38]  ( .D(n6376), .CK(CLK), .QN(n21601) );
  DFF_X1 \REGISTERS_reg[26][37]  ( .D(n6375), .CK(CLK), .QN(n21602) );
  DFF_X1 \REGISTERS_reg[26][36]  ( .D(n6374), .CK(CLK), .QN(n21603) );
  DFF_X1 \REGISTERS_reg[26][35]  ( .D(n6373), .CK(CLK), .QN(n21604) );
  DFF_X1 \REGISTERS_reg[26][34]  ( .D(n6372), .CK(CLK), .QN(n21605) );
  DFF_X1 \REGISTERS_reg[26][33]  ( .D(n6371), .CK(CLK), .QN(n21606) );
  DFF_X1 \REGISTERS_reg[26][32]  ( .D(n6370), .CK(CLK), .QN(n21607) );
  DFF_X1 \REGISTERS_reg[26][31]  ( .D(n6369), .CK(CLK), .QN(n21608) );
  DFF_X1 \REGISTERS_reg[26][30]  ( .D(n6368), .CK(CLK), .QN(n21609) );
  DFF_X1 \REGISTERS_reg[26][29]  ( .D(n6367), .CK(CLK), .QN(n21610) );
  DFF_X1 \REGISTERS_reg[26][28]  ( .D(n6366), .CK(CLK), .QN(n21611) );
  DFF_X1 \REGISTERS_reg[26][27]  ( .D(n6365), .CK(CLK), .QN(n21612) );
  DFF_X1 \REGISTERS_reg[26][26]  ( .D(n6364), .CK(CLK), .QN(n21613) );
  DFF_X1 \REGISTERS_reg[26][25]  ( .D(n6363), .CK(CLK), .QN(n21614) );
  DFF_X1 \REGISTERS_reg[26][24]  ( .D(n6362), .CK(CLK), .QN(n21615) );
  DFF_X1 \REGISTERS_reg[26][23]  ( .D(n6361), .CK(CLK), .QN(n21616) );
  DFF_X1 \REGISTERS_reg[26][22]  ( .D(n6360), .CK(CLK), .QN(n21617) );
  DFF_X1 \REGISTERS_reg[26][21]  ( .D(n6359), .CK(CLK), .QN(n21618) );
  DFF_X1 \REGISTERS_reg[26][20]  ( .D(n6358), .CK(CLK), .QN(n21619) );
  DFF_X1 \REGISTERS_reg[26][19]  ( .D(n6357), .CK(CLK), .QN(n21620) );
  DFF_X1 \REGISTERS_reg[26][18]  ( .D(n6356), .CK(CLK), .QN(n21621) );
  DFF_X1 \REGISTERS_reg[26][17]  ( .D(n6355), .CK(CLK), .QN(n21622) );
  DFF_X1 \REGISTERS_reg[26][16]  ( .D(n6354), .CK(CLK), .QN(n21623) );
  DFF_X1 \REGISTERS_reg[26][15]  ( .D(n6353), .CK(CLK), .QN(n21624) );
  DFF_X1 \REGISTERS_reg[26][14]  ( .D(n6352), .CK(CLK), .QN(n21625) );
  DFF_X1 \REGISTERS_reg[26][13]  ( .D(n6351), .CK(CLK), .QN(n21626) );
  DFF_X1 \REGISTERS_reg[26][12]  ( .D(n6350), .CK(CLK), .QN(n21627) );
  DFF_X1 \REGISTERS_reg[26][11]  ( .D(n6349), .CK(CLK), .QN(n21628) );
  DFF_X1 \REGISTERS_reg[26][10]  ( .D(n6348), .CK(CLK), .QN(n21629) );
  DFF_X1 \REGISTERS_reg[26][9]  ( .D(n6347), .CK(CLK), .QN(n21630) );
  DFF_X1 \REGISTERS_reg[26][8]  ( .D(n6346), .CK(CLK), .QN(n21631) );
  DFF_X1 \REGISTERS_reg[26][7]  ( .D(n6345), .CK(CLK), .QN(n21632) );
  DFF_X1 \REGISTERS_reg[26][6]  ( .D(n6344), .CK(CLK), .QN(n21633) );
  DFF_X1 \REGISTERS_reg[26][5]  ( .D(n6343), .CK(CLK), .QN(n21634) );
  DFF_X1 \REGISTERS_reg[26][4]  ( .D(n6342), .CK(CLK), .QN(n21635) );
  DFF_X1 \REGISTERS_reg[26][3]  ( .D(n6341), .CK(CLK), .QN(n21636) );
  DFF_X1 \REGISTERS_reg[26][2]  ( .D(n6340), .CK(CLK), .QN(n21637) );
  DFF_X1 \REGISTERS_reg[26][1]  ( .D(n6339), .CK(CLK), .QN(n21638) );
  DFF_X1 \REGISTERS_reg[26][0]  ( .D(n6338), .CK(CLK), .QN(n21639) );
  DFF_X1 \REGISTERS_reg[25][59]  ( .D(n6461), .CK(CLK), .QN(n21180) );
  DFF_X1 \REGISTERS_reg[25][58]  ( .D(n6460), .CK(CLK), .QN(n21181) );
  DFF_X1 \REGISTERS_reg[25][57]  ( .D(n6459), .CK(CLK), .QN(n21182) );
  DFF_X1 \REGISTERS_reg[25][56]  ( .D(n6458), .CK(CLK), .QN(n21183) );
  DFF_X1 \REGISTERS_reg[25][55]  ( .D(n6457), .CK(CLK), .QN(n21184) );
  DFF_X1 \REGISTERS_reg[25][54]  ( .D(n6456), .CK(CLK), .QN(n21185) );
  DFF_X1 \REGISTERS_reg[25][53]  ( .D(n6455), .CK(CLK), .QN(n21186) );
  DFF_X1 \REGISTERS_reg[25][52]  ( .D(n6454), .CK(CLK), .QN(n21187) );
  DFF_X1 \REGISTERS_reg[25][51]  ( .D(n6453), .CK(CLK), .QN(n21188) );
  DFF_X1 \REGISTERS_reg[25][50]  ( .D(n6452), .CK(CLK), .QN(n21189) );
  DFF_X1 \REGISTERS_reg[25][49]  ( .D(n6451), .CK(CLK), .QN(n21190) );
  DFF_X1 \REGISTERS_reg[25][48]  ( .D(n6450), .CK(CLK), .QN(n21191) );
  DFF_X1 \REGISTERS_reg[25][47]  ( .D(n6449), .CK(CLK), .QN(n21192) );
  DFF_X1 \REGISTERS_reg[25][46]  ( .D(n6448), .CK(CLK), .QN(n21193) );
  DFF_X1 \REGISTERS_reg[25][45]  ( .D(n6447), .CK(CLK), .QN(n21194) );
  DFF_X1 \REGISTERS_reg[25][44]  ( .D(n6446), .CK(CLK), .QN(n21195) );
  DFF_X1 \REGISTERS_reg[25][43]  ( .D(n6445), .CK(CLK), .QN(n21196) );
  DFF_X1 \REGISTERS_reg[25][42]  ( .D(n6444), .CK(CLK), .QN(n21197) );
  DFF_X1 \REGISTERS_reg[25][41]  ( .D(n6443), .CK(CLK), .QN(n21198) );
  DFF_X1 \REGISTERS_reg[25][40]  ( .D(n6442), .CK(CLK), .QN(n21199) );
  DFF_X1 \REGISTERS_reg[25][39]  ( .D(n6441), .CK(CLK), .QN(n21200) );
  DFF_X1 \REGISTERS_reg[25][38]  ( .D(n6440), .CK(CLK), .QN(n21201) );
  DFF_X1 \REGISTERS_reg[25][37]  ( .D(n6439), .CK(CLK), .QN(n21202) );
  DFF_X1 \REGISTERS_reg[25][36]  ( .D(n6438), .CK(CLK), .QN(n21203) );
  DFF_X1 \REGISTERS_reg[25][35]  ( .D(n6437), .CK(CLK), .QN(n21204) );
  DFF_X1 \REGISTERS_reg[25][34]  ( .D(n6436), .CK(CLK), .QN(n21205) );
  DFF_X1 \REGISTERS_reg[25][33]  ( .D(n6435), .CK(CLK), .QN(n21206) );
  DFF_X1 \REGISTERS_reg[25][32]  ( .D(n6434), .CK(CLK), .QN(n21207) );
  DFF_X1 \REGISTERS_reg[25][31]  ( .D(n6433), .CK(CLK), .QN(n21208) );
  DFF_X1 \REGISTERS_reg[25][30]  ( .D(n6432), .CK(CLK), .QN(n21209) );
  DFF_X1 \REGISTERS_reg[25][29]  ( .D(n6431), .CK(CLK), .QN(n21210) );
  DFF_X1 \REGISTERS_reg[25][28]  ( .D(n6430), .CK(CLK), .QN(n21211) );
  DFF_X1 \REGISTERS_reg[25][27]  ( .D(n6429), .CK(CLK), .QN(n21212) );
  DFF_X1 \REGISTERS_reg[25][26]  ( .D(n6428), .CK(CLK), .QN(n21213) );
  DFF_X1 \REGISTERS_reg[25][25]  ( .D(n6427), .CK(CLK), .QN(n21214) );
  DFF_X1 \REGISTERS_reg[25][24]  ( .D(n6426), .CK(CLK), .QN(n21215) );
  DFF_X1 \REGISTERS_reg[25][23]  ( .D(n6425), .CK(CLK), .QN(n21216) );
  DFF_X1 \REGISTERS_reg[25][22]  ( .D(n6424), .CK(CLK), .QN(n21217) );
  DFF_X1 \REGISTERS_reg[25][21]  ( .D(n6423), .CK(CLK), .QN(n21218) );
  DFF_X1 \REGISTERS_reg[25][20]  ( .D(n6422), .CK(CLK), .QN(n21219) );
  DFF_X1 \REGISTERS_reg[25][19]  ( .D(n6421), .CK(CLK), .QN(n21220) );
  DFF_X1 \REGISTERS_reg[25][18]  ( .D(n6420), .CK(CLK), .QN(n21221) );
  DFF_X1 \REGISTERS_reg[25][17]  ( .D(n6419), .CK(CLK), .QN(n21222) );
  DFF_X1 \REGISTERS_reg[25][16]  ( .D(n6418), .CK(CLK), .QN(n21223) );
  DFF_X1 \REGISTERS_reg[25][15]  ( .D(n6417), .CK(CLK), .QN(n21224) );
  DFF_X1 \REGISTERS_reg[25][14]  ( .D(n6416), .CK(CLK), .QN(n21225) );
  DFF_X1 \REGISTERS_reg[25][13]  ( .D(n6415), .CK(CLK), .QN(n21226) );
  DFF_X1 \REGISTERS_reg[25][12]  ( .D(n6414), .CK(CLK), .QN(n21227) );
  DFF_X1 \REGISTERS_reg[25][11]  ( .D(n6413), .CK(CLK), .QN(n21228) );
  DFF_X1 \REGISTERS_reg[25][10]  ( .D(n6412), .CK(CLK), .QN(n21229) );
  DFF_X1 \REGISTERS_reg[25][9]  ( .D(n6411), .CK(CLK), .QN(n21230) );
  DFF_X1 \REGISTERS_reg[25][8]  ( .D(n6410), .CK(CLK), .QN(n21231) );
  DFF_X1 \REGISTERS_reg[25][7]  ( .D(n6409), .CK(CLK), .QN(n21232) );
  DFF_X1 \REGISTERS_reg[25][6]  ( .D(n6408), .CK(CLK), .QN(n21233) );
  DFF_X1 \REGISTERS_reg[25][5]  ( .D(n6407), .CK(CLK), .QN(n21234) );
  DFF_X1 \REGISTERS_reg[25][4]  ( .D(n6406), .CK(CLK), .QN(n21235) );
  DFF_X1 \REGISTERS_reg[25][3]  ( .D(n6405), .CK(CLK), .QN(n21236) );
  DFF_X1 \REGISTERS_reg[25][2]  ( .D(n6404), .CK(CLK), .QN(n21237) );
  DFF_X1 \REGISTERS_reg[25][1]  ( .D(n6403), .CK(CLK), .QN(n21238) );
  DFF_X1 \REGISTERS_reg[25][0]  ( .D(n6402), .CK(CLK), .QN(n21239) );
  DFF_X1 \REGISTERS_reg[19][59]  ( .D(n6845), .CK(CLK), .QN(n22320) );
  DFF_X1 \REGISTERS_reg[19][58]  ( .D(n6844), .CK(CLK), .QN(n22321) );
  DFF_X1 \REGISTERS_reg[19][57]  ( .D(n6843), .CK(CLK), .QN(n22322) );
  DFF_X1 \REGISTERS_reg[19][56]  ( .D(n6842), .CK(CLK), .QN(n22323) );
  DFF_X1 \REGISTERS_reg[19][55]  ( .D(n6841), .CK(CLK), .QN(n22324) );
  DFF_X1 \REGISTERS_reg[19][54]  ( .D(n6840), .CK(CLK), .QN(n22325) );
  DFF_X1 \REGISTERS_reg[19][53]  ( .D(n6839), .CK(CLK), .QN(n22326) );
  DFF_X1 \REGISTERS_reg[19][52]  ( .D(n6838), .CK(CLK), .QN(n22327) );
  DFF_X1 \REGISTERS_reg[19][51]  ( .D(n6837), .CK(CLK), .QN(n22328) );
  DFF_X1 \REGISTERS_reg[19][50]  ( .D(n6836), .CK(CLK), .QN(n22329) );
  DFF_X1 \REGISTERS_reg[19][49]  ( .D(n6835), .CK(CLK), .QN(n22330) );
  DFF_X1 \REGISTERS_reg[19][48]  ( .D(n6834), .CK(CLK), .QN(n22331) );
  DFF_X1 \REGISTERS_reg[19][47]  ( .D(n6833), .CK(CLK), .QN(n22332) );
  DFF_X1 \REGISTERS_reg[19][46]  ( .D(n6832), .CK(CLK), .QN(n22333) );
  DFF_X1 \REGISTERS_reg[19][45]  ( .D(n6831), .CK(CLK), .QN(n22334) );
  DFF_X1 \REGISTERS_reg[19][44]  ( .D(n6830), .CK(CLK), .QN(n22335) );
  DFF_X1 \REGISTERS_reg[19][43]  ( .D(n6829), .CK(CLK), .QN(n22336) );
  DFF_X1 \REGISTERS_reg[19][42]  ( .D(n6828), .CK(CLK), .QN(n22337) );
  DFF_X1 \REGISTERS_reg[19][41]  ( .D(n6827), .CK(CLK), .QN(n22338) );
  DFF_X1 \REGISTERS_reg[19][40]  ( .D(n6826), .CK(CLK), .QN(n22339) );
  DFF_X1 \REGISTERS_reg[19][39]  ( .D(n6825), .CK(CLK), .QN(n22340) );
  DFF_X1 \REGISTERS_reg[19][38]  ( .D(n6824), .CK(CLK), .QN(n22341) );
  DFF_X1 \REGISTERS_reg[19][37]  ( .D(n6823), .CK(CLK), .QN(n22342) );
  DFF_X1 \REGISTERS_reg[19][36]  ( .D(n6822), .CK(CLK), .QN(n22343) );
  DFF_X1 \REGISTERS_reg[19][35]  ( .D(n6821), .CK(CLK), .QN(n22344) );
  DFF_X1 \REGISTERS_reg[19][34]  ( .D(n6820), .CK(CLK), .QN(n22345) );
  DFF_X1 \REGISTERS_reg[19][33]  ( .D(n6819), .CK(CLK), .QN(n22346) );
  DFF_X1 \REGISTERS_reg[19][32]  ( .D(n6818), .CK(CLK), .QN(n22347) );
  DFF_X1 \REGISTERS_reg[19][31]  ( .D(n6817), .CK(CLK), .QN(n22348) );
  DFF_X1 \REGISTERS_reg[19][30]  ( .D(n6816), .CK(CLK), .QN(n22349) );
  DFF_X1 \REGISTERS_reg[19][29]  ( .D(n6815), .CK(CLK), .QN(n22350) );
  DFF_X1 \REGISTERS_reg[19][28]  ( .D(n6814), .CK(CLK), .QN(n22351) );
  DFF_X1 \REGISTERS_reg[19][27]  ( .D(n6813), .CK(CLK), .QN(n22352) );
  DFF_X1 \REGISTERS_reg[19][26]  ( .D(n6812), .CK(CLK), .QN(n22353) );
  DFF_X1 \REGISTERS_reg[19][25]  ( .D(n6811), .CK(CLK), .QN(n22354) );
  DFF_X1 \REGISTERS_reg[19][24]  ( .D(n6810), .CK(CLK), .QN(n22355) );
  DFF_X1 \REGISTERS_reg[19][23]  ( .D(n6809), .CK(CLK), .QN(n22356) );
  DFF_X1 \REGISTERS_reg[19][22]  ( .D(n6808), .CK(CLK), .QN(n22357) );
  DFF_X1 \REGISTERS_reg[19][21]  ( .D(n6807), .CK(CLK), .QN(n22358) );
  DFF_X1 \REGISTERS_reg[19][20]  ( .D(n6806), .CK(CLK), .QN(n22359) );
  DFF_X1 \REGISTERS_reg[19][19]  ( .D(n6805), .CK(CLK), .QN(n22360) );
  DFF_X1 \REGISTERS_reg[19][18]  ( .D(n6804), .CK(CLK), .QN(n22361) );
  DFF_X1 \REGISTERS_reg[19][17]  ( .D(n6803), .CK(CLK), .QN(n22362) );
  DFF_X1 \REGISTERS_reg[19][16]  ( .D(n6802), .CK(CLK), .QN(n22363) );
  DFF_X1 \REGISTERS_reg[19][15]  ( .D(n6801), .CK(CLK), .QN(n22364) );
  DFF_X1 \REGISTERS_reg[19][14]  ( .D(n6800), .CK(CLK), .QN(n22365) );
  DFF_X1 \REGISTERS_reg[19][13]  ( .D(n6799), .CK(CLK), .QN(n22366) );
  DFF_X1 \REGISTERS_reg[19][12]  ( .D(n6798), .CK(CLK), .QN(n22367) );
  DFF_X1 \REGISTERS_reg[19][11]  ( .D(n6797), .CK(CLK), .QN(n22368) );
  DFF_X1 \REGISTERS_reg[19][10]  ( .D(n6796), .CK(CLK), .QN(n22369) );
  DFF_X1 \REGISTERS_reg[19][9]  ( .D(n6795), .CK(CLK), .QN(n22370) );
  DFF_X1 \REGISTERS_reg[19][8]  ( .D(n6794), .CK(CLK), .QN(n22371) );
  DFF_X1 \REGISTERS_reg[19][7]  ( .D(n6793), .CK(CLK), .QN(n22372) );
  DFF_X1 \REGISTERS_reg[19][6]  ( .D(n6792), .CK(CLK), .QN(n22373) );
  DFF_X1 \REGISTERS_reg[19][5]  ( .D(n6791), .CK(CLK), .QN(n22374) );
  DFF_X1 \REGISTERS_reg[19][4]  ( .D(n6790), .CK(CLK), .QN(n22375) );
  DFF_X1 \REGISTERS_reg[19][3]  ( .D(n6789), .CK(CLK), .QN(n22376) );
  DFF_X1 \REGISTERS_reg[19][2]  ( .D(n6788), .CK(CLK), .QN(n22377) );
  DFF_X1 \REGISTERS_reg[19][1]  ( .D(n6787), .CK(CLK), .QN(n22378) );
  DFF_X1 \REGISTERS_reg[19][0]  ( .D(n6786), .CK(CLK), .QN(n22379) );
  DFF_X1 \REGISTERS_reg[14][59]  ( .D(n7165), .CK(CLK), .QN(n20775) );
  DFF_X1 \REGISTERS_reg[14][58]  ( .D(n7164), .CK(CLK), .QN(n20776) );
  DFF_X1 \REGISTERS_reg[14][57]  ( .D(n7163), .CK(CLK), .QN(n20777) );
  DFF_X1 \REGISTERS_reg[14][56]  ( .D(n7162), .CK(CLK), .QN(n20778) );
  DFF_X1 \REGISTERS_reg[14][55]  ( .D(n7161), .CK(CLK), .QN(n20779) );
  DFF_X1 \REGISTERS_reg[14][54]  ( .D(n7160), .CK(CLK), .QN(n20780) );
  DFF_X1 \REGISTERS_reg[14][53]  ( .D(n7159), .CK(CLK), .QN(n20781) );
  DFF_X1 \REGISTERS_reg[14][52]  ( .D(n7158), .CK(CLK), .QN(n20782) );
  DFF_X1 \REGISTERS_reg[14][51]  ( .D(n7157), .CK(CLK), .QN(n20783) );
  DFF_X1 \REGISTERS_reg[14][50]  ( .D(n7156), .CK(CLK), .QN(n20784) );
  DFF_X1 \REGISTERS_reg[14][49]  ( .D(n7155), .CK(CLK), .QN(n20785) );
  DFF_X1 \REGISTERS_reg[14][48]  ( .D(n7154), .CK(CLK), .QN(n20786) );
  DFF_X1 \REGISTERS_reg[14][47]  ( .D(n7153), .CK(CLK), .QN(n20787) );
  DFF_X1 \REGISTERS_reg[14][46]  ( .D(n7152), .CK(CLK), .QN(n20788) );
  DFF_X1 \REGISTERS_reg[14][45]  ( .D(n7151), .CK(CLK), .QN(n20789) );
  DFF_X1 \REGISTERS_reg[14][44]  ( .D(n7150), .CK(CLK), .QN(n20790) );
  DFF_X1 \REGISTERS_reg[14][43]  ( .D(n7149), .CK(CLK), .QN(n20791) );
  DFF_X1 \REGISTERS_reg[14][42]  ( .D(n7148), .CK(CLK), .QN(n20792) );
  DFF_X1 \REGISTERS_reg[14][41]  ( .D(n7147), .CK(CLK), .QN(n20793) );
  DFF_X1 \REGISTERS_reg[14][40]  ( .D(n7146), .CK(CLK), .QN(n20794) );
  DFF_X1 \REGISTERS_reg[14][39]  ( .D(n7145), .CK(CLK), .QN(n20795) );
  DFF_X1 \REGISTERS_reg[14][38]  ( .D(n7144), .CK(CLK), .QN(n20796) );
  DFF_X1 \REGISTERS_reg[14][37]  ( .D(n7143), .CK(CLK), .QN(n20797) );
  DFF_X1 \REGISTERS_reg[14][36]  ( .D(n7142), .CK(CLK), .QN(n20798) );
  DFF_X1 \REGISTERS_reg[14][35]  ( .D(n7141), .CK(CLK), .QN(n20799) );
  DFF_X1 \REGISTERS_reg[14][34]  ( .D(n7140), .CK(CLK), .QN(n20800) );
  DFF_X1 \REGISTERS_reg[14][33]  ( .D(n7139), .CK(CLK), .QN(n20801) );
  DFF_X1 \REGISTERS_reg[14][32]  ( .D(n7138), .CK(CLK), .QN(n20802) );
  DFF_X1 \REGISTERS_reg[14][31]  ( .D(n7137), .CK(CLK), .QN(n20803) );
  DFF_X1 \REGISTERS_reg[14][30]  ( .D(n7136), .CK(CLK), .QN(n20804) );
  DFF_X1 \REGISTERS_reg[14][29]  ( .D(n7135), .CK(CLK), .QN(n20805) );
  DFF_X1 \REGISTERS_reg[14][28]  ( .D(n7134), .CK(CLK), .QN(n20806) );
  DFF_X1 \REGISTERS_reg[14][27]  ( .D(n7133), .CK(CLK), .QN(n20807) );
  DFF_X1 \REGISTERS_reg[14][26]  ( .D(n7132), .CK(CLK), .QN(n20808) );
  DFF_X1 \REGISTERS_reg[14][25]  ( .D(n7131), .CK(CLK), .QN(n20809) );
  DFF_X1 \REGISTERS_reg[14][24]  ( .D(n7130), .CK(CLK), .QN(n20810) );
  DFF_X1 \REGISTERS_reg[14][23]  ( .D(n7129), .CK(CLK), .QN(n20811) );
  DFF_X1 \REGISTERS_reg[14][22]  ( .D(n7128), .CK(CLK), .QN(n20812) );
  DFF_X1 \REGISTERS_reg[14][21]  ( .D(n7127), .CK(CLK), .QN(n20813) );
  DFF_X1 \REGISTERS_reg[14][20]  ( .D(n7126), .CK(CLK), .QN(n20814) );
  DFF_X1 \REGISTERS_reg[14][19]  ( .D(n7125), .CK(CLK), .QN(n20815) );
  DFF_X1 \REGISTERS_reg[14][18]  ( .D(n7124), .CK(CLK), .QN(n20816) );
  DFF_X1 \REGISTERS_reg[14][17]  ( .D(n7123), .CK(CLK), .QN(n20817) );
  DFF_X1 \REGISTERS_reg[14][16]  ( .D(n7122), .CK(CLK), .QN(n20818) );
  DFF_X1 \REGISTERS_reg[14][15]  ( .D(n7121), .CK(CLK), .QN(n20819) );
  DFF_X1 \REGISTERS_reg[14][14]  ( .D(n7120), .CK(CLK), .QN(n20820) );
  DFF_X1 \REGISTERS_reg[14][13]  ( .D(n7119), .CK(CLK), .QN(n20821) );
  DFF_X1 \REGISTERS_reg[14][12]  ( .D(n7118), .CK(CLK), .QN(n20822) );
  DFF_X1 \REGISTERS_reg[14][11]  ( .D(n7117), .CK(CLK), .QN(n20823) );
  DFF_X1 \REGISTERS_reg[14][10]  ( .D(n7116), .CK(CLK), .QN(n20824) );
  DFF_X1 \REGISTERS_reg[14][9]  ( .D(n7115), .CK(CLK), .QN(n20825) );
  DFF_X1 \REGISTERS_reg[14][8]  ( .D(n7114), .CK(CLK), .QN(n20826) );
  DFF_X1 \REGISTERS_reg[14][7]  ( .D(n7113), .CK(CLK), .QN(n20827) );
  DFF_X1 \REGISTERS_reg[14][6]  ( .D(n7112), .CK(CLK), .QN(n20828) );
  DFF_X1 \REGISTERS_reg[14][5]  ( .D(n7111), .CK(CLK), .QN(n20829) );
  DFF_X1 \REGISTERS_reg[14][4]  ( .D(n7110), .CK(CLK), .QN(n20830) );
  DFF_X1 \REGISTERS_reg[14][3]  ( .D(n7109), .CK(CLK), .QN(n20831) );
  DFF_X1 \REGISTERS_reg[14][2]  ( .D(n7108), .CK(CLK), .QN(n20832) );
  DFF_X1 \REGISTERS_reg[14][1]  ( .D(n7107), .CK(CLK), .QN(n20833) );
  DFF_X1 \REGISTERS_reg[14][0]  ( .D(n7106), .CK(CLK), .QN(n20834) );
  DFF_X1 \REGISTERS_reg[11][59]  ( .D(n7357), .CK(CLK), .QN(n21940) );
  DFF_X1 \REGISTERS_reg[11][58]  ( .D(n7356), .CK(CLK), .QN(n21941) );
  DFF_X1 \REGISTERS_reg[11][57]  ( .D(n7355), .CK(CLK), .QN(n21942) );
  DFF_X1 \REGISTERS_reg[11][56]  ( .D(n7354), .CK(CLK), .QN(n21943) );
  DFF_X1 \REGISTERS_reg[11][55]  ( .D(n7353), .CK(CLK), .QN(n21944) );
  DFF_X1 \REGISTERS_reg[11][54]  ( .D(n7352), .CK(CLK), .QN(n21945) );
  DFF_X1 \REGISTERS_reg[11][53]  ( .D(n7351), .CK(CLK), .QN(n21946) );
  DFF_X1 \REGISTERS_reg[11][52]  ( .D(n7350), .CK(CLK), .QN(n21947) );
  DFF_X1 \REGISTERS_reg[11][51]  ( .D(n7349), .CK(CLK), .QN(n21948) );
  DFF_X1 \REGISTERS_reg[11][50]  ( .D(n7348), .CK(CLK), .QN(n21949) );
  DFF_X1 \REGISTERS_reg[11][49]  ( .D(n7347), .CK(CLK), .QN(n21950) );
  DFF_X1 \REGISTERS_reg[11][48]  ( .D(n7346), .CK(CLK), .QN(n21951) );
  DFF_X1 \REGISTERS_reg[11][47]  ( .D(n7345), .CK(CLK), .QN(n21952) );
  DFF_X1 \REGISTERS_reg[11][46]  ( .D(n7344), .CK(CLK), .QN(n21953) );
  DFF_X1 \REGISTERS_reg[11][45]  ( .D(n7343), .CK(CLK), .QN(n21954) );
  DFF_X1 \REGISTERS_reg[11][44]  ( .D(n7342), .CK(CLK), .QN(n21955) );
  DFF_X1 \REGISTERS_reg[11][43]  ( .D(n7341), .CK(CLK), .QN(n21956) );
  DFF_X1 \REGISTERS_reg[11][42]  ( .D(n7340), .CK(CLK), .QN(n21957) );
  DFF_X1 \REGISTERS_reg[11][41]  ( .D(n7339), .CK(CLK), .QN(n21958) );
  DFF_X1 \REGISTERS_reg[11][40]  ( .D(n7338), .CK(CLK), .QN(n21959) );
  DFF_X1 \REGISTERS_reg[11][39]  ( .D(n7337), .CK(CLK), .QN(n21960) );
  DFF_X1 \REGISTERS_reg[11][38]  ( .D(n7336), .CK(CLK), .QN(n21961) );
  DFF_X1 \REGISTERS_reg[11][37]  ( .D(n7335), .CK(CLK), .QN(n21962) );
  DFF_X1 \REGISTERS_reg[11][36]  ( .D(n7334), .CK(CLK), .QN(n21963) );
  DFF_X1 \REGISTERS_reg[11][35]  ( .D(n7333), .CK(CLK), .QN(n21964) );
  DFF_X1 \REGISTERS_reg[11][34]  ( .D(n7332), .CK(CLK), .QN(n21965) );
  DFF_X1 \REGISTERS_reg[11][33]  ( .D(n7331), .CK(CLK), .QN(n21966) );
  DFF_X1 \REGISTERS_reg[11][32]  ( .D(n7330), .CK(CLK), .QN(n21967) );
  DFF_X1 \REGISTERS_reg[11][31]  ( .D(n7329), .CK(CLK), .QN(n21968) );
  DFF_X1 \REGISTERS_reg[11][30]  ( .D(n7328), .CK(CLK), .QN(n21969) );
  DFF_X1 \REGISTERS_reg[11][29]  ( .D(n7327), .CK(CLK), .QN(n21970) );
  DFF_X1 \REGISTERS_reg[11][28]  ( .D(n7326), .CK(CLK), .QN(n21971) );
  DFF_X1 \REGISTERS_reg[11][27]  ( .D(n7325), .CK(CLK), .QN(n21972) );
  DFF_X1 \REGISTERS_reg[11][26]  ( .D(n7324), .CK(CLK), .QN(n21973) );
  DFF_X1 \REGISTERS_reg[11][25]  ( .D(n7323), .CK(CLK), .QN(n21974) );
  DFF_X1 \REGISTERS_reg[11][24]  ( .D(n7322), .CK(CLK), .QN(n21975) );
  DFF_X1 \REGISTERS_reg[11][23]  ( .D(n7321), .CK(CLK), .QN(n21976) );
  DFF_X1 \REGISTERS_reg[11][22]  ( .D(n7320), .CK(CLK), .QN(n21977) );
  DFF_X1 \REGISTERS_reg[11][21]  ( .D(n7319), .CK(CLK), .QN(n21978) );
  DFF_X1 \REGISTERS_reg[11][20]  ( .D(n7318), .CK(CLK), .QN(n21979) );
  DFF_X1 \REGISTERS_reg[11][19]  ( .D(n7317), .CK(CLK), .QN(n21980) );
  DFF_X1 \REGISTERS_reg[11][18]  ( .D(n7316), .CK(CLK), .QN(n21981) );
  DFF_X1 \REGISTERS_reg[11][17]  ( .D(n7315), .CK(CLK), .QN(n21982) );
  DFF_X1 \REGISTERS_reg[11][16]  ( .D(n7314), .CK(CLK), .QN(n21983) );
  DFF_X1 \REGISTERS_reg[11][15]  ( .D(n7313), .CK(CLK), .QN(n21984) );
  DFF_X1 \REGISTERS_reg[11][14]  ( .D(n7312), .CK(CLK), .QN(n21985) );
  DFF_X1 \REGISTERS_reg[11][13]  ( .D(n7311), .CK(CLK), .QN(n21986) );
  DFF_X1 \REGISTERS_reg[11][12]  ( .D(n7310), .CK(CLK), .QN(n21987) );
  DFF_X1 \REGISTERS_reg[11][11]  ( .D(n7309), .CK(CLK), .QN(n21988) );
  DFF_X1 \REGISTERS_reg[11][10]  ( .D(n7308), .CK(CLK), .QN(n21989) );
  DFF_X1 \REGISTERS_reg[11][9]  ( .D(n7307), .CK(CLK), .QN(n21990) );
  DFF_X1 \REGISTERS_reg[11][8]  ( .D(n7306), .CK(CLK), .QN(n21991) );
  DFF_X1 \REGISTERS_reg[11][7]  ( .D(n7305), .CK(CLK), .QN(n21992) );
  DFF_X1 \REGISTERS_reg[11][6]  ( .D(n7304), .CK(CLK), .QN(n21993) );
  DFF_X1 \REGISTERS_reg[11][5]  ( .D(n7303), .CK(CLK), .QN(n21994) );
  DFF_X1 \REGISTERS_reg[11][4]  ( .D(n7302), .CK(CLK), .QN(n21995) );
  DFF_X1 \REGISTERS_reg[11][3]  ( .D(n7301), .CK(CLK), .QN(n21996) );
  DFF_X1 \REGISTERS_reg[11][2]  ( .D(n7300), .CK(CLK), .QN(n21997) );
  DFF_X1 \REGISTERS_reg[11][1]  ( .D(n7299), .CK(CLK), .QN(n21998) );
  DFF_X1 \REGISTERS_reg[11][0]  ( .D(n7298), .CK(CLK), .QN(n21999) );
  DFF_X1 \REGISTERS_reg[8][59]  ( .D(n7549), .CK(CLK), .QN(n22440) );
  DFF_X1 \REGISTERS_reg[8][58]  ( .D(n7548), .CK(CLK), .QN(n22441) );
  DFF_X1 \REGISTERS_reg[8][57]  ( .D(n7547), .CK(CLK), .QN(n22442) );
  DFF_X1 \REGISTERS_reg[8][56]  ( .D(n7546), .CK(CLK), .QN(n22443) );
  DFF_X1 \REGISTERS_reg[8][55]  ( .D(n7545), .CK(CLK), .QN(n22444) );
  DFF_X1 \REGISTERS_reg[8][54]  ( .D(n7544), .CK(CLK), .QN(n22445) );
  DFF_X1 \REGISTERS_reg[8][53]  ( .D(n7543), .CK(CLK), .QN(n22446) );
  DFF_X1 \REGISTERS_reg[8][52]  ( .D(n7542), .CK(CLK), .QN(n22447) );
  DFF_X1 \REGISTERS_reg[8][51]  ( .D(n7541), .CK(CLK), .QN(n22448) );
  DFF_X1 \REGISTERS_reg[8][50]  ( .D(n7540), .CK(CLK), .QN(n22449) );
  DFF_X1 \REGISTERS_reg[8][49]  ( .D(n7539), .CK(CLK), .QN(n22450) );
  DFF_X1 \REGISTERS_reg[8][48]  ( .D(n7538), .CK(CLK), .QN(n22451) );
  DFF_X1 \REGISTERS_reg[8][47]  ( .D(n7537), .CK(CLK), .QN(n22452) );
  DFF_X1 \REGISTERS_reg[8][46]  ( .D(n7536), .CK(CLK), .QN(n22453) );
  DFF_X1 \REGISTERS_reg[8][45]  ( .D(n7535), .CK(CLK), .QN(n22454) );
  DFF_X1 \REGISTERS_reg[8][44]  ( .D(n7534), .CK(CLK), .QN(n22455) );
  DFF_X1 \REGISTERS_reg[8][43]  ( .D(n7533), .CK(CLK), .QN(n22456) );
  DFF_X1 \REGISTERS_reg[8][42]  ( .D(n7532), .CK(CLK), .QN(n22457) );
  DFF_X1 \REGISTERS_reg[8][41]  ( .D(n7531), .CK(CLK), .QN(n22458) );
  DFF_X1 \REGISTERS_reg[8][40]  ( .D(n7530), .CK(CLK), .QN(n22459) );
  DFF_X1 \REGISTERS_reg[8][39]  ( .D(n7529), .CK(CLK), .QN(n22460) );
  DFF_X1 \REGISTERS_reg[8][38]  ( .D(n7528), .CK(CLK), .QN(n22461) );
  DFF_X1 \REGISTERS_reg[8][37]  ( .D(n7527), .CK(CLK), .QN(n22462) );
  DFF_X1 \REGISTERS_reg[8][36]  ( .D(n7526), .CK(CLK), .QN(n22463) );
  DFF_X1 \REGISTERS_reg[8][35]  ( .D(n7525), .CK(CLK), .QN(n22464) );
  DFF_X1 \REGISTERS_reg[8][34]  ( .D(n7524), .CK(CLK), .QN(n22465) );
  DFF_X1 \REGISTERS_reg[8][33]  ( .D(n7523), .CK(CLK), .QN(n22466) );
  DFF_X1 \REGISTERS_reg[8][32]  ( .D(n7522), .CK(CLK), .QN(n22467) );
  DFF_X1 \REGISTERS_reg[8][31]  ( .D(n7521), .CK(CLK), .QN(n22468) );
  DFF_X1 \REGISTERS_reg[8][30]  ( .D(n7520), .CK(CLK), .QN(n22469) );
  DFF_X1 \REGISTERS_reg[8][29]  ( .D(n7519), .CK(CLK), .QN(n22470) );
  DFF_X1 \REGISTERS_reg[8][28]  ( .D(n7518), .CK(CLK), .QN(n22471) );
  DFF_X1 \REGISTERS_reg[8][27]  ( .D(n7517), .CK(CLK), .QN(n22472) );
  DFF_X1 \REGISTERS_reg[8][26]  ( .D(n7516), .CK(CLK), .QN(n22473) );
  DFF_X1 \REGISTERS_reg[8][25]  ( .D(n7515), .CK(CLK), .QN(n22474) );
  DFF_X1 \REGISTERS_reg[8][24]  ( .D(n7514), .CK(CLK), .QN(n22475) );
  DFF_X1 \REGISTERS_reg[8][23]  ( .D(n7513), .CK(CLK), .QN(n22476) );
  DFF_X1 \REGISTERS_reg[8][22]  ( .D(n7512), .CK(CLK), .QN(n22477) );
  DFF_X1 \REGISTERS_reg[8][21]  ( .D(n7511), .CK(CLK), .QN(n22478) );
  DFF_X1 \REGISTERS_reg[8][20]  ( .D(n7510), .CK(CLK), .QN(n22479) );
  DFF_X1 \REGISTERS_reg[8][19]  ( .D(n7509), .CK(CLK), .QN(n22480) );
  DFF_X1 \REGISTERS_reg[8][18]  ( .D(n7508), .CK(CLK), .QN(n22481) );
  DFF_X1 \REGISTERS_reg[8][17]  ( .D(n7507), .CK(CLK), .QN(n22482) );
  DFF_X1 \REGISTERS_reg[8][16]  ( .D(n7506), .CK(CLK), .QN(n22483) );
  DFF_X1 \REGISTERS_reg[8][15]  ( .D(n7505), .CK(CLK), .QN(n22484) );
  DFF_X1 \REGISTERS_reg[8][14]  ( .D(n7504), .CK(CLK), .QN(n22485) );
  DFF_X1 \REGISTERS_reg[8][13]  ( .D(n7503), .CK(CLK), .QN(n22486) );
  DFF_X1 \REGISTERS_reg[8][12]  ( .D(n7502), .CK(CLK), .QN(n22487) );
  DFF_X1 \REGISTERS_reg[8][11]  ( .D(n7501), .CK(CLK), .QN(n22488) );
  DFF_X1 \REGISTERS_reg[8][10]  ( .D(n7500), .CK(CLK), .QN(n22489) );
  DFF_X1 \REGISTERS_reg[8][9]  ( .D(n7499), .CK(CLK), .QN(n22490) );
  DFF_X1 \REGISTERS_reg[8][8]  ( .D(n7498), .CK(CLK), .QN(n22491) );
  DFF_X1 \REGISTERS_reg[8][7]  ( .D(n7497), .CK(CLK), .QN(n22492) );
  DFF_X1 \REGISTERS_reg[8][6]  ( .D(n7496), .CK(CLK), .QN(n22493) );
  DFF_X1 \REGISTERS_reg[8][5]  ( .D(n7495), .CK(CLK), .QN(n22494) );
  DFF_X1 \REGISTERS_reg[8][4]  ( .D(n7494), .CK(CLK), .QN(n22495) );
  DFF_X1 \REGISTERS_reg[8][3]  ( .D(n7493), .CK(CLK), .QN(n22496) );
  DFF_X1 \REGISTERS_reg[8][2]  ( .D(n7492), .CK(CLK), .QN(n22497) );
  DFF_X1 \REGISTERS_reg[8][1]  ( .D(n7491), .CK(CLK), .QN(n22498) );
  DFF_X1 \REGISTERS_reg[8][0]  ( .D(n7490), .CK(CLK), .QN(n22499) );
  DFF_X1 \REGISTERS_reg[3][59]  ( .D(n7869), .CK(CLK), .QN(n21360) );
  DFF_X1 \REGISTERS_reg[3][58]  ( .D(n7868), .CK(CLK), .QN(n21361) );
  DFF_X1 \REGISTERS_reg[3][57]  ( .D(n7867), .CK(CLK), .QN(n21362) );
  DFF_X1 \REGISTERS_reg[3][56]  ( .D(n7866), .CK(CLK), .QN(n21363) );
  DFF_X1 \REGISTERS_reg[3][55]  ( .D(n7865), .CK(CLK), .QN(n21364) );
  DFF_X1 \REGISTERS_reg[3][54]  ( .D(n7864), .CK(CLK), .QN(n21365) );
  DFF_X1 \REGISTERS_reg[3][53]  ( .D(n7863), .CK(CLK), .QN(n21366) );
  DFF_X1 \REGISTERS_reg[3][52]  ( .D(n7862), .CK(CLK), .QN(n21367) );
  DFF_X1 \REGISTERS_reg[3][51]  ( .D(n7861), .CK(CLK), .QN(n21368) );
  DFF_X1 \REGISTERS_reg[3][50]  ( .D(n7860), .CK(CLK), .QN(n21369) );
  DFF_X1 \REGISTERS_reg[3][49]  ( .D(n7859), .CK(CLK), .QN(n21370) );
  DFF_X1 \REGISTERS_reg[3][48]  ( .D(n7858), .CK(CLK), .QN(n21371) );
  DFF_X1 \REGISTERS_reg[3][47]  ( .D(n7857), .CK(CLK), .QN(n21372) );
  DFF_X1 \REGISTERS_reg[3][46]  ( .D(n7856), .CK(CLK), .QN(n21373) );
  DFF_X1 \REGISTERS_reg[3][45]  ( .D(n7855), .CK(CLK), .QN(n21374) );
  DFF_X1 \REGISTERS_reg[3][44]  ( .D(n7854), .CK(CLK), .QN(n21375) );
  DFF_X1 \REGISTERS_reg[3][43]  ( .D(n7853), .CK(CLK), .QN(n21376) );
  DFF_X1 \REGISTERS_reg[3][42]  ( .D(n7852), .CK(CLK), .QN(n21377) );
  DFF_X1 \REGISTERS_reg[3][41]  ( .D(n7851), .CK(CLK), .QN(n21378) );
  DFF_X1 \REGISTERS_reg[3][40]  ( .D(n7850), .CK(CLK), .QN(n21379) );
  DFF_X1 \REGISTERS_reg[3][39]  ( .D(n7849), .CK(CLK), .QN(n21380) );
  DFF_X1 \REGISTERS_reg[3][38]  ( .D(n7848), .CK(CLK), .QN(n21381) );
  DFF_X1 \REGISTERS_reg[3][37]  ( .D(n7847), .CK(CLK), .QN(n21382) );
  DFF_X1 \REGISTERS_reg[3][36]  ( .D(n7846), .CK(CLK), .QN(n21383) );
  DFF_X1 \REGISTERS_reg[3][35]  ( .D(n7845), .CK(CLK), .QN(n21384) );
  DFF_X1 \REGISTERS_reg[3][34]  ( .D(n7844), .CK(CLK), .QN(n21385) );
  DFF_X1 \REGISTERS_reg[3][33]  ( .D(n7843), .CK(CLK), .QN(n21386) );
  DFF_X1 \REGISTERS_reg[3][32]  ( .D(n7842), .CK(CLK), .QN(n21387) );
  DFF_X1 \REGISTERS_reg[3][31]  ( .D(n7841), .CK(CLK), .QN(n21388) );
  DFF_X1 \REGISTERS_reg[3][30]  ( .D(n7840), .CK(CLK), .QN(n21389) );
  DFF_X1 \REGISTERS_reg[3][29]  ( .D(n7839), .CK(CLK), .QN(n21390) );
  DFF_X1 \REGISTERS_reg[3][28]  ( .D(n7838), .CK(CLK), .QN(n21391) );
  DFF_X1 \REGISTERS_reg[3][27]  ( .D(n7837), .CK(CLK), .QN(n21392) );
  DFF_X1 \REGISTERS_reg[3][26]  ( .D(n7836), .CK(CLK), .QN(n21393) );
  DFF_X1 \REGISTERS_reg[3][25]  ( .D(n7835), .CK(CLK), .QN(n21394) );
  DFF_X1 \REGISTERS_reg[3][24]  ( .D(n7834), .CK(CLK), .QN(n21395) );
  DFF_X1 \REGISTERS_reg[3][23]  ( .D(n7833), .CK(CLK), .QN(n21396) );
  DFF_X1 \REGISTERS_reg[3][22]  ( .D(n7832), .CK(CLK), .QN(n21397) );
  DFF_X1 \REGISTERS_reg[3][21]  ( .D(n7831), .CK(CLK), .QN(n21398) );
  DFF_X1 \REGISTERS_reg[3][20]  ( .D(n7830), .CK(CLK), .QN(n21399) );
  DFF_X1 \REGISTERS_reg[3][19]  ( .D(n7829), .CK(CLK), .QN(n21400) );
  DFF_X1 \REGISTERS_reg[3][18]  ( .D(n7828), .CK(CLK), .QN(n21401) );
  DFF_X1 \REGISTERS_reg[3][17]  ( .D(n7827), .CK(CLK), .QN(n21402) );
  DFF_X1 \REGISTERS_reg[3][16]  ( .D(n7826), .CK(CLK), .QN(n21403) );
  DFF_X1 \REGISTERS_reg[3][15]  ( .D(n7825), .CK(CLK), .QN(n21404) );
  DFF_X1 \REGISTERS_reg[3][14]  ( .D(n7824), .CK(CLK), .QN(n21405) );
  DFF_X1 \REGISTERS_reg[3][13]  ( .D(n7823), .CK(CLK), .QN(n21406) );
  DFF_X1 \REGISTERS_reg[3][12]  ( .D(n7822), .CK(CLK), .QN(n21407) );
  DFF_X1 \REGISTERS_reg[3][11]  ( .D(n7821), .CK(CLK), .QN(n21408) );
  DFF_X1 \REGISTERS_reg[3][10]  ( .D(n7820), .CK(CLK), .QN(n21409) );
  DFF_X1 \REGISTERS_reg[3][9]  ( .D(n7819), .CK(CLK), .QN(n21410) );
  DFF_X1 \REGISTERS_reg[3][8]  ( .D(n7818), .CK(CLK), .QN(n21411) );
  DFF_X1 \REGISTERS_reg[3][7]  ( .D(n7817), .CK(CLK), .QN(n21412) );
  DFF_X1 \REGISTERS_reg[3][6]  ( .D(n7816), .CK(CLK), .QN(n21413) );
  DFF_X1 \REGISTERS_reg[3][5]  ( .D(n7815), .CK(CLK), .QN(n21414) );
  DFF_X1 \REGISTERS_reg[3][4]  ( .D(n7814), .CK(CLK), .QN(n21415) );
  DFF_X1 \REGISTERS_reg[3][3]  ( .D(n7813), .CK(CLK), .QN(n21416) );
  DFF_X1 \REGISTERS_reg[3][2]  ( .D(n7812), .CK(CLK), .QN(n21417) );
  DFF_X1 \REGISTERS_reg[3][1]  ( .D(n7811), .CK(CLK), .QN(n21418) );
  DFF_X1 \REGISTERS_reg[3][0]  ( .D(n7810), .CK(CLK), .QN(n21419) );
  DFF_X1 \REGISTERS_reg[24][63]  ( .D(n6529), .CK(CLK), .QN(n22500) );
  DFF_X1 \REGISTERS_reg[24][62]  ( .D(n6528), .CK(CLK), .QN(n22501) );
  DFF_X1 \REGISTERS_reg[24][61]  ( .D(n6527), .CK(CLK), .QN(n22502) );
  DFF_X1 \REGISTERS_reg[24][60]  ( .D(n6526), .CK(CLK), .QN(n22503) );
  DFF_X1 \REGISTERS_reg[23][63]  ( .D(n6593), .CK(CLK), .QN(n21164) );
  DFF_X1 \REGISTERS_reg[23][62]  ( .D(n6592), .CK(CLK), .QN(n21165) );
  DFF_X1 \REGISTERS_reg[23][61]  ( .D(n6591), .CK(CLK), .QN(n21166) );
  DFF_X1 \REGISTERS_reg[23][60]  ( .D(n6590), .CK(CLK), .QN(n21167) );
  DFF_X1 \REGISTERS_reg[17][63]  ( .D(n6977), .CK(CLK), .QN(n21488) );
  DFF_X1 \REGISTERS_reg[17][62]  ( .D(n6976), .CK(CLK), .QN(n21489) );
  DFF_X1 \REGISTERS_reg[17][61]  ( .D(n6975), .CK(CLK), .QN(n21490) );
  DFF_X1 \REGISTERS_reg[17][60]  ( .D(n6974), .CK(CLK), .QN(n21491) );
  DFF_X1 \REGISTERS_reg[12][63]  ( .D(n7297), .CK(CLK), .QN(n20708) );
  DFF_X1 \REGISTERS_reg[12][62]  ( .D(n7296), .CK(CLK), .QN(n20709) );
  DFF_X1 \REGISTERS_reg[12][61]  ( .D(n7295), .CK(CLK), .QN(n20710) );
  DFF_X1 \REGISTERS_reg[12][60]  ( .D(n7294), .CK(CLK), .QN(n20711) );
  DFF_X1 \REGISTERS_reg[9][63]  ( .D(n7489), .CK(CLK), .QN(n22508) );
  DFF_X1 \REGISTERS_reg[9][62]  ( .D(n7488), .CK(CLK), .QN(n22509) );
  DFF_X1 \REGISTERS_reg[9][61]  ( .D(n7487), .CK(CLK), .QN(n22510) );
  DFF_X1 \REGISTERS_reg[9][60]  ( .D(n7486), .CK(CLK), .QN(n22511) );
  DFF_X1 \REGISTERS_reg[7][63]  ( .D(n7617), .CK(CLK), .QN(n21508) );
  DFF_X1 \REGISTERS_reg[7][62]  ( .D(n7616), .CK(CLK), .QN(n21509) );
  DFF_X1 \REGISTERS_reg[7][61]  ( .D(n7615), .CK(CLK), .QN(n21510) );
  DFF_X1 \REGISTERS_reg[7][60]  ( .D(n7614), .CK(CLK), .QN(n21511) );
  DFF_X1 \REGISTERS_reg[5][63]  ( .D(n7745), .CK(CLK), .QN(n21176) );
  DFF_X1 \REGISTERS_reg[5][62]  ( .D(n7744), .CK(CLK), .QN(n21177) );
  DFF_X1 \REGISTERS_reg[5][61]  ( .D(n7743), .CK(CLK), .QN(n21178) );
  DFF_X1 \REGISTERS_reg[5][60]  ( .D(n7742), .CK(CLK), .QN(n21179) );
  DFF_X1 \REGISTERS_reg[24][59]  ( .D(n6525), .CK(CLK), .QN(n22512) );
  DFF_X1 \REGISTERS_reg[24][58]  ( .D(n6524), .CK(CLK), .QN(n22513) );
  DFF_X1 \REGISTERS_reg[24][57]  ( .D(n6523), .CK(CLK), .QN(n22514) );
  DFF_X1 \REGISTERS_reg[24][56]  ( .D(n6522), .CK(CLK), .QN(n22515) );
  DFF_X1 \REGISTERS_reg[24][55]  ( .D(n6521), .CK(CLK), .QN(n22516) );
  DFF_X1 \REGISTERS_reg[24][54]  ( .D(n6520), .CK(CLK), .QN(n22517) );
  DFF_X1 \REGISTERS_reg[24][53]  ( .D(n6519), .CK(CLK), .QN(n22518) );
  DFF_X1 \REGISTERS_reg[24][52]  ( .D(n6518), .CK(CLK), .QN(n22519) );
  DFF_X1 \REGISTERS_reg[24][51]  ( .D(n6517), .CK(CLK), .QN(n22520) );
  DFF_X1 \REGISTERS_reg[24][50]  ( .D(n6516), .CK(CLK), .QN(n22521) );
  DFF_X1 \REGISTERS_reg[24][49]  ( .D(n6515), .CK(CLK), .QN(n22522) );
  DFF_X1 \REGISTERS_reg[24][48]  ( .D(n6514), .CK(CLK), .QN(n22523) );
  DFF_X1 \REGISTERS_reg[24][47]  ( .D(n6513), .CK(CLK), .QN(n22524) );
  DFF_X1 \REGISTERS_reg[24][46]  ( .D(n6512), .CK(CLK), .QN(n22525) );
  DFF_X1 \REGISTERS_reg[24][45]  ( .D(n6511), .CK(CLK), .QN(n22526) );
  DFF_X1 \REGISTERS_reg[24][44]  ( .D(n6510), .CK(CLK), .QN(n22527) );
  DFF_X1 \REGISTERS_reg[24][43]  ( .D(n6509), .CK(CLK), .QN(n22528) );
  DFF_X1 \REGISTERS_reg[24][42]  ( .D(n6508), .CK(CLK), .QN(n22529) );
  DFF_X1 \REGISTERS_reg[24][41]  ( .D(n6507), .CK(CLK), .QN(n22530) );
  DFF_X1 \REGISTERS_reg[24][40]  ( .D(n6506), .CK(CLK), .QN(n22531) );
  DFF_X1 \REGISTERS_reg[24][39]  ( .D(n6505), .CK(CLK), .QN(n22532) );
  DFF_X1 \REGISTERS_reg[24][38]  ( .D(n6504), .CK(CLK), .QN(n22533) );
  DFF_X1 \REGISTERS_reg[24][37]  ( .D(n6503), .CK(CLK), .QN(n22534) );
  DFF_X1 \REGISTERS_reg[24][36]  ( .D(n6502), .CK(CLK), .QN(n22535) );
  DFF_X1 \REGISTERS_reg[24][35]  ( .D(n6501), .CK(CLK), .QN(n22536) );
  DFF_X1 \REGISTERS_reg[24][34]  ( .D(n6500), .CK(CLK), .QN(n22537) );
  DFF_X1 \REGISTERS_reg[24][33]  ( .D(n6499), .CK(CLK), .QN(n22538) );
  DFF_X1 \REGISTERS_reg[24][32]  ( .D(n6498), .CK(CLK), .QN(n22539) );
  DFF_X1 \REGISTERS_reg[24][31]  ( .D(n6497), .CK(CLK), .QN(n22540) );
  DFF_X1 \REGISTERS_reg[24][30]  ( .D(n6496), .CK(CLK), .QN(n22541) );
  DFF_X1 \REGISTERS_reg[24][29]  ( .D(n6495), .CK(CLK), .QN(n22542) );
  DFF_X1 \REGISTERS_reg[24][28]  ( .D(n6494), .CK(CLK), .QN(n22543) );
  DFF_X1 \REGISTERS_reg[24][27]  ( .D(n6493), .CK(CLK), .QN(n22544) );
  DFF_X1 \REGISTERS_reg[24][26]  ( .D(n6492), .CK(CLK), .QN(n22545) );
  DFF_X1 \REGISTERS_reg[24][25]  ( .D(n6491), .CK(CLK), .QN(n22546) );
  DFF_X1 \REGISTERS_reg[24][24]  ( .D(n6490), .CK(CLK), .QN(n22547) );
  DFF_X1 \REGISTERS_reg[24][23]  ( .D(n6489), .CK(CLK), .QN(n22548) );
  DFF_X1 \REGISTERS_reg[24][22]  ( .D(n6488), .CK(CLK), .QN(n22549) );
  DFF_X1 \REGISTERS_reg[24][21]  ( .D(n6487), .CK(CLK), .QN(n22550) );
  DFF_X1 \REGISTERS_reg[24][20]  ( .D(n6486), .CK(CLK), .QN(n22551) );
  DFF_X1 \REGISTERS_reg[24][19]  ( .D(n6485), .CK(CLK), .QN(n22552) );
  DFF_X1 \REGISTERS_reg[24][18]  ( .D(n6484), .CK(CLK), .QN(n22553) );
  DFF_X1 \REGISTERS_reg[24][17]  ( .D(n6483), .CK(CLK), .QN(n22554) );
  DFF_X1 \REGISTERS_reg[24][16]  ( .D(n6482), .CK(CLK), .QN(n22555) );
  DFF_X1 \REGISTERS_reg[24][15]  ( .D(n6481), .CK(CLK), .QN(n22556) );
  DFF_X1 \REGISTERS_reg[24][14]  ( .D(n6480), .CK(CLK), .QN(n22557) );
  DFF_X1 \REGISTERS_reg[24][13]  ( .D(n6479), .CK(CLK), .QN(n22558) );
  DFF_X1 \REGISTERS_reg[24][12]  ( .D(n6478), .CK(CLK), .QN(n22559) );
  DFF_X1 \REGISTERS_reg[24][11]  ( .D(n6477), .CK(CLK), .QN(n22560) );
  DFF_X1 \REGISTERS_reg[24][10]  ( .D(n6476), .CK(CLK), .QN(n22561) );
  DFF_X1 \REGISTERS_reg[24][9]  ( .D(n6475), .CK(CLK), .QN(n22562) );
  DFF_X1 \REGISTERS_reg[24][8]  ( .D(n6474), .CK(CLK), .QN(n22563) );
  DFF_X1 \REGISTERS_reg[24][7]  ( .D(n6473), .CK(CLK), .QN(n22564) );
  DFF_X1 \REGISTERS_reg[24][6]  ( .D(n6472), .CK(CLK), .QN(n22565) );
  DFF_X1 \REGISTERS_reg[24][5]  ( .D(n6471), .CK(CLK), .QN(n22566) );
  DFF_X1 \REGISTERS_reg[24][4]  ( .D(n6470), .CK(CLK), .QN(n22567) );
  DFF_X1 \REGISTERS_reg[24][3]  ( .D(n6469), .CK(CLK), .QN(n22568) );
  DFF_X1 \REGISTERS_reg[24][2]  ( .D(n6468), .CK(CLK), .QN(n22569) );
  DFF_X1 \REGISTERS_reg[24][1]  ( .D(n6467), .CK(CLK), .QN(n22570) );
  DFF_X1 \REGISTERS_reg[24][0]  ( .D(n6466), .CK(CLK), .QN(n22571) );
  DFF_X1 \REGISTERS_reg[23][59]  ( .D(n6589), .CK(CLK), .QN(n21300) );
  DFF_X1 \REGISTERS_reg[23][58]  ( .D(n6588), .CK(CLK), .QN(n21301) );
  DFF_X1 \REGISTERS_reg[23][57]  ( .D(n6587), .CK(CLK), .QN(n21302) );
  DFF_X1 \REGISTERS_reg[23][56]  ( .D(n6586), .CK(CLK), .QN(n21303) );
  DFF_X1 \REGISTERS_reg[23][55]  ( .D(n6585), .CK(CLK), .QN(n21304) );
  DFF_X1 \REGISTERS_reg[23][54]  ( .D(n6584), .CK(CLK), .QN(n21305) );
  DFF_X1 \REGISTERS_reg[23][53]  ( .D(n6583), .CK(CLK), .QN(n21306) );
  DFF_X1 \REGISTERS_reg[23][52]  ( .D(n6582), .CK(CLK), .QN(n21307) );
  DFF_X1 \REGISTERS_reg[23][51]  ( .D(n6581), .CK(CLK), .QN(n21308) );
  DFF_X1 \REGISTERS_reg[23][50]  ( .D(n6580), .CK(CLK), .QN(n21309) );
  DFF_X1 \REGISTERS_reg[23][49]  ( .D(n6579), .CK(CLK), .QN(n21310) );
  DFF_X1 \REGISTERS_reg[23][48]  ( .D(n6578), .CK(CLK), .QN(n21311) );
  DFF_X1 \REGISTERS_reg[23][47]  ( .D(n6577), .CK(CLK), .QN(n21312) );
  DFF_X1 \REGISTERS_reg[23][46]  ( .D(n6576), .CK(CLK), .QN(n21313) );
  DFF_X1 \REGISTERS_reg[23][45]  ( .D(n6575), .CK(CLK), .QN(n21314) );
  DFF_X1 \REGISTERS_reg[23][44]  ( .D(n6574), .CK(CLK), .QN(n21315) );
  DFF_X1 \REGISTERS_reg[23][43]  ( .D(n6573), .CK(CLK), .QN(n21316) );
  DFF_X1 \REGISTERS_reg[23][42]  ( .D(n6572), .CK(CLK), .QN(n21317) );
  DFF_X1 \REGISTERS_reg[23][41]  ( .D(n6571), .CK(CLK), .QN(n21318) );
  DFF_X1 \REGISTERS_reg[23][40]  ( .D(n6570), .CK(CLK), .QN(n21319) );
  DFF_X1 \REGISTERS_reg[23][39]  ( .D(n6569), .CK(CLK), .QN(n21320) );
  DFF_X1 \REGISTERS_reg[23][38]  ( .D(n6568), .CK(CLK), .QN(n21321) );
  DFF_X1 \REGISTERS_reg[23][37]  ( .D(n6567), .CK(CLK), .QN(n21322) );
  DFF_X1 \REGISTERS_reg[23][36]  ( .D(n6566), .CK(CLK), .QN(n21323) );
  DFF_X1 \REGISTERS_reg[23][35]  ( .D(n6565), .CK(CLK), .QN(n21324) );
  DFF_X1 \REGISTERS_reg[23][34]  ( .D(n6564), .CK(CLK), .QN(n21325) );
  DFF_X1 \REGISTERS_reg[23][33]  ( .D(n6563), .CK(CLK), .QN(n21326) );
  DFF_X1 \REGISTERS_reg[23][32]  ( .D(n6562), .CK(CLK), .QN(n21327) );
  DFF_X1 \REGISTERS_reg[23][31]  ( .D(n6561), .CK(CLK), .QN(n21328) );
  DFF_X1 \REGISTERS_reg[23][30]  ( .D(n6560), .CK(CLK), .QN(n21329) );
  DFF_X1 \REGISTERS_reg[23][29]  ( .D(n6559), .CK(CLK), .QN(n21330) );
  DFF_X1 \REGISTERS_reg[23][28]  ( .D(n6558), .CK(CLK), .QN(n21331) );
  DFF_X1 \REGISTERS_reg[23][27]  ( .D(n6557), .CK(CLK), .QN(n21332) );
  DFF_X1 \REGISTERS_reg[23][26]  ( .D(n6556), .CK(CLK), .QN(n21333) );
  DFF_X1 \REGISTERS_reg[23][25]  ( .D(n6555), .CK(CLK), .QN(n21334) );
  DFF_X1 \REGISTERS_reg[23][24]  ( .D(n6554), .CK(CLK), .QN(n21335) );
  DFF_X1 \REGISTERS_reg[23][23]  ( .D(n6553), .CK(CLK), .QN(n21336) );
  DFF_X1 \REGISTERS_reg[23][22]  ( .D(n6552), .CK(CLK), .QN(n21337) );
  DFF_X1 \REGISTERS_reg[23][21]  ( .D(n6551), .CK(CLK), .QN(n21338) );
  DFF_X1 \REGISTERS_reg[23][20]  ( .D(n6550), .CK(CLK), .QN(n21339) );
  DFF_X1 \REGISTERS_reg[23][19]  ( .D(n6549), .CK(CLK), .QN(n21340) );
  DFF_X1 \REGISTERS_reg[23][18]  ( .D(n6548), .CK(CLK), .QN(n21341) );
  DFF_X1 \REGISTERS_reg[23][17]  ( .D(n6547), .CK(CLK), .QN(n21342) );
  DFF_X1 \REGISTERS_reg[23][16]  ( .D(n6546), .CK(CLK), .QN(n21343) );
  DFF_X1 \REGISTERS_reg[23][15]  ( .D(n6545), .CK(CLK), .QN(n21344) );
  DFF_X1 \REGISTERS_reg[23][14]  ( .D(n6544), .CK(CLK), .QN(n21345) );
  DFF_X1 \REGISTERS_reg[23][13]  ( .D(n6543), .CK(CLK), .QN(n21346) );
  DFF_X1 \REGISTERS_reg[23][12]  ( .D(n6542), .CK(CLK), .QN(n21347) );
  DFF_X1 \REGISTERS_reg[23][11]  ( .D(n6541), .CK(CLK), .QN(n21348) );
  DFF_X1 \REGISTERS_reg[23][10]  ( .D(n6540), .CK(CLK), .QN(n21349) );
  DFF_X1 \REGISTERS_reg[23][9]  ( .D(n6539), .CK(CLK), .QN(n21350) );
  DFF_X1 \REGISTERS_reg[23][8]  ( .D(n6538), .CK(CLK), .QN(n21351) );
  DFF_X1 \REGISTERS_reg[23][7]  ( .D(n6537), .CK(CLK), .QN(n21352) );
  DFF_X1 \REGISTERS_reg[23][6]  ( .D(n6536), .CK(CLK), .QN(n21353) );
  DFF_X1 \REGISTERS_reg[23][5]  ( .D(n6535), .CK(CLK), .QN(n21354) );
  DFF_X1 \REGISTERS_reg[23][4]  ( .D(n6534), .CK(CLK), .QN(n21355) );
  DFF_X1 \REGISTERS_reg[23][3]  ( .D(n6533), .CK(CLK), .QN(n21356) );
  DFF_X1 \REGISTERS_reg[23][2]  ( .D(n6532), .CK(CLK), .QN(n21357) );
  DFF_X1 \REGISTERS_reg[23][1]  ( .D(n6531), .CK(CLK), .QN(n21358) );
  DFF_X1 \REGISTERS_reg[23][0]  ( .D(n6530), .CK(CLK), .QN(n21359) );
  DFF_X1 \REGISTERS_reg[17][59]  ( .D(n6973), .CK(CLK), .QN(n21700) );
  DFF_X1 \REGISTERS_reg[17][58]  ( .D(n6972), .CK(CLK), .QN(n21701) );
  DFF_X1 \REGISTERS_reg[17][57]  ( .D(n6971), .CK(CLK), .QN(n21702) );
  DFF_X1 \REGISTERS_reg[17][56]  ( .D(n6970), .CK(CLK), .QN(n21703) );
  DFF_X1 \REGISTERS_reg[17][55]  ( .D(n6969), .CK(CLK), .QN(n21704) );
  DFF_X1 \REGISTERS_reg[17][54]  ( .D(n6968), .CK(CLK), .QN(n21705) );
  DFF_X1 \REGISTERS_reg[17][53]  ( .D(n6967), .CK(CLK), .QN(n21706) );
  DFF_X1 \REGISTERS_reg[17][52]  ( .D(n6966), .CK(CLK), .QN(n21707) );
  DFF_X1 \REGISTERS_reg[17][51]  ( .D(n6965), .CK(CLK), .QN(n21708) );
  DFF_X1 \REGISTERS_reg[17][50]  ( .D(n6964), .CK(CLK), .QN(n21709) );
  DFF_X1 \REGISTERS_reg[17][49]  ( .D(n6963), .CK(CLK), .QN(n21710) );
  DFF_X1 \REGISTERS_reg[17][48]  ( .D(n6962), .CK(CLK), .QN(n21711) );
  DFF_X1 \REGISTERS_reg[17][47]  ( .D(n6961), .CK(CLK), .QN(n21712) );
  DFF_X1 \REGISTERS_reg[17][46]  ( .D(n6960), .CK(CLK), .QN(n21713) );
  DFF_X1 \REGISTERS_reg[17][45]  ( .D(n6959), .CK(CLK), .QN(n21714) );
  DFF_X1 \REGISTERS_reg[17][44]  ( .D(n6958), .CK(CLK), .QN(n21715) );
  DFF_X1 \REGISTERS_reg[17][43]  ( .D(n6957), .CK(CLK), .QN(n21716) );
  DFF_X1 \REGISTERS_reg[17][42]  ( .D(n6956), .CK(CLK), .QN(n21717) );
  DFF_X1 \REGISTERS_reg[17][41]  ( .D(n6955), .CK(CLK), .QN(n21718) );
  DFF_X1 \REGISTERS_reg[17][40]  ( .D(n6954), .CK(CLK), .QN(n21719) );
  DFF_X1 \REGISTERS_reg[17][39]  ( .D(n6953), .CK(CLK), .QN(n21720) );
  DFF_X1 \REGISTERS_reg[17][38]  ( .D(n6952), .CK(CLK), .QN(n21721) );
  DFF_X1 \REGISTERS_reg[17][37]  ( .D(n6951), .CK(CLK), .QN(n21722) );
  DFF_X1 \REGISTERS_reg[17][36]  ( .D(n6950), .CK(CLK), .QN(n21723) );
  DFF_X1 \REGISTERS_reg[17][35]  ( .D(n6949), .CK(CLK), .QN(n21724) );
  DFF_X1 \REGISTERS_reg[17][34]  ( .D(n6948), .CK(CLK), .QN(n21725) );
  DFF_X1 \REGISTERS_reg[17][33]  ( .D(n6947), .CK(CLK), .QN(n21726) );
  DFF_X1 \REGISTERS_reg[17][32]  ( .D(n6946), .CK(CLK), .QN(n21727) );
  DFF_X1 \REGISTERS_reg[17][31]  ( .D(n6945), .CK(CLK), .QN(n21728) );
  DFF_X1 \REGISTERS_reg[17][30]  ( .D(n6944), .CK(CLK), .QN(n21729) );
  DFF_X1 \REGISTERS_reg[17][29]  ( .D(n6943), .CK(CLK), .QN(n21730) );
  DFF_X1 \REGISTERS_reg[17][28]  ( .D(n6942), .CK(CLK), .QN(n21731) );
  DFF_X1 \REGISTERS_reg[17][27]  ( .D(n6941), .CK(CLK), .QN(n21732) );
  DFF_X1 \REGISTERS_reg[17][26]  ( .D(n6940), .CK(CLK), .QN(n21733) );
  DFF_X1 \REGISTERS_reg[17][25]  ( .D(n6939), .CK(CLK), .QN(n21734) );
  DFF_X1 \REGISTERS_reg[17][24]  ( .D(n6938), .CK(CLK), .QN(n21735) );
  DFF_X1 \REGISTERS_reg[17][23]  ( .D(n6937), .CK(CLK), .QN(n21736) );
  DFF_X1 \REGISTERS_reg[17][22]  ( .D(n6936), .CK(CLK), .QN(n21737) );
  DFF_X1 \REGISTERS_reg[17][21]  ( .D(n6935), .CK(CLK), .QN(n21738) );
  DFF_X1 \REGISTERS_reg[17][20]  ( .D(n6934), .CK(CLK), .QN(n21739) );
  DFF_X1 \REGISTERS_reg[17][19]  ( .D(n6933), .CK(CLK), .QN(n21740) );
  DFF_X1 \REGISTERS_reg[17][18]  ( .D(n6932), .CK(CLK), .QN(n21741) );
  DFF_X1 \REGISTERS_reg[17][17]  ( .D(n6931), .CK(CLK), .QN(n21742) );
  DFF_X1 \REGISTERS_reg[17][16]  ( .D(n6930), .CK(CLK), .QN(n21743) );
  DFF_X1 \REGISTERS_reg[17][15]  ( .D(n6929), .CK(CLK), .QN(n21744) );
  DFF_X1 \REGISTERS_reg[17][14]  ( .D(n6928), .CK(CLK), .QN(n21745) );
  DFF_X1 \REGISTERS_reg[17][13]  ( .D(n6927), .CK(CLK), .QN(n21746) );
  DFF_X1 \REGISTERS_reg[17][12]  ( .D(n6926), .CK(CLK), .QN(n21747) );
  DFF_X1 \REGISTERS_reg[17][11]  ( .D(n6925), .CK(CLK), .QN(n21748) );
  DFF_X1 \REGISTERS_reg[17][10]  ( .D(n6924), .CK(CLK), .QN(n21749) );
  DFF_X1 \REGISTERS_reg[17][9]  ( .D(n6923), .CK(CLK), .QN(n21750) );
  DFF_X1 \REGISTERS_reg[17][8]  ( .D(n6922), .CK(CLK), .QN(n21751) );
  DFF_X1 \REGISTERS_reg[17][7]  ( .D(n6921), .CK(CLK), .QN(n21752) );
  DFF_X1 \REGISTERS_reg[17][6]  ( .D(n6920), .CK(CLK), .QN(n21753) );
  DFF_X1 \REGISTERS_reg[17][5]  ( .D(n6919), .CK(CLK), .QN(n21754) );
  DFF_X1 \REGISTERS_reg[17][4]  ( .D(n6918), .CK(CLK), .QN(n21755) );
  DFF_X1 \REGISTERS_reg[17][3]  ( .D(n6917), .CK(CLK), .QN(n21756) );
  DFF_X1 \REGISTERS_reg[17][2]  ( .D(n6916), .CK(CLK), .QN(n21757) );
  DFF_X1 \REGISTERS_reg[17][1]  ( .D(n6915), .CK(CLK), .QN(n21758) );
  DFF_X1 \REGISTERS_reg[17][0]  ( .D(n6914), .CK(CLK), .QN(n21759) );
  DFF_X1 \REGISTERS_reg[12][59]  ( .D(n7293), .CK(CLK), .QN(n20712) );
  DFF_X1 \REGISTERS_reg[12][58]  ( .D(n7292), .CK(CLK), .QN(n20713) );
  DFF_X1 \REGISTERS_reg[12][57]  ( .D(n7291), .CK(CLK), .QN(n20714) );
  DFF_X1 \REGISTERS_reg[12][56]  ( .D(n7290), .CK(CLK), .QN(n20715) );
  DFF_X1 \REGISTERS_reg[12][55]  ( .D(n7289), .CK(CLK), .QN(n20716) );
  DFF_X1 \REGISTERS_reg[12][54]  ( .D(n7288), .CK(CLK), .QN(n20717) );
  DFF_X1 \REGISTERS_reg[12][53]  ( .D(n7287), .CK(CLK), .QN(n20718) );
  DFF_X1 \REGISTERS_reg[12][52]  ( .D(n7286), .CK(CLK), .QN(n20719) );
  DFF_X1 \REGISTERS_reg[12][51]  ( .D(n7285), .CK(CLK), .QN(n20720) );
  DFF_X1 \REGISTERS_reg[12][50]  ( .D(n7284), .CK(CLK), .QN(n20721) );
  DFF_X1 \REGISTERS_reg[12][49]  ( .D(n7283), .CK(CLK), .QN(n20722) );
  DFF_X1 \REGISTERS_reg[12][48]  ( .D(n7282), .CK(CLK), .QN(n20723) );
  DFF_X1 \REGISTERS_reg[12][47]  ( .D(n7281), .CK(CLK), .QN(n20724) );
  DFF_X1 \REGISTERS_reg[12][46]  ( .D(n7280), .CK(CLK), .QN(n20725) );
  DFF_X1 \REGISTERS_reg[12][45]  ( .D(n7279), .CK(CLK), .QN(n20726) );
  DFF_X1 \REGISTERS_reg[12][44]  ( .D(n7278), .CK(CLK), .QN(n20727) );
  DFF_X1 \REGISTERS_reg[12][43]  ( .D(n7277), .CK(CLK), .QN(n20728) );
  DFF_X1 \REGISTERS_reg[12][42]  ( .D(n7276), .CK(CLK), .QN(n20729) );
  DFF_X1 \REGISTERS_reg[12][41]  ( .D(n7275), .CK(CLK), .QN(n20730) );
  DFF_X1 \REGISTERS_reg[12][40]  ( .D(n7274), .CK(CLK), .QN(n20731) );
  DFF_X1 \REGISTERS_reg[12][39]  ( .D(n7273), .CK(CLK), .QN(n20732) );
  DFF_X1 \REGISTERS_reg[12][38]  ( .D(n7272), .CK(CLK), .QN(n20733) );
  DFF_X1 \REGISTERS_reg[12][37]  ( .D(n7271), .CK(CLK), .QN(n20734) );
  DFF_X1 \REGISTERS_reg[12][36]  ( .D(n7270), .CK(CLK), .QN(n20735) );
  DFF_X1 \REGISTERS_reg[12][35]  ( .D(n7269), .CK(CLK), .QN(n20736) );
  DFF_X1 \REGISTERS_reg[12][34]  ( .D(n7268), .CK(CLK), .QN(n20737) );
  DFF_X1 \REGISTERS_reg[12][33]  ( .D(n7267), .CK(CLK), .QN(n20738) );
  DFF_X1 \REGISTERS_reg[12][32]  ( .D(n7266), .CK(CLK), .QN(n20739) );
  DFF_X1 \REGISTERS_reg[12][31]  ( .D(n7265), .CK(CLK), .QN(n20740) );
  DFF_X1 \REGISTERS_reg[12][30]  ( .D(n7264), .CK(CLK), .QN(n20741) );
  DFF_X1 \REGISTERS_reg[12][29]  ( .D(n7263), .CK(CLK), .QN(n20742) );
  DFF_X1 \REGISTERS_reg[12][28]  ( .D(n7262), .CK(CLK), .QN(n20743) );
  DFF_X1 \REGISTERS_reg[12][27]  ( .D(n7261), .CK(CLK), .QN(n20744) );
  DFF_X1 \REGISTERS_reg[12][26]  ( .D(n7260), .CK(CLK), .QN(n20745) );
  DFF_X1 \REGISTERS_reg[12][25]  ( .D(n7259), .CK(CLK), .QN(n20746) );
  DFF_X1 \REGISTERS_reg[12][24]  ( .D(n7258), .CK(CLK), .QN(n20747) );
  DFF_X1 \REGISTERS_reg[12][23]  ( .D(n7257), .CK(CLK), .QN(n20748) );
  DFF_X1 \REGISTERS_reg[12][22]  ( .D(n7256), .CK(CLK), .QN(n20749) );
  DFF_X1 \REGISTERS_reg[12][21]  ( .D(n7255), .CK(CLK), .QN(n20750) );
  DFF_X1 \REGISTERS_reg[12][20]  ( .D(n7254), .CK(CLK), .QN(n20751) );
  DFF_X1 \REGISTERS_reg[12][19]  ( .D(n7253), .CK(CLK), .QN(n20752) );
  DFF_X1 \REGISTERS_reg[12][18]  ( .D(n7252), .CK(CLK), .QN(n20753) );
  DFF_X1 \REGISTERS_reg[12][17]  ( .D(n7251), .CK(CLK), .QN(n20754) );
  DFF_X1 \REGISTERS_reg[12][16]  ( .D(n7250), .CK(CLK), .QN(n20755) );
  DFF_X1 \REGISTERS_reg[12][15]  ( .D(n7249), .CK(CLK), .QN(n20756) );
  DFF_X1 \REGISTERS_reg[12][14]  ( .D(n7248), .CK(CLK), .QN(n20757) );
  DFF_X1 \REGISTERS_reg[12][13]  ( .D(n7247), .CK(CLK), .QN(n20758) );
  DFF_X1 \REGISTERS_reg[12][12]  ( .D(n7246), .CK(CLK), .QN(n20759) );
  DFF_X1 \REGISTERS_reg[12][11]  ( .D(n7245), .CK(CLK), .QN(n20760) );
  DFF_X1 \REGISTERS_reg[12][10]  ( .D(n7244), .CK(CLK), .QN(n20761) );
  DFF_X1 \REGISTERS_reg[12][9]  ( .D(n7243), .CK(CLK), .QN(n20762) );
  DFF_X1 \REGISTERS_reg[12][8]  ( .D(n7242), .CK(CLK), .QN(n20763) );
  DFF_X1 \REGISTERS_reg[12][7]  ( .D(n7241), .CK(CLK), .QN(n20764) );
  DFF_X1 \REGISTERS_reg[12][6]  ( .D(n7240), .CK(CLK), .QN(n20765) );
  DFF_X1 \REGISTERS_reg[12][5]  ( .D(n7239), .CK(CLK), .QN(n20766) );
  DFF_X1 \REGISTERS_reg[12][4]  ( .D(n7238), .CK(CLK), .QN(n20767) );
  DFF_X1 \REGISTERS_reg[12][3]  ( .D(n7237), .CK(CLK), .QN(n20768) );
  DFF_X1 \REGISTERS_reg[12][2]  ( .D(n7236), .CK(CLK), .QN(n20769) );
  DFF_X1 \REGISTERS_reg[12][1]  ( .D(n7235), .CK(CLK), .QN(n20770) );
  DFF_X1 \REGISTERS_reg[12][0]  ( .D(n7234), .CK(CLK), .QN(n20771) );
  DFF_X1 \REGISTERS_reg[9][59]  ( .D(n7485), .CK(CLK), .QN(n22632) );
  DFF_X1 \REGISTERS_reg[9][58]  ( .D(n7484), .CK(CLK), .QN(n22633) );
  DFF_X1 \REGISTERS_reg[9][57]  ( .D(n7483), .CK(CLK), .QN(n22634) );
  DFF_X1 \REGISTERS_reg[9][56]  ( .D(n7482), .CK(CLK), .QN(n22635) );
  DFF_X1 \REGISTERS_reg[9][55]  ( .D(n7481), .CK(CLK), .QN(n22636) );
  DFF_X1 \REGISTERS_reg[9][54]  ( .D(n7480), .CK(CLK), .QN(n22637) );
  DFF_X1 \REGISTERS_reg[9][53]  ( .D(n7479), .CK(CLK), .QN(n22638) );
  DFF_X1 \REGISTERS_reg[9][52]  ( .D(n7478), .CK(CLK), .QN(n22639) );
  DFF_X1 \REGISTERS_reg[9][51]  ( .D(n7477), .CK(CLK), .QN(n22640) );
  DFF_X1 \REGISTERS_reg[9][50]  ( .D(n7476), .CK(CLK), .QN(n22641) );
  DFF_X1 \REGISTERS_reg[9][49]  ( .D(n7475), .CK(CLK), .QN(n22642) );
  DFF_X1 \REGISTERS_reg[9][48]  ( .D(n7474), .CK(CLK), .QN(n22643) );
  DFF_X1 \REGISTERS_reg[9][47]  ( .D(n7473), .CK(CLK), .QN(n22644) );
  DFF_X1 \REGISTERS_reg[9][46]  ( .D(n7472), .CK(CLK), .QN(n22645) );
  DFF_X1 \REGISTERS_reg[9][45]  ( .D(n7471), .CK(CLK), .QN(n22646) );
  DFF_X1 \REGISTERS_reg[9][44]  ( .D(n7470), .CK(CLK), .QN(n22647) );
  DFF_X1 \REGISTERS_reg[9][43]  ( .D(n7469), .CK(CLK), .QN(n22648) );
  DFF_X1 \REGISTERS_reg[9][42]  ( .D(n7468), .CK(CLK), .QN(n22649) );
  DFF_X1 \REGISTERS_reg[9][41]  ( .D(n7467), .CK(CLK), .QN(n22650) );
  DFF_X1 \REGISTERS_reg[9][40]  ( .D(n7466), .CK(CLK), .QN(n22651) );
  DFF_X1 \REGISTERS_reg[9][39]  ( .D(n7465), .CK(CLK), .QN(n22652) );
  DFF_X1 \REGISTERS_reg[9][38]  ( .D(n7464), .CK(CLK), .QN(n22653) );
  DFF_X1 \REGISTERS_reg[9][37]  ( .D(n7463), .CK(CLK), .QN(n22654) );
  DFF_X1 \REGISTERS_reg[9][36]  ( .D(n7462), .CK(CLK), .QN(n22655) );
  DFF_X1 \REGISTERS_reg[9][35]  ( .D(n7461), .CK(CLK), .QN(n22656) );
  DFF_X1 \REGISTERS_reg[9][34]  ( .D(n7460), .CK(CLK), .QN(n22657) );
  DFF_X1 \REGISTERS_reg[9][33]  ( .D(n7459), .CK(CLK), .QN(n22658) );
  DFF_X1 \REGISTERS_reg[9][32]  ( .D(n7458), .CK(CLK), .QN(n22659) );
  DFF_X1 \REGISTERS_reg[9][31]  ( .D(n7457), .CK(CLK), .QN(n22660) );
  DFF_X1 \REGISTERS_reg[9][30]  ( .D(n7456), .CK(CLK), .QN(n22661) );
  DFF_X1 \REGISTERS_reg[9][29]  ( .D(n7455), .CK(CLK), .QN(n22662) );
  DFF_X1 \REGISTERS_reg[9][28]  ( .D(n7454), .CK(CLK), .QN(n22663) );
  DFF_X1 \REGISTERS_reg[9][27]  ( .D(n7453), .CK(CLK), .QN(n22664) );
  DFF_X1 \REGISTERS_reg[9][26]  ( .D(n7452), .CK(CLK), .QN(n22665) );
  DFF_X1 \REGISTERS_reg[9][25]  ( .D(n7451), .CK(CLK), .QN(n22666) );
  DFF_X1 \REGISTERS_reg[9][24]  ( .D(n7450), .CK(CLK), .QN(n22667) );
  DFF_X1 \REGISTERS_reg[9][23]  ( .D(n7449), .CK(CLK), .QN(n22668) );
  DFF_X1 \REGISTERS_reg[9][22]  ( .D(n7448), .CK(CLK), .QN(n22669) );
  DFF_X1 \REGISTERS_reg[9][21]  ( .D(n7447), .CK(CLK), .QN(n22670) );
  DFF_X1 \REGISTERS_reg[9][20]  ( .D(n7446), .CK(CLK), .QN(n22671) );
  DFF_X1 \REGISTERS_reg[9][19]  ( .D(n7445), .CK(CLK), .QN(n22672) );
  DFF_X1 \REGISTERS_reg[9][18]  ( .D(n7444), .CK(CLK), .QN(n22673) );
  DFF_X1 \REGISTERS_reg[9][17]  ( .D(n7443), .CK(CLK), .QN(n22674) );
  DFF_X1 \REGISTERS_reg[9][16]  ( .D(n7442), .CK(CLK), .QN(n22675) );
  DFF_X1 \REGISTERS_reg[9][15]  ( .D(n7441), .CK(CLK), .QN(n22676) );
  DFF_X1 \REGISTERS_reg[9][14]  ( .D(n7440), .CK(CLK), .QN(n22677) );
  DFF_X1 \REGISTERS_reg[9][13]  ( .D(n7439), .CK(CLK), .QN(n22678) );
  DFF_X1 \REGISTERS_reg[9][12]  ( .D(n7438), .CK(CLK), .QN(n22679) );
  DFF_X1 \REGISTERS_reg[9][11]  ( .D(n7437), .CK(CLK), .QN(n22680) );
  DFF_X1 \REGISTERS_reg[9][10]  ( .D(n7436), .CK(CLK), .QN(n22681) );
  DFF_X1 \REGISTERS_reg[9][9]  ( .D(n7435), .CK(CLK), .QN(n22682) );
  DFF_X1 \REGISTERS_reg[9][8]  ( .D(n7434), .CK(CLK), .QN(n22683) );
  DFF_X1 \REGISTERS_reg[9][7]  ( .D(n7433), .CK(CLK), .QN(n22684) );
  DFF_X1 \REGISTERS_reg[9][6]  ( .D(n7432), .CK(CLK), .QN(n22685) );
  DFF_X1 \REGISTERS_reg[9][5]  ( .D(n7431), .CK(CLK), .QN(n22686) );
  DFF_X1 \REGISTERS_reg[9][4]  ( .D(n7430), .CK(CLK), .QN(n22687) );
  DFF_X1 \REGISTERS_reg[9][3]  ( .D(n7429), .CK(CLK), .QN(n22688) );
  DFF_X1 \REGISTERS_reg[9][2]  ( .D(n7428), .CK(CLK), .QN(n22689) );
  DFF_X1 \REGISTERS_reg[9][1]  ( .D(n7427), .CK(CLK), .QN(n22690) );
  DFF_X1 \REGISTERS_reg[9][0]  ( .D(n7426), .CK(CLK), .QN(n22691) );
  DFF_X1 \REGISTERS_reg[7][59]  ( .D(n7613), .CK(CLK), .QN(n22000) );
  DFF_X1 \REGISTERS_reg[7][58]  ( .D(n7612), .CK(CLK), .QN(n22001) );
  DFF_X1 \REGISTERS_reg[7][57]  ( .D(n7611), .CK(CLK), .QN(n22002) );
  DFF_X1 \REGISTERS_reg[7][56]  ( .D(n7610), .CK(CLK), .QN(n22003) );
  DFF_X1 \REGISTERS_reg[7][55]  ( .D(n7609), .CK(CLK), .QN(n22004) );
  DFF_X1 \REGISTERS_reg[7][54]  ( .D(n7608), .CK(CLK), .QN(n22005) );
  DFF_X1 \REGISTERS_reg[7][53]  ( .D(n7607), .CK(CLK), .QN(n22006) );
  DFF_X1 \REGISTERS_reg[7][52]  ( .D(n7606), .CK(CLK), .QN(n22007) );
  DFF_X1 \REGISTERS_reg[7][51]  ( .D(n7605), .CK(CLK), .QN(n22008) );
  DFF_X1 \REGISTERS_reg[7][50]  ( .D(n7604), .CK(CLK), .QN(n22009) );
  DFF_X1 \REGISTERS_reg[7][49]  ( .D(n7603), .CK(CLK), .QN(n22010) );
  DFF_X1 \REGISTERS_reg[7][48]  ( .D(n7602), .CK(CLK), .QN(n22011) );
  DFF_X1 \REGISTERS_reg[7][47]  ( .D(n7601), .CK(CLK), .QN(n22012) );
  DFF_X1 \REGISTERS_reg[7][46]  ( .D(n7600), .CK(CLK), .QN(n22013) );
  DFF_X1 \REGISTERS_reg[7][45]  ( .D(n7599), .CK(CLK), .QN(n22014) );
  DFF_X1 \REGISTERS_reg[7][44]  ( .D(n7598), .CK(CLK), .QN(n22015) );
  DFF_X1 \REGISTERS_reg[7][43]  ( .D(n7597), .CK(CLK), .QN(n22016) );
  DFF_X1 \REGISTERS_reg[7][42]  ( .D(n7596), .CK(CLK), .QN(n22017) );
  DFF_X1 \REGISTERS_reg[7][41]  ( .D(n7595), .CK(CLK), .QN(n22018) );
  DFF_X1 \REGISTERS_reg[7][40]  ( .D(n7594), .CK(CLK), .QN(n22019) );
  DFF_X1 \REGISTERS_reg[7][39]  ( .D(n7593), .CK(CLK), .QN(n22020) );
  DFF_X1 \REGISTERS_reg[7][38]  ( .D(n7592), .CK(CLK), .QN(n22021) );
  DFF_X1 \REGISTERS_reg[7][37]  ( .D(n7591), .CK(CLK), .QN(n22022) );
  DFF_X1 \REGISTERS_reg[7][36]  ( .D(n7590), .CK(CLK), .QN(n22023) );
  DFF_X1 \REGISTERS_reg[7][35]  ( .D(n7589), .CK(CLK), .QN(n22024) );
  DFF_X1 \REGISTERS_reg[7][34]  ( .D(n7588), .CK(CLK), .QN(n22025) );
  DFF_X1 \REGISTERS_reg[7][33]  ( .D(n7587), .CK(CLK), .QN(n22026) );
  DFF_X1 \REGISTERS_reg[7][32]  ( .D(n7586), .CK(CLK), .QN(n22027) );
  DFF_X1 \REGISTERS_reg[7][31]  ( .D(n7585), .CK(CLK), .QN(n22028) );
  DFF_X1 \REGISTERS_reg[7][30]  ( .D(n7584), .CK(CLK), .QN(n22029) );
  DFF_X1 \REGISTERS_reg[7][29]  ( .D(n7583), .CK(CLK), .QN(n22030) );
  DFF_X1 \REGISTERS_reg[7][28]  ( .D(n7582), .CK(CLK), .QN(n22031) );
  DFF_X1 \REGISTERS_reg[7][27]  ( .D(n7581), .CK(CLK), .QN(n22032) );
  DFF_X1 \REGISTERS_reg[7][26]  ( .D(n7580), .CK(CLK), .QN(n22033) );
  DFF_X1 \REGISTERS_reg[7][25]  ( .D(n7579), .CK(CLK), .QN(n22034) );
  DFF_X1 \REGISTERS_reg[7][24]  ( .D(n7578), .CK(CLK), .QN(n22035) );
  DFF_X1 \REGISTERS_reg[7][23]  ( .D(n7577), .CK(CLK), .QN(n22036) );
  DFF_X1 \REGISTERS_reg[7][22]  ( .D(n7576), .CK(CLK), .QN(n22037) );
  DFF_X1 \REGISTERS_reg[7][21]  ( .D(n7575), .CK(CLK), .QN(n22038) );
  DFF_X1 \REGISTERS_reg[7][20]  ( .D(n7574), .CK(CLK), .QN(n22039) );
  DFF_X1 \REGISTERS_reg[7][19]  ( .D(n7573), .CK(CLK), .QN(n22040) );
  DFF_X1 \REGISTERS_reg[7][18]  ( .D(n7572), .CK(CLK), .QN(n22041) );
  DFF_X1 \REGISTERS_reg[7][17]  ( .D(n7571), .CK(CLK), .QN(n22042) );
  DFF_X1 \REGISTERS_reg[7][16]  ( .D(n7570), .CK(CLK), .QN(n22043) );
  DFF_X1 \REGISTERS_reg[7][15]  ( .D(n7569), .CK(CLK), .QN(n22044) );
  DFF_X1 \REGISTERS_reg[7][14]  ( .D(n7568), .CK(CLK), .QN(n22045) );
  DFF_X1 \REGISTERS_reg[7][13]  ( .D(n7567), .CK(CLK), .QN(n22046) );
  DFF_X1 \REGISTERS_reg[7][12]  ( .D(n7566), .CK(CLK), .QN(n22047) );
  DFF_X1 \REGISTERS_reg[7][11]  ( .D(n7565), .CK(CLK), .QN(n22048) );
  DFF_X1 \REGISTERS_reg[7][10]  ( .D(n7564), .CK(CLK), .QN(n22049) );
  DFF_X1 \REGISTERS_reg[7][9]  ( .D(n7563), .CK(CLK), .QN(n22050) );
  DFF_X1 \REGISTERS_reg[7][8]  ( .D(n7562), .CK(CLK), .QN(n22051) );
  DFF_X1 \REGISTERS_reg[7][7]  ( .D(n7561), .CK(CLK), .QN(n22052) );
  DFF_X1 \REGISTERS_reg[7][6]  ( .D(n7560), .CK(CLK), .QN(n22053) );
  DFF_X1 \REGISTERS_reg[7][5]  ( .D(n7559), .CK(CLK), .QN(n22054) );
  DFF_X1 \REGISTERS_reg[7][4]  ( .D(n7558), .CK(CLK), .QN(n22055) );
  DFF_X1 \REGISTERS_reg[7][3]  ( .D(n7557), .CK(CLK), .QN(n22056) );
  DFF_X1 \REGISTERS_reg[7][2]  ( .D(n7556), .CK(CLK), .QN(n22057) );
  DFF_X1 \REGISTERS_reg[7][1]  ( .D(n7555), .CK(CLK), .QN(n22058) );
  DFF_X1 \REGISTERS_reg[7][0]  ( .D(n7554), .CK(CLK), .QN(n22059) );
  DFF_X1 \REGISTERS_reg[5][59]  ( .D(n7741), .CK(CLK), .QN(n21520) );
  DFF_X1 \REGISTERS_reg[5][58]  ( .D(n7740), .CK(CLK), .QN(n21521) );
  DFF_X1 \REGISTERS_reg[5][57]  ( .D(n7739), .CK(CLK), .QN(n21522) );
  DFF_X1 \REGISTERS_reg[5][56]  ( .D(n7738), .CK(CLK), .QN(n21523) );
  DFF_X1 \REGISTERS_reg[5][55]  ( .D(n7737), .CK(CLK), .QN(n21524) );
  DFF_X1 \REGISTERS_reg[5][54]  ( .D(n7736), .CK(CLK), .QN(n21525) );
  DFF_X1 \REGISTERS_reg[5][53]  ( .D(n7735), .CK(CLK), .QN(n21526) );
  DFF_X1 \REGISTERS_reg[5][52]  ( .D(n7734), .CK(CLK), .QN(n21527) );
  DFF_X1 \REGISTERS_reg[5][51]  ( .D(n7733), .CK(CLK), .QN(n21528) );
  DFF_X1 \REGISTERS_reg[5][50]  ( .D(n7732), .CK(CLK), .QN(n21529) );
  DFF_X1 \REGISTERS_reg[5][49]  ( .D(n7731), .CK(CLK), .QN(n21530) );
  DFF_X1 \REGISTERS_reg[5][48]  ( .D(n7730), .CK(CLK), .QN(n21531) );
  DFF_X1 \REGISTERS_reg[5][47]  ( .D(n7729), .CK(CLK), .QN(n21532) );
  DFF_X1 \REGISTERS_reg[5][46]  ( .D(n7728), .CK(CLK), .QN(n21533) );
  DFF_X1 \REGISTERS_reg[5][45]  ( .D(n7727), .CK(CLK), .QN(n21534) );
  DFF_X1 \REGISTERS_reg[5][44]  ( .D(n7726), .CK(CLK), .QN(n21535) );
  DFF_X1 \REGISTERS_reg[5][43]  ( .D(n7725), .CK(CLK), .QN(n21536) );
  DFF_X1 \REGISTERS_reg[5][42]  ( .D(n7724), .CK(CLK), .QN(n21537) );
  DFF_X1 \REGISTERS_reg[5][41]  ( .D(n7723), .CK(CLK), .QN(n21538) );
  DFF_X1 \REGISTERS_reg[5][40]  ( .D(n7722), .CK(CLK), .QN(n21539) );
  DFF_X1 \REGISTERS_reg[5][39]  ( .D(n7721), .CK(CLK), .QN(n21540) );
  DFF_X1 \REGISTERS_reg[5][38]  ( .D(n7720), .CK(CLK), .QN(n21541) );
  DFF_X1 \REGISTERS_reg[5][37]  ( .D(n7719), .CK(CLK), .QN(n21542) );
  DFF_X1 \REGISTERS_reg[5][36]  ( .D(n7718), .CK(CLK), .QN(n21543) );
  DFF_X1 \REGISTERS_reg[5][35]  ( .D(n7717), .CK(CLK), .QN(n21544) );
  DFF_X1 \REGISTERS_reg[5][34]  ( .D(n7716), .CK(CLK), .QN(n21545) );
  DFF_X1 \REGISTERS_reg[5][33]  ( .D(n7715), .CK(CLK), .QN(n21546) );
  DFF_X1 \REGISTERS_reg[5][32]  ( .D(n7714), .CK(CLK), .QN(n21547) );
  DFF_X1 \REGISTERS_reg[5][31]  ( .D(n7713), .CK(CLK), .QN(n21548) );
  DFF_X1 \REGISTERS_reg[5][30]  ( .D(n7712), .CK(CLK), .QN(n21549) );
  DFF_X1 \REGISTERS_reg[5][29]  ( .D(n7711), .CK(CLK), .QN(n21550) );
  DFF_X1 \REGISTERS_reg[5][28]  ( .D(n7710), .CK(CLK), .QN(n21551) );
  DFF_X1 \REGISTERS_reg[5][27]  ( .D(n7709), .CK(CLK), .QN(n21552) );
  DFF_X1 \REGISTERS_reg[5][26]  ( .D(n7708), .CK(CLK), .QN(n21553) );
  DFF_X1 \REGISTERS_reg[5][25]  ( .D(n7707), .CK(CLK), .QN(n21554) );
  DFF_X1 \REGISTERS_reg[5][24]  ( .D(n7706), .CK(CLK), .QN(n21555) );
  DFF_X1 \REGISTERS_reg[5][23]  ( .D(n7705), .CK(CLK), .QN(n21556) );
  DFF_X1 \REGISTERS_reg[5][22]  ( .D(n7704), .CK(CLK), .QN(n21557) );
  DFF_X1 \REGISTERS_reg[5][21]  ( .D(n7703), .CK(CLK), .QN(n21558) );
  DFF_X1 \REGISTERS_reg[5][20]  ( .D(n7702), .CK(CLK), .QN(n21559) );
  DFF_X1 \REGISTERS_reg[5][19]  ( .D(n7701), .CK(CLK), .QN(n21560) );
  DFF_X1 \REGISTERS_reg[5][18]  ( .D(n7700), .CK(CLK), .QN(n21561) );
  DFF_X1 \REGISTERS_reg[5][17]  ( .D(n7699), .CK(CLK), .QN(n21562) );
  DFF_X1 \REGISTERS_reg[5][16]  ( .D(n7698), .CK(CLK), .QN(n21563) );
  DFF_X1 \REGISTERS_reg[5][15]  ( .D(n7697), .CK(CLK), .QN(n21564) );
  DFF_X1 \REGISTERS_reg[5][14]  ( .D(n7696), .CK(CLK), .QN(n21565) );
  DFF_X1 \REGISTERS_reg[5][13]  ( .D(n7695), .CK(CLK), .QN(n21566) );
  DFF_X1 \REGISTERS_reg[5][12]  ( .D(n7694), .CK(CLK), .QN(n21567) );
  DFF_X1 \REGISTERS_reg[5][11]  ( .D(n7693), .CK(CLK), .QN(n21568) );
  DFF_X1 \REGISTERS_reg[5][10]  ( .D(n7692), .CK(CLK), .QN(n21569) );
  DFF_X1 \REGISTERS_reg[5][9]  ( .D(n7691), .CK(CLK), .QN(n21570) );
  DFF_X1 \REGISTERS_reg[5][8]  ( .D(n7690), .CK(CLK), .QN(n21571) );
  DFF_X1 \REGISTERS_reg[5][7]  ( .D(n7689), .CK(CLK), .QN(n21572) );
  DFF_X1 \REGISTERS_reg[5][6]  ( .D(n7688), .CK(CLK), .QN(n21573) );
  DFF_X1 \REGISTERS_reg[5][5]  ( .D(n7687), .CK(CLK), .QN(n21574) );
  DFF_X1 \REGISTERS_reg[5][4]  ( .D(n7686), .CK(CLK), .QN(n21575) );
  DFF_X1 \REGISTERS_reg[5][3]  ( .D(n7685), .CK(CLK), .QN(n21576) );
  DFF_X1 \REGISTERS_reg[5][2]  ( .D(n7684), .CK(CLK), .QN(n21577) );
  DFF_X1 \REGISTERS_reg[5][1]  ( .D(n7683), .CK(CLK), .QN(n21578) );
  DFF_X1 \REGISTERS_reg[5][0]  ( .D(n7682), .CK(CLK), .QN(n21579) );
  DFF_X1 \REGISTERS_reg[0][63]  ( .D(n8065), .CK(CLK), .Q(n25582), .QN(n21516)
         );
  DFF_X1 \REGISTERS_reg[0][62]  ( .D(n8064), .CK(CLK), .Q(n25581), .QN(n21517)
         );
  DFF_X1 \REGISTERS_reg[0][61]  ( .D(n8063), .CK(CLK), .Q(n25580), .QN(n21518)
         );
  DFF_X1 \REGISTERS_reg[0][60]  ( .D(n8062), .CK(CLK), .Q(n25579), .QN(n21519)
         );
  DFF_X1 \REGISTERS_reg[0][59]  ( .D(n8061), .CK(CLK), .Q(n25550), .QN(n22120)
         );
  DFF_X1 \REGISTERS_reg[0][58]  ( .D(n8060), .CK(CLK), .Q(n25549), .QN(n22121)
         );
  DFF_X1 \REGISTERS_reg[0][57]  ( .D(n8059), .CK(CLK), .Q(n25548), .QN(n22122)
         );
  DFF_X1 \REGISTERS_reg[0][56]  ( .D(n8058), .CK(CLK), .Q(n25547), .QN(n22123)
         );
  DFF_X1 \REGISTERS_reg[0][55]  ( .D(n8057), .CK(CLK), .Q(n25546), .QN(n22124)
         );
  DFF_X1 \REGISTERS_reg[0][54]  ( .D(n8056), .CK(CLK), .Q(n25545), .QN(n22125)
         );
  DFF_X1 \REGISTERS_reg[0][53]  ( .D(n8055), .CK(CLK), .Q(n25544), .QN(n22126)
         );
  DFF_X1 \REGISTERS_reg[0][52]  ( .D(n8054), .CK(CLK), .Q(n25543), .QN(n22127)
         );
  DFF_X1 \REGISTERS_reg[0][51]  ( .D(n8053), .CK(CLK), .Q(n25542), .QN(n22128)
         );
  DFF_X1 \REGISTERS_reg[0][50]  ( .D(n8052), .CK(CLK), .Q(n25541), .QN(n22129)
         );
  DFF_X1 \REGISTERS_reg[0][49]  ( .D(n8051), .CK(CLK), .Q(n25540), .QN(n22130)
         );
  DFF_X1 \REGISTERS_reg[0][48]  ( .D(n8050), .CK(CLK), .Q(n25539), .QN(n22131)
         );
  DFF_X1 \REGISTERS_reg[0][47]  ( .D(n8049), .CK(CLK), .Q(n25538), .QN(n22132)
         );
  DFF_X1 \REGISTERS_reg[0][46]  ( .D(n8048), .CK(CLK), .Q(n25537), .QN(n22133)
         );
  DFF_X1 \REGISTERS_reg[0][45]  ( .D(n8047), .CK(CLK), .Q(n25536), .QN(n22134)
         );
  DFF_X1 \REGISTERS_reg[0][44]  ( .D(n8046), .CK(CLK), .Q(n25535), .QN(n22135)
         );
  DFF_X1 \REGISTERS_reg[0][43]  ( .D(n8045), .CK(CLK), .Q(n25534), .QN(n22136)
         );
  DFF_X1 \REGISTERS_reg[0][42]  ( .D(n8044), .CK(CLK), .Q(n25533), .QN(n22137)
         );
  DFF_X1 \REGISTERS_reg[0][41]  ( .D(n8043), .CK(CLK), .Q(n25532), .QN(n22138)
         );
  DFF_X1 \REGISTERS_reg[0][40]  ( .D(n8042), .CK(CLK), .Q(n25531), .QN(n22139)
         );
  DFF_X1 \REGISTERS_reg[0][39]  ( .D(n8041), .CK(CLK), .Q(n25530), .QN(n22140)
         );
  DFF_X1 \REGISTERS_reg[0][38]  ( .D(n8040), .CK(CLK), .Q(n25529), .QN(n22141)
         );
  DFF_X1 \REGISTERS_reg[0][37]  ( .D(n8039), .CK(CLK), .Q(n25528), .QN(n22142)
         );
  DFF_X1 \REGISTERS_reg[0][36]  ( .D(n8038), .CK(CLK), .Q(n25527), .QN(n22143)
         );
  DFF_X1 \REGISTERS_reg[0][35]  ( .D(n8037), .CK(CLK), .Q(n25526), .QN(n22144)
         );
  DFF_X1 \REGISTERS_reg[0][34]  ( .D(n8036), .CK(CLK), .Q(n25525), .QN(n22145)
         );
  DFF_X1 \REGISTERS_reg[0][33]  ( .D(n8035), .CK(CLK), .Q(n25524), .QN(n22146)
         );
  DFF_X1 \REGISTERS_reg[0][32]  ( .D(n8034), .CK(CLK), .Q(n25523), .QN(n22147)
         );
  DFF_X1 \REGISTERS_reg[0][31]  ( .D(n8033), .CK(CLK), .Q(n25522), .QN(n22148)
         );
  DFF_X1 \REGISTERS_reg[0][30]  ( .D(n8032), .CK(CLK), .Q(n25521), .QN(n22149)
         );
  DFF_X1 \REGISTERS_reg[0][29]  ( .D(n8031), .CK(CLK), .Q(n25520), .QN(n22150)
         );
  DFF_X1 \REGISTERS_reg[0][28]  ( .D(n8030), .CK(CLK), .Q(n25519), .QN(n22151)
         );
  DFF_X1 \REGISTERS_reg[0][27]  ( .D(n8029), .CK(CLK), .Q(n25518), .QN(n22152)
         );
  DFF_X1 \REGISTERS_reg[0][26]  ( .D(n8028), .CK(CLK), .Q(n25517), .QN(n22153)
         );
  DFF_X1 \REGISTERS_reg[0][25]  ( .D(n8027), .CK(CLK), .Q(n25516), .QN(n22154)
         );
  DFF_X1 \REGISTERS_reg[0][24]  ( .D(n8026), .CK(CLK), .Q(n25515), .QN(n22155)
         );
  DFF_X1 \REGISTERS_reg[0][23]  ( .D(n8025), .CK(CLK), .Q(n25514), .QN(n22156)
         );
  DFF_X1 \REGISTERS_reg[0][22]  ( .D(n8024), .CK(CLK), .Q(n25513), .QN(n22157)
         );
  DFF_X1 \REGISTERS_reg[0][21]  ( .D(n8023), .CK(CLK), .Q(n25512), .QN(n22158)
         );
  DFF_X1 \REGISTERS_reg[0][20]  ( .D(n8022), .CK(CLK), .Q(n25511), .QN(n22159)
         );
  DFF_X1 \REGISTERS_reg[0][19]  ( .D(n8021), .CK(CLK), .Q(n25510), .QN(n22160)
         );
  DFF_X1 \REGISTERS_reg[0][18]  ( .D(n8020), .CK(CLK), .Q(n25509), .QN(n22161)
         );
  DFF_X1 \REGISTERS_reg[0][17]  ( .D(n8019), .CK(CLK), .Q(n25508), .QN(n22162)
         );
  DFF_X1 \REGISTERS_reg[0][16]  ( .D(n8018), .CK(CLK), .Q(n25507), .QN(n22163)
         );
  DFF_X1 \REGISTERS_reg[0][15]  ( .D(n8017), .CK(CLK), .Q(n25506), .QN(n22164)
         );
  DFF_X1 \REGISTERS_reg[0][14]  ( .D(n8016), .CK(CLK), .Q(n25505), .QN(n22165)
         );
  DFF_X1 \REGISTERS_reg[0][13]  ( .D(n8015), .CK(CLK), .Q(n25504), .QN(n22166)
         );
  DFF_X1 \REGISTERS_reg[0][12]  ( .D(n8014), .CK(CLK), .Q(n25503), .QN(n22167)
         );
  DFF_X1 \REGISTERS_reg[0][11]  ( .D(n8013), .CK(CLK), .Q(n25678), .QN(n22168)
         );
  DFF_X1 \REGISTERS_reg[0][10]  ( .D(n8012), .CK(CLK), .Q(n25677), .QN(n22169)
         );
  DFF_X1 \REGISTERS_reg[0][9]  ( .D(n8011), .CK(CLK), .Q(n25676), .QN(n22170)
         );
  DFF_X1 \REGISTERS_reg[0][8]  ( .D(n8010), .CK(CLK), .Q(n25675), .QN(n22171)
         );
  DFF_X1 \REGISTERS_reg[0][7]  ( .D(n8009), .CK(CLK), .Q(n25674), .QN(n22172)
         );
  DFF_X1 \REGISTERS_reg[0][6]  ( .D(n8008), .CK(CLK), .Q(n25673), .QN(n22173)
         );
  DFF_X1 \REGISTERS_reg[0][5]  ( .D(n8007), .CK(CLK), .Q(n25672), .QN(n22174)
         );
  DFF_X1 \REGISTERS_reg[0][4]  ( .D(n8006), .CK(CLK), .Q(n25671), .QN(n22175)
         );
  DFF_X1 \REGISTERS_reg[0][3]  ( .D(n8005), .CK(CLK), .Q(n25670), .QN(n22176)
         );
  DFF_X1 \REGISTERS_reg[0][2]  ( .D(n8004), .CK(CLK), .Q(n25669), .QN(n22177)
         );
  DFF_X1 \REGISTERS_reg[0][1]  ( .D(n8003), .CK(CLK), .Q(n25668), .QN(n22178)
         );
  DFF_X1 \REGISTERS_reg[0][0]  ( .D(n8002), .CK(CLK), .Q(n25667), .QN(n22179)
         );
  DFF_X1 \REGISTERS_reg[4][63]  ( .D(n7809), .CK(CLK), .Q(n25574), .QN(n21500)
         );
  DFF_X1 \REGISTERS_reg[4][62]  ( .D(n7808), .CK(CLK), .Q(n25573), .QN(n21501)
         );
  DFF_X1 \REGISTERS_reg[4][61]  ( .D(n7807), .CK(CLK), .Q(n25572), .QN(n21502)
         );
  DFF_X1 \REGISTERS_reg[4][60]  ( .D(n7806), .CK(CLK), .Q(n25571), .QN(n21503)
         );
  DFF_X1 \REGISTERS_reg[30][63]  ( .D(n6145), .CK(CLK), .Q(n26198), .QN(n20835) );
  DFF_X1 \REGISTERS_reg[30][62]  ( .D(n6144), .CK(CLK), .Q(n26197), .QN(n20836) );
  DFF_X1 \REGISTERS_reg[30][61]  ( .D(n6143), .CK(CLK), .Q(n26196), .QN(n20837) );
  DFF_X1 \REGISTERS_reg[30][60]  ( .D(n6142), .CK(CLK), .Q(n26195), .QN(n20838) );
  DFF_X1 \REGISTERS_reg[28][63]  ( .D(n6273), .CK(CLK), .Q(n8450), .QN(n22180)
         );
  DFF_X1 \REGISTERS_reg[28][62]  ( .D(n6272), .CK(CLK), .Q(n8453), .QN(n22181)
         );
  DFF_X1 \REGISTERS_reg[28][61]  ( .D(n6271), .CK(CLK), .Q(n8456), .QN(n22182)
         );
  DFF_X1 \REGISTERS_reg[28][60]  ( .D(n6270), .CK(CLK), .Q(n8459), .QN(n22183)
         );
  DFF_X1 \REGISTERS_reg[27][63]  ( .D(n6337), .CK(CLK), .Q(n18367), .QN(n22504) );
  DFF_X1 \REGISTERS_reg[27][62]  ( .D(n6336), .CK(CLK), .Q(n18384), .QN(n22505) );
  DFF_X1 \REGISTERS_reg[27][61]  ( .D(n6335), .CK(CLK), .Q(n18401), .QN(n22506) );
  DFF_X1 \REGISTERS_reg[27][60]  ( .D(n6334), .CK(CLK), .Q(n18418), .QN(n22507) );
  DFF_X1 \REGISTERS_reg[2][63]  ( .D(n7937), .CK(CLK), .Q(n25566), .QN(n21172)
         );
  DFF_X1 \REGISTERS_reg[2][62]  ( .D(n7936), .CK(CLK), .Q(n25565), .QN(n21173)
         );
  DFF_X1 \REGISTERS_reg[2][61]  ( .D(n7935), .CK(CLK), .Q(n25564), .QN(n21174)
         );
  DFF_X1 \REGISTERS_reg[2][60]  ( .D(n7934), .CK(CLK), .Q(n25563), .QN(n21175)
         );
  DFF_X1 \REGISTERS_reg[4][59]  ( .D(n7805), .CK(CLK), .Q(n25454), .QN(n21880)
         );
  DFF_X1 \REGISTERS_reg[4][58]  ( .D(n7804), .CK(CLK), .Q(n25453), .QN(n21881)
         );
  DFF_X1 \REGISTERS_reg[4][57]  ( .D(n7803), .CK(CLK), .Q(n25452), .QN(n21882)
         );
  DFF_X1 \REGISTERS_reg[4][56]  ( .D(n7802), .CK(CLK), .Q(n25451), .QN(n21883)
         );
  DFF_X1 \REGISTERS_reg[4][55]  ( .D(n7801), .CK(CLK), .Q(n25450), .QN(n21884)
         );
  DFF_X1 \REGISTERS_reg[4][54]  ( .D(n7800), .CK(CLK), .Q(n25449), .QN(n21885)
         );
  DFF_X1 \REGISTERS_reg[4][53]  ( .D(n7799), .CK(CLK), .Q(n25448), .QN(n21886)
         );
  DFF_X1 \REGISTERS_reg[4][52]  ( .D(n7798), .CK(CLK), .Q(n25447), .QN(n21887)
         );
  DFF_X1 \REGISTERS_reg[4][51]  ( .D(n7797), .CK(CLK), .Q(n25446), .QN(n21888)
         );
  DFF_X1 \REGISTERS_reg[4][50]  ( .D(n7796), .CK(CLK), .Q(n25445), .QN(n21889)
         );
  DFF_X1 \REGISTERS_reg[4][49]  ( .D(n7795), .CK(CLK), .Q(n25444), .QN(n21890)
         );
  DFF_X1 \REGISTERS_reg[4][48]  ( .D(n7794), .CK(CLK), .Q(n25443), .QN(n21891)
         );
  DFF_X1 \REGISTERS_reg[4][47]  ( .D(n7793), .CK(CLK), .Q(n25442), .QN(n21892)
         );
  DFF_X1 \REGISTERS_reg[4][46]  ( .D(n7792), .CK(CLK), .Q(n25441), .QN(n21893)
         );
  DFF_X1 \REGISTERS_reg[4][45]  ( .D(n7791), .CK(CLK), .Q(n25440), .QN(n21894)
         );
  DFF_X1 \REGISTERS_reg[4][44]  ( .D(n7790), .CK(CLK), .Q(n25439), .QN(n21895)
         );
  DFF_X1 \REGISTERS_reg[4][43]  ( .D(n7789), .CK(CLK), .Q(n25438), .QN(n21896)
         );
  DFF_X1 \REGISTERS_reg[4][42]  ( .D(n7788), .CK(CLK), .Q(n25437), .QN(n21897)
         );
  DFF_X1 \REGISTERS_reg[4][41]  ( .D(n7787), .CK(CLK), .Q(n25436), .QN(n21898)
         );
  DFF_X1 \REGISTERS_reg[4][40]  ( .D(n7786), .CK(CLK), .Q(n25435), .QN(n21899)
         );
  DFF_X1 \REGISTERS_reg[4][39]  ( .D(n7785), .CK(CLK), .Q(n25434), .QN(n21900)
         );
  DFF_X1 \REGISTERS_reg[4][38]  ( .D(n7784), .CK(CLK), .Q(n25433), .QN(n21901)
         );
  DFF_X1 \REGISTERS_reg[4][37]  ( .D(n7783), .CK(CLK), .Q(n25432), .QN(n21902)
         );
  DFF_X1 \REGISTERS_reg[4][36]  ( .D(n7782), .CK(CLK), .Q(n25431), .QN(n21903)
         );
  DFF_X1 \REGISTERS_reg[4][35]  ( .D(n7781), .CK(CLK), .Q(n25430), .QN(n21904)
         );
  DFF_X1 \REGISTERS_reg[4][34]  ( .D(n7780), .CK(CLK), .Q(n25429), .QN(n21905)
         );
  DFF_X1 \REGISTERS_reg[4][33]  ( .D(n7779), .CK(CLK), .Q(n25428), .QN(n21906)
         );
  DFF_X1 \REGISTERS_reg[4][32]  ( .D(n7778), .CK(CLK), .Q(n25427), .QN(n21907)
         );
  DFF_X1 \REGISTERS_reg[4][31]  ( .D(n7777), .CK(CLK), .Q(n25426), .QN(n21908)
         );
  DFF_X1 \REGISTERS_reg[4][30]  ( .D(n7776), .CK(CLK), .Q(n25425), .QN(n21909)
         );
  DFF_X1 \REGISTERS_reg[4][29]  ( .D(n7775), .CK(CLK), .Q(n25424), .QN(n21910)
         );
  DFF_X1 \REGISTERS_reg[4][28]  ( .D(n7774), .CK(CLK), .Q(n25423), .QN(n21911)
         );
  DFF_X1 \REGISTERS_reg[4][27]  ( .D(n7773), .CK(CLK), .Q(n25422), .QN(n21912)
         );
  DFF_X1 \REGISTERS_reg[4][26]  ( .D(n7772), .CK(CLK), .Q(n25421), .QN(n21913)
         );
  DFF_X1 \REGISTERS_reg[4][25]  ( .D(n7771), .CK(CLK), .Q(n25420), .QN(n21914)
         );
  DFF_X1 \REGISTERS_reg[4][24]  ( .D(n7770), .CK(CLK), .Q(n25419), .QN(n21915)
         );
  DFF_X1 \REGISTERS_reg[4][23]  ( .D(n7769), .CK(CLK), .Q(n25418), .QN(n21916)
         );
  DFF_X1 \REGISTERS_reg[4][22]  ( .D(n7768), .CK(CLK), .Q(n25417), .QN(n21917)
         );
  DFF_X1 \REGISTERS_reg[4][21]  ( .D(n7767), .CK(CLK), .Q(n25416), .QN(n21918)
         );
  DFF_X1 \REGISTERS_reg[4][20]  ( .D(n7766), .CK(CLK), .Q(n25415), .QN(n21919)
         );
  DFF_X1 \REGISTERS_reg[4][19]  ( .D(n7765), .CK(CLK), .Q(n25414), .QN(n21920)
         );
  DFF_X1 \REGISTERS_reg[4][18]  ( .D(n7764), .CK(CLK), .Q(n25413), .QN(n21921)
         );
  DFF_X1 \REGISTERS_reg[4][17]  ( .D(n7763), .CK(CLK), .Q(n25412), .QN(n21922)
         );
  DFF_X1 \REGISTERS_reg[4][16]  ( .D(n7762), .CK(CLK), .Q(n25411), .QN(n21923)
         );
  DFF_X1 \REGISTERS_reg[4][15]  ( .D(n7761), .CK(CLK), .Q(n25410), .QN(n21924)
         );
  DFF_X1 \REGISTERS_reg[4][14]  ( .D(n7760), .CK(CLK), .Q(n25409), .QN(n21925)
         );
  DFF_X1 \REGISTERS_reg[4][13]  ( .D(n7759), .CK(CLK), .Q(n25408), .QN(n21926)
         );
  DFF_X1 \REGISTERS_reg[4][12]  ( .D(n7758), .CK(CLK), .Q(n25407), .QN(n21927)
         );
  DFF_X1 \REGISTERS_reg[4][11]  ( .D(n7757), .CK(CLK), .Q(n25630), .QN(n21928)
         );
  DFF_X1 \REGISTERS_reg[4][10]  ( .D(n7756), .CK(CLK), .Q(n25629), .QN(n21929)
         );
  DFF_X1 \REGISTERS_reg[4][9]  ( .D(n7755), .CK(CLK), .Q(n25628), .QN(n21930)
         );
  DFF_X1 \REGISTERS_reg[4][8]  ( .D(n7754), .CK(CLK), .Q(n25627), .QN(n21931)
         );
  DFF_X1 \REGISTERS_reg[4][7]  ( .D(n7753), .CK(CLK), .Q(n25626), .QN(n21932)
         );
  DFF_X1 \REGISTERS_reg[4][6]  ( .D(n7752), .CK(CLK), .Q(n25625), .QN(n21933)
         );
  DFF_X1 \REGISTERS_reg[4][5]  ( .D(n7751), .CK(CLK), .Q(n25624), .QN(n21934)
         );
  DFF_X1 \REGISTERS_reg[4][4]  ( .D(n7750), .CK(CLK), .Q(n25623), .QN(n21935)
         );
  DFF_X1 \REGISTERS_reg[4][3]  ( .D(n7749), .CK(CLK), .Q(n25622), .QN(n21936)
         );
  DFF_X1 \REGISTERS_reg[4][2]  ( .D(n7748), .CK(CLK), .Q(n25621), .QN(n21937)
         );
  DFF_X1 \REGISTERS_reg[4][1]  ( .D(n7747), .CK(CLK), .Q(n25620), .QN(n21938)
         );
  DFF_X1 \REGISTERS_reg[4][0]  ( .D(n7746), .CK(CLK), .Q(n25619), .QN(n21939)
         );
  DFF_X1 \REGISTERS_reg[30][59]  ( .D(n6141), .CK(CLK), .Q(n26386), .QN(n20839) );
  DFF_X1 \REGISTERS_reg[30][58]  ( .D(n6140), .CK(CLK), .Q(n26385), .QN(n20840) );
  DFF_X1 \REGISTERS_reg[30][57]  ( .D(n6139), .CK(CLK), .Q(n26384), .QN(n20841) );
  DFF_X1 \REGISTERS_reg[30][56]  ( .D(n6138), .CK(CLK), .Q(n26383), .QN(n20842) );
  DFF_X1 \REGISTERS_reg[30][55]  ( .D(n6137), .CK(CLK), .Q(n26382), .QN(n20843) );
  DFF_X1 \REGISTERS_reg[30][54]  ( .D(n6136), .CK(CLK), .Q(n26381), .QN(n20844) );
  DFF_X1 \REGISTERS_reg[30][53]  ( .D(n6135), .CK(CLK), .Q(n26380), .QN(n20845) );
  DFF_X1 \REGISTERS_reg[30][52]  ( .D(n6134), .CK(CLK), .Q(n26379), .QN(n20846) );
  DFF_X1 \REGISTERS_reg[30][51]  ( .D(n6133), .CK(CLK), .Q(n26378), .QN(n20847) );
  DFF_X1 \REGISTERS_reg[30][50]  ( .D(n6132), .CK(CLK), .Q(n26377), .QN(n20848) );
  DFF_X1 \REGISTERS_reg[30][49]  ( .D(n6131), .CK(CLK), .Q(n26376), .QN(n20849) );
  DFF_X1 \REGISTERS_reg[30][48]  ( .D(n6130), .CK(CLK), .Q(n26375), .QN(n20850) );
  DFF_X1 \REGISTERS_reg[30][47]  ( .D(n6129), .CK(CLK), .Q(n26374), .QN(n20851) );
  DFF_X1 \REGISTERS_reg[30][46]  ( .D(n6128), .CK(CLK), .Q(n26373), .QN(n20852) );
  DFF_X1 \REGISTERS_reg[30][45]  ( .D(n6127), .CK(CLK), .Q(n26372), .QN(n20853) );
  DFF_X1 \REGISTERS_reg[30][44]  ( .D(n6126), .CK(CLK), .Q(n26371), .QN(n20854) );
  DFF_X1 \REGISTERS_reg[30][43]  ( .D(n6125), .CK(CLK), .Q(n26370), .QN(n20855) );
  DFF_X1 \REGISTERS_reg[30][42]  ( .D(n6124), .CK(CLK), .Q(n26369), .QN(n20856) );
  DFF_X1 \REGISTERS_reg[30][41]  ( .D(n6123), .CK(CLK), .Q(n26368), .QN(n20857) );
  DFF_X1 \REGISTERS_reg[30][40]  ( .D(n6122), .CK(CLK), .Q(n26367), .QN(n20858) );
  DFF_X1 \REGISTERS_reg[30][39]  ( .D(n6121), .CK(CLK), .Q(n26366), .QN(n20859) );
  DFF_X1 \REGISTERS_reg[30][38]  ( .D(n6120), .CK(CLK), .Q(n26365), .QN(n20860) );
  DFF_X1 \REGISTERS_reg[30][37]  ( .D(n6119), .CK(CLK), .Q(n26364), .QN(n20861) );
  DFF_X1 \REGISTERS_reg[30][36]  ( .D(n6118), .CK(CLK), .Q(n26363), .QN(n20862) );
  DFF_X1 \REGISTERS_reg[30][35]  ( .D(n6117), .CK(CLK), .Q(n26362), .QN(n20863) );
  DFF_X1 \REGISTERS_reg[30][34]  ( .D(n6116), .CK(CLK), .Q(n26361), .QN(n20864) );
  DFF_X1 \REGISTERS_reg[30][33]  ( .D(n6115), .CK(CLK), .Q(n26360), .QN(n20865) );
  DFF_X1 \REGISTERS_reg[30][32]  ( .D(n6114), .CK(CLK), .Q(n26359), .QN(n20866) );
  DFF_X1 \REGISTERS_reg[30][31]  ( .D(n6113), .CK(CLK), .Q(n26358), .QN(n20867) );
  DFF_X1 \REGISTERS_reg[30][30]  ( .D(n6112), .CK(CLK), .Q(n26357), .QN(n20868) );
  DFF_X1 \REGISTERS_reg[30][29]  ( .D(n6111), .CK(CLK), .Q(n26356), .QN(n20869) );
  DFF_X1 \REGISTERS_reg[30][28]  ( .D(n6110), .CK(CLK), .Q(n26355), .QN(n20870) );
  DFF_X1 \REGISTERS_reg[30][27]  ( .D(n6109), .CK(CLK), .Q(n26354), .QN(n20871) );
  DFF_X1 \REGISTERS_reg[30][26]  ( .D(n6108), .CK(CLK), .Q(n26353), .QN(n20872) );
  DFF_X1 \REGISTERS_reg[30][25]  ( .D(n6107), .CK(CLK), .Q(n26352), .QN(n20873) );
  DFF_X1 \REGISTERS_reg[30][24]  ( .D(n6106), .CK(CLK), .Q(n26351), .QN(n20874) );
  DFF_X1 \REGISTERS_reg[30][23]  ( .D(n6105), .CK(CLK), .Q(n26350), .QN(n20875) );
  DFF_X1 \REGISTERS_reg[30][22]  ( .D(n6104), .CK(CLK), .Q(n26349), .QN(n20876) );
  DFF_X1 \REGISTERS_reg[30][21]  ( .D(n6103), .CK(CLK), .Q(n26348), .QN(n20877) );
  DFF_X1 \REGISTERS_reg[30][20]  ( .D(n6102), .CK(CLK), .Q(n26347), .QN(n20878) );
  DFF_X1 \REGISTERS_reg[30][19]  ( .D(n6101), .CK(CLK), .Q(n26346), .QN(n20879) );
  DFF_X1 \REGISTERS_reg[30][18]  ( .D(n6100), .CK(CLK), .Q(n26345), .QN(n20880) );
  DFF_X1 \REGISTERS_reg[30][17]  ( .D(n6099), .CK(CLK), .Q(n26344), .QN(n20881) );
  DFF_X1 \REGISTERS_reg[30][16]  ( .D(n6098), .CK(CLK), .Q(n26343), .QN(n20882) );
  DFF_X1 \REGISTERS_reg[30][15]  ( .D(n6097), .CK(CLK), .Q(n26342), .QN(n20883) );
  DFF_X1 \REGISTERS_reg[30][14]  ( .D(n6096), .CK(CLK), .Q(n26341), .QN(n20884) );
  DFF_X1 \REGISTERS_reg[30][13]  ( .D(n6095), .CK(CLK), .Q(n26340), .QN(n20885) );
  DFF_X1 \REGISTERS_reg[30][12]  ( .D(n6094), .CK(CLK), .Q(n26339), .QN(n20886) );
  DFF_X1 \REGISTERS_reg[30][11]  ( .D(n6093), .CK(CLK), .Q(n26338), .QN(n20887) );
  DFF_X1 \REGISTERS_reg[30][10]  ( .D(n6092), .CK(CLK), .Q(n26337), .QN(n20888) );
  DFF_X1 \REGISTERS_reg[30][9]  ( .D(n6091), .CK(CLK), .Q(n26336), .QN(n20889)
         );
  DFF_X1 \REGISTERS_reg[30][8]  ( .D(n6090), .CK(CLK), .Q(n26335), .QN(n20890)
         );
  DFF_X1 \REGISTERS_reg[30][7]  ( .D(n6089), .CK(CLK), .Q(n26334), .QN(n20891)
         );
  DFF_X1 \REGISTERS_reg[30][6]  ( .D(n6088), .CK(CLK), .Q(n26333), .QN(n20892)
         );
  DFF_X1 \REGISTERS_reg[30][5]  ( .D(n6087), .CK(CLK), .Q(n26332), .QN(n20893)
         );
  DFF_X1 \REGISTERS_reg[30][4]  ( .D(n6086), .CK(CLK), .Q(n26331), .QN(n20894)
         );
  DFF_X1 \REGISTERS_reg[30][3]  ( .D(n6085), .CK(CLK), .Q(n26330), .QN(n20895)
         );
  DFF_X1 \REGISTERS_reg[30][2]  ( .D(n6084), .CK(CLK), .Q(n26329), .QN(n20896)
         );
  DFF_X1 \REGISTERS_reg[30][1]  ( .D(n6083), .CK(CLK), .Q(n26328), .QN(n20897)
         );
  DFF_X1 \REGISTERS_reg[30][0]  ( .D(n6082), .CK(CLK), .Q(n26327), .QN(n20898)
         );
  DFF_X1 \REGISTERS_reg[28][59]  ( .D(n6269), .CK(CLK), .Q(n8462), .QN(n22184)
         );
  DFF_X1 \REGISTERS_reg[28][58]  ( .D(n6268), .CK(CLK), .Q(n8465), .QN(n22185)
         );
  DFF_X1 \REGISTERS_reg[28][57]  ( .D(n6267), .CK(CLK), .Q(n8468), .QN(n22186)
         );
  DFF_X1 \REGISTERS_reg[28][56]  ( .D(n6266), .CK(CLK), .Q(n8471), .QN(n22187)
         );
  DFF_X1 \REGISTERS_reg[28][55]  ( .D(n6265), .CK(CLK), .Q(n8474), .QN(n22188)
         );
  DFF_X1 \REGISTERS_reg[28][54]  ( .D(n6264), .CK(CLK), .Q(n8477), .QN(n22189)
         );
  DFF_X1 \REGISTERS_reg[28][53]  ( .D(n6263), .CK(CLK), .Q(n8480), .QN(n22190)
         );
  DFF_X1 \REGISTERS_reg[28][52]  ( .D(n6262), .CK(CLK), .Q(n8483), .QN(n22191)
         );
  DFF_X1 \REGISTERS_reg[28][51]  ( .D(n6261), .CK(CLK), .Q(n8486), .QN(n22192)
         );
  DFF_X1 \REGISTERS_reg[28][50]  ( .D(n6260), .CK(CLK), .Q(n8489), .QN(n22193)
         );
  DFF_X1 \REGISTERS_reg[28][49]  ( .D(n6259), .CK(CLK), .Q(n8492), .QN(n22194)
         );
  DFF_X1 \REGISTERS_reg[28][48]  ( .D(n6258), .CK(CLK), .Q(n8495), .QN(n22195)
         );
  DFF_X1 \REGISTERS_reg[28][47]  ( .D(n6257), .CK(CLK), .Q(n8498), .QN(n22196)
         );
  DFF_X1 \REGISTERS_reg[28][46]  ( .D(n6256), .CK(CLK), .Q(n8501), .QN(n22197)
         );
  DFF_X1 \REGISTERS_reg[28][45]  ( .D(n6255), .CK(CLK), .Q(n8504), .QN(n22198)
         );
  DFF_X1 \REGISTERS_reg[28][44]  ( .D(n6254), .CK(CLK), .Q(n8507), .QN(n22199)
         );
  DFF_X1 \REGISTERS_reg[28][43]  ( .D(n6253), .CK(CLK), .Q(n8510), .QN(n22200)
         );
  DFF_X1 \REGISTERS_reg[28][42]  ( .D(n6252), .CK(CLK), .Q(n8513), .QN(n22201)
         );
  DFF_X1 \REGISTERS_reg[28][41]  ( .D(n6251), .CK(CLK), .Q(n8516), .QN(n22202)
         );
  DFF_X1 \REGISTERS_reg[28][40]  ( .D(n6250), .CK(CLK), .Q(n8519), .QN(n22203)
         );
  DFF_X1 \REGISTERS_reg[28][39]  ( .D(n6249), .CK(CLK), .Q(n8522), .QN(n22204)
         );
  DFF_X1 \REGISTERS_reg[28][38]  ( .D(n6248), .CK(CLK), .Q(n8525), .QN(n22205)
         );
  DFF_X1 \REGISTERS_reg[28][37]  ( .D(n6247), .CK(CLK), .Q(n8528), .QN(n22206)
         );
  DFF_X1 \REGISTERS_reg[28][36]  ( .D(n6246), .CK(CLK), .Q(n8531), .QN(n22207)
         );
  DFF_X1 \REGISTERS_reg[28][35]  ( .D(n6245), .CK(CLK), .Q(n8534), .QN(n22208)
         );
  DFF_X1 \REGISTERS_reg[28][34]  ( .D(n6244), .CK(CLK), .Q(n8537), .QN(n22209)
         );
  DFF_X1 \REGISTERS_reg[28][33]  ( .D(n6243), .CK(CLK), .Q(n8540), .QN(n22210)
         );
  DFF_X1 \REGISTERS_reg[28][32]  ( .D(n6242), .CK(CLK), .Q(n8543), .QN(n22211)
         );
  DFF_X1 \REGISTERS_reg[28][31]  ( .D(n6241), .CK(CLK), .Q(n8546), .QN(n22212)
         );
  DFF_X1 \REGISTERS_reg[28][30]  ( .D(n6240), .CK(CLK), .Q(n8549), .QN(n22213)
         );
  DFF_X1 \REGISTERS_reg[28][29]  ( .D(n6239), .CK(CLK), .Q(n8552), .QN(n22214)
         );
  DFF_X1 \REGISTERS_reg[28][28]  ( .D(n6238), .CK(CLK), .Q(n8555), .QN(n22215)
         );
  DFF_X1 \REGISTERS_reg[28][27]  ( .D(n6237), .CK(CLK), .Q(n8558), .QN(n22216)
         );
  DFF_X1 \REGISTERS_reg[28][26]  ( .D(n6236), .CK(CLK), .Q(n8561), .QN(n22217)
         );
  DFF_X1 \REGISTERS_reg[28][25]  ( .D(n6235), .CK(CLK), .Q(n8564), .QN(n22218)
         );
  DFF_X1 \REGISTERS_reg[28][24]  ( .D(n6234), .CK(CLK), .Q(n8567), .QN(n22219)
         );
  DFF_X1 \REGISTERS_reg[28][23]  ( .D(n6233), .CK(CLK), .Q(n8570), .QN(n22220)
         );
  DFF_X1 \REGISTERS_reg[28][22]  ( .D(n6232), .CK(CLK), .Q(n8573), .QN(n22221)
         );
  DFF_X1 \REGISTERS_reg[28][21]  ( .D(n6231), .CK(CLK), .Q(n8576), .QN(n22222)
         );
  DFF_X1 \REGISTERS_reg[28][20]  ( .D(n6230), .CK(CLK), .Q(n8579), .QN(n22223)
         );
  DFF_X1 \REGISTERS_reg[28][19]  ( .D(n6229), .CK(CLK), .Q(n8582), .QN(n22224)
         );
  DFF_X1 \REGISTERS_reg[28][18]  ( .D(n6228), .CK(CLK), .Q(n8585), .QN(n22225)
         );
  DFF_X1 \REGISTERS_reg[28][17]  ( .D(n6227), .CK(CLK), .Q(n8588), .QN(n22226)
         );
  DFF_X1 \REGISTERS_reg[28][16]  ( .D(n6226), .CK(CLK), .Q(n8591), .QN(n22227)
         );
  DFF_X1 \REGISTERS_reg[28][15]  ( .D(n6225), .CK(CLK), .Q(n8594), .QN(n22228)
         );
  DFF_X1 \REGISTERS_reg[28][14]  ( .D(n6224), .CK(CLK), .Q(n8597), .QN(n22229)
         );
  DFF_X1 \REGISTERS_reg[28][13]  ( .D(n6223), .CK(CLK), .Q(n8600), .QN(n22230)
         );
  DFF_X1 \REGISTERS_reg[28][12]  ( .D(n6222), .CK(CLK), .Q(n8603), .QN(n22231)
         );
  DFF_X1 \REGISTERS_reg[28][11]  ( .D(n6221), .CK(CLK), .Q(n8606), .QN(n22232)
         );
  DFF_X1 \REGISTERS_reg[28][10]  ( .D(n6220), .CK(CLK), .Q(n8609), .QN(n22233)
         );
  DFF_X1 \REGISTERS_reg[28][9]  ( .D(n6219), .CK(CLK), .Q(n8612), .QN(n22234)
         );
  DFF_X1 \REGISTERS_reg[28][8]  ( .D(n6218), .CK(CLK), .Q(n8615), .QN(n22235)
         );
  DFF_X1 \REGISTERS_reg[28][7]  ( .D(n6217), .CK(CLK), .Q(n8618), .QN(n22236)
         );
  DFF_X1 \REGISTERS_reg[28][6]  ( .D(n6216), .CK(CLK), .Q(n8621), .QN(n22237)
         );
  DFF_X1 \REGISTERS_reg[28][5]  ( .D(n6215), .CK(CLK), .Q(n8624), .QN(n22238)
         );
  DFF_X1 \REGISTERS_reg[28][4]  ( .D(n6214), .CK(CLK), .Q(n8627), .QN(n22239)
         );
  DFF_X1 \REGISTERS_reg[28][3]  ( .D(n6213), .CK(CLK), .Q(n8630), .QN(n22240)
         );
  DFF_X1 \REGISTERS_reg[28][2]  ( .D(n6212), .CK(CLK), .Q(n8633), .QN(n22241)
         );
  DFF_X1 \REGISTERS_reg[28][1]  ( .D(n6211), .CK(CLK), .Q(n8636), .QN(n22242)
         );
  DFF_X1 \REGISTERS_reg[28][0]  ( .D(n6210), .CK(CLK), .Q(n8639), .QN(n22243)
         );
  DFF_X1 \REGISTERS_reg[27][59]  ( .D(n6333), .CK(CLK), .Q(n18435), .QN(n22572) );
  DFF_X1 \REGISTERS_reg[27][58]  ( .D(n6332), .CK(CLK), .Q(n18452), .QN(n22573) );
  DFF_X1 \REGISTERS_reg[27][57]  ( .D(n6331), .CK(CLK), .Q(n18469), .QN(n22574) );
  DFF_X1 \REGISTERS_reg[27][56]  ( .D(n6330), .CK(CLK), .Q(n18486), .QN(n22575) );
  DFF_X1 \REGISTERS_reg[27][55]  ( .D(n6329), .CK(CLK), .Q(n18503), .QN(n22576) );
  DFF_X1 \REGISTERS_reg[27][54]  ( .D(n6328), .CK(CLK), .Q(n18520), .QN(n22577) );
  DFF_X1 \REGISTERS_reg[27][53]  ( .D(n6327), .CK(CLK), .Q(n18537), .QN(n22578) );
  DFF_X1 \REGISTERS_reg[27][52]  ( .D(n6326), .CK(CLK), .Q(n18554), .QN(n22579) );
  DFF_X1 \REGISTERS_reg[27][51]  ( .D(n6325), .CK(CLK), .Q(n18571), .QN(n22580) );
  DFF_X1 \REGISTERS_reg[27][50]  ( .D(n6324), .CK(CLK), .Q(n18588), .QN(n22581) );
  DFF_X1 \REGISTERS_reg[27][49]  ( .D(n6323), .CK(CLK), .Q(n18605), .QN(n22582) );
  DFF_X1 \REGISTERS_reg[27][48]  ( .D(n6322), .CK(CLK), .Q(n18622), .QN(n22583) );
  DFF_X1 \REGISTERS_reg[27][47]  ( .D(n6321), .CK(CLK), .Q(n18639), .QN(n22584) );
  DFF_X1 \REGISTERS_reg[27][46]  ( .D(n6320), .CK(CLK), .Q(n18656), .QN(n22585) );
  DFF_X1 \REGISTERS_reg[27][45]  ( .D(n6319), .CK(CLK), .Q(n18673), .QN(n22586) );
  DFF_X1 \REGISTERS_reg[27][44]  ( .D(n6318), .CK(CLK), .Q(n18690), .QN(n22587) );
  DFF_X1 \REGISTERS_reg[27][43]  ( .D(n6317), .CK(CLK), .Q(n18707), .QN(n22588) );
  DFF_X1 \REGISTERS_reg[27][42]  ( .D(n6316), .CK(CLK), .Q(n18724), .QN(n22589) );
  DFF_X1 \REGISTERS_reg[27][41]  ( .D(n6315), .CK(CLK), .Q(n18741), .QN(n22590) );
  DFF_X1 \REGISTERS_reg[27][40]  ( .D(n6314), .CK(CLK), .Q(n18758), .QN(n22591) );
  DFF_X1 \REGISTERS_reg[27][39]  ( .D(n6313), .CK(CLK), .Q(n18775), .QN(n22592) );
  DFF_X1 \REGISTERS_reg[27][38]  ( .D(n6312), .CK(CLK), .Q(n18792), .QN(n22593) );
  DFF_X1 \REGISTERS_reg[27][37]  ( .D(n6311), .CK(CLK), .Q(n18809), .QN(n22594) );
  DFF_X1 \REGISTERS_reg[27][36]  ( .D(n6310), .CK(CLK), .Q(n18826), .QN(n22595) );
  DFF_X1 \REGISTERS_reg[27][35]  ( .D(n6309), .CK(CLK), .Q(n18843), .QN(n22596) );
  DFF_X1 \REGISTERS_reg[27][34]  ( .D(n6308), .CK(CLK), .Q(n18860), .QN(n22597) );
  DFF_X1 \REGISTERS_reg[27][33]  ( .D(n6307), .CK(CLK), .Q(n18877), .QN(n22598) );
  DFF_X1 \REGISTERS_reg[27][32]  ( .D(n6306), .CK(CLK), .Q(n18894), .QN(n22599) );
  DFF_X1 \REGISTERS_reg[27][31]  ( .D(n6305), .CK(CLK), .Q(n18911), .QN(n22600) );
  DFF_X1 \REGISTERS_reg[27][30]  ( .D(n6304), .CK(CLK), .Q(n18928), .QN(n22601) );
  DFF_X1 \REGISTERS_reg[27][29]  ( .D(n6303), .CK(CLK), .Q(n18945), .QN(n22602) );
  DFF_X1 \REGISTERS_reg[27][28]  ( .D(n6302), .CK(CLK), .Q(n18962), .QN(n22603) );
  DFF_X1 \REGISTERS_reg[27][27]  ( .D(n6301), .CK(CLK), .Q(n18979), .QN(n22604) );
  DFF_X1 \REGISTERS_reg[27][26]  ( .D(n6300), .CK(CLK), .Q(n18996), .QN(n22605) );
  DFF_X1 \REGISTERS_reg[27][25]  ( .D(n6299), .CK(CLK), .Q(n19013), .QN(n22606) );
  DFF_X1 \REGISTERS_reg[27][24]  ( .D(n6298), .CK(CLK), .Q(n19030), .QN(n22607) );
  DFF_X1 \REGISTERS_reg[27][23]  ( .D(n6297), .CK(CLK), .Q(n19047), .QN(n22608) );
  DFF_X1 \REGISTERS_reg[27][22]  ( .D(n6296), .CK(CLK), .Q(n19064), .QN(n22609) );
  DFF_X1 \REGISTERS_reg[27][21]  ( .D(n6295), .CK(CLK), .Q(n19081), .QN(n22610) );
  DFF_X1 \REGISTERS_reg[27][20]  ( .D(n6294), .CK(CLK), .Q(n19098), .QN(n22611) );
  DFF_X1 \REGISTERS_reg[27][19]  ( .D(n6293), .CK(CLK), .Q(n19115), .QN(n22612) );
  DFF_X1 \REGISTERS_reg[27][18]  ( .D(n6292), .CK(CLK), .Q(n19132), .QN(n22613) );
  DFF_X1 \REGISTERS_reg[27][17]  ( .D(n6291), .CK(CLK), .Q(n19149), .QN(n22614) );
  DFF_X1 \REGISTERS_reg[27][16]  ( .D(n6290), .CK(CLK), .Q(n19166), .QN(n22615) );
  DFF_X1 \REGISTERS_reg[27][15]  ( .D(n6289), .CK(CLK), .Q(n19183), .QN(n22616) );
  DFF_X1 \REGISTERS_reg[27][14]  ( .D(n6288), .CK(CLK), .Q(n19200), .QN(n22617) );
  DFF_X1 \REGISTERS_reg[27][13]  ( .D(n6287), .CK(CLK), .Q(n19217), .QN(n22618) );
  DFF_X1 \REGISTERS_reg[27][12]  ( .D(n6286), .CK(CLK), .Q(n19234), .QN(n22619) );
  DFF_X1 \REGISTERS_reg[27][11]  ( .D(n6285), .CK(CLK), .Q(n19251), .QN(n22620) );
  DFF_X1 \REGISTERS_reg[27][10]  ( .D(n6284), .CK(CLK), .Q(n19268), .QN(n22621) );
  DFF_X1 \REGISTERS_reg[27][9]  ( .D(n6283), .CK(CLK), .Q(n19285), .QN(n22622)
         );
  DFF_X1 \REGISTERS_reg[27][8]  ( .D(n6282), .CK(CLK), .Q(n19302), .QN(n22623)
         );
  DFF_X1 \REGISTERS_reg[27][7]  ( .D(n6281), .CK(CLK), .Q(n19319), .QN(n22624)
         );
  DFF_X1 \REGISTERS_reg[27][6]  ( .D(n6280), .CK(CLK), .Q(n19336), .QN(n22625)
         );
  DFF_X1 \REGISTERS_reg[27][5]  ( .D(n6279), .CK(CLK), .Q(n19353), .QN(n22626)
         );
  DFF_X1 \REGISTERS_reg[27][4]  ( .D(n6278), .CK(CLK), .Q(n19370), .QN(n22627)
         );
  DFF_X1 \REGISTERS_reg[27][3]  ( .D(n6277), .CK(CLK), .Q(n19387), .QN(n22628)
         );
  DFF_X1 \REGISTERS_reg[27][2]  ( .D(n6276), .CK(CLK), .Q(n19404), .QN(n22629)
         );
  DFF_X1 \REGISTERS_reg[27][1]  ( .D(n6275), .CK(CLK), .Q(n19421), .QN(n22630)
         );
  DFF_X1 \REGISTERS_reg[27][0]  ( .D(n6274), .CK(CLK), .Q(n19438), .QN(n22631)
         );
  DFF_X1 \REGISTERS_reg[2][59]  ( .D(n7933), .CK(CLK), .Q(n25358), .QN(n21420)
         );
  DFF_X1 \REGISTERS_reg[2][58]  ( .D(n7932), .CK(CLK), .Q(n25357), .QN(n21421)
         );
  DFF_X1 \REGISTERS_reg[2][57]  ( .D(n7931), .CK(CLK), .Q(n25356), .QN(n21422)
         );
  DFF_X1 \REGISTERS_reg[2][56]  ( .D(n7930), .CK(CLK), .Q(n25355), .QN(n21423)
         );
  DFF_X1 \REGISTERS_reg[2][55]  ( .D(n7929), .CK(CLK), .Q(n25354), .QN(n21424)
         );
  DFF_X1 \REGISTERS_reg[2][54]  ( .D(n7928), .CK(CLK), .Q(n25353), .QN(n21425)
         );
  DFF_X1 \REGISTERS_reg[2][53]  ( .D(n7927), .CK(CLK), .Q(n25352), .QN(n21426)
         );
  DFF_X1 \REGISTERS_reg[2][52]  ( .D(n7926), .CK(CLK), .Q(n25351), .QN(n21427)
         );
  DFF_X1 \REGISTERS_reg[2][51]  ( .D(n7925), .CK(CLK), .Q(n25350), .QN(n21428)
         );
  DFF_X1 \REGISTERS_reg[2][50]  ( .D(n7924), .CK(CLK), .Q(n25349), .QN(n21429)
         );
  DFF_X1 \REGISTERS_reg[2][49]  ( .D(n7923), .CK(CLK), .Q(n25348), .QN(n21430)
         );
  DFF_X1 \REGISTERS_reg[2][48]  ( .D(n7922), .CK(CLK), .Q(n25347), .QN(n21431)
         );
  DFF_X1 \REGISTERS_reg[2][47]  ( .D(n7921), .CK(CLK), .Q(n25346), .QN(n21432)
         );
  DFF_X1 \REGISTERS_reg[2][46]  ( .D(n7920), .CK(CLK), .Q(n25345), .QN(n21433)
         );
  DFF_X1 \REGISTERS_reg[2][45]  ( .D(n7919), .CK(CLK), .Q(n25344), .QN(n21434)
         );
  DFF_X1 \REGISTERS_reg[2][44]  ( .D(n7918), .CK(CLK), .Q(n25343), .QN(n21435)
         );
  DFF_X1 \REGISTERS_reg[2][43]  ( .D(n7917), .CK(CLK), .Q(n25342), .QN(n21436)
         );
  DFF_X1 \REGISTERS_reg[2][42]  ( .D(n7916), .CK(CLK), .Q(n25341), .QN(n21437)
         );
  DFF_X1 \REGISTERS_reg[2][41]  ( .D(n7915), .CK(CLK), .Q(n25340), .QN(n21438)
         );
  DFF_X1 \REGISTERS_reg[2][40]  ( .D(n7914), .CK(CLK), .Q(n25339), .QN(n21439)
         );
  DFF_X1 \REGISTERS_reg[2][39]  ( .D(n7913), .CK(CLK), .Q(n25338), .QN(n21440)
         );
  DFF_X1 \REGISTERS_reg[2][38]  ( .D(n7912), .CK(CLK), .Q(n25337), .QN(n21441)
         );
  DFF_X1 \REGISTERS_reg[2][37]  ( .D(n7911), .CK(CLK), .Q(n25336), .QN(n21442)
         );
  DFF_X1 \REGISTERS_reg[2][36]  ( .D(n7910), .CK(CLK), .Q(n25335), .QN(n21443)
         );
  DFF_X1 \REGISTERS_reg[2][35]  ( .D(n7909), .CK(CLK), .Q(n25334), .QN(n21444)
         );
  DFF_X1 \REGISTERS_reg[2][34]  ( .D(n7908), .CK(CLK), .Q(n25333), .QN(n21445)
         );
  DFF_X1 \REGISTERS_reg[2][33]  ( .D(n7907), .CK(CLK), .Q(n25332), .QN(n21446)
         );
  DFF_X1 \REGISTERS_reg[2][32]  ( .D(n7906), .CK(CLK), .Q(n25331), .QN(n21447)
         );
  DFF_X1 \REGISTERS_reg[2][31]  ( .D(n7905), .CK(CLK), .Q(n25330), .QN(n21448)
         );
  DFF_X1 \REGISTERS_reg[2][30]  ( .D(n7904), .CK(CLK), .Q(n25329), .QN(n21449)
         );
  DFF_X1 \REGISTERS_reg[2][29]  ( .D(n7903), .CK(CLK), .Q(n25328), .QN(n21450)
         );
  DFF_X1 \REGISTERS_reg[2][28]  ( .D(n7902), .CK(CLK), .Q(n25327), .QN(n21451)
         );
  DFF_X1 \REGISTERS_reg[2][27]  ( .D(n7901), .CK(CLK), .Q(n25326), .QN(n21452)
         );
  DFF_X1 \REGISTERS_reg[2][26]  ( .D(n7900), .CK(CLK), .Q(n25325), .QN(n21453)
         );
  DFF_X1 \REGISTERS_reg[2][25]  ( .D(n7899), .CK(CLK), .Q(n25324), .QN(n21454)
         );
  DFF_X1 \REGISTERS_reg[2][24]  ( .D(n7898), .CK(CLK), .Q(n25323), .QN(n21455)
         );
  DFF_X1 \REGISTERS_reg[2][23]  ( .D(n7897), .CK(CLK), .Q(n25322), .QN(n21456)
         );
  DFF_X1 \REGISTERS_reg[2][22]  ( .D(n7896), .CK(CLK), .Q(n25321), .QN(n21457)
         );
  DFF_X1 \REGISTERS_reg[2][21]  ( .D(n7895), .CK(CLK), .Q(n25320), .QN(n21458)
         );
  DFF_X1 \REGISTERS_reg[2][20]  ( .D(n7894), .CK(CLK), .Q(n25319), .QN(n21459)
         );
  DFF_X1 \REGISTERS_reg[2][19]  ( .D(n7893), .CK(CLK), .Q(n25318), .QN(n21460)
         );
  DFF_X1 \REGISTERS_reg[2][18]  ( .D(n7892), .CK(CLK), .Q(n25317), .QN(n21461)
         );
  DFF_X1 \REGISTERS_reg[2][17]  ( .D(n7891), .CK(CLK), .Q(n25316), .QN(n21462)
         );
  DFF_X1 \REGISTERS_reg[2][16]  ( .D(n7890), .CK(CLK), .Q(n25315), .QN(n21463)
         );
  DFF_X1 \REGISTERS_reg[2][15]  ( .D(n7889), .CK(CLK), .Q(n25314), .QN(n21464)
         );
  DFF_X1 \REGISTERS_reg[2][14]  ( .D(n7888), .CK(CLK), .Q(n25313), .QN(n21465)
         );
  DFF_X1 \REGISTERS_reg[2][13]  ( .D(n7887), .CK(CLK), .Q(n25312), .QN(n21466)
         );
  DFF_X1 \REGISTERS_reg[2][12]  ( .D(n7886), .CK(CLK), .Q(n25311), .QN(n21467)
         );
  DFF_X1 \REGISTERS_reg[2][11]  ( .D(n7885), .CK(CLK), .Q(n25654), .QN(n21468)
         );
  DFF_X1 \REGISTERS_reg[2][10]  ( .D(n7884), .CK(CLK), .Q(n25653), .QN(n21469)
         );
  DFF_X1 \REGISTERS_reg[2][9]  ( .D(n7883), .CK(CLK), .Q(n25652), .QN(n21470)
         );
  DFF_X1 \REGISTERS_reg[2][8]  ( .D(n7882), .CK(CLK), .Q(n25651), .QN(n21471)
         );
  DFF_X1 \REGISTERS_reg[2][7]  ( .D(n7881), .CK(CLK), .Q(n25650), .QN(n21472)
         );
  DFF_X1 \REGISTERS_reg[2][6]  ( .D(n7880), .CK(CLK), .Q(n25649), .QN(n21473)
         );
  DFF_X1 \REGISTERS_reg[2][5]  ( .D(n7879), .CK(CLK), .Q(n25648), .QN(n21474)
         );
  DFF_X1 \REGISTERS_reg[2][4]  ( .D(n7878), .CK(CLK), .Q(n25647), .QN(n21475)
         );
  DFF_X1 \REGISTERS_reg[2][3]  ( .D(n7877), .CK(CLK), .Q(n25646), .QN(n21476)
         );
  DFF_X1 \REGISTERS_reg[2][2]  ( .D(n7876), .CK(CLK), .Q(n25645), .QN(n21477)
         );
  DFF_X1 \REGISTERS_reg[2][1]  ( .D(n7875), .CK(CLK), .Q(n25644), .QN(n21478)
         );
  DFF_X1 \REGISTERS_reg[2][0]  ( .D(n7874), .CK(CLK), .Q(n25643), .QN(n21479)
         );
  DFF_X1 \REGISTERS_reg[31][63]  ( .D(n6081), .CK(CLK), .Q(n26194), .QN(n20899) );
  DFF_X1 \REGISTERS_reg[31][62]  ( .D(n6080), .CK(CLK), .Q(n26193), .QN(n20900) );
  DFF_X1 \REGISTERS_reg[31][61]  ( .D(n6079), .CK(CLK), .Q(n26192), .QN(n20901) );
  DFF_X1 \REGISTERS_reg[31][60]  ( .D(n6078), .CK(CLK), .Q(n26191), .QN(n20902) );
  DFF_X1 \REGISTERS_reg[29][63]  ( .D(n6209), .CK(CLK), .Q(n9249), .QN(n22244)
         );
  DFF_X1 \REGISTERS_reg[29][62]  ( .D(n6208), .CK(CLK), .Q(n9252), .QN(n22245)
         );
  DFF_X1 \REGISTERS_reg[29][61]  ( .D(n6207), .CK(CLK), .Q(n9255), .QN(n22246)
         );
  DFF_X1 \REGISTERS_reg[29][60]  ( .D(n6206), .CK(CLK), .Q(n9258), .QN(n22247)
         );
  DFF_X1 \REGISTERS_reg[22][63]  ( .D(n6657), .CK(CLK), .Q(n25695), .QN(n21492) );
  DFF_X1 \REGISTERS_reg[22][62]  ( .D(n6656), .CK(CLK), .Q(n25690), .QN(n21493) );
  DFF_X1 \REGISTERS_reg[22][61]  ( .D(n6655), .CK(CLK), .Q(n25685), .QN(n21494) );
  DFF_X1 \REGISTERS_reg[22][60]  ( .D(n6654), .CK(CLK), .Q(n25680), .QN(n21495) );
  DFF_X1 \REGISTERS_reg[18][63]  ( .D(n6913), .CK(CLK), .Q(n25696), .QN(n21484) );
  DFF_X1 \REGISTERS_reg[18][62]  ( .D(n6912), .CK(CLK), .Q(n25691), .QN(n21485) );
  DFF_X1 \REGISTERS_reg[18][61]  ( .D(n6911), .CK(CLK), .Q(n25686), .QN(n21486) );
  DFF_X1 \REGISTERS_reg[18][60]  ( .D(n6910), .CK(CLK), .Q(n25681), .QN(n21487) );
  DFF_X1 \REGISTERS_reg[10][63]  ( .D(n7425), .CK(CLK), .Q(n18382), .QN(n22252) );
  DFF_X1 \REGISTERS_reg[10][62]  ( .D(n7424), .CK(CLK), .Q(n18399), .QN(n22253) );
  DFF_X1 \REGISTERS_reg[10][61]  ( .D(n7423), .CK(CLK), .Q(n18416), .QN(n22254) );
  DFF_X1 \REGISTERS_reg[10][60]  ( .D(n7422), .CK(CLK), .Q(n18433), .QN(n22255) );
  DFF_X1 \REGISTERS_reg[1][63]  ( .D(n8001), .CK(CLK), .Q(n25578), .QN(n21512)
         );
  DFF_X1 \REGISTERS_reg[1][62]  ( .D(n8000), .CK(CLK), .Q(n25577), .QN(n21513)
         );
  DFF_X1 \REGISTERS_reg[1][61]  ( .D(n7999), .CK(CLK), .Q(n25576), .QN(n21514)
         );
  DFF_X1 \REGISTERS_reg[1][60]  ( .D(n7998), .CK(CLK), .Q(n25575), .QN(n21515)
         );
  DFF_X1 \REGISTERS_reg[16][63]  ( .D(n7041), .CK(CLK), .Q(n25697), .QN(n21160) );
  DFF_X1 \REGISTERS_reg[16][62]  ( .D(n7040), .CK(CLK), .Q(n25692), .QN(n21161) );
  DFF_X1 \REGISTERS_reg[16][61]  ( .D(n7039), .CK(CLK), .Q(n25687), .QN(n21162) );
  DFF_X1 \REGISTERS_reg[16][60]  ( .D(n7038), .CK(CLK), .Q(n25682), .QN(n21163) );
  DFF_X1 \REGISTERS_reg[6][63]  ( .D(n7681), .CK(CLK), .Q(n25558), .QN(n21496)
         );
  DFF_X1 \REGISTERS_reg[6][62]  ( .D(n7680), .CK(CLK), .Q(n25557), .QN(n21497)
         );
  DFF_X1 \REGISTERS_reg[6][61]  ( .D(n7679), .CK(CLK), .Q(n25556), .QN(n21498)
         );
  DFF_X1 \REGISTERS_reg[6][60]  ( .D(n7678), .CK(CLK), .Q(n25555), .QN(n21499)
         );
  DFF_X1 \REGISTERS_reg[31][59]  ( .D(n6077), .CK(CLK), .Q(n26266), .QN(n20903) );
  DFF_X1 \REGISTERS_reg[31][58]  ( .D(n6076), .CK(CLK), .Q(n26265), .QN(n20904) );
  DFF_X1 \REGISTERS_reg[31][57]  ( .D(n6075), .CK(CLK), .Q(n26264), .QN(n20905) );
  DFF_X1 \REGISTERS_reg[31][56]  ( .D(n6074), .CK(CLK), .Q(n26263), .QN(n20906) );
  DFF_X1 \REGISTERS_reg[31][55]  ( .D(n6073), .CK(CLK), .Q(n26262), .QN(n20907) );
  DFF_X1 \REGISTERS_reg[31][54]  ( .D(n6072), .CK(CLK), .Q(n26261), .QN(n20908) );
  DFF_X1 \REGISTERS_reg[31][53]  ( .D(n6071), .CK(CLK), .Q(n26260), .QN(n20909) );
  DFF_X1 \REGISTERS_reg[31][52]  ( .D(n6070), .CK(CLK), .Q(n26259), .QN(n20910) );
  DFF_X1 \REGISTERS_reg[31][51]  ( .D(n6069), .CK(CLK), .Q(n26258), .QN(n20911) );
  DFF_X1 \REGISTERS_reg[31][50]  ( .D(n6068), .CK(CLK), .Q(n26257), .QN(n20912) );
  DFF_X1 \REGISTERS_reg[31][49]  ( .D(n6067), .CK(CLK), .Q(n26256), .QN(n20913) );
  DFF_X1 \REGISTERS_reg[31][48]  ( .D(n6066), .CK(CLK), .Q(n26255), .QN(n20914) );
  DFF_X1 \REGISTERS_reg[31][47]  ( .D(n6065), .CK(CLK), .Q(n26254), .QN(n20915) );
  DFF_X1 \REGISTERS_reg[31][46]  ( .D(n6064), .CK(CLK), .Q(n26253), .QN(n20916) );
  DFF_X1 \REGISTERS_reg[31][45]  ( .D(n6063), .CK(CLK), .Q(n26252), .QN(n20917) );
  DFF_X1 \REGISTERS_reg[31][44]  ( .D(n6062), .CK(CLK), .Q(n26251), .QN(n20918) );
  DFF_X1 \REGISTERS_reg[31][43]  ( .D(n6061), .CK(CLK), .Q(n26250), .QN(n20919) );
  DFF_X1 \REGISTERS_reg[31][42]  ( .D(n6060), .CK(CLK), .Q(n26249), .QN(n20920) );
  DFF_X1 \REGISTERS_reg[31][41]  ( .D(n6059), .CK(CLK), .Q(n26248), .QN(n20921) );
  DFF_X1 \REGISTERS_reg[31][40]  ( .D(n6058), .CK(CLK), .Q(n26247), .QN(n20922) );
  DFF_X1 \REGISTERS_reg[31][39]  ( .D(n6057), .CK(CLK), .Q(n26246), .QN(n20923) );
  DFF_X1 \REGISTERS_reg[31][38]  ( .D(n6056), .CK(CLK), .Q(n26245), .QN(n20924) );
  DFF_X1 \REGISTERS_reg[31][37]  ( .D(n6055), .CK(CLK), .Q(n26244), .QN(n20925) );
  DFF_X1 \REGISTERS_reg[31][36]  ( .D(n6054), .CK(CLK), .Q(n26243), .QN(n20926) );
  DFF_X1 \REGISTERS_reg[31][35]  ( .D(n6053), .CK(CLK), .Q(n26242), .QN(n20927) );
  DFF_X1 \REGISTERS_reg[31][34]  ( .D(n6052), .CK(CLK), .Q(n26241), .QN(n20928) );
  DFF_X1 \REGISTERS_reg[31][33]  ( .D(n6051), .CK(CLK), .Q(n26240), .QN(n20929) );
  DFF_X1 \REGISTERS_reg[31][32]  ( .D(n6050), .CK(CLK), .Q(n26239), .QN(n20930) );
  DFF_X1 \REGISTERS_reg[31][31]  ( .D(n6049), .CK(CLK), .Q(n26238), .QN(n20931) );
  DFF_X1 \REGISTERS_reg[31][30]  ( .D(n6048), .CK(CLK), .Q(n26237), .QN(n20932) );
  DFF_X1 \REGISTERS_reg[31][29]  ( .D(n6047), .CK(CLK), .Q(n26236), .QN(n20933) );
  DFF_X1 \REGISTERS_reg[31][28]  ( .D(n6046), .CK(CLK), .Q(n26235), .QN(n20934) );
  DFF_X1 \REGISTERS_reg[31][27]  ( .D(n6045), .CK(CLK), .Q(n26234), .QN(n20935) );
  DFF_X1 \REGISTERS_reg[31][26]  ( .D(n6044), .CK(CLK), .Q(n26233), .QN(n20936) );
  DFF_X1 \REGISTERS_reg[31][25]  ( .D(n6043), .CK(CLK), .Q(n26232), .QN(n20937) );
  DFF_X1 \REGISTERS_reg[31][24]  ( .D(n6042), .CK(CLK), .Q(n26231), .QN(n20938) );
  DFF_X1 \REGISTERS_reg[31][23]  ( .D(n6041), .CK(CLK), .Q(n26230), .QN(n20939) );
  DFF_X1 \REGISTERS_reg[31][22]  ( .D(n6040), .CK(CLK), .Q(n26229), .QN(n20940) );
  DFF_X1 \REGISTERS_reg[31][21]  ( .D(n6039), .CK(CLK), .Q(n26228), .QN(n20941) );
  DFF_X1 \REGISTERS_reg[31][20]  ( .D(n6038), .CK(CLK), .Q(n26227), .QN(n20942) );
  DFF_X1 \REGISTERS_reg[31][19]  ( .D(n6037), .CK(CLK), .Q(n26226), .QN(n20943) );
  DFF_X1 \REGISTERS_reg[31][18]  ( .D(n6036), .CK(CLK), .Q(n26225), .QN(n20944) );
  DFF_X1 \REGISTERS_reg[31][17]  ( .D(n6035), .CK(CLK), .Q(n26224), .QN(n20945) );
  DFF_X1 \REGISTERS_reg[31][16]  ( .D(n6034), .CK(CLK), .Q(n26223), .QN(n20946) );
  DFF_X1 \REGISTERS_reg[31][15]  ( .D(n6033), .CK(CLK), .Q(n26222), .QN(n20947) );
  DFF_X1 \REGISTERS_reg[31][14]  ( .D(n6032), .CK(CLK), .Q(n26221), .QN(n20948) );
  DFF_X1 \REGISTERS_reg[31][13]  ( .D(n6031), .CK(CLK), .Q(n26220), .QN(n20949) );
  DFF_X1 \REGISTERS_reg[31][12]  ( .D(n6030), .CK(CLK), .Q(n26219), .QN(n20950) );
  DFF_X1 \REGISTERS_reg[31][11]  ( .D(n6029), .CK(CLK), .Q(n26218), .QN(n20951) );
  DFF_X1 \REGISTERS_reg[31][10]  ( .D(n6028), .CK(CLK), .Q(n26217), .QN(n20952) );
  DFF_X1 \REGISTERS_reg[31][9]  ( .D(n6027), .CK(CLK), .Q(n26216), .QN(n20953)
         );
  DFF_X1 \REGISTERS_reg[31][8]  ( .D(n6026), .CK(CLK), .Q(n26215), .QN(n20954)
         );
  DFF_X1 \REGISTERS_reg[31][7]  ( .D(n6025), .CK(CLK), .Q(n26214), .QN(n20955)
         );
  DFF_X1 \REGISTERS_reg[31][6]  ( .D(n6024), .CK(CLK), .Q(n26213), .QN(n20956)
         );
  DFF_X1 \REGISTERS_reg[31][5]  ( .D(n6023), .CK(CLK), .Q(n26212), .QN(n20957)
         );
  DFF_X1 \REGISTERS_reg[31][4]  ( .D(n6022), .CK(CLK), .Q(n26211), .QN(n20958)
         );
  DFF_X1 \REGISTERS_reg[31][3]  ( .D(n6021), .CK(CLK), .Q(n26210), .QN(n20959)
         );
  DFF_X1 \REGISTERS_reg[31][2]  ( .D(n6020), .CK(CLK), .Q(n26209), .QN(n20960)
         );
  DFF_X1 \REGISTERS_reg[31][1]  ( .D(n6019), .CK(CLK), .Q(n26208), .QN(n20961)
         );
  DFF_X1 \REGISTERS_reg[31][0]  ( .D(n6018), .CK(CLK), .Q(n26207), .QN(n20962)
         );
  DFF_X1 \REGISTERS_reg[29][59]  ( .D(n6205), .CK(CLK), .Q(n9261), .QN(n22260)
         );
  DFF_X1 \REGISTERS_reg[29][58]  ( .D(n6204), .CK(CLK), .Q(n9264), .QN(n22261)
         );
  DFF_X1 \REGISTERS_reg[29][57]  ( .D(n6203), .CK(CLK), .Q(n9267), .QN(n22262)
         );
  DFF_X1 \REGISTERS_reg[29][56]  ( .D(n6202), .CK(CLK), .Q(n9270), .QN(n22263)
         );
  DFF_X1 \REGISTERS_reg[29][55]  ( .D(n6201), .CK(CLK), .Q(n9273), .QN(n22264)
         );
  DFF_X1 \REGISTERS_reg[29][54]  ( .D(n6200), .CK(CLK), .Q(n9276), .QN(n22265)
         );
  DFF_X1 \REGISTERS_reg[29][53]  ( .D(n6199), .CK(CLK), .Q(n9279), .QN(n22266)
         );
  DFF_X1 \REGISTERS_reg[29][52]  ( .D(n6198), .CK(CLK), .Q(n9282), .QN(n22267)
         );
  DFF_X1 \REGISTERS_reg[29][51]  ( .D(n6197), .CK(CLK), .Q(n9285), .QN(n22268)
         );
  DFF_X1 \REGISTERS_reg[29][50]  ( .D(n6196), .CK(CLK), .Q(n9288), .QN(n22269)
         );
  DFF_X1 \REGISTERS_reg[29][49]  ( .D(n6195), .CK(CLK), .Q(n9291), .QN(n22270)
         );
  DFF_X1 \REGISTERS_reg[29][48]  ( .D(n6194), .CK(CLK), .Q(n9294), .QN(n22271)
         );
  DFF_X1 \REGISTERS_reg[29][47]  ( .D(n6193), .CK(CLK), .Q(n9297), .QN(n22272)
         );
  DFF_X1 \REGISTERS_reg[29][46]  ( .D(n6192), .CK(CLK), .Q(n9300), .QN(n22273)
         );
  DFF_X1 \REGISTERS_reg[29][45]  ( .D(n6191), .CK(CLK), .Q(n9303), .QN(n22274)
         );
  DFF_X1 \REGISTERS_reg[29][44]  ( .D(n6190), .CK(CLK), .Q(n9306), .QN(n22275)
         );
  DFF_X1 \REGISTERS_reg[29][43]  ( .D(n6189), .CK(CLK), .Q(n9309), .QN(n22276)
         );
  DFF_X1 \REGISTERS_reg[29][42]  ( .D(n6188), .CK(CLK), .Q(n9312), .QN(n22277)
         );
  DFF_X1 \REGISTERS_reg[29][41]  ( .D(n6187), .CK(CLK), .Q(n9315), .QN(n22278)
         );
  DFF_X1 \REGISTERS_reg[29][40]  ( .D(n6186), .CK(CLK), .Q(n9318), .QN(n22279)
         );
  DFF_X1 \REGISTERS_reg[29][39]  ( .D(n6185), .CK(CLK), .Q(n9321), .QN(n22280)
         );
  DFF_X1 \REGISTERS_reg[29][38]  ( .D(n6184), .CK(CLK), .Q(n9324), .QN(n22281)
         );
  DFF_X1 \REGISTERS_reg[29][37]  ( .D(n6183), .CK(CLK), .Q(n9327), .QN(n22282)
         );
  DFF_X1 \REGISTERS_reg[29][36]  ( .D(n6182), .CK(CLK), .Q(n9330), .QN(n22283)
         );
  DFF_X1 \REGISTERS_reg[29][35]  ( .D(n6181), .CK(CLK), .Q(n9333), .QN(n22284)
         );
  DFF_X1 \REGISTERS_reg[29][34]  ( .D(n6180), .CK(CLK), .Q(n9336), .QN(n22285)
         );
  DFF_X1 \REGISTERS_reg[29][33]  ( .D(n6179), .CK(CLK), .Q(n9339), .QN(n22286)
         );
  DFF_X1 \REGISTERS_reg[29][32]  ( .D(n6178), .CK(CLK), .Q(n9342), .QN(n22287)
         );
  DFF_X1 \REGISTERS_reg[29][31]  ( .D(n6177), .CK(CLK), .Q(n9345), .QN(n22288)
         );
  DFF_X1 \REGISTERS_reg[29][30]  ( .D(n6176), .CK(CLK), .Q(n9348), .QN(n22289)
         );
  DFF_X1 \REGISTERS_reg[29][29]  ( .D(n6175), .CK(CLK), .Q(n9351), .QN(n22290)
         );
  DFF_X1 \REGISTERS_reg[29][28]  ( .D(n6174), .CK(CLK), .Q(n9354), .QN(n22291)
         );
  DFF_X1 \REGISTERS_reg[29][27]  ( .D(n6173), .CK(CLK), .Q(n9357), .QN(n22292)
         );
  DFF_X1 \REGISTERS_reg[29][26]  ( .D(n6172), .CK(CLK), .Q(n9360), .QN(n22293)
         );
  DFF_X1 \REGISTERS_reg[29][25]  ( .D(n6171), .CK(CLK), .Q(n9363), .QN(n22294)
         );
  DFF_X1 \REGISTERS_reg[29][24]  ( .D(n6170), .CK(CLK), .Q(n9366), .QN(n22295)
         );
  DFF_X1 \REGISTERS_reg[29][23]  ( .D(n6169), .CK(CLK), .Q(n9369), .QN(n22296)
         );
  DFF_X1 \REGISTERS_reg[29][22]  ( .D(n6168), .CK(CLK), .Q(n9372), .QN(n22297)
         );
  DFF_X1 \REGISTERS_reg[29][21]  ( .D(n6167), .CK(CLK), .Q(n9375), .QN(n22298)
         );
  DFF_X1 \REGISTERS_reg[29][20]  ( .D(n6166), .CK(CLK), .Q(n9378), .QN(n22299)
         );
  DFF_X1 \REGISTERS_reg[29][19]  ( .D(n6165), .CK(CLK), .Q(n9381), .QN(n22300)
         );
  DFF_X1 \REGISTERS_reg[29][18]  ( .D(n6164), .CK(CLK), .Q(n9384), .QN(n22301)
         );
  DFF_X1 \REGISTERS_reg[29][17]  ( .D(n6163), .CK(CLK), .Q(n9387), .QN(n22302)
         );
  DFF_X1 \REGISTERS_reg[29][16]  ( .D(n6162), .CK(CLK), .Q(n9390), .QN(n22303)
         );
  DFF_X1 \REGISTERS_reg[29][15]  ( .D(n6161), .CK(CLK), .Q(n9393), .QN(n22304)
         );
  DFF_X1 \REGISTERS_reg[29][14]  ( .D(n6160), .CK(CLK), .Q(n9396), .QN(n22305)
         );
  DFF_X1 \REGISTERS_reg[29][13]  ( .D(n6159), .CK(CLK), .Q(n9399), .QN(n22306)
         );
  DFF_X1 \REGISTERS_reg[29][12]  ( .D(n6158), .CK(CLK), .Q(n9402), .QN(n22307)
         );
  DFF_X1 \REGISTERS_reg[29][11]  ( .D(n6157), .CK(CLK), .Q(n9405), .QN(n22308)
         );
  DFF_X1 \REGISTERS_reg[29][10]  ( .D(n6156), .CK(CLK), .Q(n9408), .QN(n22309)
         );
  DFF_X1 \REGISTERS_reg[29][9]  ( .D(n6155), .CK(CLK), .Q(n9411), .QN(n22310)
         );
  DFF_X1 \REGISTERS_reg[29][8]  ( .D(n6154), .CK(CLK), .Q(n9414), .QN(n22311)
         );
  DFF_X1 \REGISTERS_reg[29][7]  ( .D(n6153), .CK(CLK), .Q(n9417), .QN(n22312)
         );
  DFF_X1 \REGISTERS_reg[29][6]  ( .D(n6152), .CK(CLK), .Q(n9420), .QN(n22313)
         );
  DFF_X1 \REGISTERS_reg[29][5]  ( .D(n6151), .CK(CLK), .Q(n9423), .QN(n22314)
         );
  DFF_X1 \REGISTERS_reg[29][4]  ( .D(n6150), .CK(CLK), .Q(n9426), .QN(n22315)
         );
  DFF_X1 \REGISTERS_reg[29][3]  ( .D(n6149), .CK(CLK), .Q(n9429), .QN(n22316)
         );
  DFF_X1 \REGISTERS_reg[29][2]  ( .D(n6148), .CK(CLK), .Q(n9432), .QN(n22317)
         );
  DFF_X1 \REGISTERS_reg[29][1]  ( .D(n6147), .CK(CLK), .Q(n9435), .QN(n22318)
         );
  DFF_X1 \REGISTERS_reg[29][0]  ( .D(n6146), .CK(CLK), .Q(n9438), .QN(n22319)
         );
  DFF_X1 \REGISTERS_reg[22][59]  ( .D(n6653), .CK(CLK), .Q(n25995), .QN(n21760) );
  DFF_X1 \REGISTERS_reg[22][58]  ( .D(n6652), .CK(CLK), .Q(n25990), .QN(n21761) );
  DFF_X1 \REGISTERS_reg[22][57]  ( .D(n6651), .CK(CLK), .Q(n25985), .QN(n21762) );
  DFF_X1 \REGISTERS_reg[22][56]  ( .D(n6650), .CK(CLK), .Q(n25980), .QN(n21763) );
  DFF_X1 \REGISTERS_reg[22][55]  ( .D(n6649), .CK(CLK), .Q(n25975), .QN(n21764) );
  DFF_X1 \REGISTERS_reg[22][54]  ( .D(n6648), .CK(CLK), .Q(n25970), .QN(n21765) );
  DFF_X1 \REGISTERS_reg[22][53]  ( .D(n6647), .CK(CLK), .Q(n25965), .QN(n21766) );
  DFF_X1 \REGISTERS_reg[22][52]  ( .D(n6646), .CK(CLK), .Q(n25960), .QN(n21767) );
  DFF_X1 \REGISTERS_reg[22][51]  ( .D(n6645), .CK(CLK), .Q(n25955), .QN(n21768) );
  DFF_X1 \REGISTERS_reg[22][50]  ( .D(n6644), .CK(CLK), .Q(n25950), .QN(n21769) );
  DFF_X1 \REGISTERS_reg[22][49]  ( .D(n6643), .CK(CLK), .Q(n25945), .QN(n21770) );
  DFF_X1 \REGISTERS_reg[22][48]  ( .D(n6642), .CK(CLK), .Q(n25940), .QN(n21771) );
  DFF_X1 \REGISTERS_reg[22][47]  ( .D(n6641), .CK(CLK), .Q(n25935), .QN(n21772) );
  DFF_X1 \REGISTERS_reg[22][46]  ( .D(n6640), .CK(CLK), .Q(n25930), .QN(n21773) );
  DFF_X1 \REGISTERS_reg[22][45]  ( .D(n6639), .CK(CLK), .Q(n25925), .QN(n21774) );
  DFF_X1 \REGISTERS_reg[22][44]  ( .D(n6638), .CK(CLK), .Q(n25920), .QN(n21775) );
  DFF_X1 \REGISTERS_reg[22][43]  ( .D(n6637), .CK(CLK), .Q(n25915), .QN(n21776) );
  DFF_X1 \REGISTERS_reg[22][42]  ( .D(n6636), .CK(CLK), .Q(n25910), .QN(n21777) );
  DFF_X1 \REGISTERS_reg[22][41]  ( .D(n6635), .CK(CLK), .Q(n25905), .QN(n21778) );
  DFF_X1 \REGISTERS_reg[22][40]  ( .D(n6634), .CK(CLK), .Q(n25900), .QN(n21779) );
  DFF_X1 \REGISTERS_reg[22][39]  ( .D(n6633), .CK(CLK), .Q(n25895), .QN(n21780) );
  DFF_X1 \REGISTERS_reg[22][38]  ( .D(n6632), .CK(CLK), .Q(n25890), .QN(n21781) );
  DFF_X1 \REGISTERS_reg[22][37]  ( .D(n6631), .CK(CLK), .Q(n25885), .QN(n21782) );
  DFF_X1 \REGISTERS_reg[22][36]  ( .D(n6630), .CK(CLK), .Q(n25880), .QN(n21783) );
  DFF_X1 \REGISTERS_reg[22][35]  ( .D(n6629), .CK(CLK), .Q(n25875), .QN(n21784) );
  DFF_X1 \REGISTERS_reg[22][34]  ( .D(n6628), .CK(CLK), .Q(n25870), .QN(n21785) );
  DFF_X1 \REGISTERS_reg[22][33]  ( .D(n6627), .CK(CLK), .Q(n25865), .QN(n21786) );
  DFF_X1 \REGISTERS_reg[22][32]  ( .D(n6626), .CK(CLK), .Q(n25860), .QN(n21787) );
  DFF_X1 \REGISTERS_reg[22][31]  ( .D(n6625), .CK(CLK), .Q(n25855), .QN(n21788) );
  DFF_X1 \REGISTERS_reg[22][30]  ( .D(n6624), .CK(CLK), .Q(n25850), .QN(n21789) );
  DFF_X1 \REGISTERS_reg[22][29]  ( .D(n6623), .CK(CLK), .Q(n25845), .QN(n21790) );
  DFF_X1 \REGISTERS_reg[22][28]  ( .D(n6622), .CK(CLK), .Q(n25840), .QN(n21791) );
  DFF_X1 \REGISTERS_reg[22][27]  ( .D(n6621), .CK(CLK), .Q(n25835), .QN(n21792) );
  DFF_X1 \REGISTERS_reg[22][26]  ( .D(n6620), .CK(CLK), .Q(n25830), .QN(n21793) );
  DFF_X1 \REGISTERS_reg[22][25]  ( .D(n6619), .CK(CLK), .Q(n25825), .QN(n21794) );
  DFF_X1 \REGISTERS_reg[22][24]  ( .D(n6618), .CK(CLK), .Q(n25820), .QN(n21795) );
  DFF_X1 \REGISTERS_reg[22][23]  ( .D(n6617), .CK(CLK), .Q(n25815), .QN(n21796) );
  DFF_X1 \REGISTERS_reg[22][22]  ( .D(n6616), .CK(CLK), .Q(n25810), .QN(n21797) );
  DFF_X1 \REGISTERS_reg[22][21]  ( .D(n6615), .CK(CLK), .Q(n25805), .QN(n21798) );
  DFF_X1 \REGISTERS_reg[22][20]  ( .D(n6614), .CK(CLK), .Q(n25800), .QN(n21799) );
  DFF_X1 \REGISTERS_reg[22][19]  ( .D(n6613), .CK(CLK), .Q(n25795), .QN(n21800) );
  DFF_X1 \REGISTERS_reg[22][18]  ( .D(n6612), .CK(CLK), .Q(n25790), .QN(n21801) );
  DFF_X1 \REGISTERS_reg[22][17]  ( .D(n6611), .CK(CLK), .Q(n25785), .QN(n21802) );
  DFF_X1 \REGISTERS_reg[22][16]  ( .D(n6610), .CK(CLK), .Q(n25780), .QN(n21803) );
  DFF_X1 \REGISTERS_reg[22][15]  ( .D(n6609), .CK(CLK), .Q(n25775), .QN(n21804) );
  DFF_X1 \REGISTERS_reg[22][14]  ( .D(n6608), .CK(CLK), .Q(n25770), .QN(n21805) );
  DFF_X1 \REGISTERS_reg[22][13]  ( .D(n6607), .CK(CLK), .Q(n25765), .QN(n21806) );
  DFF_X1 \REGISTERS_reg[22][12]  ( .D(n6606), .CK(CLK), .Q(n25760), .QN(n21807) );
  DFF_X1 \REGISTERS_reg[22][11]  ( .D(n6605), .CK(CLK), .Q(n25755), .QN(n21808) );
  DFF_X1 \REGISTERS_reg[22][10]  ( .D(n6604), .CK(CLK), .Q(n25750), .QN(n21809) );
  DFF_X1 \REGISTERS_reg[22][9]  ( .D(n6603), .CK(CLK), .Q(n25745), .QN(n21810)
         );
  DFF_X1 \REGISTERS_reg[22][8]  ( .D(n6602), .CK(CLK), .Q(n25740), .QN(n21811)
         );
  DFF_X1 \REGISTERS_reg[22][7]  ( .D(n6601), .CK(CLK), .Q(n25735), .QN(n21812)
         );
  DFF_X1 \REGISTERS_reg[22][6]  ( .D(n6600), .CK(CLK), .Q(n25730), .QN(n21813)
         );
  DFF_X1 \REGISTERS_reg[22][5]  ( .D(n6599), .CK(CLK), .Q(n25725), .QN(n21814)
         );
  DFF_X1 \REGISTERS_reg[22][4]  ( .D(n6598), .CK(CLK), .Q(n25720), .QN(n21815)
         );
  DFF_X1 \REGISTERS_reg[22][3]  ( .D(n6597), .CK(CLK), .Q(n25715), .QN(n21816)
         );
  DFF_X1 \REGISTERS_reg[22][2]  ( .D(n6596), .CK(CLK), .Q(n25710), .QN(n21817)
         );
  DFF_X1 \REGISTERS_reg[22][1]  ( .D(n6595), .CK(CLK), .Q(n25705), .QN(n21818)
         );
  DFF_X1 \REGISTERS_reg[22][0]  ( .D(n6594), .CK(CLK), .Q(n25700), .QN(n21819)
         );
  DFF_X1 \REGISTERS_reg[18][59]  ( .D(n6909), .CK(CLK), .Q(n25996), .QN(n21640) );
  DFF_X1 \REGISTERS_reg[18][58]  ( .D(n6908), .CK(CLK), .Q(n25991), .QN(n21641) );
  DFF_X1 \REGISTERS_reg[18][57]  ( .D(n6907), .CK(CLK), .Q(n25986), .QN(n21642) );
  DFF_X1 \REGISTERS_reg[18][56]  ( .D(n6906), .CK(CLK), .Q(n25981), .QN(n21643) );
  DFF_X1 \REGISTERS_reg[18][55]  ( .D(n6905), .CK(CLK), .Q(n25976), .QN(n21644) );
  DFF_X1 \REGISTERS_reg[18][54]  ( .D(n6904), .CK(CLK), .Q(n25971), .QN(n21645) );
  DFF_X1 \REGISTERS_reg[18][53]  ( .D(n6903), .CK(CLK), .Q(n25966), .QN(n21646) );
  DFF_X1 \REGISTERS_reg[18][52]  ( .D(n6902), .CK(CLK), .Q(n25961), .QN(n21647) );
  DFF_X1 \REGISTERS_reg[18][51]  ( .D(n6901), .CK(CLK), .Q(n25956), .QN(n21648) );
  DFF_X1 \REGISTERS_reg[18][50]  ( .D(n6900), .CK(CLK), .Q(n25951), .QN(n21649) );
  DFF_X1 \REGISTERS_reg[18][49]  ( .D(n6899), .CK(CLK), .Q(n25946), .QN(n21650) );
  DFF_X1 \REGISTERS_reg[18][48]  ( .D(n6898), .CK(CLK), .Q(n25941), .QN(n21651) );
  DFF_X1 \REGISTERS_reg[18][47]  ( .D(n6897), .CK(CLK), .Q(n25936), .QN(n21652) );
  DFF_X1 \REGISTERS_reg[18][46]  ( .D(n6896), .CK(CLK), .Q(n25931), .QN(n21653) );
  DFF_X1 \REGISTERS_reg[18][45]  ( .D(n6895), .CK(CLK), .Q(n25926), .QN(n21654) );
  DFF_X1 \REGISTERS_reg[18][44]  ( .D(n6894), .CK(CLK), .Q(n25921), .QN(n21655) );
  DFF_X1 \REGISTERS_reg[18][43]  ( .D(n6893), .CK(CLK), .Q(n25916), .QN(n21656) );
  DFF_X1 \REGISTERS_reg[18][42]  ( .D(n6892), .CK(CLK), .Q(n25911), .QN(n21657) );
  DFF_X1 \REGISTERS_reg[18][41]  ( .D(n6891), .CK(CLK), .Q(n25906), .QN(n21658) );
  DFF_X1 \REGISTERS_reg[18][40]  ( .D(n6890), .CK(CLK), .Q(n25901), .QN(n21659) );
  DFF_X1 \REGISTERS_reg[18][39]  ( .D(n6889), .CK(CLK), .Q(n25896), .QN(n21660) );
  DFF_X1 \REGISTERS_reg[18][38]  ( .D(n6888), .CK(CLK), .Q(n25891), .QN(n21661) );
  DFF_X1 \REGISTERS_reg[18][37]  ( .D(n6887), .CK(CLK), .Q(n25886), .QN(n21662) );
  DFF_X1 \REGISTERS_reg[18][36]  ( .D(n6886), .CK(CLK), .Q(n25881), .QN(n21663) );
  DFF_X1 \REGISTERS_reg[18][35]  ( .D(n6885), .CK(CLK), .Q(n25876), .QN(n21664) );
  DFF_X1 \REGISTERS_reg[18][34]  ( .D(n6884), .CK(CLK), .Q(n25871), .QN(n21665) );
  DFF_X1 \REGISTERS_reg[18][33]  ( .D(n6883), .CK(CLK), .Q(n25866), .QN(n21666) );
  DFF_X1 \REGISTERS_reg[18][32]  ( .D(n6882), .CK(CLK), .Q(n25861), .QN(n21667) );
  DFF_X1 \REGISTERS_reg[18][31]  ( .D(n6881), .CK(CLK), .Q(n25856), .QN(n21668) );
  DFF_X1 \REGISTERS_reg[18][30]  ( .D(n6880), .CK(CLK), .Q(n25851), .QN(n21669) );
  DFF_X1 \REGISTERS_reg[18][29]  ( .D(n6879), .CK(CLK), .Q(n25846), .QN(n21670) );
  DFF_X1 \REGISTERS_reg[18][28]  ( .D(n6878), .CK(CLK), .Q(n25841), .QN(n21671) );
  DFF_X1 \REGISTERS_reg[18][27]  ( .D(n6877), .CK(CLK), .Q(n25836), .QN(n21672) );
  DFF_X1 \REGISTERS_reg[18][26]  ( .D(n6876), .CK(CLK), .Q(n25831), .QN(n21673) );
  DFF_X1 \REGISTERS_reg[18][25]  ( .D(n6875), .CK(CLK), .Q(n25826), .QN(n21674) );
  DFF_X1 \REGISTERS_reg[18][24]  ( .D(n6874), .CK(CLK), .Q(n25821), .QN(n21675) );
  DFF_X1 \REGISTERS_reg[18][23]  ( .D(n6873), .CK(CLK), .Q(n25816), .QN(n21676) );
  DFF_X1 \REGISTERS_reg[18][22]  ( .D(n6872), .CK(CLK), .Q(n25811), .QN(n21677) );
  DFF_X1 \REGISTERS_reg[18][21]  ( .D(n6871), .CK(CLK), .Q(n25806), .QN(n21678) );
  DFF_X1 \REGISTERS_reg[18][20]  ( .D(n6870), .CK(CLK), .Q(n25801), .QN(n21679) );
  DFF_X1 \REGISTERS_reg[18][19]  ( .D(n6869), .CK(CLK), .Q(n25796), .QN(n21680) );
  DFF_X1 \REGISTERS_reg[18][18]  ( .D(n6868), .CK(CLK), .Q(n25791), .QN(n21681) );
  DFF_X1 \REGISTERS_reg[18][17]  ( .D(n6867), .CK(CLK), .Q(n25786), .QN(n21682) );
  DFF_X1 \REGISTERS_reg[18][16]  ( .D(n6866), .CK(CLK), .Q(n25781), .QN(n21683) );
  DFF_X1 \REGISTERS_reg[18][15]  ( .D(n6865), .CK(CLK), .Q(n25776), .QN(n21684) );
  DFF_X1 \REGISTERS_reg[18][14]  ( .D(n6864), .CK(CLK), .Q(n25771), .QN(n21685) );
  DFF_X1 \REGISTERS_reg[18][13]  ( .D(n6863), .CK(CLK), .Q(n25766), .QN(n21686) );
  DFF_X1 \REGISTERS_reg[18][12]  ( .D(n6862), .CK(CLK), .Q(n25761), .QN(n21687) );
  DFF_X1 \REGISTERS_reg[18][11]  ( .D(n6861), .CK(CLK), .Q(n25756), .QN(n21688) );
  DFF_X1 \REGISTERS_reg[18][10]  ( .D(n6860), .CK(CLK), .Q(n25751), .QN(n21689) );
  DFF_X1 \REGISTERS_reg[18][9]  ( .D(n6859), .CK(CLK), .Q(n25746), .QN(n21690)
         );
  DFF_X1 \REGISTERS_reg[18][8]  ( .D(n6858), .CK(CLK), .Q(n25741), .QN(n21691)
         );
  DFF_X1 \REGISTERS_reg[18][7]  ( .D(n6857), .CK(CLK), .Q(n25736), .QN(n21692)
         );
  DFF_X1 \REGISTERS_reg[18][6]  ( .D(n6856), .CK(CLK), .Q(n25731), .QN(n21693)
         );
  DFF_X1 \REGISTERS_reg[18][5]  ( .D(n6855), .CK(CLK), .Q(n25726), .QN(n21694)
         );
  DFF_X1 \REGISTERS_reg[18][4]  ( .D(n6854), .CK(CLK), .Q(n25721), .QN(n21695)
         );
  DFF_X1 \REGISTERS_reg[18][3]  ( .D(n6853), .CK(CLK), .Q(n25716), .QN(n21696)
         );
  DFF_X1 \REGISTERS_reg[18][2]  ( .D(n6852), .CK(CLK), .Q(n25711), .QN(n21697)
         );
  DFF_X1 \REGISTERS_reg[18][1]  ( .D(n6851), .CK(CLK), .Q(n25706), .QN(n21698)
         );
  DFF_X1 \REGISTERS_reg[18][0]  ( .D(n6850), .CK(CLK), .Q(n25701), .QN(n21699)
         );
  DFF_X1 \REGISTERS_reg[10][59]  ( .D(n7421), .CK(CLK), .Q(n18450), .QN(n22380) );
  DFF_X1 \REGISTERS_reg[10][58]  ( .D(n7420), .CK(CLK), .Q(n18467), .QN(n22381) );
  DFF_X1 \REGISTERS_reg[10][57]  ( .D(n7419), .CK(CLK), .Q(n18484), .QN(n22382) );
  DFF_X1 \REGISTERS_reg[10][56]  ( .D(n7418), .CK(CLK), .Q(n18501), .QN(n22383) );
  DFF_X1 \REGISTERS_reg[10][55]  ( .D(n7417), .CK(CLK), .Q(n18518), .QN(n22384) );
  DFF_X1 \REGISTERS_reg[10][54]  ( .D(n7416), .CK(CLK), .Q(n18535), .QN(n22385) );
  DFF_X1 \REGISTERS_reg[10][53]  ( .D(n7415), .CK(CLK), .Q(n18552), .QN(n22386) );
  DFF_X1 \REGISTERS_reg[10][52]  ( .D(n7414), .CK(CLK), .Q(n18569), .QN(n22387) );
  DFF_X1 \REGISTERS_reg[10][51]  ( .D(n7413), .CK(CLK), .Q(n18586), .QN(n22388) );
  DFF_X1 \REGISTERS_reg[10][50]  ( .D(n7412), .CK(CLK), .Q(n18603), .QN(n22389) );
  DFF_X1 \REGISTERS_reg[10][49]  ( .D(n7411), .CK(CLK), .Q(n18620), .QN(n22390) );
  DFF_X1 \REGISTERS_reg[10][48]  ( .D(n7410), .CK(CLK), .Q(n18637), .QN(n22391) );
  DFF_X1 \REGISTERS_reg[10][47]  ( .D(n7409), .CK(CLK), .Q(n18654), .QN(n22392) );
  DFF_X1 \REGISTERS_reg[10][46]  ( .D(n7408), .CK(CLK), .Q(n18671), .QN(n22393) );
  DFF_X1 \REGISTERS_reg[10][45]  ( .D(n7407), .CK(CLK), .Q(n18688), .QN(n22394) );
  DFF_X1 \REGISTERS_reg[10][44]  ( .D(n7406), .CK(CLK), .Q(n18705), .QN(n22395) );
  DFF_X1 \REGISTERS_reg[10][43]  ( .D(n7405), .CK(CLK), .Q(n18722), .QN(n22396) );
  DFF_X1 \REGISTERS_reg[10][42]  ( .D(n7404), .CK(CLK), .Q(n18739), .QN(n22397) );
  DFF_X1 \REGISTERS_reg[10][41]  ( .D(n7403), .CK(CLK), .Q(n18756), .QN(n22398) );
  DFF_X1 \REGISTERS_reg[10][40]  ( .D(n7402), .CK(CLK), .Q(n18773), .QN(n22399) );
  DFF_X1 \REGISTERS_reg[10][39]  ( .D(n7401), .CK(CLK), .Q(n18790), .QN(n22400) );
  DFF_X1 \REGISTERS_reg[10][38]  ( .D(n7400), .CK(CLK), .Q(n18807), .QN(n22401) );
  DFF_X1 \REGISTERS_reg[10][37]  ( .D(n7399), .CK(CLK), .Q(n18824), .QN(n22402) );
  DFF_X1 \REGISTERS_reg[10][36]  ( .D(n7398), .CK(CLK), .Q(n18841), .QN(n22403) );
  DFF_X1 \REGISTERS_reg[10][35]  ( .D(n7397), .CK(CLK), .Q(n18858), .QN(n22404) );
  DFF_X1 \REGISTERS_reg[10][34]  ( .D(n7396), .CK(CLK), .Q(n18875), .QN(n22405) );
  DFF_X1 \REGISTERS_reg[10][33]  ( .D(n7395), .CK(CLK), .Q(n18892), .QN(n22406) );
  DFF_X1 \REGISTERS_reg[10][32]  ( .D(n7394), .CK(CLK), .Q(n18909), .QN(n22407) );
  DFF_X1 \REGISTERS_reg[10][31]  ( .D(n7393), .CK(CLK), .Q(n18926), .QN(n22408) );
  DFF_X1 \REGISTERS_reg[10][30]  ( .D(n7392), .CK(CLK), .Q(n18943), .QN(n22409) );
  DFF_X1 \REGISTERS_reg[10][29]  ( .D(n7391), .CK(CLK), .Q(n18960), .QN(n22410) );
  DFF_X1 \REGISTERS_reg[10][28]  ( .D(n7390), .CK(CLK), .Q(n18977), .QN(n22411) );
  DFF_X1 \REGISTERS_reg[10][27]  ( .D(n7389), .CK(CLK), .Q(n18994), .QN(n22412) );
  DFF_X1 \REGISTERS_reg[10][26]  ( .D(n7388), .CK(CLK), .Q(n19011), .QN(n22413) );
  DFF_X1 \REGISTERS_reg[10][25]  ( .D(n7387), .CK(CLK), .Q(n19028), .QN(n22414) );
  DFF_X1 \REGISTERS_reg[10][24]  ( .D(n7386), .CK(CLK), .Q(n19045), .QN(n22415) );
  DFF_X1 \REGISTERS_reg[10][23]  ( .D(n7385), .CK(CLK), .Q(n19062), .QN(n22416) );
  DFF_X1 \REGISTERS_reg[10][22]  ( .D(n7384), .CK(CLK), .Q(n19079), .QN(n22417) );
  DFF_X1 \REGISTERS_reg[10][21]  ( .D(n7383), .CK(CLK), .Q(n19096), .QN(n22418) );
  DFF_X1 \REGISTERS_reg[10][20]  ( .D(n7382), .CK(CLK), .Q(n19113), .QN(n22419) );
  DFF_X1 \REGISTERS_reg[10][19]  ( .D(n7381), .CK(CLK), .Q(n19130), .QN(n22420) );
  DFF_X1 \REGISTERS_reg[10][18]  ( .D(n7380), .CK(CLK), .Q(n19147), .QN(n22421) );
  DFF_X1 \REGISTERS_reg[10][17]  ( .D(n7379), .CK(CLK), .Q(n19164), .QN(n22422) );
  DFF_X1 \REGISTERS_reg[10][16]  ( .D(n7378), .CK(CLK), .Q(n19181), .QN(n22423) );
  DFF_X1 \REGISTERS_reg[10][15]  ( .D(n7377), .CK(CLK), .Q(n19198), .QN(n22424) );
  DFF_X1 \REGISTERS_reg[10][14]  ( .D(n7376), .CK(CLK), .Q(n19215), .QN(n22425) );
  DFF_X1 \REGISTERS_reg[10][13]  ( .D(n7375), .CK(CLK), .Q(n19232), .QN(n22426) );
  DFF_X1 \REGISTERS_reg[10][12]  ( .D(n7374), .CK(CLK), .Q(n19249), .QN(n22427) );
  DFF_X1 \REGISTERS_reg[10][11]  ( .D(n7373), .CK(CLK), .Q(n19266), .QN(n22428) );
  DFF_X1 \REGISTERS_reg[10][10]  ( .D(n7372), .CK(CLK), .Q(n19283), .QN(n22429) );
  DFF_X1 \REGISTERS_reg[10][9]  ( .D(n7371), .CK(CLK), .Q(n19300), .QN(n22430)
         );
  DFF_X1 \REGISTERS_reg[10][8]  ( .D(n7370), .CK(CLK), .Q(n19317), .QN(n22431)
         );
  DFF_X1 \REGISTERS_reg[10][7]  ( .D(n7369), .CK(CLK), .Q(n19334), .QN(n22432)
         );
  DFF_X1 \REGISTERS_reg[10][6]  ( .D(n7368), .CK(CLK), .Q(n19351), .QN(n22433)
         );
  DFF_X1 \REGISTERS_reg[10][5]  ( .D(n7367), .CK(CLK), .Q(n19368), .QN(n22434)
         );
  DFF_X1 \REGISTERS_reg[10][4]  ( .D(n7366), .CK(CLK), .Q(n19385), .QN(n22435)
         );
  DFF_X1 \REGISTERS_reg[10][3]  ( .D(n7365), .CK(CLK), .Q(n19402), .QN(n22436)
         );
  DFF_X1 \REGISTERS_reg[10][2]  ( .D(n7364), .CK(CLK), .Q(n19419), .QN(n22437)
         );
  DFF_X1 \REGISTERS_reg[10][1]  ( .D(n7363), .CK(CLK), .Q(n19436), .QN(n22438)
         );
  DFF_X1 \REGISTERS_reg[10][0]  ( .D(n7362), .CK(CLK), .Q(n19453), .QN(n22439)
         );
  DFF_X1 \REGISTERS_reg[1][59]  ( .D(n7997), .CK(CLK), .Q(n25502), .QN(n22060)
         );
  DFF_X1 \REGISTERS_reg[1][58]  ( .D(n7996), .CK(CLK), .Q(n25501), .QN(n22061)
         );
  DFF_X1 \REGISTERS_reg[1][57]  ( .D(n7995), .CK(CLK), .Q(n25500), .QN(n22062)
         );
  DFF_X1 \REGISTERS_reg[1][56]  ( .D(n7994), .CK(CLK), .Q(n25499), .QN(n22063)
         );
  DFF_X1 \REGISTERS_reg[1][55]  ( .D(n7993), .CK(CLK), .Q(n25498), .QN(n22064)
         );
  DFF_X1 \REGISTERS_reg[1][54]  ( .D(n7992), .CK(CLK), .Q(n25497), .QN(n22065)
         );
  DFF_X1 \REGISTERS_reg[1][53]  ( .D(n7991), .CK(CLK), .Q(n25496), .QN(n22066)
         );
  DFF_X1 \REGISTERS_reg[1][52]  ( .D(n7990), .CK(CLK), .Q(n25495), .QN(n22067)
         );
  DFF_X1 \REGISTERS_reg[1][51]  ( .D(n7989), .CK(CLK), .Q(n25494), .QN(n22068)
         );
  DFF_X1 \REGISTERS_reg[1][50]  ( .D(n7988), .CK(CLK), .Q(n25493), .QN(n22069)
         );
  DFF_X1 \REGISTERS_reg[1][49]  ( .D(n7987), .CK(CLK), .Q(n25492), .QN(n22070)
         );
  DFF_X1 \REGISTERS_reg[1][48]  ( .D(n7986), .CK(CLK), .Q(n25491), .QN(n22071)
         );
  DFF_X1 \REGISTERS_reg[1][47]  ( .D(n7985), .CK(CLK), .Q(n25490), .QN(n22072)
         );
  DFF_X1 \REGISTERS_reg[1][46]  ( .D(n7984), .CK(CLK), .Q(n25489), .QN(n22073)
         );
  DFF_X1 \REGISTERS_reg[1][45]  ( .D(n7983), .CK(CLK), .Q(n25488), .QN(n22074)
         );
  DFF_X1 \REGISTERS_reg[1][44]  ( .D(n7982), .CK(CLK), .Q(n25487), .QN(n22075)
         );
  DFF_X1 \REGISTERS_reg[1][43]  ( .D(n7981), .CK(CLK), .Q(n25486), .QN(n22076)
         );
  DFF_X1 \REGISTERS_reg[1][42]  ( .D(n7980), .CK(CLK), .Q(n25485), .QN(n22077)
         );
  DFF_X1 \REGISTERS_reg[1][41]  ( .D(n7979), .CK(CLK), .Q(n25484), .QN(n22078)
         );
  DFF_X1 \REGISTERS_reg[1][40]  ( .D(n7978), .CK(CLK), .Q(n25483), .QN(n22079)
         );
  DFF_X1 \REGISTERS_reg[1][39]  ( .D(n7977), .CK(CLK), .Q(n25482), .QN(n22080)
         );
  DFF_X1 \REGISTERS_reg[1][38]  ( .D(n7976), .CK(CLK), .Q(n25481), .QN(n22081)
         );
  DFF_X1 \REGISTERS_reg[1][37]  ( .D(n7975), .CK(CLK), .Q(n25480), .QN(n22082)
         );
  DFF_X1 \REGISTERS_reg[1][36]  ( .D(n7974), .CK(CLK), .Q(n25479), .QN(n22083)
         );
  DFF_X1 \REGISTERS_reg[1][35]  ( .D(n7973), .CK(CLK), .Q(n25478), .QN(n22084)
         );
  DFF_X1 \REGISTERS_reg[1][34]  ( .D(n7972), .CK(CLK), .Q(n25477), .QN(n22085)
         );
  DFF_X1 \REGISTERS_reg[1][33]  ( .D(n7971), .CK(CLK), .Q(n25476), .QN(n22086)
         );
  DFF_X1 \REGISTERS_reg[1][32]  ( .D(n7970), .CK(CLK), .Q(n25475), .QN(n22087)
         );
  DFF_X1 \REGISTERS_reg[1][31]  ( .D(n7969), .CK(CLK), .Q(n25474), .QN(n22088)
         );
  DFF_X1 \REGISTERS_reg[1][30]  ( .D(n7968), .CK(CLK), .Q(n25473), .QN(n22089)
         );
  DFF_X1 \REGISTERS_reg[1][29]  ( .D(n7967), .CK(CLK), .Q(n25472), .QN(n22090)
         );
  DFF_X1 \REGISTERS_reg[1][28]  ( .D(n7966), .CK(CLK), .Q(n25471), .QN(n22091)
         );
  DFF_X1 \REGISTERS_reg[1][27]  ( .D(n7965), .CK(CLK), .Q(n25470), .QN(n22092)
         );
  DFF_X1 \REGISTERS_reg[1][26]  ( .D(n7964), .CK(CLK), .Q(n25469), .QN(n22093)
         );
  DFF_X1 \REGISTERS_reg[1][25]  ( .D(n7963), .CK(CLK), .Q(n25468), .QN(n22094)
         );
  DFF_X1 \REGISTERS_reg[1][24]  ( .D(n7962), .CK(CLK), .Q(n25467), .QN(n22095)
         );
  DFF_X1 \REGISTERS_reg[1][23]  ( .D(n7961), .CK(CLK), .Q(n25466), .QN(n22096)
         );
  DFF_X1 \REGISTERS_reg[1][22]  ( .D(n7960), .CK(CLK), .Q(n25465), .QN(n22097)
         );
  DFF_X1 \REGISTERS_reg[1][21]  ( .D(n7959), .CK(CLK), .Q(n25464), .QN(n22098)
         );
  DFF_X1 \REGISTERS_reg[1][20]  ( .D(n7958), .CK(CLK), .Q(n25463), .QN(n22099)
         );
  DFF_X1 \REGISTERS_reg[1][19]  ( .D(n7957), .CK(CLK), .Q(n25462), .QN(n22100)
         );
  DFF_X1 \REGISTERS_reg[1][18]  ( .D(n7956), .CK(CLK), .Q(n25461), .QN(n22101)
         );
  DFF_X1 \REGISTERS_reg[1][17]  ( .D(n7955), .CK(CLK), .Q(n25460), .QN(n22102)
         );
  DFF_X1 \REGISTERS_reg[1][16]  ( .D(n7954), .CK(CLK), .Q(n25459), .QN(n22103)
         );
  DFF_X1 \REGISTERS_reg[1][15]  ( .D(n7953), .CK(CLK), .Q(n25458), .QN(n22104)
         );
  DFF_X1 \REGISTERS_reg[1][14]  ( .D(n7952), .CK(CLK), .Q(n25457), .QN(n22105)
         );
  DFF_X1 \REGISTERS_reg[1][13]  ( .D(n7951), .CK(CLK), .Q(n25456), .QN(n22106)
         );
  DFF_X1 \REGISTERS_reg[1][12]  ( .D(n7950), .CK(CLK), .Q(n25455), .QN(n22107)
         );
  DFF_X1 \REGISTERS_reg[1][11]  ( .D(n7949), .CK(CLK), .Q(n25666), .QN(n22108)
         );
  DFF_X1 \REGISTERS_reg[1][10]  ( .D(n7948), .CK(CLK), .Q(n25665), .QN(n22109)
         );
  DFF_X1 \REGISTERS_reg[1][9]  ( .D(n7947), .CK(CLK), .Q(n25664), .QN(n22110)
         );
  DFF_X1 \REGISTERS_reg[1][8]  ( .D(n7946), .CK(CLK), .Q(n25663), .QN(n22111)
         );
  DFF_X1 \REGISTERS_reg[1][7]  ( .D(n7945), .CK(CLK), .Q(n25662), .QN(n22112)
         );
  DFF_X1 \REGISTERS_reg[1][6]  ( .D(n7944), .CK(CLK), .Q(n25661), .QN(n22113)
         );
  DFF_X1 \REGISTERS_reg[1][5]  ( .D(n7943), .CK(CLK), .Q(n25660), .QN(n22114)
         );
  DFF_X1 \REGISTERS_reg[1][4]  ( .D(n7942), .CK(CLK), .Q(n25659), .QN(n22115)
         );
  DFF_X1 \REGISTERS_reg[1][3]  ( .D(n7941), .CK(CLK), .Q(n25658), .QN(n22116)
         );
  DFF_X1 \REGISTERS_reg[1][2]  ( .D(n7940), .CK(CLK), .Q(n25657), .QN(n22117)
         );
  DFF_X1 \REGISTERS_reg[1][1]  ( .D(n7939), .CK(CLK), .Q(n25656), .QN(n22118)
         );
  DFF_X1 \REGISTERS_reg[1][0]  ( .D(n7938), .CK(CLK), .Q(n25655), .QN(n22119)
         );
  DFF_X1 \REGISTERS_reg[16][59]  ( .D(n7037), .CK(CLK), .Q(n25997), .QN(n21240) );
  DFF_X1 \REGISTERS_reg[16][58]  ( .D(n7036), .CK(CLK), .Q(n25992), .QN(n21241) );
  DFF_X1 \REGISTERS_reg[16][57]  ( .D(n7035), .CK(CLK), .Q(n25987), .QN(n21242) );
  DFF_X1 \REGISTERS_reg[16][56]  ( .D(n7034), .CK(CLK), .Q(n25982), .QN(n21243) );
  DFF_X1 \REGISTERS_reg[16][55]  ( .D(n7033), .CK(CLK), .Q(n25977), .QN(n21244) );
  DFF_X1 \REGISTERS_reg[16][54]  ( .D(n7032), .CK(CLK), .Q(n25972), .QN(n21245) );
  DFF_X1 \REGISTERS_reg[16][53]  ( .D(n7031), .CK(CLK), .Q(n25967), .QN(n21246) );
  DFF_X1 \REGISTERS_reg[16][52]  ( .D(n7030), .CK(CLK), .Q(n25962), .QN(n21247) );
  DFF_X1 \REGISTERS_reg[16][51]  ( .D(n7029), .CK(CLK), .Q(n25957), .QN(n21248) );
  DFF_X1 \REGISTERS_reg[16][50]  ( .D(n7028), .CK(CLK), .Q(n25952), .QN(n21249) );
  DFF_X1 \REGISTERS_reg[16][49]  ( .D(n7027), .CK(CLK), .Q(n25947), .QN(n21250) );
  DFF_X1 \REGISTERS_reg[16][48]  ( .D(n7026), .CK(CLK), .Q(n25942), .QN(n21251) );
  DFF_X1 \REGISTERS_reg[16][47]  ( .D(n7025), .CK(CLK), .Q(n25937), .QN(n21252) );
  DFF_X1 \REGISTERS_reg[16][46]  ( .D(n7024), .CK(CLK), .Q(n25932), .QN(n21253) );
  DFF_X1 \REGISTERS_reg[16][45]  ( .D(n7023), .CK(CLK), .Q(n25927), .QN(n21254) );
  DFF_X1 \REGISTERS_reg[16][44]  ( .D(n7022), .CK(CLK), .Q(n25922), .QN(n21255) );
  DFF_X1 \REGISTERS_reg[16][43]  ( .D(n7021), .CK(CLK), .Q(n25917), .QN(n21256) );
  DFF_X1 \REGISTERS_reg[16][42]  ( .D(n7020), .CK(CLK), .Q(n25912), .QN(n21257) );
  DFF_X1 \REGISTERS_reg[16][41]  ( .D(n7019), .CK(CLK), .Q(n25907), .QN(n21258) );
  DFF_X1 \REGISTERS_reg[16][40]  ( .D(n7018), .CK(CLK), .Q(n25902), .QN(n21259) );
  DFF_X1 \REGISTERS_reg[16][39]  ( .D(n7017), .CK(CLK), .Q(n25897), .QN(n21260) );
  DFF_X1 \REGISTERS_reg[16][38]  ( .D(n7016), .CK(CLK), .Q(n25892), .QN(n21261) );
  DFF_X1 \REGISTERS_reg[16][37]  ( .D(n7015), .CK(CLK), .Q(n25887), .QN(n21262) );
  DFF_X1 \REGISTERS_reg[16][36]  ( .D(n7014), .CK(CLK), .Q(n25882), .QN(n21263) );
  DFF_X1 \REGISTERS_reg[16][35]  ( .D(n7013), .CK(CLK), .Q(n25877), .QN(n21264) );
  DFF_X1 \REGISTERS_reg[16][34]  ( .D(n7012), .CK(CLK), .Q(n25872), .QN(n21265) );
  DFF_X1 \REGISTERS_reg[16][33]  ( .D(n7011), .CK(CLK), .Q(n25867), .QN(n21266) );
  DFF_X1 \REGISTERS_reg[16][32]  ( .D(n7010), .CK(CLK), .Q(n25862), .QN(n21267) );
  DFF_X1 \REGISTERS_reg[16][31]  ( .D(n7009), .CK(CLK), .Q(n25857), .QN(n21268) );
  DFF_X1 \REGISTERS_reg[16][30]  ( .D(n7008), .CK(CLK), .Q(n25852), .QN(n21269) );
  DFF_X1 \REGISTERS_reg[16][29]  ( .D(n7007), .CK(CLK), .Q(n25847), .QN(n21270) );
  DFF_X1 \REGISTERS_reg[16][28]  ( .D(n7006), .CK(CLK), .Q(n25842), .QN(n21271) );
  DFF_X1 \REGISTERS_reg[16][27]  ( .D(n7005), .CK(CLK), .Q(n25837), .QN(n21272) );
  DFF_X1 \REGISTERS_reg[16][26]  ( .D(n7004), .CK(CLK), .Q(n25832), .QN(n21273) );
  DFF_X1 \REGISTERS_reg[16][25]  ( .D(n7003), .CK(CLK), .Q(n25827), .QN(n21274) );
  DFF_X1 \REGISTERS_reg[16][24]  ( .D(n7002), .CK(CLK), .Q(n25822), .QN(n21275) );
  DFF_X1 \REGISTERS_reg[16][23]  ( .D(n7001), .CK(CLK), .Q(n25817), .QN(n21276) );
  DFF_X1 \REGISTERS_reg[16][22]  ( .D(n7000), .CK(CLK), .Q(n25812), .QN(n21277) );
  DFF_X1 \REGISTERS_reg[16][21]  ( .D(n6999), .CK(CLK), .Q(n25807), .QN(n21278) );
  DFF_X1 \REGISTERS_reg[16][20]  ( .D(n6998), .CK(CLK), .Q(n25802), .QN(n21279) );
  DFF_X1 \REGISTERS_reg[16][19]  ( .D(n6997), .CK(CLK), .Q(n25797), .QN(n21280) );
  DFF_X1 \REGISTERS_reg[16][18]  ( .D(n6996), .CK(CLK), .Q(n25792), .QN(n21281) );
  DFF_X1 \REGISTERS_reg[16][17]  ( .D(n6995), .CK(CLK), .Q(n25787), .QN(n21282) );
  DFF_X1 \REGISTERS_reg[16][16]  ( .D(n6994), .CK(CLK), .Q(n25782), .QN(n21283) );
  DFF_X1 \REGISTERS_reg[16][15]  ( .D(n6993), .CK(CLK), .Q(n25777), .QN(n21284) );
  DFF_X1 \REGISTERS_reg[16][14]  ( .D(n6992), .CK(CLK), .Q(n25772), .QN(n21285) );
  DFF_X1 \REGISTERS_reg[16][13]  ( .D(n6991), .CK(CLK), .Q(n25767), .QN(n21286) );
  DFF_X1 \REGISTERS_reg[16][12]  ( .D(n6990), .CK(CLK), .Q(n25762), .QN(n21287) );
  DFF_X1 \REGISTERS_reg[16][11]  ( .D(n6989), .CK(CLK), .Q(n25757), .QN(n21288) );
  DFF_X1 \REGISTERS_reg[16][10]  ( .D(n6988), .CK(CLK), .Q(n25752), .QN(n21289) );
  DFF_X1 \REGISTERS_reg[16][9]  ( .D(n6987), .CK(CLK), .Q(n25747), .QN(n21290)
         );
  DFF_X1 \REGISTERS_reg[16][8]  ( .D(n6986), .CK(CLK), .Q(n25742), .QN(n21291)
         );
  DFF_X1 \REGISTERS_reg[16][7]  ( .D(n6985), .CK(CLK), .Q(n25737), .QN(n21292)
         );
  DFF_X1 \REGISTERS_reg[16][6]  ( .D(n6984), .CK(CLK), .Q(n25732), .QN(n21293)
         );
  DFF_X1 \REGISTERS_reg[16][5]  ( .D(n6983), .CK(CLK), .Q(n25727), .QN(n21294)
         );
  DFF_X1 \REGISTERS_reg[16][4]  ( .D(n6982), .CK(CLK), .Q(n25722), .QN(n21295)
         );
  DFF_X1 \REGISTERS_reg[16][3]  ( .D(n6981), .CK(CLK), .Q(n25717), .QN(n21296)
         );
  DFF_X1 \REGISTERS_reg[16][2]  ( .D(n6980), .CK(CLK), .Q(n25712), .QN(n21297)
         );
  DFF_X1 \REGISTERS_reg[16][1]  ( .D(n6979), .CK(CLK), .Q(n25707), .QN(n21298)
         );
  DFF_X1 \REGISTERS_reg[16][0]  ( .D(n6978), .CK(CLK), .Q(n25702), .QN(n21299)
         );
  DFF_X1 \REGISTERS_reg[6][59]  ( .D(n7677), .CK(CLK), .Q(n25262), .QN(n21820)
         );
  DFF_X1 \REGISTERS_reg[6][58]  ( .D(n7676), .CK(CLK), .Q(n25261), .QN(n21821)
         );
  DFF_X1 \REGISTERS_reg[6][57]  ( .D(n7675), .CK(CLK), .Q(n25260), .QN(n21822)
         );
  DFF_X1 \REGISTERS_reg[6][56]  ( .D(n7674), .CK(CLK), .Q(n25259), .QN(n21823)
         );
  DFF_X1 \REGISTERS_reg[6][55]  ( .D(n7673), .CK(CLK), .Q(n25258), .QN(n21824)
         );
  DFF_X1 \REGISTERS_reg[6][54]  ( .D(n7672), .CK(CLK), .Q(n25257), .QN(n21825)
         );
  DFF_X1 \REGISTERS_reg[6][53]  ( .D(n7671), .CK(CLK), .Q(n25256), .QN(n21826)
         );
  DFF_X1 \REGISTERS_reg[6][52]  ( .D(n7670), .CK(CLK), .Q(n25255), .QN(n21827)
         );
  DFF_X1 \REGISTERS_reg[6][51]  ( .D(n7669), .CK(CLK), .Q(n25254), .QN(n21828)
         );
  DFF_X1 \REGISTERS_reg[6][50]  ( .D(n7668), .CK(CLK), .Q(n25253), .QN(n21829)
         );
  DFF_X1 \REGISTERS_reg[6][49]  ( .D(n7667), .CK(CLK), .Q(n25252), .QN(n21830)
         );
  DFF_X1 \REGISTERS_reg[6][48]  ( .D(n7666), .CK(CLK), .Q(n25251), .QN(n21831)
         );
  DFF_X1 \REGISTERS_reg[6][47]  ( .D(n7665), .CK(CLK), .Q(n25250), .QN(n21832)
         );
  DFF_X1 \REGISTERS_reg[6][46]  ( .D(n7664), .CK(CLK), .Q(n25249), .QN(n21833)
         );
  DFF_X1 \REGISTERS_reg[6][45]  ( .D(n7663), .CK(CLK), .Q(n25248), .QN(n21834)
         );
  DFF_X1 \REGISTERS_reg[6][44]  ( .D(n7662), .CK(CLK), .Q(n25247), .QN(n21835)
         );
  DFF_X1 \REGISTERS_reg[6][43]  ( .D(n7661), .CK(CLK), .Q(n25246), .QN(n21836)
         );
  DFF_X1 \REGISTERS_reg[6][42]  ( .D(n7660), .CK(CLK), .Q(n25245), .QN(n21837)
         );
  DFF_X1 \REGISTERS_reg[6][41]  ( .D(n7659), .CK(CLK), .Q(n25244), .QN(n21838)
         );
  DFF_X1 \REGISTERS_reg[6][40]  ( .D(n7658), .CK(CLK), .Q(n25243), .QN(n21839)
         );
  DFF_X1 \REGISTERS_reg[6][39]  ( .D(n7657), .CK(CLK), .Q(n25242), .QN(n21840)
         );
  DFF_X1 \REGISTERS_reg[6][38]  ( .D(n7656), .CK(CLK), .Q(n25241), .QN(n21841)
         );
  DFF_X1 \REGISTERS_reg[6][37]  ( .D(n7655), .CK(CLK), .Q(n25240), .QN(n21842)
         );
  DFF_X1 \REGISTERS_reg[6][36]  ( .D(n7654), .CK(CLK), .Q(n25239), .QN(n21843)
         );
  DFF_X1 \REGISTERS_reg[6][35]  ( .D(n7653), .CK(CLK), .Q(n25238), .QN(n21844)
         );
  DFF_X1 \REGISTERS_reg[6][34]  ( .D(n7652), .CK(CLK), .Q(n25237), .QN(n21845)
         );
  DFF_X1 \REGISTERS_reg[6][33]  ( .D(n7651), .CK(CLK), .Q(n25236), .QN(n21846)
         );
  DFF_X1 \REGISTERS_reg[6][32]  ( .D(n7650), .CK(CLK), .Q(n25235), .QN(n21847)
         );
  DFF_X1 \REGISTERS_reg[6][31]  ( .D(n7649), .CK(CLK), .Q(n25234), .QN(n21848)
         );
  DFF_X1 \REGISTERS_reg[6][30]  ( .D(n7648), .CK(CLK), .Q(n25233), .QN(n21849)
         );
  DFF_X1 \REGISTERS_reg[6][29]  ( .D(n7647), .CK(CLK), .Q(n25232), .QN(n21850)
         );
  DFF_X1 \REGISTERS_reg[6][28]  ( .D(n7646), .CK(CLK), .Q(n25231), .QN(n21851)
         );
  DFF_X1 \REGISTERS_reg[6][27]  ( .D(n7645), .CK(CLK), .Q(n25230), .QN(n21852)
         );
  DFF_X1 \REGISTERS_reg[6][26]  ( .D(n7644), .CK(CLK), .Q(n25229), .QN(n21853)
         );
  DFF_X1 \REGISTERS_reg[6][25]  ( .D(n7643), .CK(CLK), .Q(n25228), .QN(n21854)
         );
  DFF_X1 \REGISTERS_reg[6][24]  ( .D(n7642), .CK(CLK), .Q(n25227), .QN(n21855)
         );
  DFF_X1 \REGISTERS_reg[6][23]  ( .D(n7641), .CK(CLK), .Q(n25226), .QN(n21856)
         );
  DFF_X1 \REGISTERS_reg[6][22]  ( .D(n7640), .CK(CLK), .Q(n25225), .QN(n21857)
         );
  DFF_X1 \REGISTERS_reg[6][21]  ( .D(n7639), .CK(CLK), .Q(n25224), .QN(n21858)
         );
  DFF_X1 \REGISTERS_reg[6][20]  ( .D(n7638), .CK(CLK), .Q(n25223), .QN(n21859)
         );
  DFF_X1 \REGISTERS_reg[6][19]  ( .D(n7637), .CK(CLK), .Q(n25222), .QN(n21860)
         );
  DFF_X1 \REGISTERS_reg[6][18]  ( .D(n7636), .CK(CLK), .Q(n25221), .QN(n21861)
         );
  DFF_X1 \REGISTERS_reg[6][17]  ( .D(n7635), .CK(CLK), .Q(n25220), .QN(n21862)
         );
  DFF_X1 \REGISTERS_reg[6][16]  ( .D(n7634), .CK(CLK), .Q(n25219), .QN(n21863)
         );
  DFF_X1 \REGISTERS_reg[6][15]  ( .D(n7633), .CK(CLK), .Q(n25218), .QN(n21864)
         );
  DFF_X1 \REGISTERS_reg[6][14]  ( .D(n7632), .CK(CLK), .Q(n25217), .QN(n21865)
         );
  DFF_X1 \REGISTERS_reg[6][13]  ( .D(n7631), .CK(CLK), .Q(n25216), .QN(n21866)
         );
  DFF_X1 \REGISTERS_reg[6][12]  ( .D(n7630), .CK(CLK), .Q(n25215), .QN(n21867)
         );
  DFF_X1 \REGISTERS_reg[6][11]  ( .D(n7629), .CK(CLK), .Q(n25606), .QN(n21868)
         );
  DFF_X1 \REGISTERS_reg[6][10]  ( .D(n7628), .CK(CLK), .Q(n25605), .QN(n21869)
         );
  DFF_X1 \REGISTERS_reg[6][9]  ( .D(n7627), .CK(CLK), .Q(n25604), .QN(n21870)
         );
  DFF_X1 \REGISTERS_reg[6][8]  ( .D(n7626), .CK(CLK), .Q(n25603), .QN(n21871)
         );
  DFF_X1 \REGISTERS_reg[6][7]  ( .D(n7625), .CK(CLK), .Q(n25602), .QN(n21872)
         );
  DFF_X1 \REGISTERS_reg[6][6]  ( .D(n7624), .CK(CLK), .Q(n25601), .QN(n21873)
         );
  DFF_X1 \REGISTERS_reg[6][5]  ( .D(n7623), .CK(CLK), .Q(n25600), .QN(n21874)
         );
  DFF_X1 \REGISTERS_reg[6][4]  ( .D(n7622), .CK(CLK), .Q(n25599), .QN(n21875)
         );
  DFF_X1 \REGISTERS_reg[6][3]  ( .D(n7621), .CK(CLK), .Q(n25598), .QN(n21876)
         );
  DFF_X1 \REGISTERS_reg[6][2]  ( .D(n7620), .CK(CLK), .Q(n25597), .QN(n21877)
         );
  DFF_X1 \REGISTERS_reg[6][1]  ( .D(n7619), .CK(CLK), .Q(n25596), .QN(n21878)
         );
  DFF_X1 \REGISTERS_reg[6][0]  ( .D(n7618), .CK(CLK), .Q(n25595), .QN(n21879)
         );
  DFF_X1 \OUT2_reg[63]  ( .D(n5889), .CK(CLK), .Q(n4226) );
  INV_X1 U19266 ( .A(n26537), .ZN(n26533) );
  INV_X1 U19267 ( .A(n26762), .ZN(n26758) );
  INV_X1 U19268 ( .A(n26541), .ZN(n26535) );
  INV_X1 U19269 ( .A(n26540), .ZN(n26534) );
  INV_X1 U19270 ( .A(n26765), .ZN(n26760) );
  INV_X1 U19271 ( .A(n26763), .ZN(n26759) );
  BUF_X1 U19272 ( .A(n22722), .Z(n27162) );
  BUF_X1 U19273 ( .A(n22722), .Z(n27163) );
  BUF_X1 U19274 ( .A(n22722), .Z(n27164) );
  BUF_X1 U19275 ( .A(n22722), .Z(n27165) );
  BUF_X1 U19276 ( .A(n22760), .Z(n26946) );
  BUF_X1 U19277 ( .A(n22760), .Z(n26947) );
  BUF_X1 U19278 ( .A(n22760), .Z(n26948) );
  BUF_X1 U19279 ( .A(n22760), .Z(n26949) );
  BUF_X1 U19280 ( .A(n22753), .Z(n26982) );
  BUF_X1 U19281 ( .A(n22753), .Z(n26983) );
  BUF_X1 U19282 ( .A(n22753), .Z(n26984) );
  BUF_X1 U19283 ( .A(n22753), .Z(n26985) );
  BUF_X1 U19284 ( .A(n22719), .Z(n27174) );
  BUF_X1 U19285 ( .A(n22719), .Z(n27175) );
  BUF_X1 U19286 ( .A(n22719), .Z(n27176) );
  BUF_X1 U19287 ( .A(n22719), .Z(n27177) );
  BUF_X1 U19288 ( .A(n22724), .Z(n27150) );
  BUF_X1 U19289 ( .A(n22724), .Z(n27151) );
  BUF_X1 U19290 ( .A(n22724), .Z(n27152) );
  BUF_X1 U19291 ( .A(n22724), .Z(n27153) );
  BUF_X1 U19292 ( .A(n22743), .Z(n27042) );
  BUF_X1 U19293 ( .A(n22743), .Z(n27043) );
  BUF_X1 U19294 ( .A(n22743), .Z(n27044) );
  BUF_X1 U19295 ( .A(n22743), .Z(n27045) );
  BUF_X1 U19296 ( .A(n22764), .Z(n26922) );
  BUF_X1 U19297 ( .A(n22764), .Z(n26923) );
  BUF_X1 U19298 ( .A(n22764), .Z(n26924) );
  BUF_X1 U19299 ( .A(n22764), .Z(n26925) );
  BUF_X1 U19300 ( .A(n22762), .Z(n26934) );
  BUF_X1 U19301 ( .A(n22762), .Z(n26935) );
  BUF_X1 U19302 ( .A(n22762), .Z(n26936) );
  BUF_X1 U19303 ( .A(n22762), .Z(n26937) );
  BUF_X1 U19304 ( .A(n22693), .Z(n27270) );
  BUF_X1 U19305 ( .A(n22693), .Z(n27271) );
  BUF_X1 U19306 ( .A(n22693), .Z(n27272) );
  BUF_X1 U19307 ( .A(n22693), .Z(n27273) );
  BUF_X1 U19308 ( .A(n22697), .Z(n27258) );
  BUF_X1 U19309 ( .A(n22697), .Z(n27259) );
  BUF_X1 U19310 ( .A(n22697), .Z(n27260) );
  BUF_X1 U19311 ( .A(n22697), .Z(n27261) );
  BUF_X1 U19312 ( .A(n22715), .Z(n27186) );
  BUF_X1 U19313 ( .A(n22715), .Z(n27187) );
  BUF_X1 U19314 ( .A(n22715), .Z(n27188) );
  BUF_X1 U19315 ( .A(n22715), .Z(n27189) );
  BUF_X1 U19316 ( .A(n22726), .Z(n27138) );
  BUF_X1 U19317 ( .A(n22726), .Z(n27139) );
  BUF_X1 U19318 ( .A(n22726), .Z(n27140) );
  BUF_X1 U19319 ( .A(n22726), .Z(n27141) );
  BUF_X1 U19320 ( .A(n22706), .Z(n27222) );
  BUF_X1 U19321 ( .A(n22706), .Z(n27223) );
  BUF_X1 U19322 ( .A(n22706), .Z(n27224) );
  BUF_X1 U19323 ( .A(n22706), .Z(n27225) );
  BUF_X1 U19324 ( .A(n22712), .Z(n27198) );
  BUF_X1 U19325 ( .A(n22712), .Z(n27199) );
  BUF_X1 U19326 ( .A(n22712), .Z(n27200) );
  BUF_X1 U19327 ( .A(n22712), .Z(n27201) );
  BUF_X1 U19328 ( .A(n22749), .Z(n27006) );
  BUF_X1 U19329 ( .A(n22749), .Z(n27007) );
  BUF_X1 U19330 ( .A(n22749), .Z(n27008) );
  BUF_X1 U19331 ( .A(n22749), .Z(n27009) );
  BUF_X1 U19332 ( .A(n22739), .Z(n27066) );
  BUF_X1 U19333 ( .A(n22739), .Z(n27067) );
  BUF_X1 U19334 ( .A(n22739), .Z(n27068) );
  BUF_X1 U19335 ( .A(n22739), .Z(n27069) );
  BUF_X1 U19336 ( .A(n22741), .Z(n27054) );
  BUF_X1 U19337 ( .A(n22741), .Z(n27055) );
  BUF_X1 U19338 ( .A(n22741), .Z(n27056) );
  BUF_X1 U19339 ( .A(n22741), .Z(n27057) );
  BUF_X1 U19340 ( .A(n22758), .Z(n26958) );
  BUF_X1 U19341 ( .A(n22758), .Z(n26959) );
  BUF_X1 U19342 ( .A(n22758), .Z(n26960) );
  BUF_X1 U19343 ( .A(n22758), .Z(n26961) );
  BUF_X1 U19344 ( .A(n22709), .Z(n27210) );
  BUF_X1 U19345 ( .A(n22709), .Z(n27211) );
  BUF_X1 U19346 ( .A(n22709), .Z(n27212) );
  BUF_X1 U19347 ( .A(n22709), .Z(n27213) );
  BUF_X1 U19348 ( .A(n22700), .Z(n27246) );
  BUF_X1 U19349 ( .A(n22700), .Z(n27247) );
  BUF_X1 U19350 ( .A(n22700), .Z(n27248) );
  BUF_X1 U19351 ( .A(n22700), .Z(n27249) );
  BUF_X1 U19352 ( .A(n22703), .Z(n27234) );
  BUF_X1 U19353 ( .A(n22703), .Z(n27235) );
  BUF_X1 U19354 ( .A(n22703), .Z(n27236) );
  BUF_X1 U19355 ( .A(n22703), .Z(n27237) );
  BUF_X1 U19356 ( .A(n22751), .Z(n26994) );
  BUF_X1 U19357 ( .A(n22751), .Z(n26995) );
  BUF_X1 U19358 ( .A(n22751), .Z(n26996) );
  BUF_X1 U19359 ( .A(n22751), .Z(n26997) );
  BUF_X1 U19360 ( .A(n22736), .Z(n27078) );
  BUF_X1 U19361 ( .A(n22736), .Z(n27079) );
  BUF_X1 U19362 ( .A(n22736), .Z(n27080) );
  BUF_X1 U19363 ( .A(n22736), .Z(n27081) );
  BUF_X1 U19364 ( .A(n22756), .Z(n26970) );
  BUF_X1 U19365 ( .A(n22756), .Z(n26971) );
  BUF_X1 U19366 ( .A(n22756), .Z(n26972) );
  BUF_X1 U19367 ( .A(n22756), .Z(n26973) );
  BUF_X1 U19368 ( .A(n22768), .Z(n26898) );
  BUF_X1 U19369 ( .A(n22768), .Z(n26899) );
  BUF_X1 U19370 ( .A(n22768), .Z(n26900) );
  BUF_X1 U19371 ( .A(n22768), .Z(n26901) );
  BUF_X1 U19372 ( .A(n22766), .Z(n26910) );
  BUF_X1 U19373 ( .A(n22766), .Z(n26911) );
  BUF_X1 U19374 ( .A(n22766), .Z(n26912) );
  BUF_X1 U19375 ( .A(n22766), .Z(n26913) );
  BUF_X1 U19376 ( .A(n22732), .Z(n27102) );
  BUF_X1 U19377 ( .A(n22732), .Z(n27103) );
  BUF_X1 U19378 ( .A(n22732), .Z(n27104) );
  BUF_X1 U19379 ( .A(n22732), .Z(n27105) );
  BUF_X1 U19380 ( .A(n22728), .Z(n27126) );
  BUF_X1 U19381 ( .A(n22728), .Z(n27127) );
  BUF_X1 U19382 ( .A(n22728), .Z(n27128) );
  BUF_X1 U19383 ( .A(n22728), .Z(n27129) );
  BUF_X1 U19384 ( .A(n27275), .Z(n27277) );
  BUF_X1 U19385 ( .A(n27275), .Z(n27278) );
  BUF_X1 U19386 ( .A(n27275), .Z(n27279) );
  BUF_X1 U19387 ( .A(n27276), .Z(n27280) );
  BUF_X1 U19388 ( .A(n27276), .Z(n27281) );
  BUF_X1 U19389 ( .A(n22730), .Z(n27113) );
  BUF_X1 U19390 ( .A(n22730), .Z(n27114) );
  BUF_X1 U19391 ( .A(n22730), .Z(n27115) );
  BUF_X1 U19392 ( .A(n22730), .Z(n27116) );
  BUF_X1 U19393 ( .A(n22730), .Z(n27117) );
  BUF_X1 U19394 ( .A(n22734), .Z(n27089) );
  BUF_X1 U19395 ( .A(n22734), .Z(n27090) );
  BUF_X1 U19396 ( .A(n22734), .Z(n27091) );
  BUF_X1 U19397 ( .A(n22734), .Z(n27092) );
  BUF_X1 U19398 ( .A(n22734), .Z(n27093) );
  BUF_X1 U19399 ( .A(n22745), .Z(n27029) );
  BUF_X1 U19400 ( .A(n22745), .Z(n27030) );
  BUF_X1 U19401 ( .A(n22745), .Z(n27031) );
  BUF_X1 U19402 ( .A(n22745), .Z(n27032) );
  BUF_X1 U19403 ( .A(n22745), .Z(n27033) );
  BUF_X1 U19404 ( .A(n22747), .Z(n27017) );
  BUF_X1 U19405 ( .A(n22747), .Z(n27018) );
  BUF_X1 U19406 ( .A(n22747), .Z(n27019) );
  BUF_X1 U19407 ( .A(n22747), .Z(n27020) );
  BUF_X1 U19408 ( .A(n22747), .Z(n27021) );
  BUF_X1 U19409 ( .A(n23980), .Z(n26636) );
  BUF_X1 U19410 ( .A(n23980), .Z(n26637) );
  BUF_X1 U19411 ( .A(n23980), .Z(n26638) );
  BUF_X1 U19412 ( .A(n23980), .Z(n26639) );
  BUF_X1 U19413 ( .A(n23980), .Z(n26640) );
  BUF_X1 U19414 ( .A(n22781), .Z(n26861) );
  BUF_X1 U19415 ( .A(n22781), .Z(n26862) );
  BUF_X1 U19416 ( .A(n22781), .Z(n26863) );
  BUF_X1 U19417 ( .A(n22781), .Z(n26864) );
  BUF_X1 U19418 ( .A(n22781), .Z(n26865) );
  BUF_X1 U19419 ( .A(n22760), .Z(n26945) );
  BUF_X1 U19420 ( .A(n22753), .Z(n26981) );
  BUF_X1 U19421 ( .A(n22764), .Z(n26921) );
  BUF_X1 U19422 ( .A(n22762), .Z(n26933) );
  BUF_X1 U19423 ( .A(n22758), .Z(n26957) );
  BUF_X1 U19424 ( .A(n22756), .Z(n26969) );
  BUF_X1 U19425 ( .A(n22768), .Z(n26897) );
  BUF_X1 U19426 ( .A(n22766), .Z(n26909) );
  BUF_X1 U19427 ( .A(n22722), .Z(n27161) );
  BUF_X1 U19428 ( .A(n22719), .Z(n27173) );
  BUF_X1 U19429 ( .A(n22724), .Z(n27149) );
  BUF_X1 U19430 ( .A(n22743), .Z(n27041) );
  BUF_X1 U19431 ( .A(n22693), .Z(n27269) );
  BUF_X1 U19432 ( .A(n22697), .Z(n27257) );
  BUF_X1 U19433 ( .A(n22715), .Z(n27185) );
  BUF_X1 U19434 ( .A(n22726), .Z(n27137) );
  BUF_X1 U19435 ( .A(n22706), .Z(n27221) );
  BUF_X1 U19436 ( .A(n22712), .Z(n27197) );
  BUF_X1 U19437 ( .A(n22749), .Z(n27005) );
  BUF_X1 U19438 ( .A(n22739), .Z(n27065) );
  BUF_X1 U19439 ( .A(n22741), .Z(n27053) );
  BUF_X1 U19440 ( .A(n22709), .Z(n27209) );
  BUF_X1 U19441 ( .A(n22700), .Z(n27245) );
  BUF_X1 U19442 ( .A(n22703), .Z(n27233) );
  BUF_X1 U19443 ( .A(n22751), .Z(n26993) );
  BUF_X1 U19444 ( .A(n22736), .Z(n27077) );
  BUF_X1 U19445 ( .A(n22732), .Z(n27101) );
  BUF_X1 U19446 ( .A(n22728), .Z(n27125) );
  BUF_X1 U19447 ( .A(n26526), .Z(n26541) );
  BUF_X1 U19448 ( .A(n26526), .Z(n26540) );
  BUF_X1 U19449 ( .A(n26526), .Z(n26539) );
  BUF_X1 U19450 ( .A(n26525), .Z(n26538) );
  BUF_X1 U19451 ( .A(n26525), .Z(n26537) );
  BUF_X1 U19452 ( .A(n26751), .Z(n26766) );
  BUF_X1 U19453 ( .A(n26751), .Z(n26765) );
  BUF_X1 U19454 ( .A(n26751), .Z(n26764) );
  BUF_X1 U19455 ( .A(n26750), .Z(n26763) );
  BUF_X1 U19456 ( .A(n26750), .Z(n26762) );
  BUF_X1 U19457 ( .A(n26525), .Z(n26536) );
  BUF_X1 U19458 ( .A(n26750), .Z(n26761) );
  BUF_X1 U19459 ( .A(n26529), .Z(n26550) );
  BUF_X1 U19460 ( .A(n26529), .Z(n26549) );
  BUF_X1 U19461 ( .A(n26529), .Z(n26548) );
  BUF_X1 U19462 ( .A(n26528), .Z(n26547) );
  BUF_X1 U19463 ( .A(n26528), .Z(n26546) );
  BUF_X1 U19464 ( .A(n26528), .Z(n26545) );
  BUF_X1 U19465 ( .A(n26527), .Z(n26544) );
  BUF_X1 U19466 ( .A(n26527), .Z(n26543) );
  BUF_X1 U19467 ( .A(n26527), .Z(n26542) );
  BUF_X1 U19468 ( .A(n26754), .Z(n26775) );
  BUF_X1 U19469 ( .A(n26754), .Z(n26774) );
  BUF_X1 U19470 ( .A(n26754), .Z(n26773) );
  BUF_X1 U19471 ( .A(n26753), .Z(n26772) );
  BUF_X1 U19472 ( .A(n26753), .Z(n26771) );
  BUF_X1 U19473 ( .A(n26753), .Z(n26770) );
  BUF_X1 U19474 ( .A(n26752), .Z(n26768) );
  BUF_X1 U19475 ( .A(n26752), .Z(n26767) );
  BUF_X1 U19476 ( .A(n26752), .Z(n26769) );
  BUF_X1 U19477 ( .A(n26530), .Z(n26551) );
  BUF_X1 U19478 ( .A(n26755), .Z(n26776) );
  BUF_X1 U19479 ( .A(n23992), .Z(n26582) );
  BUF_X1 U19480 ( .A(n24017), .Z(n26459) );
  BUF_X1 U19481 ( .A(n23992), .Z(n26583) );
  BUF_X1 U19482 ( .A(n24017), .Z(n26460) );
  BUF_X1 U19483 ( .A(n23992), .Z(n26584) );
  BUF_X1 U19484 ( .A(n24017), .Z(n26461) );
  BUF_X1 U19485 ( .A(n23992), .Z(n26585) );
  BUF_X1 U19486 ( .A(n24017), .Z(n26462) );
  BUF_X1 U19487 ( .A(n23992), .Z(n26586) );
  BUF_X1 U19488 ( .A(n24017), .Z(n26463) );
  BUF_X1 U19489 ( .A(n22793), .Z(n26807) );
  BUF_X1 U19490 ( .A(n22818), .Z(n26684) );
  BUF_X1 U19491 ( .A(n22793), .Z(n26808) );
  BUF_X1 U19492 ( .A(n22818), .Z(n26685) );
  BUF_X1 U19493 ( .A(n22793), .Z(n26809) );
  BUF_X1 U19494 ( .A(n22818), .Z(n26686) );
  BUF_X1 U19495 ( .A(n22793), .Z(n26810) );
  BUF_X1 U19496 ( .A(n22818), .Z(n26687) );
  BUF_X1 U19497 ( .A(n22793), .Z(n26811) );
  BUF_X1 U19498 ( .A(n22818), .Z(n26688) );
  BUF_X1 U19499 ( .A(n24012), .Z(n26483) );
  BUF_X1 U19500 ( .A(n24012), .Z(n26484) );
  BUF_X1 U19501 ( .A(n24012), .Z(n26485) );
  BUF_X1 U19502 ( .A(n24012), .Z(n26486) );
  BUF_X1 U19503 ( .A(n24012), .Z(n26487) );
  BUF_X1 U19504 ( .A(n22813), .Z(n26708) );
  BUF_X1 U19505 ( .A(n22813), .Z(n26709) );
  BUF_X1 U19506 ( .A(n22813), .Z(n26710) );
  BUF_X1 U19507 ( .A(n22813), .Z(n26711) );
  BUF_X1 U19508 ( .A(n22813), .Z(n26712) );
  BUF_X1 U19509 ( .A(n23987), .Z(n26606) );
  BUF_X1 U19510 ( .A(n23977), .Z(n26654) );
  BUF_X1 U19511 ( .A(n23982), .Z(n26630) );
  BUF_X1 U19512 ( .A(n24007), .Z(n26507) );
  BUF_X1 U19513 ( .A(n24002), .Z(n26552) );
  BUF_X1 U19514 ( .A(n23987), .Z(n26607) );
  BUF_X1 U19515 ( .A(n23977), .Z(n26655) );
  BUF_X1 U19516 ( .A(n23982), .Z(n26631) );
  BUF_X1 U19517 ( .A(n24007), .Z(n26508) );
  BUF_X1 U19518 ( .A(n24002), .Z(n26553) );
  BUF_X1 U19519 ( .A(n23987), .Z(n26608) );
  BUF_X1 U19520 ( .A(n23977), .Z(n26656) );
  BUF_X1 U19521 ( .A(n23982), .Z(n26632) );
  BUF_X1 U19522 ( .A(n24007), .Z(n26509) );
  BUF_X1 U19523 ( .A(n24002), .Z(n26554) );
  BUF_X1 U19524 ( .A(n23987), .Z(n26609) );
  BUF_X1 U19525 ( .A(n23977), .Z(n26657) );
  BUF_X1 U19526 ( .A(n23982), .Z(n26633) );
  BUF_X1 U19527 ( .A(n24007), .Z(n26510) );
  BUF_X1 U19528 ( .A(n24002), .Z(n26555) );
  BUF_X1 U19529 ( .A(n23987), .Z(n26610) );
  BUF_X1 U19530 ( .A(n23977), .Z(n26658) );
  BUF_X1 U19531 ( .A(n23982), .Z(n26634) );
  BUF_X1 U19532 ( .A(n24007), .Z(n26511) );
  BUF_X1 U19533 ( .A(n24002), .Z(n26556) );
  BUF_X1 U19534 ( .A(n22788), .Z(n26831) );
  BUF_X1 U19535 ( .A(n22778), .Z(n26879) );
  BUF_X1 U19536 ( .A(n22783), .Z(n26855) );
  BUF_X1 U19537 ( .A(n22808), .Z(n26732) );
  BUF_X1 U19538 ( .A(n22803), .Z(n26777) );
  BUF_X1 U19539 ( .A(n22788), .Z(n26832) );
  BUF_X1 U19540 ( .A(n22778), .Z(n26880) );
  BUF_X1 U19541 ( .A(n22783), .Z(n26856) );
  BUF_X1 U19542 ( .A(n22808), .Z(n26733) );
  BUF_X1 U19543 ( .A(n22803), .Z(n26778) );
  BUF_X1 U19544 ( .A(n22788), .Z(n26833) );
  BUF_X1 U19545 ( .A(n22778), .Z(n26881) );
  BUF_X1 U19546 ( .A(n22783), .Z(n26857) );
  BUF_X1 U19547 ( .A(n22808), .Z(n26734) );
  BUF_X1 U19548 ( .A(n22803), .Z(n26779) );
  BUF_X1 U19549 ( .A(n22788), .Z(n26834) );
  BUF_X1 U19550 ( .A(n22778), .Z(n26882) );
  BUF_X1 U19551 ( .A(n22783), .Z(n26858) );
  BUF_X1 U19552 ( .A(n22808), .Z(n26735) );
  BUF_X1 U19553 ( .A(n22803), .Z(n26780) );
  BUF_X1 U19554 ( .A(n22788), .Z(n26835) );
  BUF_X1 U19555 ( .A(n22778), .Z(n26883) );
  BUF_X1 U19556 ( .A(n22783), .Z(n26859) );
  BUF_X1 U19557 ( .A(n22808), .Z(n26736) );
  BUF_X1 U19558 ( .A(n22803), .Z(n26781) );
  BUF_X1 U19559 ( .A(n23989), .Z(n26595) );
  BUF_X1 U19560 ( .A(n23984), .Z(n26619) );
  BUF_X1 U19561 ( .A(n23974), .Z(n26667) );
  BUF_X1 U19562 ( .A(n23979), .Z(n26643) );
  BUF_X1 U19563 ( .A(n24004), .Z(n26520) );
  BUF_X1 U19564 ( .A(n23999), .Z(n26565) );
  BUF_X1 U19565 ( .A(n23989), .Z(n26596) );
  BUF_X1 U19566 ( .A(n23984), .Z(n26620) );
  BUF_X1 U19567 ( .A(n23974), .Z(n26668) );
  BUF_X1 U19568 ( .A(n23979), .Z(n26644) );
  BUF_X1 U19569 ( .A(n24004), .Z(n26521) );
  BUF_X1 U19570 ( .A(n23999), .Z(n26566) );
  BUF_X1 U19571 ( .A(n23989), .Z(n26597) );
  BUF_X1 U19572 ( .A(n23984), .Z(n26621) );
  BUF_X1 U19573 ( .A(n23974), .Z(n26669) );
  BUF_X1 U19574 ( .A(n23979), .Z(n26645) );
  BUF_X1 U19575 ( .A(n24004), .Z(n26522) );
  BUF_X1 U19576 ( .A(n23999), .Z(n26567) );
  BUF_X1 U19577 ( .A(n23989), .Z(n26598) );
  BUF_X1 U19578 ( .A(n23984), .Z(n26622) );
  BUF_X1 U19579 ( .A(n23974), .Z(n26670) );
  BUF_X1 U19580 ( .A(n23979), .Z(n26646) );
  BUF_X1 U19581 ( .A(n24004), .Z(n26523) );
  BUF_X1 U19582 ( .A(n23999), .Z(n26568) );
  BUF_X1 U19583 ( .A(n22790), .Z(n26820) );
  BUF_X1 U19584 ( .A(n22785), .Z(n26844) );
  BUF_X1 U19585 ( .A(n22775), .Z(n26892) );
  BUF_X1 U19586 ( .A(n22780), .Z(n26868) );
  BUF_X1 U19587 ( .A(n22805), .Z(n26745) );
  BUF_X1 U19588 ( .A(n22800), .Z(n26790) );
  BUF_X1 U19589 ( .A(n22790), .Z(n26821) );
  BUF_X1 U19590 ( .A(n22785), .Z(n26845) );
  BUF_X1 U19591 ( .A(n22775), .Z(n26893) );
  BUF_X1 U19592 ( .A(n22780), .Z(n26869) );
  BUF_X1 U19593 ( .A(n22805), .Z(n26746) );
  BUF_X1 U19594 ( .A(n22800), .Z(n26791) );
  BUF_X1 U19595 ( .A(n22790), .Z(n26822) );
  BUF_X1 U19596 ( .A(n22785), .Z(n26846) );
  BUF_X1 U19597 ( .A(n22775), .Z(n26894) );
  BUF_X1 U19598 ( .A(n22780), .Z(n26870) );
  BUF_X1 U19599 ( .A(n22805), .Z(n26747) );
  BUF_X1 U19600 ( .A(n22800), .Z(n26792) );
  BUF_X1 U19601 ( .A(n22790), .Z(n26823) );
  BUF_X1 U19602 ( .A(n22785), .Z(n26847) );
  BUF_X1 U19603 ( .A(n22775), .Z(n26895) );
  BUF_X1 U19604 ( .A(n22780), .Z(n26871) );
  BUF_X1 U19605 ( .A(n22805), .Z(n26748) );
  BUF_X1 U19606 ( .A(n22800), .Z(n26793) );
  BUF_X1 U19607 ( .A(n23993), .Z(n26576) );
  BUF_X1 U19608 ( .A(n24018), .Z(n26453) );
  BUF_X1 U19609 ( .A(n23993), .Z(n26577) );
  BUF_X1 U19610 ( .A(n24018), .Z(n26454) );
  BUF_X1 U19611 ( .A(n23993), .Z(n26578) );
  BUF_X1 U19612 ( .A(n24018), .Z(n26455) );
  BUF_X1 U19613 ( .A(n23993), .Z(n26579) );
  BUF_X1 U19614 ( .A(n24018), .Z(n26456) );
  BUF_X1 U19615 ( .A(n23993), .Z(n26580) );
  BUF_X1 U19616 ( .A(n24018), .Z(n26457) );
  BUF_X1 U19617 ( .A(n22794), .Z(n26801) );
  BUF_X1 U19618 ( .A(n22819), .Z(n26678) );
  BUF_X1 U19619 ( .A(n22794), .Z(n26802) );
  BUF_X1 U19620 ( .A(n22819), .Z(n26679) );
  BUF_X1 U19621 ( .A(n22794), .Z(n26803) );
  BUF_X1 U19622 ( .A(n22819), .Z(n26680) );
  BUF_X1 U19623 ( .A(n22794), .Z(n26804) );
  BUF_X1 U19624 ( .A(n22819), .Z(n26681) );
  BUF_X1 U19625 ( .A(n22794), .Z(n26805) );
  BUF_X1 U19626 ( .A(n22819), .Z(n26682) );
  BUF_X1 U19627 ( .A(n23988), .Z(n26600) );
  BUF_X1 U19628 ( .A(n23978), .Z(n26648) );
  BUF_X1 U19629 ( .A(n23983), .Z(n26624) );
  BUF_X1 U19630 ( .A(n24008), .Z(n26501) );
  BUF_X1 U19631 ( .A(n24013), .Z(n26477) );
  BUF_X1 U19632 ( .A(n23988), .Z(n26601) );
  BUF_X1 U19633 ( .A(n23978), .Z(n26649) );
  BUF_X1 U19634 ( .A(n23983), .Z(n26625) );
  BUF_X1 U19635 ( .A(n24008), .Z(n26502) );
  BUF_X1 U19636 ( .A(n24013), .Z(n26478) );
  BUF_X1 U19637 ( .A(n23988), .Z(n26602) );
  BUF_X1 U19638 ( .A(n23978), .Z(n26650) );
  BUF_X1 U19639 ( .A(n23983), .Z(n26626) );
  BUF_X1 U19640 ( .A(n24008), .Z(n26503) );
  BUF_X1 U19641 ( .A(n24013), .Z(n26479) );
  BUF_X1 U19642 ( .A(n23988), .Z(n26603) );
  BUF_X1 U19643 ( .A(n23978), .Z(n26651) );
  BUF_X1 U19644 ( .A(n23983), .Z(n26627) );
  BUF_X1 U19645 ( .A(n24008), .Z(n26504) );
  BUF_X1 U19646 ( .A(n24013), .Z(n26480) );
  BUF_X1 U19647 ( .A(n23988), .Z(n26604) );
  BUF_X1 U19648 ( .A(n23978), .Z(n26652) );
  BUF_X1 U19649 ( .A(n23983), .Z(n26628) );
  BUF_X1 U19650 ( .A(n24008), .Z(n26505) );
  BUF_X1 U19651 ( .A(n24013), .Z(n26481) );
  BUF_X1 U19652 ( .A(n22789), .Z(n26825) );
  BUF_X1 U19653 ( .A(n22779), .Z(n26873) );
  BUF_X1 U19654 ( .A(n22784), .Z(n26849) );
  BUF_X1 U19655 ( .A(n22809), .Z(n26726) );
  BUF_X1 U19656 ( .A(n22814), .Z(n26702) );
  BUF_X1 U19657 ( .A(n22789), .Z(n26826) );
  BUF_X1 U19658 ( .A(n22779), .Z(n26874) );
  BUF_X1 U19659 ( .A(n22784), .Z(n26850) );
  BUF_X1 U19660 ( .A(n22809), .Z(n26727) );
  BUF_X1 U19661 ( .A(n22814), .Z(n26703) );
  BUF_X1 U19662 ( .A(n22789), .Z(n26827) );
  BUF_X1 U19663 ( .A(n22779), .Z(n26875) );
  BUF_X1 U19664 ( .A(n22784), .Z(n26851) );
  BUF_X1 U19665 ( .A(n22809), .Z(n26728) );
  BUF_X1 U19666 ( .A(n22814), .Z(n26704) );
  BUF_X1 U19667 ( .A(n22789), .Z(n26828) );
  BUF_X1 U19668 ( .A(n22779), .Z(n26876) );
  BUF_X1 U19669 ( .A(n22784), .Z(n26852) );
  BUF_X1 U19670 ( .A(n22809), .Z(n26729) );
  BUF_X1 U19671 ( .A(n22814), .Z(n26705) );
  BUF_X1 U19672 ( .A(n22789), .Z(n26829) );
  BUF_X1 U19673 ( .A(n22779), .Z(n26877) );
  BUF_X1 U19674 ( .A(n22784), .Z(n26853) );
  BUF_X1 U19675 ( .A(n22809), .Z(n26730) );
  BUF_X1 U19676 ( .A(n22814), .Z(n26706) );
  BUF_X1 U19677 ( .A(n23994), .Z(n26570) );
  BUF_X1 U19678 ( .A(n24019), .Z(n26447) );
  BUF_X1 U19679 ( .A(n23994), .Z(n26571) );
  BUF_X1 U19680 ( .A(n24019), .Z(n26448) );
  BUF_X1 U19681 ( .A(n23994), .Z(n26572) );
  BUF_X1 U19682 ( .A(n24019), .Z(n26449) );
  BUF_X1 U19683 ( .A(n23994), .Z(n26573) );
  BUF_X1 U19684 ( .A(n24019), .Z(n26450) );
  BUF_X1 U19685 ( .A(n23994), .Z(n26574) );
  BUF_X1 U19686 ( .A(n24019), .Z(n26451) );
  BUF_X1 U19687 ( .A(n22795), .Z(n26795) );
  BUF_X1 U19688 ( .A(n22820), .Z(n26672) );
  BUF_X1 U19689 ( .A(n22795), .Z(n26796) );
  BUF_X1 U19690 ( .A(n22820), .Z(n26673) );
  BUF_X1 U19691 ( .A(n22795), .Z(n26797) );
  BUF_X1 U19692 ( .A(n22820), .Z(n26674) );
  BUF_X1 U19693 ( .A(n22795), .Z(n26798) );
  BUF_X1 U19694 ( .A(n22820), .Z(n26675) );
  BUF_X1 U19695 ( .A(n22795), .Z(n26799) );
  BUF_X1 U19696 ( .A(n22820), .Z(n26676) );
  BUF_X1 U19697 ( .A(n22696), .Z(n27263) );
  BUF_X1 U19698 ( .A(n22714), .Z(n27191) );
  BUF_X1 U19699 ( .A(n22705), .Z(n27227) );
  BUF_X1 U19700 ( .A(n22711), .Z(n27203) );
  BUF_X1 U19701 ( .A(n22708), .Z(n27215) );
  BUF_X1 U19702 ( .A(n22699), .Z(n27251) );
  BUF_X1 U19703 ( .A(n22702), .Z(n27239) );
  BUF_X1 U19704 ( .A(n22721), .Z(n27167) );
  BUF_X1 U19705 ( .A(n22759), .Z(n26951) );
  BUF_X1 U19706 ( .A(n22752), .Z(n26987) );
  BUF_X1 U19707 ( .A(n22718), .Z(n27179) );
  BUF_X1 U19708 ( .A(n22723), .Z(n27155) );
  BUF_X1 U19709 ( .A(n22742), .Z(n27047) );
  BUF_X1 U19710 ( .A(n22763), .Z(n26927) );
  BUF_X1 U19711 ( .A(n22761), .Z(n26939) );
  BUF_X1 U19712 ( .A(n22725), .Z(n27143) );
  BUF_X1 U19713 ( .A(n22748), .Z(n27011) );
  BUF_X1 U19714 ( .A(n22738), .Z(n27071) );
  BUF_X1 U19715 ( .A(n22740), .Z(n27059) );
  BUF_X1 U19716 ( .A(n22757), .Z(n26963) );
  BUF_X1 U19717 ( .A(n22750), .Z(n26999) );
  BUF_X1 U19718 ( .A(n22735), .Z(n27083) );
  BUF_X1 U19719 ( .A(n22755), .Z(n26975) );
  BUF_X1 U19720 ( .A(n22729), .Z(n27119) );
  BUF_X1 U19721 ( .A(n22733), .Z(n27095) );
  BUF_X1 U19722 ( .A(n22744), .Z(n27035) );
  BUF_X1 U19723 ( .A(n22746), .Z(n27023) );
  BUF_X1 U19724 ( .A(n22767), .Z(n26903) );
  BUF_X1 U19725 ( .A(n22765), .Z(n26915) );
  BUF_X1 U19726 ( .A(n22731), .Z(n27107) );
  BUF_X1 U19727 ( .A(n22727), .Z(n27131) );
  BUF_X1 U19728 ( .A(n22696), .Z(n27264) );
  BUF_X1 U19729 ( .A(n22696), .Z(n27265) );
  BUF_X1 U19730 ( .A(n22696), .Z(n27266) );
  BUF_X1 U19731 ( .A(n22696), .Z(n27267) );
  BUF_X1 U19732 ( .A(n22714), .Z(n27192) );
  BUF_X1 U19733 ( .A(n22714), .Z(n27193) );
  BUF_X1 U19734 ( .A(n22714), .Z(n27194) );
  BUF_X1 U19735 ( .A(n22714), .Z(n27195) );
  BUF_X1 U19736 ( .A(n22705), .Z(n27228) );
  BUF_X1 U19737 ( .A(n22705), .Z(n27229) );
  BUF_X1 U19738 ( .A(n22705), .Z(n27230) );
  BUF_X1 U19739 ( .A(n22705), .Z(n27231) );
  BUF_X1 U19740 ( .A(n22711), .Z(n27204) );
  BUF_X1 U19741 ( .A(n22711), .Z(n27205) );
  BUF_X1 U19742 ( .A(n22711), .Z(n27206) );
  BUF_X1 U19743 ( .A(n22711), .Z(n27207) );
  BUF_X1 U19744 ( .A(n22708), .Z(n27216) );
  BUF_X1 U19745 ( .A(n22708), .Z(n27217) );
  BUF_X1 U19746 ( .A(n22708), .Z(n27218) );
  BUF_X1 U19747 ( .A(n22708), .Z(n27219) );
  BUF_X1 U19748 ( .A(n22699), .Z(n27252) );
  BUF_X1 U19749 ( .A(n22699), .Z(n27253) );
  BUF_X1 U19750 ( .A(n22699), .Z(n27254) );
  BUF_X1 U19751 ( .A(n22699), .Z(n27255) );
  BUF_X1 U19752 ( .A(n22702), .Z(n27240) );
  BUF_X1 U19753 ( .A(n22702), .Z(n27241) );
  BUF_X1 U19754 ( .A(n22702), .Z(n27242) );
  BUF_X1 U19755 ( .A(n22702), .Z(n27243) );
  BUF_X1 U19756 ( .A(n22721), .Z(n27168) );
  BUF_X1 U19757 ( .A(n22721), .Z(n27169) );
  BUF_X1 U19758 ( .A(n22721), .Z(n27170) );
  BUF_X1 U19759 ( .A(n22721), .Z(n27171) );
  BUF_X1 U19760 ( .A(n22759), .Z(n26952) );
  BUF_X1 U19761 ( .A(n22759), .Z(n26953) );
  BUF_X1 U19762 ( .A(n22759), .Z(n26954) );
  BUF_X1 U19763 ( .A(n22759), .Z(n26955) );
  BUF_X1 U19764 ( .A(n22752), .Z(n26988) );
  BUF_X1 U19765 ( .A(n22752), .Z(n26989) );
  BUF_X1 U19766 ( .A(n22752), .Z(n26990) );
  BUF_X1 U19767 ( .A(n22752), .Z(n26991) );
  BUF_X1 U19768 ( .A(n22718), .Z(n27180) );
  BUF_X1 U19769 ( .A(n22718), .Z(n27181) );
  BUF_X1 U19770 ( .A(n22718), .Z(n27182) );
  BUF_X1 U19771 ( .A(n22718), .Z(n27183) );
  BUF_X1 U19772 ( .A(n22723), .Z(n27156) );
  BUF_X1 U19773 ( .A(n22723), .Z(n27157) );
  BUF_X1 U19774 ( .A(n22723), .Z(n27158) );
  BUF_X1 U19775 ( .A(n22723), .Z(n27159) );
  BUF_X1 U19776 ( .A(n22742), .Z(n27048) );
  BUF_X1 U19777 ( .A(n22742), .Z(n27049) );
  BUF_X1 U19778 ( .A(n22742), .Z(n27050) );
  BUF_X1 U19779 ( .A(n22742), .Z(n27051) );
  BUF_X1 U19780 ( .A(n22763), .Z(n26928) );
  BUF_X1 U19781 ( .A(n22763), .Z(n26929) );
  BUF_X1 U19782 ( .A(n22763), .Z(n26930) );
  BUF_X1 U19783 ( .A(n22763), .Z(n26931) );
  BUF_X1 U19784 ( .A(n22761), .Z(n26940) );
  BUF_X1 U19785 ( .A(n22761), .Z(n26941) );
  BUF_X1 U19786 ( .A(n22761), .Z(n26942) );
  BUF_X1 U19787 ( .A(n22761), .Z(n26943) );
  BUF_X1 U19788 ( .A(n22725), .Z(n27144) );
  BUF_X1 U19789 ( .A(n22725), .Z(n27145) );
  BUF_X1 U19790 ( .A(n22725), .Z(n27146) );
  BUF_X1 U19791 ( .A(n22725), .Z(n27147) );
  BUF_X1 U19792 ( .A(n22748), .Z(n27012) );
  BUF_X1 U19793 ( .A(n22748), .Z(n27013) );
  BUF_X1 U19794 ( .A(n22748), .Z(n27014) );
  BUF_X1 U19795 ( .A(n22748), .Z(n27015) );
  BUF_X1 U19796 ( .A(n22738), .Z(n27072) );
  BUF_X1 U19797 ( .A(n22738), .Z(n27073) );
  BUF_X1 U19798 ( .A(n22738), .Z(n27074) );
  BUF_X1 U19799 ( .A(n22738), .Z(n27075) );
  BUF_X1 U19800 ( .A(n22740), .Z(n27060) );
  BUF_X1 U19801 ( .A(n22740), .Z(n27061) );
  BUF_X1 U19802 ( .A(n22740), .Z(n27062) );
  BUF_X1 U19803 ( .A(n22740), .Z(n27063) );
  BUF_X1 U19804 ( .A(n22757), .Z(n26964) );
  BUF_X1 U19805 ( .A(n22757), .Z(n26965) );
  BUF_X1 U19806 ( .A(n22757), .Z(n26966) );
  BUF_X1 U19807 ( .A(n22757), .Z(n26967) );
  BUF_X1 U19808 ( .A(n22750), .Z(n27000) );
  BUF_X1 U19809 ( .A(n22750), .Z(n27001) );
  BUF_X1 U19810 ( .A(n22750), .Z(n27002) );
  BUF_X1 U19811 ( .A(n22750), .Z(n27003) );
  BUF_X1 U19812 ( .A(n22735), .Z(n27084) );
  BUF_X1 U19813 ( .A(n22735), .Z(n27085) );
  BUF_X1 U19814 ( .A(n22735), .Z(n27086) );
  BUF_X1 U19815 ( .A(n22735), .Z(n27087) );
  BUF_X1 U19816 ( .A(n22755), .Z(n26976) );
  BUF_X1 U19817 ( .A(n22755), .Z(n26977) );
  BUF_X1 U19818 ( .A(n22755), .Z(n26978) );
  BUF_X1 U19819 ( .A(n22755), .Z(n26979) );
  BUF_X1 U19820 ( .A(n22729), .Z(n27120) );
  BUF_X1 U19821 ( .A(n22729), .Z(n27121) );
  BUF_X1 U19822 ( .A(n22729), .Z(n27122) );
  BUF_X1 U19823 ( .A(n22729), .Z(n27123) );
  BUF_X1 U19824 ( .A(n22733), .Z(n27096) );
  BUF_X1 U19825 ( .A(n22733), .Z(n27097) );
  BUF_X1 U19826 ( .A(n22733), .Z(n27098) );
  BUF_X1 U19827 ( .A(n22733), .Z(n27099) );
  BUF_X1 U19828 ( .A(n22744), .Z(n27036) );
  BUF_X1 U19829 ( .A(n22744), .Z(n27037) );
  BUF_X1 U19830 ( .A(n22744), .Z(n27038) );
  BUF_X1 U19831 ( .A(n22744), .Z(n27039) );
  BUF_X1 U19832 ( .A(n22746), .Z(n27024) );
  BUF_X1 U19833 ( .A(n22746), .Z(n27025) );
  BUF_X1 U19834 ( .A(n22746), .Z(n27026) );
  BUF_X1 U19835 ( .A(n22746), .Z(n27027) );
  BUF_X1 U19836 ( .A(n22767), .Z(n26904) );
  BUF_X1 U19837 ( .A(n22767), .Z(n26905) );
  BUF_X1 U19838 ( .A(n22767), .Z(n26906) );
  BUF_X1 U19839 ( .A(n22767), .Z(n26907) );
  BUF_X1 U19840 ( .A(n22765), .Z(n26916) );
  BUF_X1 U19841 ( .A(n22765), .Z(n26917) );
  BUF_X1 U19842 ( .A(n22765), .Z(n26918) );
  BUF_X1 U19843 ( .A(n22765), .Z(n26919) );
  BUF_X1 U19844 ( .A(n22731), .Z(n27108) );
  BUF_X1 U19845 ( .A(n22731), .Z(n27109) );
  BUF_X1 U19846 ( .A(n22731), .Z(n27110) );
  BUF_X1 U19847 ( .A(n22731), .Z(n27111) );
  BUF_X1 U19848 ( .A(n22727), .Z(n27132) );
  BUF_X1 U19849 ( .A(n22727), .Z(n27133) );
  BUF_X1 U19850 ( .A(n22727), .Z(n27134) );
  BUF_X1 U19851 ( .A(n22727), .Z(n27135) );
  NAND2_X1 U19852 ( .A1(n25143), .A2(n25151), .ZN(n23980) );
  NAND2_X1 U19853 ( .A1(n23944), .A2(n23952), .ZN(n22781) );
  NAND2_X1 U19854 ( .A1(n27475), .A2(n27119), .ZN(n22730) );
  NAND2_X1 U19855 ( .A1(n27475), .A2(n27095), .ZN(n22734) );
  NAND2_X1 U19856 ( .A1(n27475), .A2(n27035), .ZN(n22745) );
  NAND2_X1 U19857 ( .A1(n27475), .A2(n27023), .ZN(n22747) );
  BUF_X1 U19858 ( .A(n23990), .Z(n26588) );
  BUF_X1 U19859 ( .A(n23985), .Z(n26612) );
  BUF_X1 U19860 ( .A(n23975), .Z(n26660) );
  BUF_X1 U19861 ( .A(n24005), .Z(n26513) );
  BUF_X1 U19862 ( .A(n24000), .Z(n26558) );
  BUF_X1 U19863 ( .A(n23990), .Z(n26589) );
  BUF_X1 U19864 ( .A(n23985), .Z(n26613) );
  BUF_X1 U19865 ( .A(n23975), .Z(n26661) );
  BUF_X1 U19866 ( .A(n24005), .Z(n26514) );
  BUF_X1 U19867 ( .A(n24000), .Z(n26559) );
  BUF_X1 U19868 ( .A(n23990), .Z(n26590) );
  BUF_X1 U19869 ( .A(n23985), .Z(n26614) );
  BUF_X1 U19870 ( .A(n23975), .Z(n26662) );
  BUF_X1 U19871 ( .A(n24005), .Z(n26515) );
  BUF_X1 U19872 ( .A(n24000), .Z(n26560) );
  BUF_X1 U19873 ( .A(n23990), .Z(n26591) );
  BUF_X1 U19874 ( .A(n23985), .Z(n26615) );
  BUF_X1 U19875 ( .A(n23975), .Z(n26663) );
  BUF_X1 U19876 ( .A(n24005), .Z(n26516) );
  BUF_X1 U19877 ( .A(n24000), .Z(n26561) );
  BUF_X1 U19878 ( .A(n23990), .Z(n26592) );
  BUF_X1 U19879 ( .A(n23985), .Z(n26616) );
  BUF_X1 U19880 ( .A(n23975), .Z(n26664) );
  BUF_X1 U19881 ( .A(n24005), .Z(n26517) );
  BUF_X1 U19882 ( .A(n24000), .Z(n26562) );
  BUF_X1 U19883 ( .A(n22791), .Z(n26813) );
  BUF_X1 U19884 ( .A(n22786), .Z(n26837) );
  BUF_X1 U19885 ( .A(n22776), .Z(n26885) );
  BUF_X1 U19886 ( .A(n22806), .Z(n26738) );
  BUF_X1 U19887 ( .A(n22801), .Z(n26783) );
  BUF_X1 U19888 ( .A(n22791), .Z(n26814) );
  BUF_X1 U19889 ( .A(n22786), .Z(n26838) );
  BUF_X1 U19890 ( .A(n22776), .Z(n26886) );
  BUF_X1 U19891 ( .A(n22806), .Z(n26739) );
  BUF_X1 U19892 ( .A(n22801), .Z(n26784) );
  BUF_X1 U19893 ( .A(n22791), .Z(n26815) );
  BUF_X1 U19894 ( .A(n22786), .Z(n26839) );
  BUF_X1 U19895 ( .A(n22776), .Z(n26887) );
  BUF_X1 U19896 ( .A(n22806), .Z(n26740) );
  BUF_X1 U19897 ( .A(n22801), .Z(n26785) );
  BUF_X1 U19898 ( .A(n22791), .Z(n26816) );
  BUF_X1 U19899 ( .A(n22786), .Z(n26840) );
  BUF_X1 U19900 ( .A(n22776), .Z(n26888) );
  BUF_X1 U19901 ( .A(n22806), .Z(n26741) );
  BUF_X1 U19902 ( .A(n22801), .Z(n26786) );
  BUF_X1 U19903 ( .A(n22791), .Z(n26817) );
  BUF_X1 U19904 ( .A(n22786), .Z(n26841) );
  BUF_X1 U19905 ( .A(n22776), .Z(n26889) );
  BUF_X1 U19906 ( .A(n22806), .Z(n26742) );
  BUF_X1 U19907 ( .A(n22801), .Z(n26787) );
  BUF_X1 U19908 ( .A(n23989), .Z(n26594) );
  BUF_X1 U19909 ( .A(n23984), .Z(n26618) );
  BUF_X1 U19910 ( .A(n23974), .Z(n26666) );
  BUF_X1 U19911 ( .A(n23979), .Z(n26642) );
  BUF_X1 U19912 ( .A(n24004), .Z(n26519) );
  BUF_X1 U19913 ( .A(n23999), .Z(n26564) );
  BUF_X1 U19914 ( .A(n22790), .Z(n26819) );
  BUF_X1 U19915 ( .A(n22785), .Z(n26843) );
  BUF_X1 U19916 ( .A(n22775), .Z(n26891) );
  BUF_X1 U19917 ( .A(n22780), .Z(n26867) );
  BUF_X1 U19918 ( .A(n22805), .Z(n26744) );
  BUF_X1 U19919 ( .A(n22800), .Z(n26789) );
  NAND2_X1 U19920 ( .A1(n27476), .A2(n26951), .ZN(n22760) );
  NAND2_X1 U19921 ( .A1(n27476), .A2(n26987), .ZN(n22753) );
  NAND2_X1 U19922 ( .A1(n27476), .A2(n26927), .ZN(n22764) );
  NAND2_X1 U19923 ( .A1(n27476), .A2(n26939), .ZN(n22762) );
  NAND2_X1 U19924 ( .A1(n27476), .A2(n26963), .ZN(n22758) );
  NAND2_X1 U19925 ( .A1(n27476), .A2(n26975), .ZN(n22756) );
  NAND2_X1 U19926 ( .A1(n27476), .A2(n26903), .ZN(n22768) );
  NAND2_X1 U19927 ( .A1(n27476), .A2(n26915), .ZN(n22766) );
  NAND2_X1 U19928 ( .A1(n27474), .A2(n27263), .ZN(n22697) );
  NAND2_X1 U19929 ( .A1(n27474), .A2(n27251), .ZN(n22700) );
  NAND2_X1 U19930 ( .A1(n27474), .A2(n27239), .ZN(n22703) );
  NAND2_X1 U19931 ( .A1(n27474), .A2(n27167), .ZN(n22722) );
  NAND2_X1 U19932 ( .A1(n27474), .A2(n27179), .ZN(n22719) );
  NAND2_X1 U19933 ( .A1(n27474), .A2(n27155), .ZN(n22724) );
  NAND2_X1 U19934 ( .A1(n27475), .A2(n27047), .ZN(n22743) );
  NAND2_X1 U19935 ( .A1(n27474), .A2(n27277), .ZN(n22693) );
  NAND2_X1 U19936 ( .A1(n27474), .A2(n27143), .ZN(n22726) );
  NAND2_X1 U19937 ( .A1(n27475), .A2(n27011), .ZN(n22749) );
  NAND2_X1 U19938 ( .A1(n27475), .A2(n27071), .ZN(n22739) );
  NAND2_X1 U19939 ( .A1(n27475), .A2(n27059), .ZN(n22741) );
  NAND2_X1 U19940 ( .A1(n27475), .A2(n26999), .ZN(n22751) );
  NAND2_X1 U19941 ( .A1(n27475), .A2(n27083), .ZN(n22736) );
  NAND2_X1 U19942 ( .A1(n27474), .A2(n27191), .ZN(n22715) );
  NAND2_X1 U19943 ( .A1(n27474), .A2(n27227), .ZN(n22706) );
  NAND2_X1 U19944 ( .A1(n27474), .A2(n27203), .ZN(n22712) );
  NAND2_X1 U19945 ( .A1(n27474), .A2(n27215), .ZN(n22709) );
  NAND2_X1 U19946 ( .A1(n27475), .A2(n27107), .ZN(n22732) );
  NAND2_X1 U19947 ( .A1(n27475), .A2(n27131), .ZN(n22728) );
  BUF_X1 U19948 ( .A(n22692), .Z(n27275) );
  BUF_X1 U19949 ( .A(n22692), .Z(n27276) );
  BUF_X1 U19950 ( .A(n26531), .Z(n26529) );
  BUF_X1 U19951 ( .A(n26531), .Z(n26528) );
  BUF_X1 U19952 ( .A(n26532), .Z(n26527) );
  BUF_X1 U19953 ( .A(n26532), .Z(n26526) );
  BUF_X1 U19954 ( .A(n26532), .Z(n26525) );
  BUF_X1 U19955 ( .A(n26756), .Z(n26754) );
  BUF_X1 U19956 ( .A(n26756), .Z(n26753) );
  BUF_X1 U19957 ( .A(n26757), .Z(n26751) );
  BUF_X1 U19958 ( .A(n26757), .Z(n26750) );
  BUF_X1 U19959 ( .A(n26757), .Z(n26752) );
  BUF_X1 U19960 ( .A(n26531), .Z(n26530) );
  BUF_X1 U19961 ( .A(n26756), .Z(n26755) );
  OAI22_X1 U19962 ( .A1(n27318), .A2(n27168), .B1(n27162), .B2(n22679), .ZN(
        n7438) );
  OAI22_X1 U19963 ( .A1(n27321), .A2(n27168), .B1(n27162), .B2(n22678), .ZN(
        n7439) );
  OAI22_X1 U19964 ( .A1(n27324), .A2(n27168), .B1(n27162), .B2(n22677), .ZN(
        n7440) );
  OAI22_X1 U19965 ( .A1(n27327), .A2(n27168), .B1(n27162), .B2(n22676), .ZN(
        n7441) );
  OAI22_X1 U19966 ( .A1(n27330), .A2(n27168), .B1(n27162), .B2(n22675), .ZN(
        n7442) );
  OAI22_X1 U19967 ( .A1(n27333), .A2(n27168), .B1(n27162), .B2(n22674), .ZN(
        n7443) );
  OAI22_X1 U19968 ( .A1(n27336), .A2(n27168), .B1(n27162), .B2(n22673), .ZN(
        n7444) );
  OAI22_X1 U19969 ( .A1(n27339), .A2(n27168), .B1(n27162), .B2(n22672), .ZN(
        n7445) );
  OAI22_X1 U19970 ( .A1(n27342), .A2(n27168), .B1(n27162), .B2(n22671), .ZN(
        n7446) );
  OAI22_X1 U19971 ( .A1(n27345), .A2(n27168), .B1(n27162), .B2(n22670), .ZN(
        n7447) );
  OAI22_X1 U19972 ( .A1(n27348), .A2(n27168), .B1(n27162), .B2(n22669), .ZN(
        n7448) );
  OAI22_X1 U19973 ( .A1(n27351), .A2(n27169), .B1(n27162), .B2(n22668), .ZN(
        n7449) );
  OAI22_X1 U19974 ( .A1(n27354), .A2(n27169), .B1(n27163), .B2(n22667), .ZN(
        n7450) );
  OAI22_X1 U19975 ( .A1(n27357), .A2(n27169), .B1(n27163), .B2(n22666), .ZN(
        n7451) );
  OAI22_X1 U19976 ( .A1(n27360), .A2(n27169), .B1(n27163), .B2(n22665), .ZN(
        n7452) );
  OAI22_X1 U19977 ( .A1(n27363), .A2(n27169), .B1(n27163), .B2(n22664), .ZN(
        n7453) );
  OAI22_X1 U19978 ( .A1(n27366), .A2(n27169), .B1(n27163), .B2(n22663), .ZN(
        n7454) );
  OAI22_X1 U19979 ( .A1(n27369), .A2(n27169), .B1(n27163), .B2(n22662), .ZN(
        n7455) );
  OAI22_X1 U19980 ( .A1(n27372), .A2(n27169), .B1(n27163), .B2(n22661), .ZN(
        n7456) );
  OAI22_X1 U19981 ( .A1(n27375), .A2(n27169), .B1(n27163), .B2(n22660), .ZN(
        n7457) );
  OAI22_X1 U19982 ( .A1(n27378), .A2(n27169), .B1(n27163), .B2(n22659), .ZN(
        n7458) );
  OAI22_X1 U19983 ( .A1(n27381), .A2(n27169), .B1(n27163), .B2(n22658), .ZN(
        n7459) );
  OAI22_X1 U19984 ( .A1(n27384), .A2(n27169), .B1(n27163), .B2(n22657), .ZN(
        n7460) );
  OAI22_X1 U19985 ( .A1(n27387), .A2(n27170), .B1(n27163), .B2(n22656), .ZN(
        n7461) );
  OAI22_X1 U19986 ( .A1(n27390), .A2(n27170), .B1(n27164), .B2(n22655), .ZN(
        n7462) );
  OAI22_X1 U19987 ( .A1(n27393), .A2(n27170), .B1(n27164), .B2(n22654), .ZN(
        n7463) );
  OAI22_X1 U19988 ( .A1(n27396), .A2(n27170), .B1(n27164), .B2(n22653), .ZN(
        n7464) );
  OAI22_X1 U19989 ( .A1(n27399), .A2(n27170), .B1(n27164), .B2(n22652), .ZN(
        n7465) );
  OAI22_X1 U19990 ( .A1(n27402), .A2(n27170), .B1(n27164), .B2(n22651), .ZN(
        n7466) );
  OAI22_X1 U19991 ( .A1(n27405), .A2(n27170), .B1(n27164), .B2(n22650), .ZN(
        n7467) );
  OAI22_X1 U19992 ( .A1(n27408), .A2(n27170), .B1(n27164), .B2(n22649), .ZN(
        n7468) );
  OAI22_X1 U19993 ( .A1(n27411), .A2(n27170), .B1(n27164), .B2(n22648), .ZN(
        n7469) );
  OAI22_X1 U19994 ( .A1(n27414), .A2(n27170), .B1(n27164), .B2(n22647), .ZN(
        n7470) );
  OAI22_X1 U19995 ( .A1(n27417), .A2(n27170), .B1(n27164), .B2(n22646), .ZN(
        n7471) );
  OAI22_X1 U19996 ( .A1(n27420), .A2(n27170), .B1(n27164), .B2(n22645), .ZN(
        n7472) );
  OAI22_X1 U19997 ( .A1(n27423), .A2(n27171), .B1(n27164), .B2(n22644), .ZN(
        n7473) );
  OAI22_X1 U19998 ( .A1(n27426), .A2(n27171), .B1(n27165), .B2(n22643), .ZN(
        n7474) );
  OAI22_X1 U19999 ( .A1(n27429), .A2(n27171), .B1(n27165), .B2(n22642), .ZN(
        n7475) );
  OAI22_X1 U20000 ( .A1(n27432), .A2(n27171), .B1(n27165), .B2(n22641), .ZN(
        n7476) );
  OAI22_X1 U20001 ( .A1(n27435), .A2(n27171), .B1(n27165), .B2(n22640), .ZN(
        n7477) );
  OAI22_X1 U20002 ( .A1(n27438), .A2(n27171), .B1(n27165), .B2(n22639), .ZN(
        n7478) );
  OAI22_X1 U20003 ( .A1(n27441), .A2(n27171), .B1(n27165), .B2(n22638), .ZN(
        n7479) );
  OAI22_X1 U20004 ( .A1(n27444), .A2(n27171), .B1(n27165), .B2(n22637), .ZN(
        n7480) );
  OAI22_X1 U20005 ( .A1(n27447), .A2(n27171), .B1(n27165), .B2(n22636), .ZN(
        n7481) );
  OAI22_X1 U20006 ( .A1(n27450), .A2(n27171), .B1(n27165), .B2(n22635), .ZN(
        n7482) );
  OAI22_X1 U20007 ( .A1(n27453), .A2(n27171), .B1(n27165), .B2(n22634), .ZN(
        n7483) );
  OAI22_X1 U20008 ( .A1(n27456), .A2(n27171), .B1(n27165), .B2(n22633), .ZN(
        n7484) );
  OAI22_X1 U20009 ( .A1(n27459), .A2(n27172), .B1(n27165), .B2(n22632), .ZN(
        n7485) );
  OAI22_X1 U20010 ( .A1(n27319), .A2(n26988), .B1(n26982), .B2(n22559), .ZN(
        n6478) );
  OAI22_X1 U20011 ( .A1(n27322), .A2(n26988), .B1(n26982), .B2(n22558), .ZN(
        n6479) );
  OAI22_X1 U20012 ( .A1(n27325), .A2(n26988), .B1(n26982), .B2(n22557), .ZN(
        n6480) );
  OAI22_X1 U20013 ( .A1(n27328), .A2(n26988), .B1(n26982), .B2(n22556), .ZN(
        n6481) );
  OAI22_X1 U20014 ( .A1(n27331), .A2(n26988), .B1(n26982), .B2(n22555), .ZN(
        n6482) );
  OAI22_X1 U20015 ( .A1(n27334), .A2(n26988), .B1(n26982), .B2(n22554), .ZN(
        n6483) );
  OAI22_X1 U20016 ( .A1(n27337), .A2(n26988), .B1(n26982), .B2(n22553), .ZN(
        n6484) );
  OAI22_X1 U20017 ( .A1(n27340), .A2(n26988), .B1(n26982), .B2(n22552), .ZN(
        n6485) );
  OAI22_X1 U20018 ( .A1(n27343), .A2(n26988), .B1(n26982), .B2(n22551), .ZN(
        n6486) );
  OAI22_X1 U20019 ( .A1(n27346), .A2(n26988), .B1(n26982), .B2(n22550), .ZN(
        n6487) );
  OAI22_X1 U20020 ( .A1(n27349), .A2(n26988), .B1(n26982), .B2(n22549), .ZN(
        n6488) );
  OAI22_X1 U20021 ( .A1(n27352), .A2(n26989), .B1(n26982), .B2(n22548), .ZN(
        n6489) );
  OAI22_X1 U20022 ( .A1(n27355), .A2(n26989), .B1(n26983), .B2(n22547), .ZN(
        n6490) );
  OAI22_X1 U20023 ( .A1(n27358), .A2(n26989), .B1(n26983), .B2(n22546), .ZN(
        n6491) );
  OAI22_X1 U20024 ( .A1(n27361), .A2(n26989), .B1(n26983), .B2(n22545), .ZN(
        n6492) );
  OAI22_X1 U20025 ( .A1(n27364), .A2(n26989), .B1(n26983), .B2(n22544), .ZN(
        n6493) );
  OAI22_X1 U20026 ( .A1(n27367), .A2(n26989), .B1(n26983), .B2(n22543), .ZN(
        n6494) );
  OAI22_X1 U20027 ( .A1(n27370), .A2(n26989), .B1(n26983), .B2(n22542), .ZN(
        n6495) );
  OAI22_X1 U20028 ( .A1(n27373), .A2(n26989), .B1(n26983), .B2(n22541), .ZN(
        n6496) );
  OAI22_X1 U20029 ( .A1(n27376), .A2(n26989), .B1(n26983), .B2(n22540), .ZN(
        n6497) );
  OAI22_X1 U20030 ( .A1(n27379), .A2(n26989), .B1(n26983), .B2(n22539), .ZN(
        n6498) );
  OAI22_X1 U20031 ( .A1(n27382), .A2(n26989), .B1(n26983), .B2(n22538), .ZN(
        n6499) );
  OAI22_X1 U20032 ( .A1(n27385), .A2(n26989), .B1(n26983), .B2(n22537), .ZN(
        n6500) );
  OAI22_X1 U20033 ( .A1(n27388), .A2(n26990), .B1(n26983), .B2(n22536), .ZN(
        n6501) );
  OAI22_X1 U20034 ( .A1(n27391), .A2(n26990), .B1(n26984), .B2(n22535), .ZN(
        n6502) );
  OAI22_X1 U20035 ( .A1(n27394), .A2(n26990), .B1(n26984), .B2(n22534), .ZN(
        n6503) );
  OAI22_X1 U20036 ( .A1(n27397), .A2(n26990), .B1(n26984), .B2(n22533), .ZN(
        n6504) );
  OAI22_X1 U20037 ( .A1(n27400), .A2(n26990), .B1(n26984), .B2(n22532), .ZN(
        n6505) );
  OAI22_X1 U20038 ( .A1(n27403), .A2(n26990), .B1(n26984), .B2(n22531), .ZN(
        n6506) );
  OAI22_X1 U20039 ( .A1(n27406), .A2(n26990), .B1(n26984), .B2(n22530), .ZN(
        n6507) );
  OAI22_X1 U20040 ( .A1(n27409), .A2(n26990), .B1(n26984), .B2(n22529), .ZN(
        n6508) );
  OAI22_X1 U20041 ( .A1(n27412), .A2(n26990), .B1(n26984), .B2(n22528), .ZN(
        n6509) );
  OAI22_X1 U20042 ( .A1(n27415), .A2(n26990), .B1(n26984), .B2(n22527), .ZN(
        n6510) );
  OAI22_X1 U20043 ( .A1(n27418), .A2(n26990), .B1(n26984), .B2(n22526), .ZN(
        n6511) );
  OAI22_X1 U20044 ( .A1(n27421), .A2(n26990), .B1(n26984), .B2(n22525), .ZN(
        n6512) );
  OAI22_X1 U20045 ( .A1(n27424), .A2(n26991), .B1(n26984), .B2(n22524), .ZN(
        n6513) );
  OAI22_X1 U20046 ( .A1(n27427), .A2(n26991), .B1(n26985), .B2(n22523), .ZN(
        n6514) );
  OAI22_X1 U20047 ( .A1(n27430), .A2(n26991), .B1(n26985), .B2(n22522), .ZN(
        n6515) );
  OAI22_X1 U20048 ( .A1(n27433), .A2(n26991), .B1(n26985), .B2(n22521), .ZN(
        n6516) );
  OAI22_X1 U20049 ( .A1(n27436), .A2(n26991), .B1(n26985), .B2(n22520), .ZN(
        n6517) );
  OAI22_X1 U20050 ( .A1(n27439), .A2(n26991), .B1(n26985), .B2(n22519), .ZN(
        n6518) );
  OAI22_X1 U20051 ( .A1(n27442), .A2(n26991), .B1(n26985), .B2(n22518), .ZN(
        n6519) );
  OAI22_X1 U20052 ( .A1(n27445), .A2(n26991), .B1(n26985), .B2(n22517), .ZN(
        n6520) );
  OAI22_X1 U20053 ( .A1(n27448), .A2(n26991), .B1(n26985), .B2(n22516), .ZN(
        n6521) );
  OAI22_X1 U20054 ( .A1(n27451), .A2(n26991), .B1(n26985), .B2(n22515), .ZN(
        n6522) );
  OAI22_X1 U20055 ( .A1(n27454), .A2(n26991), .B1(n26985), .B2(n22514), .ZN(
        n6523) );
  OAI22_X1 U20056 ( .A1(n27457), .A2(n26991), .B1(n26985), .B2(n22513), .ZN(
        n6524) );
  OAI22_X1 U20057 ( .A1(n27460), .A2(n26992), .B1(n26985), .B2(n22512), .ZN(
        n6525) );
  OAI22_X1 U20058 ( .A1(n27318), .A2(n27180), .B1(n27174), .B2(n22487), .ZN(
        n7502) );
  OAI22_X1 U20059 ( .A1(n27321), .A2(n27180), .B1(n27174), .B2(n22486), .ZN(
        n7503) );
  OAI22_X1 U20060 ( .A1(n27324), .A2(n27180), .B1(n27174), .B2(n22485), .ZN(
        n7504) );
  OAI22_X1 U20061 ( .A1(n27327), .A2(n27180), .B1(n27174), .B2(n22484), .ZN(
        n7505) );
  OAI22_X1 U20062 ( .A1(n27330), .A2(n27180), .B1(n27174), .B2(n22483), .ZN(
        n7506) );
  OAI22_X1 U20063 ( .A1(n27333), .A2(n27180), .B1(n27174), .B2(n22482), .ZN(
        n7507) );
  OAI22_X1 U20064 ( .A1(n27336), .A2(n27180), .B1(n27174), .B2(n22481), .ZN(
        n7508) );
  OAI22_X1 U20065 ( .A1(n27339), .A2(n27180), .B1(n27174), .B2(n22480), .ZN(
        n7509) );
  OAI22_X1 U20066 ( .A1(n27342), .A2(n27180), .B1(n27174), .B2(n22479), .ZN(
        n7510) );
  OAI22_X1 U20067 ( .A1(n27345), .A2(n27180), .B1(n27174), .B2(n22478), .ZN(
        n7511) );
  OAI22_X1 U20068 ( .A1(n27348), .A2(n27180), .B1(n27174), .B2(n22477), .ZN(
        n7512) );
  OAI22_X1 U20069 ( .A1(n27351), .A2(n27181), .B1(n27174), .B2(n22476), .ZN(
        n7513) );
  OAI22_X1 U20070 ( .A1(n27354), .A2(n27181), .B1(n27175), .B2(n22475), .ZN(
        n7514) );
  OAI22_X1 U20071 ( .A1(n27357), .A2(n27181), .B1(n27175), .B2(n22474), .ZN(
        n7515) );
  OAI22_X1 U20072 ( .A1(n27360), .A2(n27181), .B1(n27175), .B2(n22473), .ZN(
        n7516) );
  OAI22_X1 U20073 ( .A1(n27363), .A2(n27181), .B1(n27175), .B2(n22472), .ZN(
        n7517) );
  OAI22_X1 U20074 ( .A1(n27366), .A2(n27181), .B1(n27175), .B2(n22471), .ZN(
        n7518) );
  OAI22_X1 U20075 ( .A1(n27369), .A2(n27181), .B1(n27175), .B2(n22470), .ZN(
        n7519) );
  OAI22_X1 U20076 ( .A1(n27372), .A2(n27181), .B1(n27175), .B2(n22469), .ZN(
        n7520) );
  OAI22_X1 U20077 ( .A1(n27375), .A2(n27181), .B1(n27175), .B2(n22468), .ZN(
        n7521) );
  OAI22_X1 U20078 ( .A1(n27378), .A2(n27181), .B1(n27175), .B2(n22467), .ZN(
        n7522) );
  OAI22_X1 U20079 ( .A1(n27381), .A2(n27181), .B1(n27175), .B2(n22466), .ZN(
        n7523) );
  OAI22_X1 U20080 ( .A1(n27384), .A2(n27181), .B1(n27175), .B2(n22465), .ZN(
        n7524) );
  OAI22_X1 U20081 ( .A1(n27387), .A2(n27182), .B1(n27175), .B2(n22464), .ZN(
        n7525) );
  OAI22_X1 U20082 ( .A1(n27390), .A2(n27182), .B1(n27176), .B2(n22463), .ZN(
        n7526) );
  OAI22_X1 U20083 ( .A1(n27393), .A2(n27182), .B1(n27176), .B2(n22462), .ZN(
        n7527) );
  OAI22_X1 U20084 ( .A1(n27396), .A2(n27182), .B1(n27176), .B2(n22461), .ZN(
        n7528) );
  OAI22_X1 U20085 ( .A1(n27399), .A2(n27182), .B1(n27176), .B2(n22460), .ZN(
        n7529) );
  OAI22_X1 U20086 ( .A1(n27402), .A2(n27182), .B1(n27176), .B2(n22459), .ZN(
        n7530) );
  OAI22_X1 U20087 ( .A1(n27405), .A2(n27182), .B1(n27176), .B2(n22458), .ZN(
        n7531) );
  OAI22_X1 U20088 ( .A1(n27408), .A2(n27182), .B1(n27176), .B2(n22457), .ZN(
        n7532) );
  OAI22_X1 U20089 ( .A1(n27411), .A2(n27182), .B1(n27176), .B2(n22456), .ZN(
        n7533) );
  OAI22_X1 U20090 ( .A1(n27414), .A2(n27182), .B1(n27176), .B2(n22455), .ZN(
        n7534) );
  OAI22_X1 U20091 ( .A1(n27417), .A2(n27182), .B1(n27176), .B2(n22454), .ZN(
        n7535) );
  OAI22_X1 U20092 ( .A1(n27420), .A2(n27182), .B1(n27176), .B2(n22453), .ZN(
        n7536) );
  OAI22_X1 U20093 ( .A1(n27423), .A2(n27183), .B1(n27176), .B2(n22452), .ZN(
        n7537) );
  OAI22_X1 U20094 ( .A1(n27426), .A2(n27183), .B1(n27177), .B2(n22451), .ZN(
        n7538) );
  OAI22_X1 U20095 ( .A1(n27429), .A2(n27183), .B1(n27177), .B2(n22450), .ZN(
        n7539) );
  OAI22_X1 U20096 ( .A1(n27432), .A2(n27183), .B1(n27177), .B2(n22449), .ZN(
        n7540) );
  OAI22_X1 U20097 ( .A1(n27435), .A2(n27183), .B1(n27177), .B2(n22448), .ZN(
        n7541) );
  OAI22_X1 U20098 ( .A1(n27438), .A2(n27183), .B1(n27177), .B2(n22447), .ZN(
        n7542) );
  OAI22_X1 U20099 ( .A1(n27441), .A2(n27183), .B1(n27177), .B2(n22446), .ZN(
        n7543) );
  OAI22_X1 U20100 ( .A1(n27444), .A2(n27183), .B1(n27177), .B2(n22445), .ZN(
        n7544) );
  OAI22_X1 U20101 ( .A1(n27447), .A2(n27183), .B1(n27177), .B2(n22444), .ZN(
        n7545) );
  OAI22_X1 U20102 ( .A1(n27450), .A2(n27183), .B1(n27177), .B2(n22443), .ZN(
        n7546) );
  OAI22_X1 U20103 ( .A1(n27453), .A2(n27183), .B1(n27177), .B2(n22442), .ZN(
        n7547) );
  OAI22_X1 U20104 ( .A1(n27456), .A2(n27183), .B1(n27177), .B2(n22441), .ZN(
        n7548) );
  OAI22_X1 U20105 ( .A1(n27459), .A2(n27184), .B1(n27177), .B2(n22440), .ZN(
        n7549) );
  OAI22_X1 U20106 ( .A1(n27319), .A2(n27048), .B1(n27042), .B2(n22367), .ZN(
        n6798) );
  OAI22_X1 U20107 ( .A1(n27322), .A2(n27048), .B1(n27042), .B2(n22366), .ZN(
        n6799) );
  OAI22_X1 U20108 ( .A1(n27325), .A2(n27048), .B1(n27042), .B2(n22365), .ZN(
        n6800) );
  OAI22_X1 U20109 ( .A1(n27328), .A2(n27048), .B1(n27042), .B2(n22364), .ZN(
        n6801) );
  OAI22_X1 U20110 ( .A1(n27331), .A2(n27048), .B1(n27042), .B2(n22363), .ZN(
        n6802) );
  OAI22_X1 U20111 ( .A1(n27334), .A2(n27048), .B1(n27042), .B2(n22362), .ZN(
        n6803) );
  OAI22_X1 U20112 ( .A1(n27337), .A2(n27048), .B1(n27042), .B2(n22361), .ZN(
        n6804) );
  OAI22_X1 U20113 ( .A1(n27340), .A2(n27048), .B1(n27042), .B2(n22360), .ZN(
        n6805) );
  OAI22_X1 U20114 ( .A1(n27343), .A2(n27048), .B1(n27042), .B2(n22359), .ZN(
        n6806) );
  OAI22_X1 U20115 ( .A1(n27346), .A2(n27048), .B1(n27042), .B2(n22358), .ZN(
        n6807) );
  OAI22_X1 U20116 ( .A1(n27349), .A2(n27048), .B1(n27042), .B2(n22357), .ZN(
        n6808) );
  OAI22_X1 U20117 ( .A1(n27352), .A2(n27049), .B1(n27042), .B2(n22356), .ZN(
        n6809) );
  OAI22_X1 U20118 ( .A1(n27355), .A2(n27049), .B1(n27043), .B2(n22355), .ZN(
        n6810) );
  OAI22_X1 U20119 ( .A1(n27358), .A2(n27049), .B1(n27043), .B2(n22354), .ZN(
        n6811) );
  OAI22_X1 U20120 ( .A1(n27361), .A2(n27049), .B1(n27043), .B2(n22353), .ZN(
        n6812) );
  OAI22_X1 U20121 ( .A1(n27364), .A2(n27049), .B1(n27043), .B2(n22352), .ZN(
        n6813) );
  OAI22_X1 U20122 ( .A1(n27367), .A2(n27049), .B1(n27043), .B2(n22351), .ZN(
        n6814) );
  OAI22_X1 U20123 ( .A1(n27370), .A2(n27049), .B1(n27043), .B2(n22350), .ZN(
        n6815) );
  OAI22_X1 U20124 ( .A1(n27373), .A2(n27049), .B1(n27043), .B2(n22349), .ZN(
        n6816) );
  OAI22_X1 U20125 ( .A1(n27376), .A2(n27049), .B1(n27043), .B2(n22348), .ZN(
        n6817) );
  OAI22_X1 U20126 ( .A1(n27379), .A2(n27049), .B1(n27043), .B2(n22347), .ZN(
        n6818) );
  OAI22_X1 U20127 ( .A1(n27382), .A2(n27049), .B1(n27043), .B2(n22346), .ZN(
        n6819) );
  OAI22_X1 U20128 ( .A1(n27385), .A2(n27049), .B1(n27043), .B2(n22345), .ZN(
        n6820) );
  OAI22_X1 U20129 ( .A1(n27388), .A2(n27050), .B1(n27043), .B2(n22344), .ZN(
        n6821) );
  OAI22_X1 U20130 ( .A1(n27391), .A2(n27050), .B1(n27044), .B2(n22343), .ZN(
        n6822) );
  OAI22_X1 U20131 ( .A1(n27394), .A2(n27050), .B1(n27044), .B2(n22342), .ZN(
        n6823) );
  OAI22_X1 U20132 ( .A1(n27397), .A2(n27050), .B1(n27044), .B2(n22341), .ZN(
        n6824) );
  OAI22_X1 U20133 ( .A1(n27400), .A2(n27050), .B1(n27044), .B2(n22340), .ZN(
        n6825) );
  OAI22_X1 U20134 ( .A1(n27403), .A2(n27050), .B1(n27044), .B2(n22339), .ZN(
        n6826) );
  OAI22_X1 U20135 ( .A1(n27406), .A2(n27050), .B1(n27044), .B2(n22338), .ZN(
        n6827) );
  OAI22_X1 U20136 ( .A1(n27409), .A2(n27050), .B1(n27044), .B2(n22337), .ZN(
        n6828) );
  OAI22_X1 U20137 ( .A1(n27412), .A2(n27050), .B1(n27044), .B2(n22336), .ZN(
        n6829) );
  OAI22_X1 U20138 ( .A1(n27415), .A2(n27050), .B1(n27044), .B2(n22335), .ZN(
        n6830) );
  OAI22_X1 U20139 ( .A1(n27418), .A2(n27050), .B1(n27044), .B2(n22334), .ZN(
        n6831) );
  OAI22_X1 U20140 ( .A1(n27421), .A2(n27050), .B1(n27044), .B2(n22333), .ZN(
        n6832) );
  OAI22_X1 U20141 ( .A1(n27424), .A2(n27051), .B1(n27044), .B2(n22332), .ZN(
        n6833) );
  OAI22_X1 U20142 ( .A1(n27427), .A2(n27051), .B1(n27045), .B2(n22331), .ZN(
        n6834) );
  OAI22_X1 U20143 ( .A1(n27430), .A2(n27051), .B1(n27045), .B2(n22330), .ZN(
        n6835) );
  OAI22_X1 U20144 ( .A1(n27433), .A2(n27051), .B1(n27045), .B2(n22329), .ZN(
        n6836) );
  OAI22_X1 U20145 ( .A1(n27436), .A2(n27051), .B1(n27045), .B2(n22328), .ZN(
        n6837) );
  OAI22_X1 U20146 ( .A1(n27439), .A2(n27051), .B1(n27045), .B2(n22327), .ZN(
        n6838) );
  OAI22_X1 U20147 ( .A1(n27442), .A2(n27051), .B1(n27045), .B2(n22326), .ZN(
        n6839) );
  OAI22_X1 U20148 ( .A1(n27445), .A2(n27051), .B1(n27045), .B2(n22325), .ZN(
        n6840) );
  OAI22_X1 U20149 ( .A1(n27448), .A2(n27051), .B1(n27045), .B2(n22324), .ZN(
        n6841) );
  OAI22_X1 U20150 ( .A1(n27451), .A2(n27051), .B1(n27045), .B2(n22323), .ZN(
        n6842) );
  OAI22_X1 U20151 ( .A1(n27454), .A2(n27051), .B1(n27045), .B2(n22322), .ZN(
        n6843) );
  OAI22_X1 U20152 ( .A1(n27457), .A2(n27051), .B1(n27045), .B2(n22321), .ZN(
        n6844) );
  OAI22_X1 U20153 ( .A1(n27460), .A2(n27052), .B1(n27045), .B2(n22320), .ZN(
        n6845) );
  OAI22_X1 U20154 ( .A1(n27318), .A2(n27192), .B1(n27186), .B2(n22047), .ZN(
        n7566) );
  OAI22_X1 U20155 ( .A1(n27321), .A2(n27192), .B1(n27186), .B2(n22046), .ZN(
        n7567) );
  OAI22_X1 U20156 ( .A1(n27324), .A2(n27192), .B1(n27186), .B2(n22045), .ZN(
        n7568) );
  OAI22_X1 U20157 ( .A1(n27327), .A2(n27192), .B1(n27186), .B2(n22044), .ZN(
        n7569) );
  OAI22_X1 U20158 ( .A1(n27330), .A2(n27192), .B1(n27186), .B2(n22043), .ZN(
        n7570) );
  OAI22_X1 U20159 ( .A1(n27333), .A2(n27192), .B1(n27186), .B2(n22042), .ZN(
        n7571) );
  OAI22_X1 U20160 ( .A1(n27336), .A2(n27192), .B1(n27186), .B2(n22041), .ZN(
        n7572) );
  OAI22_X1 U20161 ( .A1(n27339), .A2(n27192), .B1(n27186), .B2(n22040), .ZN(
        n7573) );
  OAI22_X1 U20162 ( .A1(n27342), .A2(n27192), .B1(n27186), .B2(n22039), .ZN(
        n7574) );
  OAI22_X1 U20163 ( .A1(n27345), .A2(n27192), .B1(n27186), .B2(n22038), .ZN(
        n7575) );
  OAI22_X1 U20164 ( .A1(n27348), .A2(n27192), .B1(n27186), .B2(n22037), .ZN(
        n7576) );
  OAI22_X1 U20165 ( .A1(n27351), .A2(n27193), .B1(n27186), .B2(n22036), .ZN(
        n7577) );
  OAI22_X1 U20166 ( .A1(n27354), .A2(n27193), .B1(n27187), .B2(n22035), .ZN(
        n7578) );
  OAI22_X1 U20167 ( .A1(n27357), .A2(n27193), .B1(n27187), .B2(n22034), .ZN(
        n7579) );
  OAI22_X1 U20168 ( .A1(n27360), .A2(n27193), .B1(n27187), .B2(n22033), .ZN(
        n7580) );
  OAI22_X1 U20169 ( .A1(n27363), .A2(n27193), .B1(n27187), .B2(n22032), .ZN(
        n7581) );
  OAI22_X1 U20170 ( .A1(n27366), .A2(n27193), .B1(n27187), .B2(n22031), .ZN(
        n7582) );
  OAI22_X1 U20171 ( .A1(n27369), .A2(n27193), .B1(n27187), .B2(n22030), .ZN(
        n7583) );
  OAI22_X1 U20172 ( .A1(n27372), .A2(n27193), .B1(n27187), .B2(n22029), .ZN(
        n7584) );
  OAI22_X1 U20173 ( .A1(n27375), .A2(n27193), .B1(n27187), .B2(n22028), .ZN(
        n7585) );
  OAI22_X1 U20174 ( .A1(n27378), .A2(n27193), .B1(n27187), .B2(n22027), .ZN(
        n7586) );
  OAI22_X1 U20175 ( .A1(n27381), .A2(n27193), .B1(n27187), .B2(n22026), .ZN(
        n7587) );
  OAI22_X1 U20176 ( .A1(n27384), .A2(n27193), .B1(n27187), .B2(n22025), .ZN(
        n7588) );
  OAI22_X1 U20177 ( .A1(n27387), .A2(n27194), .B1(n27187), .B2(n22024), .ZN(
        n7589) );
  OAI22_X1 U20178 ( .A1(n27390), .A2(n27194), .B1(n27188), .B2(n22023), .ZN(
        n7590) );
  OAI22_X1 U20179 ( .A1(n27393), .A2(n27194), .B1(n27188), .B2(n22022), .ZN(
        n7591) );
  OAI22_X1 U20180 ( .A1(n27396), .A2(n27194), .B1(n27188), .B2(n22021), .ZN(
        n7592) );
  OAI22_X1 U20181 ( .A1(n27399), .A2(n27194), .B1(n27188), .B2(n22020), .ZN(
        n7593) );
  OAI22_X1 U20182 ( .A1(n27402), .A2(n27194), .B1(n27188), .B2(n22019), .ZN(
        n7594) );
  OAI22_X1 U20183 ( .A1(n27405), .A2(n27194), .B1(n27188), .B2(n22018), .ZN(
        n7595) );
  OAI22_X1 U20184 ( .A1(n27408), .A2(n27194), .B1(n27188), .B2(n22017), .ZN(
        n7596) );
  OAI22_X1 U20185 ( .A1(n27411), .A2(n27194), .B1(n27188), .B2(n22016), .ZN(
        n7597) );
  OAI22_X1 U20186 ( .A1(n27414), .A2(n27194), .B1(n27188), .B2(n22015), .ZN(
        n7598) );
  OAI22_X1 U20187 ( .A1(n27417), .A2(n27194), .B1(n27188), .B2(n22014), .ZN(
        n7599) );
  OAI22_X1 U20188 ( .A1(n27420), .A2(n27194), .B1(n27188), .B2(n22013), .ZN(
        n7600) );
  OAI22_X1 U20189 ( .A1(n27423), .A2(n27195), .B1(n27188), .B2(n22012), .ZN(
        n7601) );
  OAI22_X1 U20190 ( .A1(n27426), .A2(n27195), .B1(n27189), .B2(n22011), .ZN(
        n7602) );
  OAI22_X1 U20191 ( .A1(n27429), .A2(n27195), .B1(n27189), .B2(n22010), .ZN(
        n7603) );
  OAI22_X1 U20192 ( .A1(n27432), .A2(n27195), .B1(n27189), .B2(n22009), .ZN(
        n7604) );
  OAI22_X1 U20193 ( .A1(n27435), .A2(n27195), .B1(n27189), .B2(n22008), .ZN(
        n7605) );
  OAI22_X1 U20194 ( .A1(n27438), .A2(n27195), .B1(n27189), .B2(n22007), .ZN(
        n7606) );
  OAI22_X1 U20195 ( .A1(n27441), .A2(n27195), .B1(n27189), .B2(n22006), .ZN(
        n7607) );
  OAI22_X1 U20196 ( .A1(n27444), .A2(n27195), .B1(n27189), .B2(n22005), .ZN(
        n7608) );
  OAI22_X1 U20197 ( .A1(n27447), .A2(n27195), .B1(n27189), .B2(n22004), .ZN(
        n7609) );
  OAI22_X1 U20198 ( .A1(n27450), .A2(n27195), .B1(n27189), .B2(n22003), .ZN(
        n7610) );
  OAI22_X1 U20199 ( .A1(n27453), .A2(n27195), .B1(n27189), .B2(n22002), .ZN(
        n7611) );
  OAI22_X1 U20200 ( .A1(n27456), .A2(n27195), .B1(n27189), .B2(n22001), .ZN(
        n7612) );
  OAI22_X1 U20201 ( .A1(n27459), .A2(n27196), .B1(n27189), .B2(n22000), .ZN(
        n7613) );
  OAI22_X1 U20202 ( .A1(n27318), .A2(n27144), .B1(n27138), .B2(n21987), .ZN(
        n7310) );
  OAI22_X1 U20203 ( .A1(n27321), .A2(n27144), .B1(n27138), .B2(n21986), .ZN(
        n7311) );
  OAI22_X1 U20204 ( .A1(n27324), .A2(n27144), .B1(n27138), .B2(n21985), .ZN(
        n7312) );
  OAI22_X1 U20205 ( .A1(n27327), .A2(n27144), .B1(n27138), .B2(n21984), .ZN(
        n7313) );
  OAI22_X1 U20206 ( .A1(n27330), .A2(n27144), .B1(n27138), .B2(n21983), .ZN(
        n7314) );
  OAI22_X1 U20207 ( .A1(n27333), .A2(n27144), .B1(n27138), .B2(n21982), .ZN(
        n7315) );
  OAI22_X1 U20208 ( .A1(n27336), .A2(n27144), .B1(n27138), .B2(n21981), .ZN(
        n7316) );
  OAI22_X1 U20209 ( .A1(n27339), .A2(n27144), .B1(n27138), .B2(n21980), .ZN(
        n7317) );
  OAI22_X1 U20210 ( .A1(n27342), .A2(n27144), .B1(n27138), .B2(n21979), .ZN(
        n7318) );
  OAI22_X1 U20211 ( .A1(n27345), .A2(n27144), .B1(n27138), .B2(n21978), .ZN(
        n7319) );
  OAI22_X1 U20212 ( .A1(n27348), .A2(n27144), .B1(n27138), .B2(n21977), .ZN(
        n7320) );
  OAI22_X1 U20213 ( .A1(n27351), .A2(n27145), .B1(n27138), .B2(n21976), .ZN(
        n7321) );
  OAI22_X1 U20214 ( .A1(n27354), .A2(n27145), .B1(n27139), .B2(n21975), .ZN(
        n7322) );
  OAI22_X1 U20215 ( .A1(n27357), .A2(n27145), .B1(n27139), .B2(n21974), .ZN(
        n7323) );
  OAI22_X1 U20216 ( .A1(n27360), .A2(n27145), .B1(n27139), .B2(n21973), .ZN(
        n7324) );
  OAI22_X1 U20217 ( .A1(n27363), .A2(n27145), .B1(n27139), .B2(n21972), .ZN(
        n7325) );
  OAI22_X1 U20218 ( .A1(n27366), .A2(n27145), .B1(n27139), .B2(n21971), .ZN(
        n7326) );
  OAI22_X1 U20219 ( .A1(n27369), .A2(n27145), .B1(n27139), .B2(n21970), .ZN(
        n7327) );
  OAI22_X1 U20220 ( .A1(n27372), .A2(n27145), .B1(n27139), .B2(n21969), .ZN(
        n7328) );
  OAI22_X1 U20221 ( .A1(n27375), .A2(n27145), .B1(n27139), .B2(n21968), .ZN(
        n7329) );
  OAI22_X1 U20222 ( .A1(n27378), .A2(n27145), .B1(n27139), .B2(n21967), .ZN(
        n7330) );
  OAI22_X1 U20223 ( .A1(n27381), .A2(n27145), .B1(n27139), .B2(n21966), .ZN(
        n7331) );
  OAI22_X1 U20224 ( .A1(n27384), .A2(n27145), .B1(n27139), .B2(n21965), .ZN(
        n7332) );
  OAI22_X1 U20225 ( .A1(n27387), .A2(n27146), .B1(n27139), .B2(n21964), .ZN(
        n7333) );
  OAI22_X1 U20226 ( .A1(n27390), .A2(n27146), .B1(n27140), .B2(n21963), .ZN(
        n7334) );
  OAI22_X1 U20227 ( .A1(n27393), .A2(n27146), .B1(n27140), .B2(n21962), .ZN(
        n7335) );
  OAI22_X1 U20228 ( .A1(n27396), .A2(n27146), .B1(n27140), .B2(n21961), .ZN(
        n7336) );
  OAI22_X1 U20229 ( .A1(n27399), .A2(n27146), .B1(n27140), .B2(n21960), .ZN(
        n7337) );
  OAI22_X1 U20230 ( .A1(n27402), .A2(n27146), .B1(n27140), .B2(n21959), .ZN(
        n7338) );
  OAI22_X1 U20231 ( .A1(n27405), .A2(n27146), .B1(n27140), .B2(n21958), .ZN(
        n7339) );
  OAI22_X1 U20232 ( .A1(n27408), .A2(n27146), .B1(n27140), .B2(n21957), .ZN(
        n7340) );
  OAI22_X1 U20233 ( .A1(n27411), .A2(n27146), .B1(n27140), .B2(n21956), .ZN(
        n7341) );
  OAI22_X1 U20234 ( .A1(n27414), .A2(n27146), .B1(n27140), .B2(n21955), .ZN(
        n7342) );
  OAI22_X1 U20235 ( .A1(n27417), .A2(n27146), .B1(n27140), .B2(n21954), .ZN(
        n7343) );
  OAI22_X1 U20236 ( .A1(n27420), .A2(n27146), .B1(n27140), .B2(n21953), .ZN(
        n7344) );
  OAI22_X1 U20237 ( .A1(n27423), .A2(n27147), .B1(n27140), .B2(n21952), .ZN(
        n7345) );
  OAI22_X1 U20238 ( .A1(n27426), .A2(n27147), .B1(n27141), .B2(n21951), .ZN(
        n7346) );
  OAI22_X1 U20239 ( .A1(n27429), .A2(n27147), .B1(n27141), .B2(n21950), .ZN(
        n7347) );
  OAI22_X1 U20240 ( .A1(n27432), .A2(n27147), .B1(n27141), .B2(n21949), .ZN(
        n7348) );
  OAI22_X1 U20241 ( .A1(n27435), .A2(n27147), .B1(n27141), .B2(n21948), .ZN(
        n7349) );
  OAI22_X1 U20242 ( .A1(n27438), .A2(n27147), .B1(n27141), .B2(n21947), .ZN(
        n7350) );
  OAI22_X1 U20243 ( .A1(n27441), .A2(n27147), .B1(n27141), .B2(n21946), .ZN(
        n7351) );
  OAI22_X1 U20244 ( .A1(n27444), .A2(n27147), .B1(n27141), .B2(n21945), .ZN(
        n7352) );
  OAI22_X1 U20245 ( .A1(n27447), .A2(n27147), .B1(n27141), .B2(n21944), .ZN(
        n7353) );
  OAI22_X1 U20246 ( .A1(n27450), .A2(n27147), .B1(n27141), .B2(n21943), .ZN(
        n7354) );
  OAI22_X1 U20247 ( .A1(n27453), .A2(n27147), .B1(n27141), .B2(n21942), .ZN(
        n7355) );
  OAI22_X1 U20248 ( .A1(n27456), .A2(n27147), .B1(n27141), .B2(n21941), .ZN(
        n7356) );
  OAI22_X1 U20249 ( .A1(n27459), .A2(n27148), .B1(n27141), .B2(n21940), .ZN(
        n7357) );
  OAI22_X1 U20250 ( .A1(n27319), .A2(n27072), .B1(n27066), .B2(n21747), .ZN(
        n6926) );
  OAI22_X1 U20251 ( .A1(n27322), .A2(n27072), .B1(n27066), .B2(n21746), .ZN(
        n6927) );
  OAI22_X1 U20252 ( .A1(n27325), .A2(n27072), .B1(n27066), .B2(n21745), .ZN(
        n6928) );
  OAI22_X1 U20253 ( .A1(n27328), .A2(n27072), .B1(n27066), .B2(n21744), .ZN(
        n6929) );
  OAI22_X1 U20254 ( .A1(n27331), .A2(n27072), .B1(n27066), .B2(n21743), .ZN(
        n6930) );
  OAI22_X1 U20255 ( .A1(n27334), .A2(n27072), .B1(n27066), .B2(n21742), .ZN(
        n6931) );
  OAI22_X1 U20256 ( .A1(n27337), .A2(n27072), .B1(n27066), .B2(n21741), .ZN(
        n6932) );
  OAI22_X1 U20257 ( .A1(n27340), .A2(n27072), .B1(n27066), .B2(n21740), .ZN(
        n6933) );
  OAI22_X1 U20258 ( .A1(n27343), .A2(n27072), .B1(n27066), .B2(n21739), .ZN(
        n6934) );
  OAI22_X1 U20259 ( .A1(n27346), .A2(n27072), .B1(n27066), .B2(n21738), .ZN(
        n6935) );
  OAI22_X1 U20260 ( .A1(n27349), .A2(n27072), .B1(n27066), .B2(n21737), .ZN(
        n6936) );
  OAI22_X1 U20261 ( .A1(n27352), .A2(n27073), .B1(n27066), .B2(n21736), .ZN(
        n6937) );
  OAI22_X1 U20262 ( .A1(n27355), .A2(n27073), .B1(n27067), .B2(n21735), .ZN(
        n6938) );
  OAI22_X1 U20263 ( .A1(n27358), .A2(n27073), .B1(n27067), .B2(n21734), .ZN(
        n6939) );
  OAI22_X1 U20264 ( .A1(n27361), .A2(n27073), .B1(n27067), .B2(n21733), .ZN(
        n6940) );
  OAI22_X1 U20265 ( .A1(n27364), .A2(n27073), .B1(n27067), .B2(n21732), .ZN(
        n6941) );
  OAI22_X1 U20266 ( .A1(n27367), .A2(n27073), .B1(n27067), .B2(n21731), .ZN(
        n6942) );
  OAI22_X1 U20267 ( .A1(n27370), .A2(n27073), .B1(n27067), .B2(n21730), .ZN(
        n6943) );
  OAI22_X1 U20268 ( .A1(n27373), .A2(n27073), .B1(n27067), .B2(n21729), .ZN(
        n6944) );
  OAI22_X1 U20269 ( .A1(n27376), .A2(n27073), .B1(n27067), .B2(n21728), .ZN(
        n6945) );
  OAI22_X1 U20270 ( .A1(n27379), .A2(n27073), .B1(n27067), .B2(n21727), .ZN(
        n6946) );
  OAI22_X1 U20271 ( .A1(n27382), .A2(n27073), .B1(n27067), .B2(n21726), .ZN(
        n6947) );
  OAI22_X1 U20272 ( .A1(n27385), .A2(n27073), .B1(n27067), .B2(n21725), .ZN(
        n6948) );
  OAI22_X1 U20273 ( .A1(n27388), .A2(n27074), .B1(n27067), .B2(n21724), .ZN(
        n6949) );
  OAI22_X1 U20274 ( .A1(n27391), .A2(n27074), .B1(n27068), .B2(n21723), .ZN(
        n6950) );
  OAI22_X1 U20275 ( .A1(n27394), .A2(n27074), .B1(n27068), .B2(n21722), .ZN(
        n6951) );
  OAI22_X1 U20276 ( .A1(n27397), .A2(n27074), .B1(n27068), .B2(n21721), .ZN(
        n6952) );
  OAI22_X1 U20277 ( .A1(n27400), .A2(n27074), .B1(n27068), .B2(n21720), .ZN(
        n6953) );
  OAI22_X1 U20278 ( .A1(n27403), .A2(n27074), .B1(n27068), .B2(n21719), .ZN(
        n6954) );
  OAI22_X1 U20279 ( .A1(n27406), .A2(n27074), .B1(n27068), .B2(n21718), .ZN(
        n6955) );
  OAI22_X1 U20280 ( .A1(n27409), .A2(n27074), .B1(n27068), .B2(n21717), .ZN(
        n6956) );
  OAI22_X1 U20281 ( .A1(n27412), .A2(n27074), .B1(n27068), .B2(n21716), .ZN(
        n6957) );
  OAI22_X1 U20282 ( .A1(n27415), .A2(n27074), .B1(n27068), .B2(n21715), .ZN(
        n6958) );
  OAI22_X1 U20283 ( .A1(n27418), .A2(n27074), .B1(n27068), .B2(n21714), .ZN(
        n6959) );
  OAI22_X1 U20284 ( .A1(n27421), .A2(n27074), .B1(n27068), .B2(n21713), .ZN(
        n6960) );
  OAI22_X1 U20285 ( .A1(n27424), .A2(n27075), .B1(n27068), .B2(n21712), .ZN(
        n6961) );
  OAI22_X1 U20286 ( .A1(n27427), .A2(n27075), .B1(n27069), .B2(n21711), .ZN(
        n6962) );
  OAI22_X1 U20287 ( .A1(n27430), .A2(n27075), .B1(n27069), .B2(n21710), .ZN(
        n6963) );
  OAI22_X1 U20288 ( .A1(n27433), .A2(n27075), .B1(n27069), .B2(n21709), .ZN(
        n6964) );
  OAI22_X1 U20289 ( .A1(n27436), .A2(n27075), .B1(n27069), .B2(n21708), .ZN(
        n6965) );
  OAI22_X1 U20290 ( .A1(n27439), .A2(n27075), .B1(n27069), .B2(n21707), .ZN(
        n6966) );
  OAI22_X1 U20291 ( .A1(n27442), .A2(n27075), .B1(n27069), .B2(n21706), .ZN(
        n6967) );
  OAI22_X1 U20292 ( .A1(n27445), .A2(n27075), .B1(n27069), .B2(n21705), .ZN(
        n6968) );
  OAI22_X1 U20293 ( .A1(n27448), .A2(n27075), .B1(n27069), .B2(n21704), .ZN(
        n6969) );
  OAI22_X1 U20294 ( .A1(n27451), .A2(n27075), .B1(n27069), .B2(n21703), .ZN(
        n6970) );
  OAI22_X1 U20295 ( .A1(n27454), .A2(n27075), .B1(n27069), .B2(n21702), .ZN(
        n6971) );
  OAI22_X1 U20296 ( .A1(n27457), .A2(n27075), .B1(n27069), .B2(n21701), .ZN(
        n6972) );
  OAI22_X1 U20297 ( .A1(n27460), .A2(n27076), .B1(n27069), .B2(n21700), .ZN(
        n6973) );
  OAI22_X1 U20298 ( .A1(n27320), .A2(n26964), .B1(n26958), .B2(n21627), .ZN(
        n6350) );
  OAI22_X1 U20299 ( .A1(n27323), .A2(n26964), .B1(n26958), .B2(n21626), .ZN(
        n6351) );
  OAI22_X1 U20300 ( .A1(n27326), .A2(n26964), .B1(n26958), .B2(n21625), .ZN(
        n6352) );
  OAI22_X1 U20301 ( .A1(n27329), .A2(n26964), .B1(n26958), .B2(n21624), .ZN(
        n6353) );
  OAI22_X1 U20302 ( .A1(n27332), .A2(n26964), .B1(n26958), .B2(n21623), .ZN(
        n6354) );
  OAI22_X1 U20303 ( .A1(n27335), .A2(n26964), .B1(n26958), .B2(n21622), .ZN(
        n6355) );
  OAI22_X1 U20304 ( .A1(n27338), .A2(n26964), .B1(n26958), .B2(n21621), .ZN(
        n6356) );
  OAI22_X1 U20305 ( .A1(n27341), .A2(n26964), .B1(n26958), .B2(n21620), .ZN(
        n6357) );
  OAI22_X1 U20306 ( .A1(n27344), .A2(n26964), .B1(n26958), .B2(n21619), .ZN(
        n6358) );
  OAI22_X1 U20307 ( .A1(n27347), .A2(n26964), .B1(n26958), .B2(n21618), .ZN(
        n6359) );
  OAI22_X1 U20308 ( .A1(n27350), .A2(n26964), .B1(n26958), .B2(n21617), .ZN(
        n6360) );
  OAI22_X1 U20309 ( .A1(n27353), .A2(n26965), .B1(n26958), .B2(n21616), .ZN(
        n6361) );
  OAI22_X1 U20310 ( .A1(n27356), .A2(n26965), .B1(n26959), .B2(n21615), .ZN(
        n6362) );
  OAI22_X1 U20311 ( .A1(n27359), .A2(n26965), .B1(n26959), .B2(n21614), .ZN(
        n6363) );
  OAI22_X1 U20312 ( .A1(n27362), .A2(n26965), .B1(n26959), .B2(n21613), .ZN(
        n6364) );
  OAI22_X1 U20313 ( .A1(n27365), .A2(n26965), .B1(n26959), .B2(n21612), .ZN(
        n6365) );
  OAI22_X1 U20314 ( .A1(n27368), .A2(n26965), .B1(n26959), .B2(n21611), .ZN(
        n6366) );
  OAI22_X1 U20315 ( .A1(n27371), .A2(n26965), .B1(n26959), .B2(n21610), .ZN(
        n6367) );
  OAI22_X1 U20316 ( .A1(n27374), .A2(n26965), .B1(n26959), .B2(n21609), .ZN(
        n6368) );
  OAI22_X1 U20317 ( .A1(n27377), .A2(n26965), .B1(n26959), .B2(n21608), .ZN(
        n6369) );
  OAI22_X1 U20318 ( .A1(n27380), .A2(n26965), .B1(n26959), .B2(n21607), .ZN(
        n6370) );
  OAI22_X1 U20319 ( .A1(n27383), .A2(n26965), .B1(n26959), .B2(n21606), .ZN(
        n6371) );
  OAI22_X1 U20320 ( .A1(n27386), .A2(n26965), .B1(n26959), .B2(n21605), .ZN(
        n6372) );
  OAI22_X1 U20321 ( .A1(n27389), .A2(n26966), .B1(n26959), .B2(n21604), .ZN(
        n6373) );
  OAI22_X1 U20322 ( .A1(n27392), .A2(n26966), .B1(n26960), .B2(n21603), .ZN(
        n6374) );
  OAI22_X1 U20323 ( .A1(n27395), .A2(n26966), .B1(n26960), .B2(n21602), .ZN(
        n6375) );
  OAI22_X1 U20324 ( .A1(n27398), .A2(n26966), .B1(n26960), .B2(n21601), .ZN(
        n6376) );
  OAI22_X1 U20325 ( .A1(n27401), .A2(n26966), .B1(n26960), .B2(n21600), .ZN(
        n6377) );
  OAI22_X1 U20326 ( .A1(n27404), .A2(n26966), .B1(n26960), .B2(n21599), .ZN(
        n6378) );
  OAI22_X1 U20327 ( .A1(n27407), .A2(n26966), .B1(n26960), .B2(n21598), .ZN(
        n6379) );
  OAI22_X1 U20328 ( .A1(n27410), .A2(n26966), .B1(n26960), .B2(n21597), .ZN(
        n6380) );
  OAI22_X1 U20329 ( .A1(n27413), .A2(n26966), .B1(n26960), .B2(n21596), .ZN(
        n6381) );
  OAI22_X1 U20330 ( .A1(n27416), .A2(n26966), .B1(n26960), .B2(n21595), .ZN(
        n6382) );
  OAI22_X1 U20331 ( .A1(n27419), .A2(n26966), .B1(n26960), .B2(n21594), .ZN(
        n6383) );
  OAI22_X1 U20332 ( .A1(n27422), .A2(n26966), .B1(n26960), .B2(n21593), .ZN(
        n6384) );
  OAI22_X1 U20333 ( .A1(n27425), .A2(n26967), .B1(n26960), .B2(n21592), .ZN(
        n6385) );
  OAI22_X1 U20334 ( .A1(n27428), .A2(n26967), .B1(n26961), .B2(n21591), .ZN(
        n6386) );
  OAI22_X1 U20335 ( .A1(n27431), .A2(n26967), .B1(n26961), .B2(n21590), .ZN(
        n6387) );
  OAI22_X1 U20336 ( .A1(n27434), .A2(n26967), .B1(n26961), .B2(n21589), .ZN(
        n6388) );
  OAI22_X1 U20337 ( .A1(n27437), .A2(n26967), .B1(n26961), .B2(n21588), .ZN(
        n6389) );
  OAI22_X1 U20338 ( .A1(n27440), .A2(n26967), .B1(n26961), .B2(n21587), .ZN(
        n6390) );
  OAI22_X1 U20339 ( .A1(n27443), .A2(n26967), .B1(n26961), .B2(n21586), .ZN(
        n6391) );
  OAI22_X1 U20340 ( .A1(n27446), .A2(n26967), .B1(n26961), .B2(n21585), .ZN(
        n6392) );
  OAI22_X1 U20341 ( .A1(n27449), .A2(n26967), .B1(n26961), .B2(n21584), .ZN(
        n6393) );
  OAI22_X1 U20342 ( .A1(n27452), .A2(n26967), .B1(n26961), .B2(n21583), .ZN(
        n6394) );
  OAI22_X1 U20343 ( .A1(n27455), .A2(n26967), .B1(n26961), .B2(n21582), .ZN(
        n6395) );
  OAI22_X1 U20344 ( .A1(n27458), .A2(n26967), .B1(n26961), .B2(n21581), .ZN(
        n6396) );
  OAI22_X1 U20345 ( .A1(n27461), .A2(n26968), .B1(n26961), .B2(n21580), .ZN(
        n6397) );
  OAI22_X1 U20346 ( .A1(n27318), .A2(n27216), .B1(n27210), .B2(n21567), .ZN(
        n7694) );
  OAI22_X1 U20347 ( .A1(n27321), .A2(n27216), .B1(n27210), .B2(n21566), .ZN(
        n7695) );
  OAI22_X1 U20348 ( .A1(n27324), .A2(n27216), .B1(n27210), .B2(n21565), .ZN(
        n7696) );
  OAI22_X1 U20349 ( .A1(n27327), .A2(n27216), .B1(n27210), .B2(n21564), .ZN(
        n7697) );
  OAI22_X1 U20350 ( .A1(n27330), .A2(n27216), .B1(n27210), .B2(n21563), .ZN(
        n7698) );
  OAI22_X1 U20351 ( .A1(n27333), .A2(n27216), .B1(n27210), .B2(n21562), .ZN(
        n7699) );
  OAI22_X1 U20352 ( .A1(n27336), .A2(n27216), .B1(n27210), .B2(n21561), .ZN(
        n7700) );
  OAI22_X1 U20353 ( .A1(n27339), .A2(n27216), .B1(n27210), .B2(n21560), .ZN(
        n7701) );
  OAI22_X1 U20354 ( .A1(n27342), .A2(n27216), .B1(n27210), .B2(n21559), .ZN(
        n7702) );
  OAI22_X1 U20355 ( .A1(n27345), .A2(n27216), .B1(n27210), .B2(n21558), .ZN(
        n7703) );
  OAI22_X1 U20356 ( .A1(n27348), .A2(n27216), .B1(n27210), .B2(n21557), .ZN(
        n7704) );
  OAI22_X1 U20357 ( .A1(n27351), .A2(n27217), .B1(n27210), .B2(n21556), .ZN(
        n7705) );
  OAI22_X1 U20358 ( .A1(n27354), .A2(n27217), .B1(n27211), .B2(n21555), .ZN(
        n7706) );
  OAI22_X1 U20359 ( .A1(n27357), .A2(n27217), .B1(n27211), .B2(n21554), .ZN(
        n7707) );
  OAI22_X1 U20360 ( .A1(n27360), .A2(n27217), .B1(n27211), .B2(n21553), .ZN(
        n7708) );
  OAI22_X1 U20361 ( .A1(n27363), .A2(n27217), .B1(n27211), .B2(n21552), .ZN(
        n7709) );
  OAI22_X1 U20362 ( .A1(n27366), .A2(n27217), .B1(n27211), .B2(n21551), .ZN(
        n7710) );
  OAI22_X1 U20363 ( .A1(n27369), .A2(n27217), .B1(n27211), .B2(n21550), .ZN(
        n7711) );
  OAI22_X1 U20364 ( .A1(n27372), .A2(n27217), .B1(n27211), .B2(n21549), .ZN(
        n7712) );
  OAI22_X1 U20365 ( .A1(n27375), .A2(n27217), .B1(n27211), .B2(n21548), .ZN(
        n7713) );
  OAI22_X1 U20366 ( .A1(n27378), .A2(n27217), .B1(n27211), .B2(n21547), .ZN(
        n7714) );
  OAI22_X1 U20367 ( .A1(n27381), .A2(n27217), .B1(n27211), .B2(n21546), .ZN(
        n7715) );
  OAI22_X1 U20368 ( .A1(n27384), .A2(n27217), .B1(n27211), .B2(n21545), .ZN(
        n7716) );
  OAI22_X1 U20369 ( .A1(n27387), .A2(n27218), .B1(n27211), .B2(n21544), .ZN(
        n7717) );
  OAI22_X1 U20370 ( .A1(n27390), .A2(n27218), .B1(n27212), .B2(n21543), .ZN(
        n7718) );
  OAI22_X1 U20371 ( .A1(n27393), .A2(n27218), .B1(n27212), .B2(n21542), .ZN(
        n7719) );
  OAI22_X1 U20372 ( .A1(n27396), .A2(n27218), .B1(n27212), .B2(n21541), .ZN(
        n7720) );
  OAI22_X1 U20373 ( .A1(n27399), .A2(n27218), .B1(n27212), .B2(n21540), .ZN(
        n7721) );
  OAI22_X1 U20374 ( .A1(n27402), .A2(n27218), .B1(n27212), .B2(n21539), .ZN(
        n7722) );
  OAI22_X1 U20375 ( .A1(n27405), .A2(n27218), .B1(n27212), .B2(n21538), .ZN(
        n7723) );
  OAI22_X1 U20376 ( .A1(n27408), .A2(n27218), .B1(n27212), .B2(n21537), .ZN(
        n7724) );
  OAI22_X1 U20377 ( .A1(n27411), .A2(n27218), .B1(n27212), .B2(n21536), .ZN(
        n7725) );
  OAI22_X1 U20378 ( .A1(n27414), .A2(n27218), .B1(n27212), .B2(n21535), .ZN(
        n7726) );
  OAI22_X1 U20379 ( .A1(n27417), .A2(n27218), .B1(n27212), .B2(n21534), .ZN(
        n7727) );
  OAI22_X1 U20380 ( .A1(n27420), .A2(n27218), .B1(n27212), .B2(n21533), .ZN(
        n7728) );
  OAI22_X1 U20381 ( .A1(n27423), .A2(n27219), .B1(n27212), .B2(n21532), .ZN(
        n7729) );
  OAI22_X1 U20382 ( .A1(n27426), .A2(n27219), .B1(n27213), .B2(n21531), .ZN(
        n7730) );
  OAI22_X1 U20383 ( .A1(n27429), .A2(n27219), .B1(n27213), .B2(n21530), .ZN(
        n7731) );
  OAI22_X1 U20384 ( .A1(n27432), .A2(n27219), .B1(n27213), .B2(n21529), .ZN(
        n7732) );
  OAI22_X1 U20385 ( .A1(n27435), .A2(n27219), .B1(n27213), .B2(n21528), .ZN(
        n7733) );
  OAI22_X1 U20386 ( .A1(n27438), .A2(n27219), .B1(n27213), .B2(n21527), .ZN(
        n7734) );
  OAI22_X1 U20387 ( .A1(n27441), .A2(n27219), .B1(n27213), .B2(n21526), .ZN(
        n7735) );
  OAI22_X1 U20388 ( .A1(n27444), .A2(n27219), .B1(n27213), .B2(n21525), .ZN(
        n7736) );
  OAI22_X1 U20389 ( .A1(n27447), .A2(n27219), .B1(n27213), .B2(n21524), .ZN(
        n7737) );
  OAI22_X1 U20390 ( .A1(n27450), .A2(n27219), .B1(n27213), .B2(n21523), .ZN(
        n7738) );
  OAI22_X1 U20391 ( .A1(n27453), .A2(n27219), .B1(n27213), .B2(n21522), .ZN(
        n7739) );
  OAI22_X1 U20392 ( .A1(n27456), .A2(n27219), .B1(n27213), .B2(n21521), .ZN(
        n7740) );
  OAI22_X1 U20393 ( .A1(n27459), .A2(n27220), .B1(n27213), .B2(n21520), .ZN(
        n7741) );
  OAI22_X1 U20394 ( .A1(n27318), .A2(n27240), .B1(n27234), .B2(n21407), .ZN(
        n7822) );
  OAI22_X1 U20395 ( .A1(n27321), .A2(n27240), .B1(n27234), .B2(n21406), .ZN(
        n7823) );
  OAI22_X1 U20396 ( .A1(n27324), .A2(n27240), .B1(n27234), .B2(n21405), .ZN(
        n7824) );
  OAI22_X1 U20397 ( .A1(n27327), .A2(n27240), .B1(n27234), .B2(n21404), .ZN(
        n7825) );
  OAI22_X1 U20398 ( .A1(n27330), .A2(n27240), .B1(n27234), .B2(n21403), .ZN(
        n7826) );
  OAI22_X1 U20399 ( .A1(n27333), .A2(n27240), .B1(n27234), .B2(n21402), .ZN(
        n7827) );
  OAI22_X1 U20400 ( .A1(n27336), .A2(n27240), .B1(n27234), .B2(n21401), .ZN(
        n7828) );
  OAI22_X1 U20401 ( .A1(n27339), .A2(n27240), .B1(n27234), .B2(n21400), .ZN(
        n7829) );
  OAI22_X1 U20402 ( .A1(n27342), .A2(n27240), .B1(n27234), .B2(n21399), .ZN(
        n7830) );
  OAI22_X1 U20403 ( .A1(n27345), .A2(n27240), .B1(n27234), .B2(n21398), .ZN(
        n7831) );
  OAI22_X1 U20404 ( .A1(n27348), .A2(n27240), .B1(n27234), .B2(n21397), .ZN(
        n7832) );
  OAI22_X1 U20405 ( .A1(n27351), .A2(n27241), .B1(n27234), .B2(n21396), .ZN(
        n7833) );
  OAI22_X1 U20406 ( .A1(n27354), .A2(n27241), .B1(n27235), .B2(n21395), .ZN(
        n7834) );
  OAI22_X1 U20407 ( .A1(n27357), .A2(n27241), .B1(n27235), .B2(n21394), .ZN(
        n7835) );
  OAI22_X1 U20408 ( .A1(n27360), .A2(n27241), .B1(n27235), .B2(n21393), .ZN(
        n7836) );
  OAI22_X1 U20409 ( .A1(n27363), .A2(n27241), .B1(n27235), .B2(n21392), .ZN(
        n7837) );
  OAI22_X1 U20410 ( .A1(n27366), .A2(n27241), .B1(n27235), .B2(n21391), .ZN(
        n7838) );
  OAI22_X1 U20411 ( .A1(n27369), .A2(n27241), .B1(n27235), .B2(n21390), .ZN(
        n7839) );
  OAI22_X1 U20412 ( .A1(n27372), .A2(n27241), .B1(n27235), .B2(n21389), .ZN(
        n7840) );
  OAI22_X1 U20413 ( .A1(n27375), .A2(n27241), .B1(n27235), .B2(n21388), .ZN(
        n7841) );
  OAI22_X1 U20414 ( .A1(n27378), .A2(n27241), .B1(n27235), .B2(n21387), .ZN(
        n7842) );
  OAI22_X1 U20415 ( .A1(n27381), .A2(n27241), .B1(n27235), .B2(n21386), .ZN(
        n7843) );
  OAI22_X1 U20416 ( .A1(n27384), .A2(n27241), .B1(n27235), .B2(n21385), .ZN(
        n7844) );
  OAI22_X1 U20417 ( .A1(n27387), .A2(n27242), .B1(n27235), .B2(n21384), .ZN(
        n7845) );
  OAI22_X1 U20418 ( .A1(n27390), .A2(n27242), .B1(n27236), .B2(n21383), .ZN(
        n7846) );
  OAI22_X1 U20419 ( .A1(n27393), .A2(n27242), .B1(n27236), .B2(n21382), .ZN(
        n7847) );
  OAI22_X1 U20420 ( .A1(n27396), .A2(n27242), .B1(n27236), .B2(n21381), .ZN(
        n7848) );
  OAI22_X1 U20421 ( .A1(n27399), .A2(n27242), .B1(n27236), .B2(n21380), .ZN(
        n7849) );
  OAI22_X1 U20422 ( .A1(n27402), .A2(n27242), .B1(n27236), .B2(n21379), .ZN(
        n7850) );
  OAI22_X1 U20423 ( .A1(n27405), .A2(n27242), .B1(n27236), .B2(n21378), .ZN(
        n7851) );
  OAI22_X1 U20424 ( .A1(n27408), .A2(n27242), .B1(n27236), .B2(n21377), .ZN(
        n7852) );
  OAI22_X1 U20425 ( .A1(n27411), .A2(n27242), .B1(n27236), .B2(n21376), .ZN(
        n7853) );
  OAI22_X1 U20426 ( .A1(n27414), .A2(n27242), .B1(n27236), .B2(n21375), .ZN(
        n7854) );
  OAI22_X1 U20427 ( .A1(n27417), .A2(n27242), .B1(n27236), .B2(n21374), .ZN(
        n7855) );
  OAI22_X1 U20428 ( .A1(n27420), .A2(n27242), .B1(n27236), .B2(n21373), .ZN(
        n7856) );
  OAI22_X1 U20429 ( .A1(n27423), .A2(n27243), .B1(n27236), .B2(n21372), .ZN(
        n7857) );
  OAI22_X1 U20430 ( .A1(n27426), .A2(n27243), .B1(n27237), .B2(n21371), .ZN(
        n7858) );
  OAI22_X1 U20431 ( .A1(n27429), .A2(n27243), .B1(n27237), .B2(n21370), .ZN(
        n7859) );
  OAI22_X1 U20432 ( .A1(n27432), .A2(n27243), .B1(n27237), .B2(n21369), .ZN(
        n7860) );
  OAI22_X1 U20433 ( .A1(n27435), .A2(n27243), .B1(n27237), .B2(n21368), .ZN(
        n7861) );
  OAI22_X1 U20434 ( .A1(n27438), .A2(n27243), .B1(n27237), .B2(n21367), .ZN(
        n7862) );
  OAI22_X1 U20435 ( .A1(n27441), .A2(n27243), .B1(n27237), .B2(n21366), .ZN(
        n7863) );
  OAI22_X1 U20436 ( .A1(n27444), .A2(n27243), .B1(n27237), .B2(n21365), .ZN(
        n7864) );
  OAI22_X1 U20437 ( .A1(n27447), .A2(n27243), .B1(n27237), .B2(n21364), .ZN(
        n7865) );
  OAI22_X1 U20438 ( .A1(n27450), .A2(n27243), .B1(n27237), .B2(n21363), .ZN(
        n7866) );
  OAI22_X1 U20439 ( .A1(n27453), .A2(n27243), .B1(n27237), .B2(n21362), .ZN(
        n7867) );
  OAI22_X1 U20440 ( .A1(n27456), .A2(n27243), .B1(n27237), .B2(n21361), .ZN(
        n7868) );
  OAI22_X1 U20441 ( .A1(n27459), .A2(n27244), .B1(n27237), .B2(n21360), .ZN(
        n7869) );
  OAI22_X1 U20442 ( .A1(n27319), .A2(n27000), .B1(n26994), .B2(n21347), .ZN(
        n6542) );
  OAI22_X1 U20443 ( .A1(n27322), .A2(n27000), .B1(n26994), .B2(n21346), .ZN(
        n6543) );
  OAI22_X1 U20444 ( .A1(n27325), .A2(n27000), .B1(n26994), .B2(n21345), .ZN(
        n6544) );
  OAI22_X1 U20445 ( .A1(n27328), .A2(n27000), .B1(n26994), .B2(n21344), .ZN(
        n6545) );
  OAI22_X1 U20446 ( .A1(n27331), .A2(n27000), .B1(n26994), .B2(n21343), .ZN(
        n6546) );
  OAI22_X1 U20447 ( .A1(n27334), .A2(n27000), .B1(n26994), .B2(n21342), .ZN(
        n6547) );
  OAI22_X1 U20448 ( .A1(n27337), .A2(n27000), .B1(n26994), .B2(n21341), .ZN(
        n6548) );
  OAI22_X1 U20449 ( .A1(n27340), .A2(n27000), .B1(n26994), .B2(n21340), .ZN(
        n6549) );
  OAI22_X1 U20450 ( .A1(n27343), .A2(n27000), .B1(n26994), .B2(n21339), .ZN(
        n6550) );
  OAI22_X1 U20451 ( .A1(n27346), .A2(n27000), .B1(n26994), .B2(n21338), .ZN(
        n6551) );
  OAI22_X1 U20452 ( .A1(n27349), .A2(n27000), .B1(n26994), .B2(n21337), .ZN(
        n6552) );
  OAI22_X1 U20453 ( .A1(n27352), .A2(n27001), .B1(n26994), .B2(n21336), .ZN(
        n6553) );
  OAI22_X1 U20454 ( .A1(n27355), .A2(n27001), .B1(n26995), .B2(n21335), .ZN(
        n6554) );
  OAI22_X1 U20455 ( .A1(n27358), .A2(n27001), .B1(n26995), .B2(n21334), .ZN(
        n6555) );
  OAI22_X1 U20456 ( .A1(n27361), .A2(n27001), .B1(n26995), .B2(n21333), .ZN(
        n6556) );
  OAI22_X1 U20457 ( .A1(n27364), .A2(n27001), .B1(n26995), .B2(n21332), .ZN(
        n6557) );
  OAI22_X1 U20458 ( .A1(n27367), .A2(n27001), .B1(n26995), .B2(n21331), .ZN(
        n6558) );
  OAI22_X1 U20459 ( .A1(n27370), .A2(n27001), .B1(n26995), .B2(n21330), .ZN(
        n6559) );
  OAI22_X1 U20460 ( .A1(n27373), .A2(n27001), .B1(n26995), .B2(n21329), .ZN(
        n6560) );
  OAI22_X1 U20461 ( .A1(n27376), .A2(n27001), .B1(n26995), .B2(n21328), .ZN(
        n6561) );
  OAI22_X1 U20462 ( .A1(n27379), .A2(n27001), .B1(n26995), .B2(n21327), .ZN(
        n6562) );
  OAI22_X1 U20463 ( .A1(n27382), .A2(n27001), .B1(n26995), .B2(n21326), .ZN(
        n6563) );
  OAI22_X1 U20464 ( .A1(n27385), .A2(n27001), .B1(n26995), .B2(n21325), .ZN(
        n6564) );
  OAI22_X1 U20465 ( .A1(n27388), .A2(n27002), .B1(n26995), .B2(n21324), .ZN(
        n6565) );
  OAI22_X1 U20466 ( .A1(n27391), .A2(n27002), .B1(n26996), .B2(n21323), .ZN(
        n6566) );
  OAI22_X1 U20467 ( .A1(n27394), .A2(n27002), .B1(n26996), .B2(n21322), .ZN(
        n6567) );
  OAI22_X1 U20468 ( .A1(n27397), .A2(n27002), .B1(n26996), .B2(n21321), .ZN(
        n6568) );
  OAI22_X1 U20469 ( .A1(n27400), .A2(n27002), .B1(n26996), .B2(n21320), .ZN(
        n6569) );
  OAI22_X1 U20470 ( .A1(n27403), .A2(n27002), .B1(n26996), .B2(n21319), .ZN(
        n6570) );
  OAI22_X1 U20471 ( .A1(n27406), .A2(n27002), .B1(n26996), .B2(n21318), .ZN(
        n6571) );
  OAI22_X1 U20472 ( .A1(n27409), .A2(n27002), .B1(n26996), .B2(n21317), .ZN(
        n6572) );
  OAI22_X1 U20473 ( .A1(n27412), .A2(n27002), .B1(n26996), .B2(n21316), .ZN(
        n6573) );
  OAI22_X1 U20474 ( .A1(n27415), .A2(n27002), .B1(n26996), .B2(n21315), .ZN(
        n6574) );
  OAI22_X1 U20475 ( .A1(n27418), .A2(n27002), .B1(n26996), .B2(n21314), .ZN(
        n6575) );
  OAI22_X1 U20476 ( .A1(n27421), .A2(n27002), .B1(n26996), .B2(n21313), .ZN(
        n6576) );
  OAI22_X1 U20477 ( .A1(n27424), .A2(n27003), .B1(n26996), .B2(n21312), .ZN(
        n6577) );
  OAI22_X1 U20478 ( .A1(n27427), .A2(n27003), .B1(n26997), .B2(n21311), .ZN(
        n6578) );
  OAI22_X1 U20479 ( .A1(n27430), .A2(n27003), .B1(n26997), .B2(n21310), .ZN(
        n6579) );
  OAI22_X1 U20480 ( .A1(n27433), .A2(n27003), .B1(n26997), .B2(n21309), .ZN(
        n6580) );
  OAI22_X1 U20481 ( .A1(n27436), .A2(n27003), .B1(n26997), .B2(n21308), .ZN(
        n6581) );
  OAI22_X1 U20482 ( .A1(n27439), .A2(n27003), .B1(n26997), .B2(n21307), .ZN(
        n6582) );
  OAI22_X1 U20483 ( .A1(n27442), .A2(n27003), .B1(n26997), .B2(n21306), .ZN(
        n6583) );
  OAI22_X1 U20484 ( .A1(n27445), .A2(n27003), .B1(n26997), .B2(n21305), .ZN(
        n6584) );
  OAI22_X1 U20485 ( .A1(n27448), .A2(n27003), .B1(n26997), .B2(n21304), .ZN(
        n6585) );
  OAI22_X1 U20486 ( .A1(n27451), .A2(n27003), .B1(n26997), .B2(n21303), .ZN(
        n6586) );
  OAI22_X1 U20487 ( .A1(n27454), .A2(n27003), .B1(n26997), .B2(n21302), .ZN(
        n6587) );
  OAI22_X1 U20488 ( .A1(n27457), .A2(n27003), .B1(n26997), .B2(n21301), .ZN(
        n6588) );
  OAI22_X1 U20489 ( .A1(n27460), .A2(n27004), .B1(n26997), .B2(n21300), .ZN(
        n6589) );
  OAI22_X1 U20490 ( .A1(n27319), .A2(n26976), .B1(n26970), .B2(n21227), .ZN(
        n6414) );
  OAI22_X1 U20491 ( .A1(n27322), .A2(n26976), .B1(n26970), .B2(n21226), .ZN(
        n6415) );
  OAI22_X1 U20492 ( .A1(n27325), .A2(n26976), .B1(n26970), .B2(n21225), .ZN(
        n6416) );
  OAI22_X1 U20493 ( .A1(n27328), .A2(n26976), .B1(n26970), .B2(n21224), .ZN(
        n6417) );
  OAI22_X1 U20494 ( .A1(n27331), .A2(n26976), .B1(n26970), .B2(n21223), .ZN(
        n6418) );
  OAI22_X1 U20495 ( .A1(n27334), .A2(n26976), .B1(n26970), .B2(n21222), .ZN(
        n6419) );
  OAI22_X1 U20496 ( .A1(n27337), .A2(n26976), .B1(n26970), .B2(n21221), .ZN(
        n6420) );
  OAI22_X1 U20497 ( .A1(n27340), .A2(n26976), .B1(n26970), .B2(n21220), .ZN(
        n6421) );
  OAI22_X1 U20498 ( .A1(n27343), .A2(n26976), .B1(n26970), .B2(n21219), .ZN(
        n6422) );
  OAI22_X1 U20499 ( .A1(n27346), .A2(n26976), .B1(n26970), .B2(n21218), .ZN(
        n6423) );
  OAI22_X1 U20500 ( .A1(n27349), .A2(n26976), .B1(n26970), .B2(n21217), .ZN(
        n6424) );
  OAI22_X1 U20501 ( .A1(n27352), .A2(n26977), .B1(n26970), .B2(n21216), .ZN(
        n6425) );
  OAI22_X1 U20502 ( .A1(n27355), .A2(n26977), .B1(n26971), .B2(n21215), .ZN(
        n6426) );
  OAI22_X1 U20503 ( .A1(n27358), .A2(n26977), .B1(n26971), .B2(n21214), .ZN(
        n6427) );
  OAI22_X1 U20504 ( .A1(n27361), .A2(n26977), .B1(n26971), .B2(n21213), .ZN(
        n6428) );
  OAI22_X1 U20505 ( .A1(n27364), .A2(n26977), .B1(n26971), .B2(n21212), .ZN(
        n6429) );
  OAI22_X1 U20506 ( .A1(n27367), .A2(n26977), .B1(n26971), .B2(n21211), .ZN(
        n6430) );
  OAI22_X1 U20507 ( .A1(n27370), .A2(n26977), .B1(n26971), .B2(n21210), .ZN(
        n6431) );
  OAI22_X1 U20508 ( .A1(n27373), .A2(n26977), .B1(n26971), .B2(n21209), .ZN(
        n6432) );
  OAI22_X1 U20509 ( .A1(n27376), .A2(n26977), .B1(n26971), .B2(n21208), .ZN(
        n6433) );
  OAI22_X1 U20510 ( .A1(n27379), .A2(n26977), .B1(n26971), .B2(n21207), .ZN(
        n6434) );
  OAI22_X1 U20511 ( .A1(n27382), .A2(n26977), .B1(n26971), .B2(n21206), .ZN(
        n6435) );
  OAI22_X1 U20512 ( .A1(n27385), .A2(n26977), .B1(n26971), .B2(n21205), .ZN(
        n6436) );
  OAI22_X1 U20513 ( .A1(n27388), .A2(n26978), .B1(n26971), .B2(n21204), .ZN(
        n6437) );
  OAI22_X1 U20514 ( .A1(n27391), .A2(n26978), .B1(n26972), .B2(n21203), .ZN(
        n6438) );
  OAI22_X1 U20515 ( .A1(n27394), .A2(n26978), .B1(n26972), .B2(n21202), .ZN(
        n6439) );
  OAI22_X1 U20516 ( .A1(n27397), .A2(n26978), .B1(n26972), .B2(n21201), .ZN(
        n6440) );
  OAI22_X1 U20517 ( .A1(n27400), .A2(n26978), .B1(n26972), .B2(n21200), .ZN(
        n6441) );
  OAI22_X1 U20518 ( .A1(n27403), .A2(n26978), .B1(n26972), .B2(n21199), .ZN(
        n6442) );
  OAI22_X1 U20519 ( .A1(n27406), .A2(n26978), .B1(n26972), .B2(n21198), .ZN(
        n6443) );
  OAI22_X1 U20520 ( .A1(n27409), .A2(n26978), .B1(n26972), .B2(n21197), .ZN(
        n6444) );
  OAI22_X1 U20521 ( .A1(n27412), .A2(n26978), .B1(n26972), .B2(n21196), .ZN(
        n6445) );
  OAI22_X1 U20522 ( .A1(n27415), .A2(n26978), .B1(n26972), .B2(n21195), .ZN(
        n6446) );
  OAI22_X1 U20523 ( .A1(n27418), .A2(n26978), .B1(n26972), .B2(n21194), .ZN(
        n6447) );
  OAI22_X1 U20524 ( .A1(n27421), .A2(n26978), .B1(n26972), .B2(n21193), .ZN(
        n6448) );
  OAI22_X1 U20525 ( .A1(n27424), .A2(n26979), .B1(n26972), .B2(n21192), .ZN(
        n6449) );
  OAI22_X1 U20526 ( .A1(n27427), .A2(n26979), .B1(n26973), .B2(n21191), .ZN(
        n6450) );
  OAI22_X1 U20527 ( .A1(n27430), .A2(n26979), .B1(n26973), .B2(n21190), .ZN(
        n6451) );
  OAI22_X1 U20528 ( .A1(n27433), .A2(n26979), .B1(n26973), .B2(n21189), .ZN(
        n6452) );
  OAI22_X1 U20529 ( .A1(n27436), .A2(n26979), .B1(n26973), .B2(n21188), .ZN(
        n6453) );
  OAI22_X1 U20530 ( .A1(n27439), .A2(n26979), .B1(n26973), .B2(n21187), .ZN(
        n6454) );
  OAI22_X1 U20531 ( .A1(n27442), .A2(n26979), .B1(n26973), .B2(n21186), .ZN(
        n6455) );
  OAI22_X1 U20532 ( .A1(n27445), .A2(n26979), .B1(n26973), .B2(n21185), .ZN(
        n6456) );
  OAI22_X1 U20533 ( .A1(n27448), .A2(n26979), .B1(n26973), .B2(n21184), .ZN(
        n6457) );
  OAI22_X1 U20534 ( .A1(n27451), .A2(n26979), .B1(n26973), .B2(n21183), .ZN(
        n6458) );
  OAI22_X1 U20535 ( .A1(n27454), .A2(n26979), .B1(n26973), .B2(n21182), .ZN(
        n6459) );
  OAI22_X1 U20536 ( .A1(n27457), .A2(n26979), .B1(n26973), .B2(n21181), .ZN(
        n6460) );
  OAI22_X1 U20537 ( .A1(n27460), .A2(n26980), .B1(n26973), .B2(n21180), .ZN(
        n6461) );
  OAI22_X1 U20538 ( .A1(n27319), .A2(n27108), .B1(n27102), .B2(n20822), .ZN(
        n7118) );
  OAI22_X1 U20539 ( .A1(n27322), .A2(n27108), .B1(n27102), .B2(n20821), .ZN(
        n7119) );
  OAI22_X1 U20540 ( .A1(n27325), .A2(n27108), .B1(n27102), .B2(n20820), .ZN(
        n7120) );
  OAI22_X1 U20541 ( .A1(n27328), .A2(n27108), .B1(n27102), .B2(n20819), .ZN(
        n7121) );
  OAI22_X1 U20542 ( .A1(n27331), .A2(n27108), .B1(n27102), .B2(n20818), .ZN(
        n7122) );
  OAI22_X1 U20543 ( .A1(n27334), .A2(n27108), .B1(n27102), .B2(n20817), .ZN(
        n7123) );
  OAI22_X1 U20544 ( .A1(n27337), .A2(n27108), .B1(n27102), .B2(n20816), .ZN(
        n7124) );
  OAI22_X1 U20545 ( .A1(n27340), .A2(n27108), .B1(n27102), .B2(n20815), .ZN(
        n7125) );
  OAI22_X1 U20546 ( .A1(n27343), .A2(n27108), .B1(n27102), .B2(n20814), .ZN(
        n7126) );
  OAI22_X1 U20547 ( .A1(n27346), .A2(n27108), .B1(n27102), .B2(n20813), .ZN(
        n7127) );
  OAI22_X1 U20548 ( .A1(n27349), .A2(n27108), .B1(n27102), .B2(n20812), .ZN(
        n7128) );
  OAI22_X1 U20549 ( .A1(n27352), .A2(n27109), .B1(n27102), .B2(n20811), .ZN(
        n7129) );
  OAI22_X1 U20550 ( .A1(n27355), .A2(n27109), .B1(n27103), .B2(n20810), .ZN(
        n7130) );
  OAI22_X1 U20551 ( .A1(n27358), .A2(n27109), .B1(n27103), .B2(n20809), .ZN(
        n7131) );
  OAI22_X1 U20552 ( .A1(n27361), .A2(n27109), .B1(n27103), .B2(n20808), .ZN(
        n7132) );
  OAI22_X1 U20553 ( .A1(n27364), .A2(n27109), .B1(n27103), .B2(n20807), .ZN(
        n7133) );
  OAI22_X1 U20554 ( .A1(n27367), .A2(n27109), .B1(n27103), .B2(n20806), .ZN(
        n7134) );
  OAI22_X1 U20555 ( .A1(n27370), .A2(n27109), .B1(n27103), .B2(n20805), .ZN(
        n7135) );
  OAI22_X1 U20556 ( .A1(n27373), .A2(n27109), .B1(n27103), .B2(n20804), .ZN(
        n7136) );
  OAI22_X1 U20557 ( .A1(n27376), .A2(n27109), .B1(n27103), .B2(n20803), .ZN(
        n7137) );
  OAI22_X1 U20558 ( .A1(n27379), .A2(n27109), .B1(n27103), .B2(n20802), .ZN(
        n7138) );
  OAI22_X1 U20559 ( .A1(n27382), .A2(n27109), .B1(n27103), .B2(n20801), .ZN(
        n7139) );
  OAI22_X1 U20560 ( .A1(n27385), .A2(n27109), .B1(n27103), .B2(n20800), .ZN(
        n7140) );
  OAI22_X1 U20561 ( .A1(n27388), .A2(n27110), .B1(n27103), .B2(n20799), .ZN(
        n7141) );
  OAI22_X1 U20562 ( .A1(n27391), .A2(n27110), .B1(n27104), .B2(n20798), .ZN(
        n7142) );
  OAI22_X1 U20563 ( .A1(n27394), .A2(n27110), .B1(n27104), .B2(n20797), .ZN(
        n7143) );
  OAI22_X1 U20564 ( .A1(n27397), .A2(n27110), .B1(n27104), .B2(n20796), .ZN(
        n7144) );
  OAI22_X1 U20565 ( .A1(n27400), .A2(n27110), .B1(n27104), .B2(n20795), .ZN(
        n7145) );
  OAI22_X1 U20566 ( .A1(n27403), .A2(n27110), .B1(n27104), .B2(n20794), .ZN(
        n7146) );
  OAI22_X1 U20567 ( .A1(n27406), .A2(n27110), .B1(n27104), .B2(n20793), .ZN(
        n7147) );
  OAI22_X1 U20568 ( .A1(n27409), .A2(n27110), .B1(n27104), .B2(n20792), .ZN(
        n7148) );
  OAI22_X1 U20569 ( .A1(n27412), .A2(n27110), .B1(n27104), .B2(n20791), .ZN(
        n7149) );
  OAI22_X1 U20570 ( .A1(n27415), .A2(n27110), .B1(n27104), .B2(n20790), .ZN(
        n7150) );
  OAI22_X1 U20571 ( .A1(n27418), .A2(n27110), .B1(n27104), .B2(n20789), .ZN(
        n7151) );
  OAI22_X1 U20572 ( .A1(n27421), .A2(n27110), .B1(n27104), .B2(n20788), .ZN(
        n7152) );
  OAI22_X1 U20573 ( .A1(n27424), .A2(n27111), .B1(n27104), .B2(n20787), .ZN(
        n7153) );
  OAI22_X1 U20574 ( .A1(n27427), .A2(n27111), .B1(n27105), .B2(n20786), .ZN(
        n7154) );
  OAI22_X1 U20575 ( .A1(n27430), .A2(n27111), .B1(n27105), .B2(n20785), .ZN(
        n7155) );
  OAI22_X1 U20576 ( .A1(n27433), .A2(n27111), .B1(n27105), .B2(n20784), .ZN(
        n7156) );
  OAI22_X1 U20577 ( .A1(n27436), .A2(n27111), .B1(n27105), .B2(n20783), .ZN(
        n7157) );
  OAI22_X1 U20578 ( .A1(n27439), .A2(n27111), .B1(n27105), .B2(n20782), .ZN(
        n7158) );
  OAI22_X1 U20579 ( .A1(n27442), .A2(n27111), .B1(n27105), .B2(n20781), .ZN(
        n7159) );
  OAI22_X1 U20580 ( .A1(n27445), .A2(n27111), .B1(n27105), .B2(n20780), .ZN(
        n7160) );
  OAI22_X1 U20581 ( .A1(n27448), .A2(n27111), .B1(n27105), .B2(n20779), .ZN(
        n7161) );
  OAI22_X1 U20582 ( .A1(n27451), .A2(n27111), .B1(n27105), .B2(n20778), .ZN(
        n7162) );
  OAI22_X1 U20583 ( .A1(n27454), .A2(n27111), .B1(n27105), .B2(n20777), .ZN(
        n7163) );
  OAI22_X1 U20584 ( .A1(n27457), .A2(n27111), .B1(n27105), .B2(n20776), .ZN(
        n7164) );
  OAI22_X1 U20585 ( .A1(n27460), .A2(n27112), .B1(n27105), .B2(n20775), .ZN(
        n7165) );
  OAI22_X1 U20586 ( .A1(n27318), .A2(n27132), .B1(n27126), .B2(n20759), .ZN(
        n7246) );
  OAI22_X1 U20587 ( .A1(n27321), .A2(n27132), .B1(n27126), .B2(n20758), .ZN(
        n7247) );
  OAI22_X1 U20588 ( .A1(n27324), .A2(n27132), .B1(n27126), .B2(n20757), .ZN(
        n7248) );
  OAI22_X1 U20589 ( .A1(n27327), .A2(n27132), .B1(n27126), .B2(n20756), .ZN(
        n7249) );
  OAI22_X1 U20590 ( .A1(n27330), .A2(n27132), .B1(n27126), .B2(n20755), .ZN(
        n7250) );
  OAI22_X1 U20591 ( .A1(n27333), .A2(n27132), .B1(n27126), .B2(n20754), .ZN(
        n7251) );
  OAI22_X1 U20592 ( .A1(n27336), .A2(n27132), .B1(n27126), .B2(n20753), .ZN(
        n7252) );
  OAI22_X1 U20593 ( .A1(n27339), .A2(n27132), .B1(n27126), .B2(n20752), .ZN(
        n7253) );
  OAI22_X1 U20594 ( .A1(n27342), .A2(n27132), .B1(n27126), .B2(n20751), .ZN(
        n7254) );
  OAI22_X1 U20595 ( .A1(n27345), .A2(n27132), .B1(n27126), .B2(n20750), .ZN(
        n7255) );
  OAI22_X1 U20596 ( .A1(n27348), .A2(n27132), .B1(n27126), .B2(n20749), .ZN(
        n7256) );
  OAI22_X1 U20597 ( .A1(n27351), .A2(n27133), .B1(n27126), .B2(n20748), .ZN(
        n7257) );
  OAI22_X1 U20598 ( .A1(n27354), .A2(n27133), .B1(n27127), .B2(n20747), .ZN(
        n7258) );
  OAI22_X1 U20599 ( .A1(n27357), .A2(n27133), .B1(n27127), .B2(n20746), .ZN(
        n7259) );
  OAI22_X1 U20600 ( .A1(n27360), .A2(n27133), .B1(n27127), .B2(n20745), .ZN(
        n7260) );
  OAI22_X1 U20601 ( .A1(n27363), .A2(n27133), .B1(n27127), .B2(n20744), .ZN(
        n7261) );
  OAI22_X1 U20602 ( .A1(n27366), .A2(n27133), .B1(n27127), .B2(n20743), .ZN(
        n7262) );
  OAI22_X1 U20603 ( .A1(n27369), .A2(n27133), .B1(n27127), .B2(n20742), .ZN(
        n7263) );
  OAI22_X1 U20604 ( .A1(n27372), .A2(n27133), .B1(n27127), .B2(n20741), .ZN(
        n7264) );
  OAI22_X1 U20605 ( .A1(n27375), .A2(n27133), .B1(n27127), .B2(n20740), .ZN(
        n7265) );
  OAI22_X1 U20606 ( .A1(n27378), .A2(n27133), .B1(n27127), .B2(n20739), .ZN(
        n7266) );
  OAI22_X1 U20607 ( .A1(n27381), .A2(n27133), .B1(n27127), .B2(n20738), .ZN(
        n7267) );
  OAI22_X1 U20608 ( .A1(n27384), .A2(n27133), .B1(n27127), .B2(n20737), .ZN(
        n7268) );
  OAI22_X1 U20609 ( .A1(n27387), .A2(n27134), .B1(n27127), .B2(n20736), .ZN(
        n7269) );
  OAI22_X1 U20610 ( .A1(n27390), .A2(n27134), .B1(n27128), .B2(n20735), .ZN(
        n7270) );
  OAI22_X1 U20611 ( .A1(n27393), .A2(n27134), .B1(n27128), .B2(n20734), .ZN(
        n7271) );
  OAI22_X1 U20612 ( .A1(n27396), .A2(n27134), .B1(n27128), .B2(n20733), .ZN(
        n7272) );
  OAI22_X1 U20613 ( .A1(n27399), .A2(n27134), .B1(n27128), .B2(n20732), .ZN(
        n7273) );
  OAI22_X1 U20614 ( .A1(n27402), .A2(n27134), .B1(n27128), .B2(n20731), .ZN(
        n7274) );
  OAI22_X1 U20615 ( .A1(n27405), .A2(n27134), .B1(n27128), .B2(n20730), .ZN(
        n7275) );
  OAI22_X1 U20616 ( .A1(n27408), .A2(n27134), .B1(n27128), .B2(n20729), .ZN(
        n7276) );
  OAI22_X1 U20617 ( .A1(n27411), .A2(n27134), .B1(n27128), .B2(n20728), .ZN(
        n7277) );
  OAI22_X1 U20618 ( .A1(n27414), .A2(n27134), .B1(n27128), .B2(n20727), .ZN(
        n7278) );
  OAI22_X1 U20619 ( .A1(n27417), .A2(n27134), .B1(n27128), .B2(n20726), .ZN(
        n7279) );
  OAI22_X1 U20620 ( .A1(n27420), .A2(n27134), .B1(n27128), .B2(n20725), .ZN(
        n7280) );
  OAI22_X1 U20621 ( .A1(n27423), .A2(n27135), .B1(n27128), .B2(n20724), .ZN(
        n7281) );
  OAI22_X1 U20622 ( .A1(n27426), .A2(n27135), .B1(n27129), .B2(n20723), .ZN(
        n7282) );
  OAI22_X1 U20623 ( .A1(n27429), .A2(n27135), .B1(n27129), .B2(n20722), .ZN(
        n7283) );
  OAI22_X1 U20624 ( .A1(n27432), .A2(n27135), .B1(n27129), .B2(n20721), .ZN(
        n7284) );
  OAI22_X1 U20625 ( .A1(n27435), .A2(n27135), .B1(n27129), .B2(n20720), .ZN(
        n7285) );
  OAI22_X1 U20626 ( .A1(n27438), .A2(n27135), .B1(n27129), .B2(n20719), .ZN(
        n7286) );
  OAI22_X1 U20627 ( .A1(n27441), .A2(n27135), .B1(n27129), .B2(n20718), .ZN(
        n7287) );
  OAI22_X1 U20628 ( .A1(n27444), .A2(n27135), .B1(n27129), .B2(n20717), .ZN(
        n7288) );
  OAI22_X1 U20629 ( .A1(n27447), .A2(n27135), .B1(n27129), .B2(n20716), .ZN(
        n7289) );
  OAI22_X1 U20630 ( .A1(n27450), .A2(n27135), .B1(n27129), .B2(n20715), .ZN(
        n7290) );
  OAI22_X1 U20631 ( .A1(n27453), .A2(n27135), .B1(n27129), .B2(n20714), .ZN(
        n7291) );
  OAI22_X1 U20632 ( .A1(n27456), .A2(n27135), .B1(n27129), .B2(n20713), .ZN(
        n7292) );
  OAI22_X1 U20633 ( .A1(n27459), .A2(n27136), .B1(n27129), .B2(n20712), .ZN(
        n7293) );
  OAI22_X1 U20634 ( .A1(n27462), .A2(n27172), .B1(n27166), .B2(n22511), .ZN(
        n7486) );
  OAI22_X1 U20635 ( .A1(n27465), .A2(n27172), .B1(n27166), .B2(n22510), .ZN(
        n7487) );
  OAI22_X1 U20636 ( .A1(n27468), .A2(n27172), .B1(n27166), .B2(n22509), .ZN(
        n7488) );
  OAI22_X1 U20637 ( .A1(n27471), .A2(n27172), .B1(n27166), .B2(n22508), .ZN(
        n7489) );
  OAI22_X1 U20638 ( .A1(n27463), .A2(n26992), .B1(n26986), .B2(n22503), .ZN(
        n6526) );
  OAI22_X1 U20639 ( .A1(n27466), .A2(n26992), .B1(n26986), .B2(n22502), .ZN(
        n6527) );
  OAI22_X1 U20640 ( .A1(n27469), .A2(n26992), .B1(n26986), .B2(n22501), .ZN(
        n6528) );
  OAI22_X1 U20641 ( .A1(n27472), .A2(n26992), .B1(n26986), .B2(n22500), .ZN(
        n6529) );
  OAI22_X1 U20642 ( .A1(n27462), .A2(n27184), .B1(n27178), .B2(n22259), .ZN(
        n7550) );
  OAI22_X1 U20643 ( .A1(n27465), .A2(n27184), .B1(n27178), .B2(n22258), .ZN(
        n7551) );
  OAI22_X1 U20644 ( .A1(n27468), .A2(n27184), .B1(n27178), .B2(n22257), .ZN(
        n7552) );
  OAI22_X1 U20645 ( .A1(n27471), .A2(n27184), .B1(n27178), .B2(n22256), .ZN(
        n7553) );
  OAI22_X1 U20646 ( .A1(n27463), .A2(n27052), .B1(n27046), .B2(n22251), .ZN(
        n6846) );
  OAI22_X1 U20647 ( .A1(n27466), .A2(n27052), .B1(n27046), .B2(n22250), .ZN(
        n6847) );
  OAI22_X1 U20648 ( .A1(n27469), .A2(n27052), .B1(n27046), .B2(n22249), .ZN(
        n6848) );
  OAI22_X1 U20649 ( .A1(n27472), .A2(n27052), .B1(n27046), .B2(n22248), .ZN(
        n6849) );
  OAI22_X1 U20650 ( .A1(n27462), .A2(n27196), .B1(n27190), .B2(n21511), .ZN(
        n7614) );
  OAI22_X1 U20651 ( .A1(n27465), .A2(n27196), .B1(n27190), .B2(n21510), .ZN(
        n7615) );
  OAI22_X1 U20652 ( .A1(n27468), .A2(n27196), .B1(n27190), .B2(n21509), .ZN(
        n7616) );
  OAI22_X1 U20653 ( .A1(n27471), .A2(n27196), .B1(n27190), .B2(n21508), .ZN(
        n7617) );
  OAI22_X1 U20654 ( .A1(n27462), .A2(n27148), .B1(n27142), .B2(n21507), .ZN(
        n7358) );
  OAI22_X1 U20655 ( .A1(n27465), .A2(n27148), .B1(n27142), .B2(n21506), .ZN(
        n7359) );
  OAI22_X1 U20656 ( .A1(n27468), .A2(n27148), .B1(n27142), .B2(n21505), .ZN(
        n7360) );
  OAI22_X1 U20657 ( .A1(n27471), .A2(n27148), .B1(n27142), .B2(n21504), .ZN(
        n7361) );
  OAI22_X1 U20658 ( .A1(n27463), .A2(n27076), .B1(n27070), .B2(n21491), .ZN(
        n6974) );
  OAI22_X1 U20659 ( .A1(n27466), .A2(n27076), .B1(n27070), .B2(n21490), .ZN(
        n6975) );
  OAI22_X1 U20660 ( .A1(n27469), .A2(n27076), .B1(n27070), .B2(n21489), .ZN(
        n6976) );
  OAI22_X1 U20661 ( .A1(n27472), .A2(n27076), .B1(n27070), .B2(n21488), .ZN(
        n6977) );
  OAI22_X1 U20662 ( .A1(n27464), .A2(n26968), .B1(n26962), .B2(n21483), .ZN(
        n6398) );
  OAI22_X1 U20663 ( .A1(n27467), .A2(n26968), .B1(n26962), .B2(n21482), .ZN(
        n6399) );
  OAI22_X1 U20664 ( .A1(n27470), .A2(n26968), .B1(n26962), .B2(n21481), .ZN(
        n6400) );
  OAI22_X1 U20665 ( .A1(n27473), .A2(n26968), .B1(n26962), .B2(n21480), .ZN(
        n6401) );
  OAI22_X1 U20666 ( .A1(n27462), .A2(n27220), .B1(n27214), .B2(n21179), .ZN(
        n7742) );
  OAI22_X1 U20667 ( .A1(n27465), .A2(n27220), .B1(n27214), .B2(n21178), .ZN(
        n7743) );
  OAI22_X1 U20668 ( .A1(n27468), .A2(n27220), .B1(n27214), .B2(n21177), .ZN(
        n7744) );
  OAI22_X1 U20669 ( .A1(n27471), .A2(n27220), .B1(n27214), .B2(n21176), .ZN(
        n7745) );
  OAI22_X1 U20670 ( .A1(n27462), .A2(n27244), .B1(n27238), .B2(n21171), .ZN(
        n7870) );
  OAI22_X1 U20671 ( .A1(n27465), .A2(n27244), .B1(n27238), .B2(n21170), .ZN(
        n7871) );
  OAI22_X1 U20672 ( .A1(n27468), .A2(n27244), .B1(n27238), .B2(n21169), .ZN(
        n7872) );
  OAI22_X1 U20673 ( .A1(n27471), .A2(n27244), .B1(n27238), .B2(n21168), .ZN(
        n7873) );
  OAI22_X1 U20674 ( .A1(n27463), .A2(n27004), .B1(n26998), .B2(n21167), .ZN(
        n6590) );
  OAI22_X1 U20675 ( .A1(n27466), .A2(n27004), .B1(n26998), .B2(n21166), .ZN(
        n6591) );
  OAI22_X1 U20676 ( .A1(n27469), .A2(n27004), .B1(n26998), .B2(n21165), .ZN(
        n6592) );
  OAI22_X1 U20677 ( .A1(n27472), .A2(n27004), .B1(n26998), .B2(n21164), .ZN(
        n6593) );
  OAI22_X1 U20678 ( .A1(n27463), .A2(n26980), .B1(n26974), .B2(n21159), .ZN(
        n6462) );
  OAI22_X1 U20679 ( .A1(n27466), .A2(n26980), .B1(n26974), .B2(n21158), .ZN(
        n6463) );
  OAI22_X1 U20680 ( .A1(n27469), .A2(n26980), .B1(n26974), .B2(n21157), .ZN(
        n6464) );
  OAI22_X1 U20681 ( .A1(n27472), .A2(n26980), .B1(n26974), .B2(n21156), .ZN(
        n6465) );
  OAI22_X1 U20682 ( .A1(n27472), .A2(n27112), .B1(n27106), .B2(n21155), .ZN(
        n7169) );
  OAI22_X1 U20683 ( .A1(n27463), .A2(n27112), .B1(n27106), .B2(n20774), .ZN(
        n7166) );
  OAI22_X1 U20684 ( .A1(n27466), .A2(n27112), .B1(n27106), .B2(n20773), .ZN(
        n7167) );
  OAI22_X1 U20685 ( .A1(n27469), .A2(n27112), .B1(n27106), .B2(n20772), .ZN(
        n7168) );
  OAI22_X1 U20686 ( .A1(n27462), .A2(n27136), .B1(n27130), .B2(n20711), .ZN(
        n7294) );
  OAI22_X1 U20687 ( .A1(n27465), .A2(n27136), .B1(n27130), .B2(n20710), .ZN(
        n7295) );
  OAI22_X1 U20688 ( .A1(n27468), .A2(n27136), .B1(n27130), .B2(n20709), .ZN(
        n7296) );
  OAI22_X1 U20689 ( .A1(n27471), .A2(n27136), .B1(n27130), .B2(n20708), .ZN(
        n7297) );
  OAI22_X1 U20690 ( .A1(n27282), .A2(n27167), .B1(n27161), .B2(n22691), .ZN(
        n7426) );
  OAI22_X1 U20691 ( .A1(n27285), .A2(n27167), .B1(n27161), .B2(n22690), .ZN(
        n7427) );
  OAI22_X1 U20692 ( .A1(n27288), .A2(n27167), .B1(n27161), .B2(n22689), .ZN(
        n7428) );
  OAI22_X1 U20693 ( .A1(n27291), .A2(n27167), .B1(n27161), .B2(n22688), .ZN(
        n7429) );
  OAI22_X1 U20694 ( .A1(n27294), .A2(n27167), .B1(n27161), .B2(n22687), .ZN(
        n7430) );
  OAI22_X1 U20695 ( .A1(n27297), .A2(n27167), .B1(n27161), .B2(n22686), .ZN(
        n7431) );
  OAI22_X1 U20696 ( .A1(n27300), .A2(n27167), .B1(n27161), .B2(n22685), .ZN(
        n7432) );
  OAI22_X1 U20697 ( .A1(n27303), .A2(n27167), .B1(n27161), .B2(n22684), .ZN(
        n7433) );
  OAI22_X1 U20698 ( .A1(n27306), .A2(n27167), .B1(n27161), .B2(n22683), .ZN(
        n7434) );
  OAI22_X1 U20699 ( .A1(n27309), .A2(n27167), .B1(n27161), .B2(n22682), .ZN(
        n7435) );
  OAI22_X1 U20700 ( .A1(n27312), .A2(n27167), .B1(n27161), .B2(n22681), .ZN(
        n7436) );
  OAI22_X1 U20701 ( .A1(n27315), .A2(n27168), .B1(n27161), .B2(n22680), .ZN(
        n7437) );
  OAI22_X1 U20702 ( .A1(n27283), .A2(n26987), .B1(n26981), .B2(n22571), .ZN(
        n6466) );
  OAI22_X1 U20703 ( .A1(n27286), .A2(n26987), .B1(n26981), .B2(n22570), .ZN(
        n6467) );
  OAI22_X1 U20704 ( .A1(n27289), .A2(n26987), .B1(n26981), .B2(n22569), .ZN(
        n6468) );
  OAI22_X1 U20705 ( .A1(n27292), .A2(n26987), .B1(n26981), .B2(n22568), .ZN(
        n6469) );
  OAI22_X1 U20706 ( .A1(n27295), .A2(n26987), .B1(n26981), .B2(n22567), .ZN(
        n6470) );
  OAI22_X1 U20707 ( .A1(n27298), .A2(n26987), .B1(n26981), .B2(n22566), .ZN(
        n6471) );
  OAI22_X1 U20708 ( .A1(n27301), .A2(n26987), .B1(n26981), .B2(n22565), .ZN(
        n6472) );
  OAI22_X1 U20709 ( .A1(n27304), .A2(n26987), .B1(n26981), .B2(n22564), .ZN(
        n6473) );
  OAI22_X1 U20710 ( .A1(n27307), .A2(n26987), .B1(n26981), .B2(n22563), .ZN(
        n6474) );
  OAI22_X1 U20711 ( .A1(n27310), .A2(n26987), .B1(n26981), .B2(n22562), .ZN(
        n6475) );
  OAI22_X1 U20712 ( .A1(n27313), .A2(n26987), .B1(n26981), .B2(n22561), .ZN(
        n6476) );
  OAI22_X1 U20713 ( .A1(n27316), .A2(n26988), .B1(n26981), .B2(n22560), .ZN(
        n6477) );
  OAI22_X1 U20714 ( .A1(n27282), .A2(n27179), .B1(n27173), .B2(n22499), .ZN(
        n7490) );
  OAI22_X1 U20715 ( .A1(n27285), .A2(n27179), .B1(n27173), .B2(n22498), .ZN(
        n7491) );
  OAI22_X1 U20716 ( .A1(n27288), .A2(n27179), .B1(n27173), .B2(n22497), .ZN(
        n7492) );
  OAI22_X1 U20717 ( .A1(n27291), .A2(n27179), .B1(n27173), .B2(n22496), .ZN(
        n7493) );
  OAI22_X1 U20718 ( .A1(n27294), .A2(n27179), .B1(n27173), .B2(n22495), .ZN(
        n7494) );
  OAI22_X1 U20719 ( .A1(n27297), .A2(n27179), .B1(n27173), .B2(n22494), .ZN(
        n7495) );
  OAI22_X1 U20720 ( .A1(n27300), .A2(n27179), .B1(n27173), .B2(n22493), .ZN(
        n7496) );
  OAI22_X1 U20721 ( .A1(n27303), .A2(n27179), .B1(n27173), .B2(n22492), .ZN(
        n7497) );
  OAI22_X1 U20722 ( .A1(n27306), .A2(n27179), .B1(n27173), .B2(n22491), .ZN(
        n7498) );
  OAI22_X1 U20723 ( .A1(n27309), .A2(n27179), .B1(n27173), .B2(n22490), .ZN(
        n7499) );
  OAI22_X1 U20724 ( .A1(n27312), .A2(n27179), .B1(n27173), .B2(n22489), .ZN(
        n7500) );
  OAI22_X1 U20725 ( .A1(n27315), .A2(n27180), .B1(n27173), .B2(n22488), .ZN(
        n7501) );
  OAI22_X1 U20726 ( .A1(n27283), .A2(n27047), .B1(n27041), .B2(n22379), .ZN(
        n6786) );
  OAI22_X1 U20727 ( .A1(n27286), .A2(n27047), .B1(n27041), .B2(n22378), .ZN(
        n6787) );
  OAI22_X1 U20728 ( .A1(n27289), .A2(n27047), .B1(n27041), .B2(n22377), .ZN(
        n6788) );
  OAI22_X1 U20729 ( .A1(n27292), .A2(n27047), .B1(n27041), .B2(n22376), .ZN(
        n6789) );
  OAI22_X1 U20730 ( .A1(n27295), .A2(n27047), .B1(n27041), .B2(n22375), .ZN(
        n6790) );
  OAI22_X1 U20731 ( .A1(n27298), .A2(n27047), .B1(n27041), .B2(n22374), .ZN(
        n6791) );
  OAI22_X1 U20732 ( .A1(n27301), .A2(n27047), .B1(n27041), .B2(n22373), .ZN(
        n6792) );
  OAI22_X1 U20733 ( .A1(n27304), .A2(n27047), .B1(n27041), .B2(n22372), .ZN(
        n6793) );
  OAI22_X1 U20734 ( .A1(n27307), .A2(n27047), .B1(n27041), .B2(n22371), .ZN(
        n6794) );
  OAI22_X1 U20735 ( .A1(n27310), .A2(n27047), .B1(n27041), .B2(n22370), .ZN(
        n6795) );
  OAI22_X1 U20736 ( .A1(n27313), .A2(n27047), .B1(n27041), .B2(n22369), .ZN(
        n6796) );
  OAI22_X1 U20737 ( .A1(n27316), .A2(n27048), .B1(n27041), .B2(n22368), .ZN(
        n6797) );
  OAI22_X1 U20738 ( .A1(n27282), .A2(n27191), .B1(n27185), .B2(n22059), .ZN(
        n7554) );
  OAI22_X1 U20739 ( .A1(n27285), .A2(n27191), .B1(n27185), .B2(n22058), .ZN(
        n7555) );
  OAI22_X1 U20740 ( .A1(n27288), .A2(n27191), .B1(n27185), .B2(n22057), .ZN(
        n7556) );
  OAI22_X1 U20741 ( .A1(n27291), .A2(n27191), .B1(n27185), .B2(n22056), .ZN(
        n7557) );
  OAI22_X1 U20742 ( .A1(n27294), .A2(n27191), .B1(n27185), .B2(n22055), .ZN(
        n7558) );
  OAI22_X1 U20743 ( .A1(n27297), .A2(n27191), .B1(n27185), .B2(n22054), .ZN(
        n7559) );
  OAI22_X1 U20744 ( .A1(n27300), .A2(n27191), .B1(n27185), .B2(n22053), .ZN(
        n7560) );
  OAI22_X1 U20745 ( .A1(n27303), .A2(n27191), .B1(n27185), .B2(n22052), .ZN(
        n7561) );
  OAI22_X1 U20746 ( .A1(n27306), .A2(n27191), .B1(n27185), .B2(n22051), .ZN(
        n7562) );
  OAI22_X1 U20747 ( .A1(n27309), .A2(n27191), .B1(n27185), .B2(n22050), .ZN(
        n7563) );
  OAI22_X1 U20748 ( .A1(n27312), .A2(n27191), .B1(n27185), .B2(n22049), .ZN(
        n7564) );
  OAI22_X1 U20749 ( .A1(n27315), .A2(n27192), .B1(n27185), .B2(n22048), .ZN(
        n7565) );
  OAI22_X1 U20750 ( .A1(n27282), .A2(n27143), .B1(n27137), .B2(n21999), .ZN(
        n7298) );
  OAI22_X1 U20751 ( .A1(n27285), .A2(n27143), .B1(n27137), .B2(n21998), .ZN(
        n7299) );
  OAI22_X1 U20752 ( .A1(n27288), .A2(n27143), .B1(n27137), .B2(n21997), .ZN(
        n7300) );
  OAI22_X1 U20753 ( .A1(n27291), .A2(n27143), .B1(n27137), .B2(n21996), .ZN(
        n7301) );
  OAI22_X1 U20754 ( .A1(n27294), .A2(n27143), .B1(n27137), .B2(n21995), .ZN(
        n7302) );
  OAI22_X1 U20755 ( .A1(n27297), .A2(n27143), .B1(n27137), .B2(n21994), .ZN(
        n7303) );
  OAI22_X1 U20756 ( .A1(n27300), .A2(n27143), .B1(n27137), .B2(n21993), .ZN(
        n7304) );
  OAI22_X1 U20757 ( .A1(n27303), .A2(n27143), .B1(n27137), .B2(n21992), .ZN(
        n7305) );
  OAI22_X1 U20758 ( .A1(n27306), .A2(n27143), .B1(n27137), .B2(n21991), .ZN(
        n7306) );
  OAI22_X1 U20759 ( .A1(n27309), .A2(n27143), .B1(n27137), .B2(n21990), .ZN(
        n7307) );
  OAI22_X1 U20760 ( .A1(n27312), .A2(n27143), .B1(n27137), .B2(n21989), .ZN(
        n7308) );
  OAI22_X1 U20761 ( .A1(n27315), .A2(n27144), .B1(n27137), .B2(n21988), .ZN(
        n7309) );
  OAI22_X1 U20762 ( .A1(n27283), .A2(n27071), .B1(n27065), .B2(n21759), .ZN(
        n6914) );
  OAI22_X1 U20763 ( .A1(n27286), .A2(n27071), .B1(n27065), .B2(n21758), .ZN(
        n6915) );
  OAI22_X1 U20764 ( .A1(n27289), .A2(n27071), .B1(n27065), .B2(n21757), .ZN(
        n6916) );
  OAI22_X1 U20765 ( .A1(n27292), .A2(n27071), .B1(n27065), .B2(n21756), .ZN(
        n6917) );
  OAI22_X1 U20766 ( .A1(n27295), .A2(n27071), .B1(n27065), .B2(n21755), .ZN(
        n6918) );
  OAI22_X1 U20767 ( .A1(n27298), .A2(n27071), .B1(n27065), .B2(n21754), .ZN(
        n6919) );
  OAI22_X1 U20768 ( .A1(n27301), .A2(n27071), .B1(n27065), .B2(n21753), .ZN(
        n6920) );
  OAI22_X1 U20769 ( .A1(n27304), .A2(n27071), .B1(n27065), .B2(n21752), .ZN(
        n6921) );
  OAI22_X1 U20770 ( .A1(n27307), .A2(n27071), .B1(n27065), .B2(n21751), .ZN(
        n6922) );
  OAI22_X1 U20771 ( .A1(n27310), .A2(n27071), .B1(n27065), .B2(n21750), .ZN(
        n6923) );
  OAI22_X1 U20772 ( .A1(n27313), .A2(n27071), .B1(n27065), .B2(n21749), .ZN(
        n6924) );
  OAI22_X1 U20773 ( .A1(n27316), .A2(n27072), .B1(n27065), .B2(n21748), .ZN(
        n6925) );
  OAI22_X1 U20774 ( .A1(n27284), .A2(n26963), .B1(n26957), .B2(n21639), .ZN(
        n6338) );
  OAI22_X1 U20775 ( .A1(n27287), .A2(n26963), .B1(n26957), .B2(n21638), .ZN(
        n6339) );
  OAI22_X1 U20776 ( .A1(n27290), .A2(n26963), .B1(n26957), .B2(n21637), .ZN(
        n6340) );
  OAI22_X1 U20777 ( .A1(n27293), .A2(n26963), .B1(n26957), .B2(n21636), .ZN(
        n6341) );
  OAI22_X1 U20778 ( .A1(n27296), .A2(n26963), .B1(n26957), .B2(n21635), .ZN(
        n6342) );
  OAI22_X1 U20779 ( .A1(n27299), .A2(n26963), .B1(n26957), .B2(n21634), .ZN(
        n6343) );
  OAI22_X1 U20780 ( .A1(n27302), .A2(n26963), .B1(n26957), .B2(n21633), .ZN(
        n6344) );
  OAI22_X1 U20781 ( .A1(n27305), .A2(n26963), .B1(n26957), .B2(n21632), .ZN(
        n6345) );
  OAI22_X1 U20782 ( .A1(n27308), .A2(n26963), .B1(n26957), .B2(n21631), .ZN(
        n6346) );
  OAI22_X1 U20783 ( .A1(n27311), .A2(n26963), .B1(n26957), .B2(n21630), .ZN(
        n6347) );
  OAI22_X1 U20784 ( .A1(n27314), .A2(n26963), .B1(n26957), .B2(n21629), .ZN(
        n6348) );
  OAI22_X1 U20785 ( .A1(n27317), .A2(n26964), .B1(n26957), .B2(n21628), .ZN(
        n6349) );
  OAI22_X1 U20786 ( .A1(n27282), .A2(n27215), .B1(n27209), .B2(n21579), .ZN(
        n7682) );
  OAI22_X1 U20787 ( .A1(n27285), .A2(n27215), .B1(n27209), .B2(n21578), .ZN(
        n7683) );
  OAI22_X1 U20788 ( .A1(n27288), .A2(n27215), .B1(n27209), .B2(n21577), .ZN(
        n7684) );
  OAI22_X1 U20789 ( .A1(n27291), .A2(n27215), .B1(n27209), .B2(n21576), .ZN(
        n7685) );
  OAI22_X1 U20790 ( .A1(n27294), .A2(n27215), .B1(n27209), .B2(n21575), .ZN(
        n7686) );
  OAI22_X1 U20791 ( .A1(n27297), .A2(n27215), .B1(n27209), .B2(n21574), .ZN(
        n7687) );
  OAI22_X1 U20792 ( .A1(n27300), .A2(n27215), .B1(n27209), .B2(n21573), .ZN(
        n7688) );
  OAI22_X1 U20793 ( .A1(n27303), .A2(n27215), .B1(n27209), .B2(n21572), .ZN(
        n7689) );
  OAI22_X1 U20794 ( .A1(n27306), .A2(n27215), .B1(n27209), .B2(n21571), .ZN(
        n7690) );
  OAI22_X1 U20795 ( .A1(n27309), .A2(n27215), .B1(n27209), .B2(n21570), .ZN(
        n7691) );
  OAI22_X1 U20796 ( .A1(n27312), .A2(n27215), .B1(n27209), .B2(n21569), .ZN(
        n7692) );
  OAI22_X1 U20797 ( .A1(n27315), .A2(n27216), .B1(n27209), .B2(n21568), .ZN(
        n7693) );
  OAI22_X1 U20798 ( .A1(n27282), .A2(n27239), .B1(n27233), .B2(n21419), .ZN(
        n7810) );
  OAI22_X1 U20799 ( .A1(n27285), .A2(n27239), .B1(n27233), .B2(n21418), .ZN(
        n7811) );
  OAI22_X1 U20800 ( .A1(n27288), .A2(n27239), .B1(n27233), .B2(n21417), .ZN(
        n7812) );
  OAI22_X1 U20801 ( .A1(n27291), .A2(n27239), .B1(n27233), .B2(n21416), .ZN(
        n7813) );
  OAI22_X1 U20802 ( .A1(n27294), .A2(n27239), .B1(n27233), .B2(n21415), .ZN(
        n7814) );
  OAI22_X1 U20803 ( .A1(n27297), .A2(n27239), .B1(n27233), .B2(n21414), .ZN(
        n7815) );
  OAI22_X1 U20804 ( .A1(n27300), .A2(n27239), .B1(n27233), .B2(n21413), .ZN(
        n7816) );
  OAI22_X1 U20805 ( .A1(n27303), .A2(n27239), .B1(n27233), .B2(n21412), .ZN(
        n7817) );
  OAI22_X1 U20806 ( .A1(n27306), .A2(n27239), .B1(n27233), .B2(n21411), .ZN(
        n7818) );
  OAI22_X1 U20807 ( .A1(n27309), .A2(n27239), .B1(n27233), .B2(n21410), .ZN(
        n7819) );
  OAI22_X1 U20808 ( .A1(n27312), .A2(n27239), .B1(n27233), .B2(n21409), .ZN(
        n7820) );
  OAI22_X1 U20809 ( .A1(n27315), .A2(n27240), .B1(n27233), .B2(n21408), .ZN(
        n7821) );
  OAI22_X1 U20810 ( .A1(n27283), .A2(n26999), .B1(n26993), .B2(n21359), .ZN(
        n6530) );
  OAI22_X1 U20811 ( .A1(n27286), .A2(n26999), .B1(n26993), .B2(n21358), .ZN(
        n6531) );
  OAI22_X1 U20812 ( .A1(n27289), .A2(n26999), .B1(n26993), .B2(n21357), .ZN(
        n6532) );
  OAI22_X1 U20813 ( .A1(n27292), .A2(n26999), .B1(n26993), .B2(n21356), .ZN(
        n6533) );
  OAI22_X1 U20814 ( .A1(n27295), .A2(n26999), .B1(n26993), .B2(n21355), .ZN(
        n6534) );
  OAI22_X1 U20815 ( .A1(n27298), .A2(n26999), .B1(n26993), .B2(n21354), .ZN(
        n6535) );
  OAI22_X1 U20816 ( .A1(n27301), .A2(n26999), .B1(n26993), .B2(n21353), .ZN(
        n6536) );
  OAI22_X1 U20817 ( .A1(n27304), .A2(n26999), .B1(n26993), .B2(n21352), .ZN(
        n6537) );
  OAI22_X1 U20818 ( .A1(n27307), .A2(n26999), .B1(n26993), .B2(n21351), .ZN(
        n6538) );
  OAI22_X1 U20819 ( .A1(n27310), .A2(n26999), .B1(n26993), .B2(n21350), .ZN(
        n6539) );
  OAI22_X1 U20820 ( .A1(n27313), .A2(n26999), .B1(n26993), .B2(n21349), .ZN(
        n6540) );
  OAI22_X1 U20821 ( .A1(n27316), .A2(n27000), .B1(n26993), .B2(n21348), .ZN(
        n6541) );
  OAI22_X1 U20822 ( .A1(n27283), .A2(n26975), .B1(n26969), .B2(n21239), .ZN(
        n6402) );
  OAI22_X1 U20823 ( .A1(n27286), .A2(n26975), .B1(n26969), .B2(n21238), .ZN(
        n6403) );
  OAI22_X1 U20824 ( .A1(n27289), .A2(n26975), .B1(n26969), .B2(n21237), .ZN(
        n6404) );
  OAI22_X1 U20825 ( .A1(n27292), .A2(n26975), .B1(n26969), .B2(n21236), .ZN(
        n6405) );
  OAI22_X1 U20826 ( .A1(n27295), .A2(n26975), .B1(n26969), .B2(n21235), .ZN(
        n6406) );
  OAI22_X1 U20827 ( .A1(n27298), .A2(n26975), .B1(n26969), .B2(n21234), .ZN(
        n6407) );
  OAI22_X1 U20828 ( .A1(n27301), .A2(n26975), .B1(n26969), .B2(n21233), .ZN(
        n6408) );
  OAI22_X1 U20829 ( .A1(n27304), .A2(n26975), .B1(n26969), .B2(n21232), .ZN(
        n6409) );
  OAI22_X1 U20830 ( .A1(n27307), .A2(n26975), .B1(n26969), .B2(n21231), .ZN(
        n6410) );
  OAI22_X1 U20831 ( .A1(n27310), .A2(n26975), .B1(n26969), .B2(n21230), .ZN(
        n6411) );
  OAI22_X1 U20832 ( .A1(n27313), .A2(n26975), .B1(n26969), .B2(n21229), .ZN(
        n6412) );
  OAI22_X1 U20833 ( .A1(n27316), .A2(n26976), .B1(n26969), .B2(n21228), .ZN(
        n6413) );
  OAI22_X1 U20834 ( .A1(n27283), .A2(n27107), .B1(n27101), .B2(n20834), .ZN(
        n7106) );
  OAI22_X1 U20835 ( .A1(n27286), .A2(n27107), .B1(n27101), .B2(n20833), .ZN(
        n7107) );
  OAI22_X1 U20836 ( .A1(n27289), .A2(n27107), .B1(n27101), .B2(n20832), .ZN(
        n7108) );
  OAI22_X1 U20837 ( .A1(n27292), .A2(n27107), .B1(n27101), .B2(n20831), .ZN(
        n7109) );
  OAI22_X1 U20838 ( .A1(n27295), .A2(n27107), .B1(n27101), .B2(n20830), .ZN(
        n7110) );
  OAI22_X1 U20839 ( .A1(n27298), .A2(n27107), .B1(n27101), .B2(n20829), .ZN(
        n7111) );
  OAI22_X1 U20840 ( .A1(n27301), .A2(n27107), .B1(n27101), .B2(n20828), .ZN(
        n7112) );
  OAI22_X1 U20841 ( .A1(n27304), .A2(n27107), .B1(n27101), .B2(n20827), .ZN(
        n7113) );
  OAI22_X1 U20842 ( .A1(n27307), .A2(n27107), .B1(n27101), .B2(n20826), .ZN(
        n7114) );
  OAI22_X1 U20843 ( .A1(n27310), .A2(n27107), .B1(n27101), .B2(n20825), .ZN(
        n7115) );
  OAI22_X1 U20844 ( .A1(n27313), .A2(n27107), .B1(n27101), .B2(n20824), .ZN(
        n7116) );
  OAI22_X1 U20845 ( .A1(n27316), .A2(n27108), .B1(n27101), .B2(n20823), .ZN(
        n7117) );
  OAI22_X1 U20846 ( .A1(n27282), .A2(n27131), .B1(n27125), .B2(n20771), .ZN(
        n7234) );
  OAI22_X1 U20847 ( .A1(n27285), .A2(n27131), .B1(n27125), .B2(n20770), .ZN(
        n7235) );
  OAI22_X1 U20848 ( .A1(n27288), .A2(n27131), .B1(n27125), .B2(n20769), .ZN(
        n7236) );
  OAI22_X1 U20849 ( .A1(n27291), .A2(n27131), .B1(n27125), .B2(n20768), .ZN(
        n7237) );
  OAI22_X1 U20850 ( .A1(n27294), .A2(n27131), .B1(n27125), .B2(n20767), .ZN(
        n7238) );
  OAI22_X1 U20851 ( .A1(n27297), .A2(n27131), .B1(n27125), .B2(n20766), .ZN(
        n7239) );
  OAI22_X1 U20852 ( .A1(n27300), .A2(n27131), .B1(n27125), .B2(n20765), .ZN(
        n7240) );
  OAI22_X1 U20853 ( .A1(n27303), .A2(n27131), .B1(n27125), .B2(n20764), .ZN(
        n7241) );
  OAI22_X1 U20854 ( .A1(n27306), .A2(n27131), .B1(n27125), .B2(n20763), .ZN(
        n7242) );
  OAI22_X1 U20855 ( .A1(n27309), .A2(n27131), .B1(n27125), .B2(n20762), .ZN(
        n7243) );
  OAI22_X1 U20856 ( .A1(n27312), .A2(n27131), .B1(n27125), .B2(n20761), .ZN(
        n7244) );
  OAI22_X1 U20857 ( .A1(n27315), .A2(n27132), .B1(n27125), .B2(n20760), .ZN(
        n7245) );
  NAND2_X1 U20858 ( .A1(n25136), .A2(n25137), .ZN(n5763) );
  NOR4_X1 U20859 ( .A1(n25156), .A2(n25157), .A3(n25158), .A4(n25159), .ZN(
        n25136) );
  NOR4_X1 U20860 ( .A1(n25138), .A2(n25139), .A3(n25140), .A4(n25141), .ZN(
        n25137) );
  OAI221_X1 U20861 ( .B1(n21579), .B2(n26495), .C1(n21419), .C2(n26489), .A(
        n25162), .ZN(n25157) );
  NAND2_X1 U20862 ( .A1(n25118), .A2(n25119), .ZN(n5765) );
  NOR4_X1 U20863 ( .A1(n25128), .A2(n25129), .A3(n25130), .A4(n25131), .ZN(
        n25118) );
  NOR4_X1 U20864 ( .A1(n25120), .A2(n25121), .A3(n25122), .A4(n25123), .ZN(
        n25119) );
  OAI221_X1 U20865 ( .B1(n21578), .B2(n26495), .C1(n21418), .C2(n26489), .A(
        n25134), .ZN(n25129) );
  NAND2_X1 U20866 ( .A1(n25100), .A2(n25101), .ZN(n5767) );
  NOR4_X1 U20867 ( .A1(n25110), .A2(n25111), .A3(n25112), .A4(n25113), .ZN(
        n25100) );
  NOR4_X1 U20868 ( .A1(n25102), .A2(n25103), .A3(n25104), .A4(n25105), .ZN(
        n25101) );
  OAI221_X1 U20869 ( .B1(n21577), .B2(n26495), .C1(n21417), .C2(n26489), .A(
        n25116), .ZN(n25111) );
  NAND2_X1 U20870 ( .A1(n25082), .A2(n25083), .ZN(n5769) );
  NOR4_X1 U20871 ( .A1(n25092), .A2(n25093), .A3(n25094), .A4(n25095), .ZN(
        n25082) );
  NOR4_X1 U20872 ( .A1(n25084), .A2(n25085), .A3(n25086), .A4(n25087), .ZN(
        n25083) );
  OAI221_X1 U20873 ( .B1(n21576), .B2(n26495), .C1(n21416), .C2(n26489), .A(
        n25098), .ZN(n25093) );
  NAND2_X1 U20874 ( .A1(n25064), .A2(n25065), .ZN(n5771) );
  NOR4_X1 U20875 ( .A1(n25074), .A2(n25075), .A3(n25076), .A4(n25077), .ZN(
        n25064) );
  NOR4_X1 U20876 ( .A1(n25066), .A2(n25067), .A3(n25068), .A4(n25069), .ZN(
        n25065) );
  OAI221_X1 U20877 ( .B1(n21575), .B2(n26495), .C1(n21415), .C2(n26489), .A(
        n25080), .ZN(n25075) );
  NAND2_X1 U20878 ( .A1(n25046), .A2(n25047), .ZN(n5773) );
  NOR4_X1 U20879 ( .A1(n25056), .A2(n25057), .A3(n25058), .A4(n25059), .ZN(
        n25046) );
  NOR4_X1 U20880 ( .A1(n25048), .A2(n25049), .A3(n25050), .A4(n25051), .ZN(
        n25047) );
  OAI221_X1 U20881 ( .B1(n21574), .B2(n26495), .C1(n21414), .C2(n26489), .A(
        n25062), .ZN(n25057) );
  NAND2_X1 U20882 ( .A1(n25028), .A2(n25029), .ZN(n5775) );
  NOR4_X1 U20883 ( .A1(n25038), .A2(n25039), .A3(n25040), .A4(n25041), .ZN(
        n25028) );
  NOR4_X1 U20884 ( .A1(n25030), .A2(n25031), .A3(n25032), .A4(n25033), .ZN(
        n25029) );
  OAI221_X1 U20885 ( .B1(n21573), .B2(n26495), .C1(n21413), .C2(n26489), .A(
        n25044), .ZN(n25039) );
  NAND2_X1 U20886 ( .A1(n25010), .A2(n25011), .ZN(n5777) );
  NOR4_X1 U20887 ( .A1(n25020), .A2(n25021), .A3(n25022), .A4(n25023), .ZN(
        n25010) );
  NOR4_X1 U20888 ( .A1(n25012), .A2(n25013), .A3(n25014), .A4(n25015), .ZN(
        n25011) );
  OAI221_X1 U20889 ( .B1(n21572), .B2(n26495), .C1(n21412), .C2(n26489), .A(
        n25026), .ZN(n25021) );
  NAND2_X1 U20890 ( .A1(n24992), .A2(n24993), .ZN(n5779) );
  NOR4_X1 U20891 ( .A1(n25002), .A2(n25003), .A3(n25004), .A4(n25005), .ZN(
        n24992) );
  NOR4_X1 U20892 ( .A1(n24994), .A2(n24995), .A3(n24996), .A4(n24997), .ZN(
        n24993) );
  OAI221_X1 U20893 ( .B1(n21571), .B2(n26495), .C1(n21411), .C2(n26489), .A(
        n25008), .ZN(n25003) );
  NAND2_X1 U20894 ( .A1(n24974), .A2(n24975), .ZN(n5781) );
  NOR4_X1 U20895 ( .A1(n24984), .A2(n24985), .A3(n24986), .A4(n24987), .ZN(
        n24974) );
  NOR4_X1 U20896 ( .A1(n24976), .A2(n24977), .A3(n24978), .A4(n24979), .ZN(
        n24975) );
  OAI221_X1 U20897 ( .B1(n21570), .B2(n26495), .C1(n21410), .C2(n26489), .A(
        n24990), .ZN(n24985) );
  NAND2_X1 U20898 ( .A1(n24956), .A2(n24957), .ZN(n5783) );
  NOR4_X1 U20899 ( .A1(n24966), .A2(n24967), .A3(n24968), .A4(n24969), .ZN(
        n24956) );
  NOR4_X1 U20900 ( .A1(n24958), .A2(n24959), .A3(n24960), .A4(n24961), .ZN(
        n24957) );
  OAI221_X1 U20901 ( .B1(n21569), .B2(n26495), .C1(n21409), .C2(n26489), .A(
        n24972), .ZN(n24967) );
  NAND2_X1 U20902 ( .A1(n24938), .A2(n24939), .ZN(n5785) );
  NOR4_X1 U20903 ( .A1(n24948), .A2(n24949), .A3(n24950), .A4(n24951), .ZN(
        n24938) );
  NOR4_X1 U20904 ( .A1(n24940), .A2(n24941), .A3(n24942), .A4(n24943), .ZN(
        n24939) );
  OAI221_X1 U20905 ( .B1(n21568), .B2(n26495), .C1(n21408), .C2(n26489), .A(
        n24954), .ZN(n24949) );
  NAND2_X1 U20906 ( .A1(n24920), .A2(n24921), .ZN(n5787) );
  NOR4_X1 U20907 ( .A1(n24930), .A2(n24931), .A3(n24932), .A4(n24933), .ZN(
        n24920) );
  NOR4_X1 U20908 ( .A1(n24922), .A2(n24923), .A3(n24924), .A4(n24925), .ZN(
        n24921) );
  OAI221_X1 U20909 ( .B1(n21567), .B2(n26496), .C1(n21407), .C2(n26490), .A(
        n24936), .ZN(n24931) );
  NAND2_X1 U20910 ( .A1(n24902), .A2(n24903), .ZN(n5789) );
  NOR4_X1 U20911 ( .A1(n24912), .A2(n24913), .A3(n24914), .A4(n24915), .ZN(
        n24902) );
  NOR4_X1 U20912 ( .A1(n24904), .A2(n24905), .A3(n24906), .A4(n24907), .ZN(
        n24903) );
  OAI221_X1 U20913 ( .B1(n21566), .B2(n26496), .C1(n21406), .C2(n26490), .A(
        n24918), .ZN(n24913) );
  NAND2_X1 U20914 ( .A1(n24884), .A2(n24885), .ZN(n5791) );
  NOR4_X1 U20915 ( .A1(n24894), .A2(n24895), .A3(n24896), .A4(n24897), .ZN(
        n24884) );
  NOR4_X1 U20916 ( .A1(n24886), .A2(n24887), .A3(n24888), .A4(n24889), .ZN(
        n24885) );
  OAI221_X1 U20917 ( .B1(n21565), .B2(n26496), .C1(n21405), .C2(n26490), .A(
        n24900), .ZN(n24895) );
  NAND2_X1 U20918 ( .A1(n24866), .A2(n24867), .ZN(n5793) );
  NOR4_X1 U20919 ( .A1(n24876), .A2(n24877), .A3(n24878), .A4(n24879), .ZN(
        n24866) );
  NOR4_X1 U20920 ( .A1(n24868), .A2(n24869), .A3(n24870), .A4(n24871), .ZN(
        n24867) );
  OAI221_X1 U20921 ( .B1(n21564), .B2(n26496), .C1(n21404), .C2(n26490), .A(
        n24882), .ZN(n24877) );
  NAND2_X1 U20922 ( .A1(n24848), .A2(n24849), .ZN(n5795) );
  NOR4_X1 U20923 ( .A1(n24858), .A2(n24859), .A3(n24860), .A4(n24861), .ZN(
        n24848) );
  NOR4_X1 U20924 ( .A1(n24850), .A2(n24851), .A3(n24852), .A4(n24853), .ZN(
        n24849) );
  OAI221_X1 U20925 ( .B1(n21563), .B2(n26496), .C1(n21403), .C2(n26490), .A(
        n24864), .ZN(n24859) );
  NAND2_X1 U20926 ( .A1(n24830), .A2(n24831), .ZN(n5797) );
  NOR4_X1 U20927 ( .A1(n24840), .A2(n24841), .A3(n24842), .A4(n24843), .ZN(
        n24830) );
  NOR4_X1 U20928 ( .A1(n24832), .A2(n24833), .A3(n24834), .A4(n24835), .ZN(
        n24831) );
  OAI221_X1 U20929 ( .B1(n21562), .B2(n26496), .C1(n21402), .C2(n26490), .A(
        n24846), .ZN(n24841) );
  NAND2_X1 U20930 ( .A1(n24812), .A2(n24813), .ZN(n5799) );
  NOR4_X1 U20931 ( .A1(n24822), .A2(n24823), .A3(n24824), .A4(n24825), .ZN(
        n24812) );
  NOR4_X1 U20932 ( .A1(n24814), .A2(n24815), .A3(n24816), .A4(n24817), .ZN(
        n24813) );
  OAI221_X1 U20933 ( .B1(n21561), .B2(n26496), .C1(n21401), .C2(n26490), .A(
        n24828), .ZN(n24823) );
  NAND2_X1 U20934 ( .A1(n24794), .A2(n24795), .ZN(n5801) );
  NOR4_X1 U20935 ( .A1(n24804), .A2(n24805), .A3(n24806), .A4(n24807), .ZN(
        n24794) );
  NOR4_X1 U20936 ( .A1(n24796), .A2(n24797), .A3(n24798), .A4(n24799), .ZN(
        n24795) );
  OAI221_X1 U20937 ( .B1(n21560), .B2(n26496), .C1(n21400), .C2(n26490), .A(
        n24810), .ZN(n24805) );
  NAND2_X1 U20938 ( .A1(n24776), .A2(n24777), .ZN(n5803) );
  NOR4_X1 U20939 ( .A1(n24786), .A2(n24787), .A3(n24788), .A4(n24789), .ZN(
        n24776) );
  NOR4_X1 U20940 ( .A1(n24778), .A2(n24779), .A3(n24780), .A4(n24781), .ZN(
        n24777) );
  OAI221_X1 U20941 ( .B1(n21559), .B2(n26496), .C1(n21399), .C2(n26490), .A(
        n24792), .ZN(n24787) );
  NAND2_X1 U20942 ( .A1(n24758), .A2(n24759), .ZN(n5805) );
  NOR4_X1 U20943 ( .A1(n24768), .A2(n24769), .A3(n24770), .A4(n24771), .ZN(
        n24758) );
  NOR4_X1 U20944 ( .A1(n24760), .A2(n24761), .A3(n24762), .A4(n24763), .ZN(
        n24759) );
  OAI221_X1 U20945 ( .B1(n21558), .B2(n26496), .C1(n21398), .C2(n26490), .A(
        n24774), .ZN(n24769) );
  NAND2_X1 U20946 ( .A1(n24740), .A2(n24741), .ZN(n5807) );
  NOR4_X1 U20947 ( .A1(n24750), .A2(n24751), .A3(n24752), .A4(n24753), .ZN(
        n24740) );
  NOR4_X1 U20948 ( .A1(n24742), .A2(n24743), .A3(n24744), .A4(n24745), .ZN(
        n24741) );
  OAI221_X1 U20949 ( .B1(n21557), .B2(n26496), .C1(n21397), .C2(n26490), .A(
        n24756), .ZN(n24751) );
  NAND2_X1 U20950 ( .A1(n24722), .A2(n24723), .ZN(n5809) );
  NOR4_X1 U20951 ( .A1(n24732), .A2(n24733), .A3(n24734), .A4(n24735), .ZN(
        n24722) );
  NOR4_X1 U20952 ( .A1(n24724), .A2(n24725), .A3(n24726), .A4(n24727), .ZN(
        n24723) );
  OAI221_X1 U20953 ( .B1(n21556), .B2(n26496), .C1(n21396), .C2(n26490), .A(
        n24738), .ZN(n24733) );
  NAND2_X1 U20954 ( .A1(n24704), .A2(n24705), .ZN(n5811) );
  NOR4_X1 U20955 ( .A1(n24714), .A2(n24715), .A3(n24716), .A4(n24717), .ZN(
        n24704) );
  NOR4_X1 U20956 ( .A1(n24706), .A2(n24707), .A3(n24708), .A4(n24709), .ZN(
        n24705) );
  OAI221_X1 U20957 ( .B1(n21555), .B2(n26497), .C1(n21395), .C2(n26491), .A(
        n24720), .ZN(n24715) );
  NAND2_X1 U20958 ( .A1(n24686), .A2(n24687), .ZN(n5813) );
  NOR4_X1 U20959 ( .A1(n24696), .A2(n24697), .A3(n24698), .A4(n24699), .ZN(
        n24686) );
  NOR4_X1 U20960 ( .A1(n24688), .A2(n24689), .A3(n24690), .A4(n24691), .ZN(
        n24687) );
  OAI221_X1 U20961 ( .B1(n21554), .B2(n26497), .C1(n21394), .C2(n26491), .A(
        n24702), .ZN(n24697) );
  NAND2_X1 U20962 ( .A1(n24668), .A2(n24669), .ZN(n5815) );
  NOR4_X1 U20963 ( .A1(n24678), .A2(n24679), .A3(n24680), .A4(n24681), .ZN(
        n24668) );
  NOR4_X1 U20964 ( .A1(n24670), .A2(n24671), .A3(n24672), .A4(n24673), .ZN(
        n24669) );
  OAI221_X1 U20965 ( .B1(n21553), .B2(n26497), .C1(n21393), .C2(n26491), .A(
        n24684), .ZN(n24679) );
  NAND2_X1 U20966 ( .A1(n24650), .A2(n24651), .ZN(n5817) );
  NOR4_X1 U20967 ( .A1(n24660), .A2(n24661), .A3(n24662), .A4(n24663), .ZN(
        n24650) );
  NOR4_X1 U20968 ( .A1(n24652), .A2(n24653), .A3(n24654), .A4(n24655), .ZN(
        n24651) );
  OAI221_X1 U20969 ( .B1(n21552), .B2(n26497), .C1(n21392), .C2(n26491), .A(
        n24666), .ZN(n24661) );
  NAND2_X1 U20970 ( .A1(n24632), .A2(n24633), .ZN(n5819) );
  NOR4_X1 U20971 ( .A1(n24642), .A2(n24643), .A3(n24644), .A4(n24645), .ZN(
        n24632) );
  NOR4_X1 U20972 ( .A1(n24634), .A2(n24635), .A3(n24636), .A4(n24637), .ZN(
        n24633) );
  OAI221_X1 U20973 ( .B1(n21551), .B2(n26497), .C1(n21391), .C2(n26491), .A(
        n24648), .ZN(n24643) );
  NAND2_X1 U20974 ( .A1(n24614), .A2(n24615), .ZN(n5821) );
  NOR4_X1 U20975 ( .A1(n24624), .A2(n24625), .A3(n24626), .A4(n24627), .ZN(
        n24614) );
  NOR4_X1 U20976 ( .A1(n24616), .A2(n24617), .A3(n24618), .A4(n24619), .ZN(
        n24615) );
  OAI221_X1 U20977 ( .B1(n21550), .B2(n26497), .C1(n21390), .C2(n26491), .A(
        n24630), .ZN(n24625) );
  NAND2_X1 U20978 ( .A1(n24596), .A2(n24597), .ZN(n5823) );
  NOR4_X1 U20979 ( .A1(n24606), .A2(n24607), .A3(n24608), .A4(n24609), .ZN(
        n24596) );
  NOR4_X1 U20980 ( .A1(n24598), .A2(n24599), .A3(n24600), .A4(n24601), .ZN(
        n24597) );
  OAI221_X1 U20981 ( .B1(n21549), .B2(n26497), .C1(n21389), .C2(n26491), .A(
        n24612), .ZN(n24607) );
  NAND2_X1 U20982 ( .A1(n24578), .A2(n24579), .ZN(n5825) );
  NOR4_X1 U20983 ( .A1(n24588), .A2(n24589), .A3(n24590), .A4(n24591), .ZN(
        n24578) );
  NOR4_X1 U20984 ( .A1(n24580), .A2(n24581), .A3(n24582), .A4(n24583), .ZN(
        n24579) );
  OAI221_X1 U20985 ( .B1(n21548), .B2(n26497), .C1(n21388), .C2(n26491), .A(
        n24594), .ZN(n24589) );
  NAND2_X1 U20986 ( .A1(n24560), .A2(n24561), .ZN(n5827) );
  NOR4_X1 U20987 ( .A1(n24570), .A2(n24571), .A3(n24572), .A4(n24573), .ZN(
        n24560) );
  NOR4_X1 U20988 ( .A1(n24562), .A2(n24563), .A3(n24564), .A4(n24565), .ZN(
        n24561) );
  OAI221_X1 U20989 ( .B1(n21547), .B2(n26497), .C1(n21387), .C2(n26491), .A(
        n24576), .ZN(n24571) );
  NAND2_X1 U20990 ( .A1(n24542), .A2(n24543), .ZN(n5829) );
  NOR4_X1 U20991 ( .A1(n24552), .A2(n24553), .A3(n24554), .A4(n24555), .ZN(
        n24542) );
  NOR4_X1 U20992 ( .A1(n24544), .A2(n24545), .A3(n24546), .A4(n24547), .ZN(
        n24543) );
  OAI221_X1 U20993 ( .B1(n21546), .B2(n26497), .C1(n21386), .C2(n26491), .A(
        n24558), .ZN(n24553) );
  NAND2_X1 U20994 ( .A1(n24524), .A2(n24525), .ZN(n5831) );
  NOR4_X1 U20995 ( .A1(n24534), .A2(n24535), .A3(n24536), .A4(n24537), .ZN(
        n24524) );
  NOR4_X1 U20996 ( .A1(n24526), .A2(n24527), .A3(n24528), .A4(n24529), .ZN(
        n24525) );
  OAI221_X1 U20997 ( .B1(n21545), .B2(n26497), .C1(n21385), .C2(n26491), .A(
        n24540), .ZN(n24535) );
  NAND2_X1 U20998 ( .A1(n24506), .A2(n24507), .ZN(n5833) );
  NOR4_X1 U20999 ( .A1(n24516), .A2(n24517), .A3(n24518), .A4(n24519), .ZN(
        n24506) );
  NOR4_X1 U21000 ( .A1(n24508), .A2(n24509), .A3(n24510), .A4(n24511), .ZN(
        n24507) );
  OAI221_X1 U21001 ( .B1(n21544), .B2(n26497), .C1(n21384), .C2(n26491), .A(
        n24522), .ZN(n24517) );
  NAND2_X1 U21002 ( .A1(n24488), .A2(n24489), .ZN(n5835) );
  NOR4_X1 U21003 ( .A1(n24498), .A2(n24499), .A3(n24500), .A4(n24501), .ZN(
        n24488) );
  NOR4_X1 U21004 ( .A1(n24490), .A2(n24491), .A3(n24492), .A4(n24493), .ZN(
        n24489) );
  OAI221_X1 U21005 ( .B1(n21543), .B2(n26498), .C1(n21383), .C2(n26492), .A(
        n24504), .ZN(n24499) );
  NAND2_X1 U21006 ( .A1(n24470), .A2(n24471), .ZN(n5837) );
  NOR4_X1 U21007 ( .A1(n24480), .A2(n24481), .A3(n24482), .A4(n24483), .ZN(
        n24470) );
  NOR4_X1 U21008 ( .A1(n24472), .A2(n24473), .A3(n24474), .A4(n24475), .ZN(
        n24471) );
  OAI221_X1 U21009 ( .B1(n21542), .B2(n26498), .C1(n21382), .C2(n26492), .A(
        n24486), .ZN(n24481) );
  NAND2_X1 U21010 ( .A1(n24452), .A2(n24453), .ZN(n5839) );
  NOR4_X1 U21011 ( .A1(n24462), .A2(n24463), .A3(n24464), .A4(n24465), .ZN(
        n24452) );
  NOR4_X1 U21012 ( .A1(n24454), .A2(n24455), .A3(n24456), .A4(n24457), .ZN(
        n24453) );
  OAI221_X1 U21013 ( .B1(n21541), .B2(n26498), .C1(n21381), .C2(n26492), .A(
        n24468), .ZN(n24463) );
  NAND2_X1 U21014 ( .A1(n24434), .A2(n24435), .ZN(n5841) );
  NOR4_X1 U21015 ( .A1(n24444), .A2(n24445), .A3(n24446), .A4(n24447), .ZN(
        n24434) );
  NOR4_X1 U21016 ( .A1(n24436), .A2(n24437), .A3(n24438), .A4(n24439), .ZN(
        n24435) );
  OAI221_X1 U21017 ( .B1(n21540), .B2(n26498), .C1(n21380), .C2(n26492), .A(
        n24450), .ZN(n24445) );
  NAND2_X1 U21018 ( .A1(n24416), .A2(n24417), .ZN(n5843) );
  NOR4_X1 U21019 ( .A1(n24426), .A2(n24427), .A3(n24428), .A4(n24429), .ZN(
        n24416) );
  NOR4_X1 U21020 ( .A1(n24418), .A2(n24419), .A3(n24420), .A4(n24421), .ZN(
        n24417) );
  OAI221_X1 U21021 ( .B1(n21539), .B2(n26498), .C1(n21379), .C2(n26492), .A(
        n24432), .ZN(n24427) );
  NAND2_X1 U21022 ( .A1(n24398), .A2(n24399), .ZN(n5845) );
  NOR4_X1 U21023 ( .A1(n24408), .A2(n24409), .A3(n24410), .A4(n24411), .ZN(
        n24398) );
  NOR4_X1 U21024 ( .A1(n24400), .A2(n24401), .A3(n24402), .A4(n24403), .ZN(
        n24399) );
  OAI221_X1 U21025 ( .B1(n21538), .B2(n26498), .C1(n21378), .C2(n26492), .A(
        n24414), .ZN(n24409) );
  NAND2_X1 U21026 ( .A1(n24380), .A2(n24381), .ZN(n5847) );
  NOR4_X1 U21027 ( .A1(n24390), .A2(n24391), .A3(n24392), .A4(n24393), .ZN(
        n24380) );
  NOR4_X1 U21028 ( .A1(n24382), .A2(n24383), .A3(n24384), .A4(n24385), .ZN(
        n24381) );
  OAI221_X1 U21029 ( .B1(n21537), .B2(n26498), .C1(n21377), .C2(n26492), .A(
        n24396), .ZN(n24391) );
  NAND2_X1 U21030 ( .A1(n24362), .A2(n24363), .ZN(n5849) );
  NOR4_X1 U21031 ( .A1(n24372), .A2(n24373), .A3(n24374), .A4(n24375), .ZN(
        n24362) );
  NOR4_X1 U21032 ( .A1(n24364), .A2(n24365), .A3(n24366), .A4(n24367), .ZN(
        n24363) );
  OAI221_X1 U21033 ( .B1(n21536), .B2(n26498), .C1(n21376), .C2(n26492), .A(
        n24378), .ZN(n24373) );
  NAND2_X1 U21034 ( .A1(n24344), .A2(n24345), .ZN(n5851) );
  NOR4_X1 U21035 ( .A1(n24354), .A2(n24355), .A3(n24356), .A4(n24357), .ZN(
        n24344) );
  NOR4_X1 U21036 ( .A1(n24346), .A2(n24347), .A3(n24348), .A4(n24349), .ZN(
        n24345) );
  OAI221_X1 U21037 ( .B1(n21535), .B2(n26498), .C1(n21375), .C2(n26492), .A(
        n24360), .ZN(n24355) );
  NAND2_X1 U21038 ( .A1(n24326), .A2(n24327), .ZN(n5853) );
  NOR4_X1 U21039 ( .A1(n24336), .A2(n24337), .A3(n24338), .A4(n24339), .ZN(
        n24326) );
  NOR4_X1 U21040 ( .A1(n24328), .A2(n24329), .A3(n24330), .A4(n24331), .ZN(
        n24327) );
  OAI221_X1 U21041 ( .B1(n21534), .B2(n26498), .C1(n21374), .C2(n26492), .A(
        n24342), .ZN(n24337) );
  NAND2_X1 U21042 ( .A1(n24308), .A2(n24309), .ZN(n5855) );
  NOR4_X1 U21043 ( .A1(n24318), .A2(n24319), .A3(n24320), .A4(n24321), .ZN(
        n24308) );
  NOR4_X1 U21044 ( .A1(n24310), .A2(n24311), .A3(n24312), .A4(n24313), .ZN(
        n24309) );
  OAI221_X1 U21045 ( .B1(n21533), .B2(n26498), .C1(n21373), .C2(n26492), .A(
        n24324), .ZN(n24319) );
  NAND2_X1 U21046 ( .A1(n24290), .A2(n24291), .ZN(n5857) );
  NOR4_X1 U21047 ( .A1(n24300), .A2(n24301), .A3(n24302), .A4(n24303), .ZN(
        n24290) );
  NOR4_X1 U21048 ( .A1(n24292), .A2(n24293), .A3(n24294), .A4(n24295), .ZN(
        n24291) );
  OAI221_X1 U21049 ( .B1(n21532), .B2(n26498), .C1(n21372), .C2(n26492), .A(
        n24306), .ZN(n24301) );
  NAND2_X1 U21050 ( .A1(n23937), .A2(n23938), .ZN(n5891) );
  NOR4_X1 U21051 ( .A1(n23957), .A2(n23958), .A3(n23959), .A4(n23960), .ZN(
        n23937) );
  NOR4_X1 U21052 ( .A1(n23939), .A2(n23940), .A3(n23941), .A4(n23942), .ZN(
        n23938) );
  OAI221_X1 U21053 ( .B1(n21579), .B2(n26720), .C1(n21419), .C2(n26714), .A(
        n23963), .ZN(n23958) );
  NAND2_X1 U21054 ( .A1(n23919), .A2(n23920), .ZN(n5893) );
  NOR4_X1 U21055 ( .A1(n23929), .A2(n23930), .A3(n23931), .A4(n23932), .ZN(
        n23919) );
  NOR4_X1 U21056 ( .A1(n23921), .A2(n23922), .A3(n23923), .A4(n23924), .ZN(
        n23920) );
  OAI221_X1 U21057 ( .B1(n21578), .B2(n26720), .C1(n21418), .C2(n26714), .A(
        n23935), .ZN(n23930) );
  NAND2_X1 U21058 ( .A1(n23901), .A2(n23902), .ZN(n5895) );
  NOR4_X1 U21059 ( .A1(n23911), .A2(n23912), .A3(n23913), .A4(n23914), .ZN(
        n23901) );
  NOR4_X1 U21060 ( .A1(n23903), .A2(n23904), .A3(n23905), .A4(n23906), .ZN(
        n23902) );
  OAI221_X1 U21061 ( .B1(n21577), .B2(n26720), .C1(n21417), .C2(n26714), .A(
        n23917), .ZN(n23912) );
  NAND2_X1 U21062 ( .A1(n23883), .A2(n23884), .ZN(n5897) );
  NOR4_X1 U21063 ( .A1(n23893), .A2(n23894), .A3(n23895), .A4(n23896), .ZN(
        n23883) );
  NOR4_X1 U21064 ( .A1(n23885), .A2(n23886), .A3(n23887), .A4(n23888), .ZN(
        n23884) );
  OAI221_X1 U21065 ( .B1(n21576), .B2(n26720), .C1(n21416), .C2(n26714), .A(
        n23899), .ZN(n23894) );
  NAND2_X1 U21066 ( .A1(n23865), .A2(n23866), .ZN(n5899) );
  NOR4_X1 U21067 ( .A1(n23875), .A2(n23876), .A3(n23877), .A4(n23878), .ZN(
        n23865) );
  NOR4_X1 U21068 ( .A1(n23867), .A2(n23868), .A3(n23869), .A4(n23870), .ZN(
        n23866) );
  OAI221_X1 U21069 ( .B1(n21575), .B2(n26720), .C1(n21415), .C2(n26714), .A(
        n23881), .ZN(n23876) );
  NAND2_X1 U21070 ( .A1(n23847), .A2(n23848), .ZN(n5901) );
  NOR4_X1 U21071 ( .A1(n23857), .A2(n23858), .A3(n23859), .A4(n23860), .ZN(
        n23847) );
  NOR4_X1 U21072 ( .A1(n23849), .A2(n23850), .A3(n23851), .A4(n23852), .ZN(
        n23848) );
  OAI221_X1 U21073 ( .B1(n21574), .B2(n26720), .C1(n21414), .C2(n26714), .A(
        n23863), .ZN(n23858) );
  NAND2_X1 U21074 ( .A1(n23829), .A2(n23830), .ZN(n5903) );
  NOR4_X1 U21075 ( .A1(n23839), .A2(n23840), .A3(n23841), .A4(n23842), .ZN(
        n23829) );
  NOR4_X1 U21076 ( .A1(n23831), .A2(n23832), .A3(n23833), .A4(n23834), .ZN(
        n23830) );
  OAI221_X1 U21077 ( .B1(n21573), .B2(n26720), .C1(n21413), .C2(n26714), .A(
        n23845), .ZN(n23840) );
  NAND2_X1 U21078 ( .A1(n23811), .A2(n23812), .ZN(n5905) );
  NOR4_X1 U21079 ( .A1(n23821), .A2(n23822), .A3(n23823), .A4(n23824), .ZN(
        n23811) );
  NOR4_X1 U21080 ( .A1(n23813), .A2(n23814), .A3(n23815), .A4(n23816), .ZN(
        n23812) );
  OAI221_X1 U21081 ( .B1(n21572), .B2(n26720), .C1(n21412), .C2(n26714), .A(
        n23827), .ZN(n23822) );
  NAND2_X1 U21082 ( .A1(n23793), .A2(n23794), .ZN(n5907) );
  NOR4_X1 U21083 ( .A1(n23803), .A2(n23804), .A3(n23805), .A4(n23806), .ZN(
        n23793) );
  NOR4_X1 U21084 ( .A1(n23795), .A2(n23796), .A3(n23797), .A4(n23798), .ZN(
        n23794) );
  OAI221_X1 U21085 ( .B1(n21571), .B2(n26720), .C1(n21411), .C2(n26714), .A(
        n23809), .ZN(n23804) );
  NAND2_X1 U21086 ( .A1(n23775), .A2(n23776), .ZN(n5909) );
  NOR4_X1 U21087 ( .A1(n23785), .A2(n23786), .A3(n23787), .A4(n23788), .ZN(
        n23775) );
  NOR4_X1 U21088 ( .A1(n23777), .A2(n23778), .A3(n23779), .A4(n23780), .ZN(
        n23776) );
  OAI221_X1 U21089 ( .B1(n21570), .B2(n26720), .C1(n21410), .C2(n26714), .A(
        n23791), .ZN(n23786) );
  NAND2_X1 U21090 ( .A1(n23757), .A2(n23758), .ZN(n5911) );
  NOR4_X1 U21091 ( .A1(n23767), .A2(n23768), .A3(n23769), .A4(n23770), .ZN(
        n23757) );
  NOR4_X1 U21092 ( .A1(n23759), .A2(n23760), .A3(n23761), .A4(n23762), .ZN(
        n23758) );
  OAI221_X1 U21093 ( .B1(n21569), .B2(n26720), .C1(n21409), .C2(n26714), .A(
        n23773), .ZN(n23768) );
  NAND2_X1 U21094 ( .A1(n23739), .A2(n23740), .ZN(n5913) );
  NOR4_X1 U21095 ( .A1(n23749), .A2(n23750), .A3(n23751), .A4(n23752), .ZN(
        n23739) );
  NOR4_X1 U21096 ( .A1(n23741), .A2(n23742), .A3(n23743), .A4(n23744), .ZN(
        n23740) );
  OAI221_X1 U21097 ( .B1(n21568), .B2(n26720), .C1(n21408), .C2(n26714), .A(
        n23755), .ZN(n23750) );
  NAND2_X1 U21098 ( .A1(n23721), .A2(n23722), .ZN(n5915) );
  NOR4_X1 U21099 ( .A1(n23731), .A2(n23732), .A3(n23733), .A4(n23734), .ZN(
        n23721) );
  NOR4_X1 U21100 ( .A1(n23723), .A2(n23724), .A3(n23725), .A4(n23726), .ZN(
        n23722) );
  OAI221_X1 U21101 ( .B1(n21567), .B2(n26721), .C1(n21407), .C2(n26715), .A(
        n23737), .ZN(n23732) );
  NAND2_X1 U21102 ( .A1(n23703), .A2(n23704), .ZN(n5917) );
  NOR4_X1 U21103 ( .A1(n23713), .A2(n23714), .A3(n23715), .A4(n23716), .ZN(
        n23703) );
  NOR4_X1 U21104 ( .A1(n23705), .A2(n23706), .A3(n23707), .A4(n23708), .ZN(
        n23704) );
  OAI221_X1 U21105 ( .B1(n21566), .B2(n26721), .C1(n21406), .C2(n26715), .A(
        n23719), .ZN(n23714) );
  NAND2_X1 U21106 ( .A1(n23685), .A2(n23686), .ZN(n5919) );
  NOR4_X1 U21107 ( .A1(n23695), .A2(n23696), .A3(n23697), .A4(n23698), .ZN(
        n23685) );
  NOR4_X1 U21108 ( .A1(n23687), .A2(n23688), .A3(n23689), .A4(n23690), .ZN(
        n23686) );
  OAI221_X1 U21109 ( .B1(n21565), .B2(n26721), .C1(n21405), .C2(n26715), .A(
        n23701), .ZN(n23696) );
  NAND2_X1 U21110 ( .A1(n23667), .A2(n23668), .ZN(n5921) );
  NOR4_X1 U21111 ( .A1(n23677), .A2(n23678), .A3(n23679), .A4(n23680), .ZN(
        n23667) );
  NOR4_X1 U21112 ( .A1(n23669), .A2(n23670), .A3(n23671), .A4(n23672), .ZN(
        n23668) );
  OAI221_X1 U21113 ( .B1(n21564), .B2(n26721), .C1(n21404), .C2(n26715), .A(
        n23683), .ZN(n23678) );
  NAND2_X1 U21114 ( .A1(n23649), .A2(n23650), .ZN(n5923) );
  NOR4_X1 U21115 ( .A1(n23659), .A2(n23660), .A3(n23661), .A4(n23662), .ZN(
        n23649) );
  NOR4_X1 U21116 ( .A1(n23651), .A2(n23652), .A3(n23653), .A4(n23654), .ZN(
        n23650) );
  OAI221_X1 U21117 ( .B1(n21563), .B2(n26721), .C1(n21403), .C2(n26715), .A(
        n23665), .ZN(n23660) );
  NAND2_X1 U21118 ( .A1(n23631), .A2(n23632), .ZN(n5925) );
  NOR4_X1 U21119 ( .A1(n23641), .A2(n23642), .A3(n23643), .A4(n23644), .ZN(
        n23631) );
  NOR4_X1 U21120 ( .A1(n23633), .A2(n23634), .A3(n23635), .A4(n23636), .ZN(
        n23632) );
  OAI221_X1 U21121 ( .B1(n21562), .B2(n26721), .C1(n21402), .C2(n26715), .A(
        n23647), .ZN(n23642) );
  NAND2_X1 U21122 ( .A1(n23613), .A2(n23614), .ZN(n5927) );
  NOR4_X1 U21123 ( .A1(n23623), .A2(n23624), .A3(n23625), .A4(n23626), .ZN(
        n23613) );
  NOR4_X1 U21124 ( .A1(n23615), .A2(n23616), .A3(n23617), .A4(n23618), .ZN(
        n23614) );
  OAI221_X1 U21125 ( .B1(n21561), .B2(n26721), .C1(n21401), .C2(n26715), .A(
        n23629), .ZN(n23624) );
  NAND2_X1 U21126 ( .A1(n23595), .A2(n23596), .ZN(n5929) );
  NOR4_X1 U21127 ( .A1(n23605), .A2(n23606), .A3(n23607), .A4(n23608), .ZN(
        n23595) );
  NOR4_X1 U21128 ( .A1(n23597), .A2(n23598), .A3(n23599), .A4(n23600), .ZN(
        n23596) );
  OAI221_X1 U21129 ( .B1(n21560), .B2(n26721), .C1(n21400), .C2(n26715), .A(
        n23611), .ZN(n23606) );
  NAND2_X1 U21130 ( .A1(n23577), .A2(n23578), .ZN(n5931) );
  NOR4_X1 U21131 ( .A1(n23587), .A2(n23588), .A3(n23589), .A4(n23590), .ZN(
        n23577) );
  NOR4_X1 U21132 ( .A1(n23579), .A2(n23580), .A3(n23581), .A4(n23582), .ZN(
        n23578) );
  OAI221_X1 U21133 ( .B1(n21559), .B2(n26721), .C1(n21399), .C2(n26715), .A(
        n23593), .ZN(n23588) );
  NAND2_X1 U21134 ( .A1(n23559), .A2(n23560), .ZN(n5933) );
  NOR4_X1 U21135 ( .A1(n23569), .A2(n23570), .A3(n23571), .A4(n23572), .ZN(
        n23559) );
  NOR4_X1 U21136 ( .A1(n23561), .A2(n23562), .A3(n23563), .A4(n23564), .ZN(
        n23560) );
  OAI221_X1 U21137 ( .B1(n21558), .B2(n26721), .C1(n21398), .C2(n26715), .A(
        n23575), .ZN(n23570) );
  NAND2_X1 U21138 ( .A1(n23541), .A2(n23542), .ZN(n5935) );
  NOR4_X1 U21139 ( .A1(n23551), .A2(n23552), .A3(n23553), .A4(n23554), .ZN(
        n23541) );
  NOR4_X1 U21140 ( .A1(n23543), .A2(n23544), .A3(n23545), .A4(n23546), .ZN(
        n23542) );
  OAI221_X1 U21141 ( .B1(n21557), .B2(n26721), .C1(n21397), .C2(n26715), .A(
        n23557), .ZN(n23552) );
  NAND2_X1 U21142 ( .A1(n23523), .A2(n23524), .ZN(n5937) );
  NOR4_X1 U21143 ( .A1(n23533), .A2(n23534), .A3(n23535), .A4(n23536), .ZN(
        n23523) );
  NOR4_X1 U21144 ( .A1(n23525), .A2(n23526), .A3(n23527), .A4(n23528), .ZN(
        n23524) );
  OAI221_X1 U21145 ( .B1(n21556), .B2(n26721), .C1(n21396), .C2(n26715), .A(
        n23539), .ZN(n23534) );
  NAND2_X1 U21146 ( .A1(n23505), .A2(n23506), .ZN(n5939) );
  NOR4_X1 U21147 ( .A1(n23515), .A2(n23516), .A3(n23517), .A4(n23518), .ZN(
        n23505) );
  NOR4_X1 U21148 ( .A1(n23507), .A2(n23508), .A3(n23509), .A4(n23510), .ZN(
        n23506) );
  OAI221_X1 U21149 ( .B1(n21555), .B2(n26722), .C1(n21395), .C2(n26716), .A(
        n23521), .ZN(n23516) );
  NAND2_X1 U21150 ( .A1(n23487), .A2(n23488), .ZN(n5941) );
  NOR4_X1 U21151 ( .A1(n23497), .A2(n23498), .A3(n23499), .A4(n23500), .ZN(
        n23487) );
  NOR4_X1 U21152 ( .A1(n23489), .A2(n23490), .A3(n23491), .A4(n23492), .ZN(
        n23488) );
  OAI221_X1 U21153 ( .B1(n21554), .B2(n26722), .C1(n21394), .C2(n26716), .A(
        n23503), .ZN(n23498) );
  NAND2_X1 U21154 ( .A1(n23469), .A2(n23470), .ZN(n5943) );
  NOR4_X1 U21155 ( .A1(n23479), .A2(n23480), .A3(n23481), .A4(n23482), .ZN(
        n23469) );
  NOR4_X1 U21156 ( .A1(n23471), .A2(n23472), .A3(n23473), .A4(n23474), .ZN(
        n23470) );
  OAI221_X1 U21157 ( .B1(n21553), .B2(n26722), .C1(n21393), .C2(n26716), .A(
        n23485), .ZN(n23480) );
  NAND2_X1 U21158 ( .A1(n23451), .A2(n23452), .ZN(n5945) );
  NOR4_X1 U21159 ( .A1(n23461), .A2(n23462), .A3(n23463), .A4(n23464), .ZN(
        n23451) );
  NOR4_X1 U21160 ( .A1(n23453), .A2(n23454), .A3(n23455), .A4(n23456), .ZN(
        n23452) );
  OAI221_X1 U21161 ( .B1(n21552), .B2(n26722), .C1(n21392), .C2(n26716), .A(
        n23467), .ZN(n23462) );
  NAND2_X1 U21162 ( .A1(n23433), .A2(n23434), .ZN(n5947) );
  NOR4_X1 U21163 ( .A1(n23443), .A2(n23444), .A3(n23445), .A4(n23446), .ZN(
        n23433) );
  NOR4_X1 U21164 ( .A1(n23435), .A2(n23436), .A3(n23437), .A4(n23438), .ZN(
        n23434) );
  OAI221_X1 U21165 ( .B1(n21551), .B2(n26722), .C1(n21391), .C2(n26716), .A(
        n23449), .ZN(n23444) );
  NAND2_X1 U21166 ( .A1(n23415), .A2(n23416), .ZN(n5949) );
  NOR4_X1 U21167 ( .A1(n23425), .A2(n23426), .A3(n23427), .A4(n23428), .ZN(
        n23415) );
  NOR4_X1 U21168 ( .A1(n23417), .A2(n23418), .A3(n23419), .A4(n23420), .ZN(
        n23416) );
  OAI221_X1 U21169 ( .B1(n21550), .B2(n26722), .C1(n21390), .C2(n26716), .A(
        n23431), .ZN(n23426) );
  NAND2_X1 U21170 ( .A1(n23397), .A2(n23398), .ZN(n5951) );
  NOR4_X1 U21171 ( .A1(n23407), .A2(n23408), .A3(n23409), .A4(n23410), .ZN(
        n23397) );
  NOR4_X1 U21172 ( .A1(n23399), .A2(n23400), .A3(n23401), .A4(n23402), .ZN(
        n23398) );
  OAI221_X1 U21173 ( .B1(n21549), .B2(n26722), .C1(n21389), .C2(n26716), .A(
        n23413), .ZN(n23408) );
  NAND2_X1 U21174 ( .A1(n23379), .A2(n23380), .ZN(n5953) );
  NOR4_X1 U21175 ( .A1(n23389), .A2(n23390), .A3(n23391), .A4(n23392), .ZN(
        n23379) );
  NOR4_X1 U21176 ( .A1(n23381), .A2(n23382), .A3(n23383), .A4(n23384), .ZN(
        n23380) );
  OAI221_X1 U21177 ( .B1(n21548), .B2(n26722), .C1(n21388), .C2(n26716), .A(
        n23395), .ZN(n23390) );
  NAND2_X1 U21178 ( .A1(n23361), .A2(n23362), .ZN(n5955) );
  NOR4_X1 U21179 ( .A1(n23371), .A2(n23372), .A3(n23373), .A4(n23374), .ZN(
        n23361) );
  NOR4_X1 U21180 ( .A1(n23363), .A2(n23364), .A3(n23365), .A4(n23366), .ZN(
        n23362) );
  OAI221_X1 U21181 ( .B1(n21547), .B2(n26722), .C1(n21387), .C2(n26716), .A(
        n23377), .ZN(n23372) );
  NAND2_X1 U21182 ( .A1(n23343), .A2(n23344), .ZN(n5957) );
  NOR4_X1 U21183 ( .A1(n23353), .A2(n23354), .A3(n23355), .A4(n23356), .ZN(
        n23343) );
  NOR4_X1 U21184 ( .A1(n23345), .A2(n23346), .A3(n23347), .A4(n23348), .ZN(
        n23344) );
  OAI221_X1 U21185 ( .B1(n21546), .B2(n26722), .C1(n21386), .C2(n26716), .A(
        n23359), .ZN(n23354) );
  NAND2_X1 U21186 ( .A1(n23325), .A2(n23326), .ZN(n5959) );
  NOR4_X1 U21187 ( .A1(n23335), .A2(n23336), .A3(n23337), .A4(n23338), .ZN(
        n23325) );
  NOR4_X1 U21188 ( .A1(n23327), .A2(n23328), .A3(n23329), .A4(n23330), .ZN(
        n23326) );
  OAI221_X1 U21189 ( .B1(n21545), .B2(n26722), .C1(n21385), .C2(n26716), .A(
        n23341), .ZN(n23336) );
  NAND2_X1 U21190 ( .A1(n23307), .A2(n23308), .ZN(n5961) );
  NOR4_X1 U21191 ( .A1(n23317), .A2(n23318), .A3(n23319), .A4(n23320), .ZN(
        n23307) );
  NOR4_X1 U21192 ( .A1(n23309), .A2(n23310), .A3(n23311), .A4(n23312), .ZN(
        n23308) );
  OAI221_X1 U21193 ( .B1(n21544), .B2(n26722), .C1(n21384), .C2(n26716), .A(
        n23323), .ZN(n23318) );
  NAND2_X1 U21194 ( .A1(n23289), .A2(n23290), .ZN(n5963) );
  NOR4_X1 U21195 ( .A1(n23299), .A2(n23300), .A3(n23301), .A4(n23302), .ZN(
        n23289) );
  NOR4_X1 U21196 ( .A1(n23291), .A2(n23292), .A3(n23293), .A4(n23294), .ZN(
        n23290) );
  OAI221_X1 U21197 ( .B1(n21543), .B2(n26723), .C1(n21383), .C2(n26717), .A(
        n23305), .ZN(n23300) );
  NAND2_X1 U21198 ( .A1(n23271), .A2(n23272), .ZN(n5965) );
  NOR4_X1 U21199 ( .A1(n23281), .A2(n23282), .A3(n23283), .A4(n23284), .ZN(
        n23271) );
  NOR4_X1 U21200 ( .A1(n23273), .A2(n23274), .A3(n23275), .A4(n23276), .ZN(
        n23272) );
  OAI221_X1 U21201 ( .B1(n21542), .B2(n26723), .C1(n21382), .C2(n26717), .A(
        n23287), .ZN(n23282) );
  NAND2_X1 U21202 ( .A1(n23253), .A2(n23254), .ZN(n5967) );
  NOR4_X1 U21203 ( .A1(n23263), .A2(n23264), .A3(n23265), .A4(n23266), .ZN(
        n23253) );
  NOR4_X1 U21204 ( .A1(n23255), .A2(n23256), .A3(n23257), .A4(n23258), .ZN(
        n23254) );
  OAI221_X1 U21205 ( .B1(n21541), .B2(n26723), .C1(n21381), .C2(n26717), .A(
        n23269), .ZN(n23264) );
  NAND2_X1 U21206 ( .A1(n23235), .A2(n23236), .ZN(n5969) );
  NOR4_X1 U21207 ( .A1(n23245), .A2(n23246), .A3(n23247), .A4(n23248), .ZN(
        n23235) );
  NOR4_X1 U21208 ( .A1(n23237), .A2(n23238), .A3(n23239), .A4(n23240), .ZN(
        n23236) );
  OAI221_X1 U21209 ( .B1(n21540), .B2(n26723), .C1(n21380), .C2(n26717), .A(
        n23251), .ZN(n23246) );
  NAND2_X1 U21210 ( .A1(n23217), .A2(n23218), .ZN(n5971) );
  NOR4_X1 U21211 ( .A1(n23227), .A2(n23228), .A3(n23229), .A4(n23230), .ZN(
        n23217) );
  NOR4_X1 U21212 ( .A1(n23219), .A2(n23220), .A3(n23221), .A4(n23222), .ZN(
        n23218) );
  OAI221_X1 U21213 ( .B1(n21539), .B2(n26723), .C1(n21379), .C2(n26717), .A(
        n23233), .ZN(n23228) );
  NAND2_X1 U21214 ( .A1(n23199), .A2(n23200), .ZN(n5973) );
  NOR4_X1 U21215 ( .A1(n23209), .A2(n23210), .A3(n23211), .A4(n23212), .ZN(
        n23199) );
  NOR4_X1 U21216 ( .A1(n23201), .A2(n23202), .A3(n23203), .A4(n23204), .ZN(
        n23200) );
  OAI221_X1 U21217 ( .B1(n21538), .B2(n26723), .C1(n21378), .C2(n26717), .A(
        n23215), .ZN(n23210) );
  NAND2_X1 U21218 ( .A1(n23181), .A2(n23182), .ZN(n5975) );
  NOR4_X1 U21219 ( .A1(n23191), .A2(n23192), .A3(n23193), .A4(n23194), .ZN(
        n23181) );
  NOR4_X1 U21220 ( .A1(n23183), .A2(n23184), .A3(n23185), .A4(n23186), .ZN(
        n23182) );
  OAI221_X1 U21221 ( .B1(n21537), .B2(n26723), .C1(n21377), .C2(n26717), .A(
        n23197), .ZN(n23192) );
  NAND2_X1 U21222 ( .A1(n23163), .A2(n23164), .ZN(n5977) );
  NOR4_X1 U21223 ( .A1(n23173), .A2(n23174), .A3(n23175), .A4(n23176), .ZN(
        n23163) );
  NOR4_X1 U21224 ( .A1(n23165), .A2(n23166), .A3(n23167), .A4(n23168), .ZN(
        n23164) );
  OAI221_X1 U21225 ( .B1(n21536), .B2(n26723), .C1(n21376), .C2(n26717), .A(
        n23179), .ZN(n23174) );
  NAND2_X1 U21226 ( .A1(n23145), .A2(n23146), .ZN(n5979) );
  NOR4_X1 U21227 ( .A1(n23155), .A2(n23156), .A3(n23157), .A4(n23158), .ZN(
        n23145) );
  NOR4_X1 U21228 ( .A1(n23147), .A2(n23148), .A3(n23149), .A4(n23150), .ZN(
        n23146) );
  OAI221_X1 U21229 ( .B1(n21535), .B2(n26723), .C1(n21375), .C2(n26717), .A(
        n23161), .ZN(n23156) );
  NAND2_X1 U21230 ( .A1(n23127), .A2(n23128), .ZN(n5981) );
  NOR4_X1 U21231 ( .A1(n23137), .A2(n23138), .A3(n23139), .A4(n23140), .ZN(
        n23127) );
  NOR4_X1 U21232 ( .A1(n23129), .A2(n23130), .A3(n23131), .A4(n23132), .ZN(
        n23128) );
  OAI221_X1 U21233 ( .B1(n21534), .B2(n26723), .C1(n21374), .C2(n26717), .A(
        n23143), .ZN(n23138) );
  NAND2_X1 U21234 ( .A1(n23109), .A2(n23110), .ZN(n5983) );
  NOR4_X1 U21235 ( .A1(n23119), .A2(n23120), .A3(n23121), .A4(n23122), .ZN(
        n23109) );
  NOR4_X1 U21236 ( .A1(n23111), .A2(n23112), .A3(n23113), .A4(n23114), .ZN(
        n23110) );
  OAI221_X1 U21237 ( .B1(n21533), .B2(n26723), .C1(n21373), .C2(n26717), .A(
        n23125), .ZN(n23120) );
  NAND2_X1 U21238 ( .A1(n23091), .A2(n23092), .ZN(n5985) );
  NOR4_X1 U21239 ( .A1(n23101), .A2(n23102), .A3(n23103), .A4(n23104), .ZN(
        n23091) );
  NOR4_X1 U21240 ( .A1(n23093), .A2(n23094), .A3(n23095), .A4(n23096), .ZN(
        n23092) );
  OAI221_X1 U21241 ( .B1(n21532), .B2(n26723), .C1(n21372), .C2(n26717), .A(
        n23107), .ZN(n23102) );
  NAND2_X1 U21242 ( .A1(n23968), .A2(n23969), .ZN(n5889) );
  NOR4_X1 U21243 ( .A1(n23995), .A2(n23996), .A3(n23997), .A4(n23998), .ZN(
        n23968) );
  NOR4_X1 U21244 ( .A1(n23970), .A2(n23971), .A3(n23972), .A4(n23973), .ZN(
        n23969) );
  OAI221_X1 U21245 ( .B1(n21176), .B2(n26500), .C1(n21168), .C2(n26494), .A(
        n24011), .ZN(n23996) );
  NAND2_X1 U21246 ( .A1(n24056), .A2(n24057), .ZN(n5883) );
  NOR4_X1 U21247 ( .A1(n24066), .A2(n24067), .A3(n24068), .A4(n24069), .ZN(
        n24056) );
  NOR4_X1 U21248 ( .A1(n24058), .A2(n24059), .A3(n24060), .A4(n24061), .ZN(
        n24057) );
  OAI221_X1 U21249 ( .B1(n21179), .B2(n26500), .C1(n21171), .C2(n26494), .A(
        n24072), .ZN(n24067) );
  NAND2_X1 U21250 ( .A1(n24038), .A2(n24039), .ZN(n5885) );
  NOR4_X1 U21251 ( .A1(n24048), .A2(n24049), .A3(n24050), .A4(n24051), .ZN(
        n24038) );
  NOR4_X1 U21252 ( .A1(n24040), .A2(n24041), .A3(n24042), .A4(n24043), .ZN(
        n24039) );
  OAI221_X1 U21253 ( .B1(n21178), .B2(n26500), .C1(n21170), .C2(n26494), .A(
        n24054), .ZN(n24049) );
  NAND2_X1 U21254 ( .A1(n24020), .A2(n24021), .ZN(n5887) );
  NOR4_X1 U21255 ( .A1(n24030), .A2(n24031), .A3(n24032), .A4(n24033), .ZN(
        n24020) );
  NOR4_X1 U21256 ( .A1(n24022), .A2(n24023), .A3(n24024), .A4(n24025), .ZN(
        n24021) );
  OAI221_X1 U21257 ( .B1(n21177), .B2(n26500), .C1(n21169), .C2(n26494), .A(
        n24036), .ZN(n24031) );
  NAND2_X1 U21258 ( .A1(n22857), .A2(n22858), .ZN(n6011) );
  NOR4_X1 U21259 ( .A1(n22867), .A2(n22868), .A3(n22869), .A4(n22870), .ZN(
        n22857) );
  NOR4_X1 U21260 ( .A1(n22859), .A2(n22860), .A3(n22861), .A4(n22862), .ZN(
        n22858) );
  OAI221_X1 U21261 ( .B1(n21179), .B2(n26725), .C1(n21171), .C2(n26719), .A(
        n22873), .ZN(n22868) );
  NAND2_X1 U21262 ( .A1(n22839), .A2(n22840), .ZN(n6013) );
  NOR4_X1 U21263 ( .A1(n22849), .A2(n22850), .A3(n22851), .A4(n22852), .ZN(
        n22839) );
  NOR4_X1 U21264 ( .A1(n22841), .A2(n22842), .A3(n22843), .A4(n22844), .ZN(
        n22840) );
  OAI221_X1 U21265 ( .B1(n21178), .B2(n26725), .C1(n21170), .C2(n26719), .A(
        n22855), .ZN(n22850) );
  NAND2_X1 U21266 ( .A1(n22821), .A2(n22822), .ZN(n6015) );
  NOR4_X1 U21267 ( .A1(n22831), .A2(n22832), .A3(n22833), .A4(n22834), .ZN(
        n22821) );
  NOR4_X1 U21268 ( .A1(n22823), .A2(n22824), .A3(n22825), .A4(n22826), .ZN(
        n22822) );
  OAI221_X1 U21269 ( .B1(n21177), .B2(n26725), .C1(n21169), .C2(n26719), .A(
        n22837), .ZN(n22832) );
  NAND2_X1 U21270 ( .A1(n22769), .A2(n22770), .ZN(n6017) );
  NOR4_X1 U21271 ( .A1(n22796), .A2(n22797), .A3(n22798), .A4(n22799), .ZN(
        n22769) );
  NOR4_X1 U21272 ( .A1(n22771), .A2(n22772), .A3(n22773), .A4(n22774), .ZN(
        n22770) );
  OAI221_X1 U21273 ( .B1(n21176), .B2(n26725), .C1(n21168), .C2(n26719), .A(
        n22812), .ZN(n22797) );
  NAND2_X1 U21274 ( .A1(n24272), .A2(n24273), .ZN(n5859) );
  NOR4_X1 U21275 ( .A1(n24282), .A2(n24283), .A3(n24284), .A4(n24285), .ZN(
        n24272) );
  NOR4_X1 U21276 ( .A1(n24274), .A2(n24275), .A3(n24276), .A4(n24277), .ZN(
        n24273) );
  OAI221_X1 U21277 ( .B1(n21531), .B2(n26499), .C1(n21371), .C2(n26493), .A(
        n24288), .ZN(n24283) );
  NAND2_X1 U21278 ( .A1(n24254), .A2(n24255), .ZN(n5861) );
  NOR4_X1 U21279 ( .A1(n24264), .A2(n24265), .A3(n24266), .A4(n24267), .ZN(
        n24254) );
  NOR4_X1 U21280 ( .A1(n24256), .A2(n24257), .A3(n24258), .A4(n24259), .ZN(
        n24255) );
  OAI221_X1 U21281 ( .B1(n21530), .B2(n26499), .C1(n21370), .C2(n26493), .A(
        n24270), .ZN(n24265) );
  NAND2_X1 U21282 ( .A1(n24236), .A2(n24237), .ZN(n5863) );
  NOR4_X1 U21283 ( .A1(n24246), .A2(n24247), .A3(n24248), .A4(n24249), .ZN(
        n24236) );
  NOR4_X1 U21284 ( .A1(n24238), .A2(n24239), .A3(n24240), .A4(n24241), .ZN(
        n24237) );
  OAI221_X1 U21285 ( .B1(n21529), .B2(n26499), .C1(n21369), .C2(n26493), .A(
        n24252), .ZN(n24247) );
  NAND2_X1 U21286 ( .A1(n24218), .A2(n24219), .ZN(n5865) );
  NOR4_X1 U21287 ( .A1(n24228), .A2(n24229), .A3(n24230), .A4(n24231), .ZN(
        n24218) );
  NOR4_X1 U21288 ( .A1(n24220), .A2(n24221), .A3(n24222), .A4(n24223), .ZN(
        n24219) );
  OAI221_X1 U21289 ( .B1(n21528), .B2(n26499), .C1(n21368), .C2(n26493), .A(
        n24234), .ZN(n24229) );
  NAND2_X1 U21290 ( .A1(n24200), .A2(n24201), .ZN(n5867) );
  NOR4_X1 U21291 ( .A1(n24210), .A2(n24211), .A3(n24212), .A4(n24213), .ZN(
        n24200) );
  NOR4_X1 U21292 ( .A1(n24202), .A2(n24203), .A3(n24204), .A4(n24205), .ZN(
        n24201) );
  OAI221_X1 U21293 ( .B1(n21527), .B2(n26499), .C1(n21367), .C2(n26493), .A(
        n24216), .ZN(n24211) );
  NAND2_X1 U21294 ( .A1(n24182), .A2(n24183), .ZN(n5869) );
  NOR4_X1 U21295 ( .A1(n24192), .A2(n24193), .A3(n24194), .A4(n24195), .ZN(
        n24182) );
  NOR4_X1 U21296 ( .A1(n24184), .A2(n24185), .A3(n24186), .A4(n24187), .ZN(
        n24183) );
  OAI221_X1 U21297 ( .B1(n21526), .B2(n26499), .C1(n21366), .C2(n26493), .A(
        n24198), .ZN(n24193) );
  NAND2_X1 U21298 ( .A1(n24164), .A2(n24165), .ZN(n5871) );
  NOR4_X1 U21299 ( .A1(n24174), .A2(n24175), .A3(n24176), .A4(n24177), .ZN(
        n24164) );
  NOR4_X1 U21300 ( .A1(n24166), .A2(n24167), .A3(n24168), .A4(n24169), .ZN(
        n24165) );
  OAI221_X1 U21301 ( .B1(n21525), .B2(n26499), .C1(n21365), .C2(n26493), .A(
        n24180), .ZN(n24175) );
  NAND2_X1 U21302 ( .A1(n24146), .A2(n24147), .ZN(n5873) );
  NOR4_X1 U21303 ( .A1(n24156), .A2(n24157), .A3(n24158), .A4(n24159), .ZN(
        n24146) );
  NOR4_X1 U21304 ( .A1(n24148), .A2(n24149), .A3(n24150), .A4(n24151), .ZN(
        n24147) );
  OAI221_X1 U21305 ( .B1(n21524), .B2(n26499), .C1(n21364), .C2(n26493), .A(
        n24162), .ZN(n24157) );
  NAND2_X1 U21306 ( .A1(n24128), .A2(n24129), .ZN(n5875) );
  NOR4_X1 U21307 ( .A1(n24138), .A2(n24139), .A3(n24140), .A4(n24141), .ZN(
        n24128) );
  NOR4_X1 U21308 ( .A1(n24130), .A2(n24131), .A3(n24132), .A4(n24133), .ZN(
        n24129) );
  OAI221_X1 U21309 ( .B1(n21523), .B2(n26499), .C1(n21363), .C2(n26493), .A(
        n24144), .ZN(n24139) );
  NAND2_X1 U21310 ( .A1(n24110), .A2(n24111), .ZN(n5877) );
  NOR4_X1 U21311 ( .A1(n24120), .A2(n24121), .A3(n24122), .A4(n24123), .ZN(
        n24110) );
  NOR4_X1 U21312 ( .A1(n24112), .A2(n24113), .A3(n24114), .A4(n24115), .ZN(
        n24111) );
  OAI221_X1 U21313 ( .B1(n21522), .B2(n26499), .C1(n21362), .C2(n26493), .A(
        n24126), .ZN(n24121) );
  NAND2_X1 U21314 ( .A1(n24092), .A2(n24093), .ZN(n5879) );
  NOR4_X1 U21315 ( .A1(n24102), .A2(n24103), .A3(n24104), .A4(n24105), .ZN(
        n24092) );
  NOR4_X1 U21316 ( .A1(n24094), .A2(n24095), .A3(n24096), .A4(n24097), .ZN(
        n24093) );
  OAI221_X1 U21317 ( .B1(n21521), .B2(n26499), .C1(n21361), .C2(n26493), .A(
        n24108), .ZN(n24103) );
  NAND2_X1 U21318 ( .A1(n24074), .A2(n24075), .ZN(n5881) );
  NOR4_X1 U21319 ( .A1(n24084), .A2(n24085), .A3(n24086), .A4(n24087), .ZN(
        n24074) );
  NOR4_X1 U21320 ( .A1(n24076), .A2(n24077), .A3(n24078), .A4(n24079), .ZN(
        n24075) );
  OAI221_X1 U21321 ( .B1(n21520), .B2(n26499), .C1(n21360), .C2(n26493), .A(
        n24090), .ZN(n24085) );
  NAND2_X1 U21322 ( .A1(n23073), .A2(n23074), .ZN(n5987) );
  NOR4_X1 U21323 ( .A1(n23083), .A2(n23084), .A3(n23085), .A4(n23086), .ZN(
        n23073) );
  NOR4_X1 U21324 ( .A1(n23075), .A2(n23076), .A3(n23077), .A4(n23078), .ZN(
        n23074) );
  OAI221_X1 U21325 ( .B1(n21531), .B2(n26724), .C1(n21371), .C2(n26718), .A(
        n23089), .ZN(n23084) );
  NAND2_X1 U21326 ( .A1(n23055), .A2(n23056), .ZN(n5989) );
  NOR4_X1 U21327 ( .A1(n23065), .A2(n23066), .A3(n23067), .A4(n23068), .ZN(
        n23055) );
  NOR4_X1 U21328 ( .A1(n23057), .A2(n23058), .A3(n23059), .A4(n23060), .ZN(
        n23056) );
  OAI221_X1 U21329 ( .B1(n21530), .B2(n26724), .C1(n21370), .C2(n26718), .A(
        n23071), .ZN(n23066) );
  NAND2_X1 U21330 ( .A1(n23037), .A2(n23038), .ZN(n5991) );
  NOR4_X1 U21331 ( .A1(n23047), .A2(n23048), .A3(n23049), .A4(n23050), .ZN(
        n23037) );
  NOR4_X1 U21332 ( .A1(n23039), .A2(n23040), .A3(n23041), .A4(n23042), .ZN(
        n23038) );
  OAI221_X1 U21333 ( .B1(n21529), .B2(n26724), .C1(n21369), .C2(n26718), .A(
        n23053), .ZN(n23048) );
  NAND2_X1 U21334 ( .A1(n23019), .A2(n23020), .ZN(n5993) );
  NOR4_X1 U21335 ( .A1(n23029), .A2(n23030), .A3(n23031), .A4(n23032), .ZN(
        n23019) );
  NOR4_X1 U21336 ( .A1(n23021), .A2(n23022), .A3(n23023), .A4(n23024), .ZN(
        n23020) );
  OAI221_X1 U21337 ( .B1(n21528), .B2(n26724), .C1(n21368), .C2(n26718), .A(
        n23035), .ZN(n23030) );
  NAND2_X1 U21338 ( .A1(n23001), .A2(n23002), .ZN(n5995) );
  NOR4_X1 U21339 ( .A1(n23011), .A2(n23012), .A3(n23013), .A4(n23014), .ZN(
        n23001) );
  NOR4_X1 U21340 ( .A1(n23003), .A2(n23004), .A3(n23005), .A4(n23006), .ZN(
        n23002) );
  OAI221_X1 U21341 ( .B1(n21527), .B2(n26724), .C1(n21367), .C2(n26718), .A(
        n23017), .ZN(n23012) );
  NAND2_X1 U21342 ( .A1(n22983), .A2(n22984), .ZN(n5997) );
  NOR4_X1 U21343 ( .A1(n22993), .A2(n22994), .A3(n22995), .A4(n22996), .ZN(
        n22983) );
  NOR4_X1 U21344 ( .A1(n22985), .A2(n22986), .A3(n22987), .A4(n22988), .ZN(
        n22984) );
  OAI221_X1 U21345 ( .B1(n21526), .B2(n26724), .C1(n21366), .C2(n26718), .A(
        n22999), .ZN(n22994) );
  NAND2_X1 U21346 ( .A1(n22965), .A2(n22966), .ZN(n5999) );
  NOR4_X1 U21347 ( .A1(n22975), .A2(n22976), .A3(n22977), .A4(n22978), .ZN(
        n22965) );
  NOR4_X1 U21348 ( .A1(n22967), .A2(n22968), .A3(n22969), .A4(n22970), .ZN(
        n22966) );
  OAI221_X1 U21349 ( .B1(n21525), .B2(n26724), .C1(n21365), .C2(n26718), .A(
        n22981), .ZN(n22976) );
  NAND2_X1 U21350 ( .A1(n22947), .A2(n22948), .ZN(n6001) );
  NOR4_X1 U21351 ( .A1(n22957), .A2(n22958), .A3(n22959), .A4(n22960), .ZN(
        n22947) );
  NOR4_X1 U21352 ( .A1(n22949), .A2(n22950), .A3(n22951), .A4(n22952), .ZN(
        n22948) );
  OAI221_X1 U21353 ( .B1(n21524), .B2(n26724), .C1(n21364), .C2(n26718), .A(
        n22963), .ZN(n22958) );
  NAND2_X1 U21354 ( .A1(n22929), .A2(n22930), .ZN(n6003) );
  NOR4_X1 U21355 ( .A1(n22939), .A2(n22940), .A3(n22941), .A4(n22942), .ZN(
        n22929) );
  NOR4_X1 U21356 ( .A1(n22931), .A2(n22932), .A3(n22933), .A4(n22934), .ZN(
        n22930) );
  OAI221_X1 U21357 ( .B1(n21523), .B2(n26724), .C1(n21363), .C2(n26718), .A(
        n22945), .ZN(n22940) );
  NAND2_X1 U21358 ( .A1(n22911), .A2(n22912), .ZN(n6005) );
  NOR4_X1 U21359 ( .A1(n22921), .A2(n22922), .A3(n22923), .A4(n22924), .ZN(
        n22911) );
  NOR4_X1 U21360 ( .A1(n22913), .A2(n22914), .A3(n22915), .A4(n22916), .ZN(
        n22912) );
  OAI221_X1 U21361 ( .B1(n21522), .B2(n26724), .C1(n21362), .C2(n26718), .A(
        n22927), .ZN(n22922) );
  NAND2_X1 U21362 ( .A1(n22893), .A2(n22894), .ZN(n6007) );
  NOR4_X1 U21363 ( .A1(n22903), .A2(n22904), .A3(n22905), .A4(n22906), .ZN(
        n22893) );
  NOR4_X1 U21364 ( .A1(n22895), .A2(n22896), .A3(n22897), .A4(n22898), .ZN(
        n22894) );
  OAI221_X1 U21365 ( .B1(n21521), .B2(n26724), .C1(n21361), .C2(n26718), .A(
        n22909), .ZN(n22904) );
  NAND2_X1 U21366 ( .A1(n22875), .A2(n22876), .ZN(n6009) );
  NOR4_X1 U21367 ( .A1(n22885), .A2(n22886), .A3(n22887), .A4(n22888), .ZN(
        n22875) );
  NOR4_X1 U21368 ( .A1(n22877), .A2(n22878), .A3(n22879), .A4(n22880), .ZN(
        n22876) );
  OAI221_X1 U21369 ( .B1(n21520), .B2(n26724), .C1(n21360), .C2(n26718), .A(
        n22891), .ZN(n22886) );
  BUF_X1 U21370 ( .A(n24010), .Z(n26489) );
  BUF_X1 U21371 ( .A(n24010), .Z(n26490) );
  BUF_X1 U21372 ( .A(n24010), .Z(n26491) );
  BUF_X1 U21373 ( .A(n24010), .Z(n26492) );
  BUF_X1 U21374 ( .A(n22811), .Z(n26714) );
  BUF_X1 U21375 ( .A(n22811), .Z(n26715) );
  BUF_X1 U21376 ( .A(n22811), .Z(n26716) );
  BUF_X1 U21377 ( .A(n22811), .Z(n26717) );
  INV_X1 U21378 ( .A(n27487), .ZN(n27477) );
  INV_X1 U21379 ( .A(n27487), .ZN(n27478) );
  INV_X1 U21380 ( .A(n27487), .ZN(n27479) );
  INV_X1 U21381 ( .A(n27487), .ZN(n27480) );
  INV_X1 U21382 ( .A(n27487), .ZN(n27481) );
  INV_X1 U21383 ( .A(n27487), .ZN(n27483) );
  INV_X1 U21384 ( .A(n27487), .ZN(n27482) );
  INV_X1 U21385 ( .A(n27487), .ZN(n27485) );
  INV_X1 U21386 ( .A(n27487), .ZN(n27486) );
  INV_X1 U21387 ( .A(n27487), .ZN(n27484) );
  BUF_X1 U21388 ( .A(n24014), .Z(n26471) );
  BUF_X1 U21389 ( .A(n24009), .Z(n26495) );
  BUF_X1 U21390 ( .A(n24014), .Z(n26472) );
  BUF_X1 U21391 ( .A(n24009), .Z(n26496) );
  BUF_X1 U21392 ( .A(n24014), .Z(n26473) );
  BUF_X1 U21393 ( .A(n24009), .Z(n26497) );
  BUF_X1 U21394 ( .A(n24014), .Z(n26474) );
  BUF_X1 U21395 ( .A(n24009), .Z(n26498) );
  BUF_X1 U21396 ( .A(n22815), .Z(n26696) );
  BUF_X1 U21397 ( .A(n22810), .Z(n26720) );
  BUF_X1 U21398 ( .A(n22815), .Z(n26697) );
  BUF_X1 U21399 ( .A(n22810), .Z(n26721) );
  BUF_X1 U21400 ( .A(n22815), .Z(n26698) );
  BUF_X1 U21401 ( .A(n22810), .Z(n26722) );
  BUF_X1 U21402 ( .A(n22815), .Z(n26699) );
  BUF_X1 U21403 ( .A(n22810), .Z(n26723) );
  NOR3_X1 U21404 ( .A1(n20640), .A2(n20643), .A3(n20639), .ZN(n25143) );
  NOR3_X1 U21405 ( .A1(n20635), .A2(n20638), .A3(n20634), .ZN(n23944) );
  AND3_X1 U21406 ( .A1(n20631), .A2(n20630), .A3(n22717), .ZN(n22695) );
  NAND2_X1 U21407 ( .A1(n22704), .A2(n22695), .ZN(n22702) );
  NAND2_X1 U21408 ( .A1(n22698), .A2(n22695), .ZN(n22696) );
  NAND2_X1 U21409 ( .A1(n22701), .A2(n22695), .ZN(n22699) );
  AND3_X1 U21410 ( .A1(n20642), .A2(n20641), .A3(n25164), .ZN(n25151) );
  AND3_X1 U21411 ( .A1(n20637), .A2(n20636), .A3(n23965), .ZN(n23952) );
  BUF_X1 U21412 ( .A(n20707), .Z(n27282) );
  BUF_X1 U21413 ( .A(n20706), .Z(n27285) );
  BUF_X1 U21414 ( .A(n20705), .Z(n27288) );
  BUF_X1 U21415 ( .A(n20704), .Z(n27291) );
  BUF_X1 U21416 ( .A(n20703), .Z(n27294) );
  BUF_X1 U21417 ( .A(n20702), .Z(n27297) );
  BUF_X1 U21418 ( .A(n20701), .Z(n27300) );
  BUF_X1 U21419 ( .A(n20700), .Z(n27303) );
  BUF_X1 U21420 ( .A(n20699), .Z(n27306) );
  BUF_X1 U21421 ( .A(n20698), .Z(n27309) );
  BUF_X1 U21422 ( .A(n20697), .Z(n27312) );
  BUF_X1 U21423 ( .A(n20696), .Z(n27315) );
  BUF_X1 U21424 ( .A(n20695), .Z(n27318) );
  BUF_X1 U21425 ( .A(n20694), .Z(n27321) );
  BUF_X1 U21426 ( .A(n20693), .Z(n27324) );
  BUF_X1 U21427 ( .A(n20692), .Z(n27327) );
  BUF_X1 U21428 ( .A(n20691), .Z(n27330) );
  BUF_X1 U21429 ( .A(n20690), .Z(n27333) );
  BUF_X1 U21430 ( .A(n20689), .Z(n27336) );
  BUF_X1 U21431 ( .A(n20688), .Z(n27339) );
  BUF_X1 U21432 ( .A(n20687), .Z(n27342) );
  BUF_X1 U21433 ( .A(n20686), .Z(n27345) );
  BUF_X1 U21434 ( .A(n20685), .Z(n27348) );
  BUF_X1 U21435 ( .A(n20684), .Z(n27351) );
  BUF_X1 U21436 ( .A(n20683), .Z(n27354) );
  BUF_X1 U21437 ( .A(n20682), .Z(n27357) );
  BUF_X1 U21438 ( .A(n20681), .Z(n27360) );
  BUF_X1 U21439 ( .A(n20680), .Z(n27363) );
  BUF_X1 U21440 ( .A(n20679), .Z(n27366) );
  BUF_X1 U21441 ( .A(n20678), .Z(n27369) );
  BUF_X1 U21442 ( .A(n20677), .Z(n27372) );
  BUF_X1 U21443 ( .A(n20676), .Z(n27375) );
  BUF_X1 U21444 ( .A(n20675), .Z(n27378) );
  BUF_X1 U21445 ( .A(n20674), .Z(n27381) );
  BUF_X1 U21446 ( .A(n20673), .Z(n27384) );
  BUF_X1 U21447 ( .A(n20672), .Z(n27387) );
  BUF_X1 U21448 ( .A(n20671), .Z(n27390) );
  BUF_X1 U21449 ( .A(n20670), .Z(n27393) );
  BUF_X1 U21450 ( .A(n20669), .Z(n27396) );
  BUF_X1 U21451 ( .A(n20668), .Z(n27399) );
  BUF_X1 U21452 ( .A(n20667), .Z(n27402) );
  BUF_X1 U21453 ( .A(n20666), .Z(n27405) );
  BUF_X1 U21454 ( .A(n20665), .Z(n27408) );
  BUF_X1 U21455 ( .A(n20664), .Z(n27411) );
  BUF_X1 U21456 ( .A(n20663), .Z(n27414) );
  BUF_X1 U21457 ( .A(n20662), .Z(n27417) );
  BUF_X1 U21458 ( .A(n20661), .Z(n27420) );
  BUF_X1 U21459 ( .A(n20660), .Z(n27423) );
  BUF_X1 U21460 ( .A(n20659), .Z(n27426) );
  BUF_X1 U21461 ( .A(n20658), .Z(n27429) );
  BUF_X1 U21462 ( .A(n20657), .Z(n27432) );
  BUF_X1 U21463 ( .A(n20656), .Z(n27435) );
  BUF_X1 U21464 ( .A(n20655), .Z(n27438) );
  BUF_X1 U21465 ( .A(n20654), .Z(n27441) );
  BUF_X1 U21466 ( .A(n20653), .Z(n27444) );
  BUF_X1 U21467 ( .A(n20652), .Z(n27447) );
  BUF_X1 U21468 ( .A(n20651), .Z(n27450) );
  BUF_X1 U21469 ( .A(n20650), .Z(n27453) );
  BUF_X1 U21470 ( .A(n20649), .Z(n27456) );
  BUF_X1 U21471 ( .A(n20648), .Z(n27459) );
  BUF_X1 U21472 ( .A(n20647), .Z(n27462) );
  BUF_X1 U21473 ( .A(n20646), .Z(n27465) );
  BUF_X1 U21474 ( .A(n20645), .Z(n27468) );
  BUF_X1 U21475 ( .A(n20644), .Z(n27471) );
  BUF_X1 U21476 ( .A(n20644), .Z(n27472) );
  BUF_X1 U21477 ( .A(n20707), .Z(n27283) );
  BUF_X1 U21478 ( .A(n20706), .Z(n27286) );
  BUF_X1 U21479 ( .A(n20705), .Z(n27289) );
  BUF_X1 U21480 ( .A(n20704), .Z(n27292) );
  BUF_X1 U21481 ( .A(n20703), .Z(n27295) );
  BUF_X1 U21482 ( .A(n20702), .Z(n27298) );
  BUF_X1 U21483 ( .A(n20701), .Z(n27301) );
  BUF_X1 U21484 ( .A(n20700), .Z(n27304) );
  BUF_X1 U21485 ( .A(n20699), .Z(n27307) );
  BUF_X1 U21486 ( .A(n20698), .Z(n27310) );
  BUF_X1 U21487 ( .A(n20697), .Z(n27313) );
  BUF_X1 U21488 ( .A(n20696), .Z(n27316) );
  BUF_X1 U21489 ( .A(n20695), .Z(n27319) );
  BUF_X1 U21490 ( .A(n20694), .Z(n27322) );
  BUF_X1 U21491 ( .A(n20693), .Z(n27325) );
  BUF_X1 U21492 ( .A(n20692), .Z(n27328) );
  BUF_X1 U21493 ( .A(n20691), .Z(n27331) );
  BUF_X1 U21494 ( .A(n20690), .Z(n27334) );
  BUF_X1 U21495 ( .A(n20689), .Z(n27337) );
  BUF_X1 U21496 ( .A(n20688), .Z(n27340) );
  BUF_X1 U21497 ( .A(n20687), .Z(n27343) );
  BUF_X1 U21498 ( .A(n20686), .Z(n27346) );
  BUF_X1 U21499 ( .A(n20685), .Z(n27349) );
  BUF_X1 U21500 ( .A(n20684), .Z(n27352) );
  BUF_X1 U21501 ( .A(n20683), .Z(n27355) );
  BUF_X1 U21502 ( .A(n20682), .Z(n27358) );
  BUF_X1 U21503 ( .A(n20681), .Z(n27361) );
  BUF_X1 U21504 ( .A(n20680), .Z(n27364) );
  BUF_X1 U21505 ( .A(n20679), .Z(n27367) );
  BUF_X1 U21506 ( .A(n20678), .Z(n27370) );
  BUF_X1 U21507 ( .A(n20677), .Z(n27373) );
  BUF_X1 U21508 ( .A(n20676), .Z(n27376) );
  BUF_X1 U21509 ( .A(n20675), .Z(n27379) );
  BUF_X1 U21510 ( .A(n20674), .Z(n27382) );
  BUF_X1 U21511 ( .A(n20673), .Z(n27385) );
  BUF_X1 U21512 ( .A(n20672), .Z(n27388) );
  BUF_X1 U21513 ( .A(n20671), .Z(n27391) );
  BUF_X1 U21514 ( .A(n20670), .Z(n27394) );
  BUF_X1 U21515 ( .A(n20669), .Z(n27397) );
  BUF_X1 U21516 ( .A(n20668), .Z(n27400) );
  BUF_X1 U21517 ( .A(n20667), .Z(n27403) );
  BUF_X1 U21518 ( .A(n20666), .Z(n27406) );
  BUF_X1 U21519 ( .A(n20665), .Z(n27409) );
  BUF_X1 U21520 ( .A(n20664), .Z(n27412) );
  BUF_X1 U21521 ( .A(n20663), .Z(n27415) );
  BUF_X1 U21522 ( .A(n20662), .Z(n27418) );
  BUF_X1 U21523 ( .A(n20661), .Z(n27421) );
  BUF_X1 U21524 ( .A(n20660), .Z(n27424) );
  BUF_X1 U21525 ( .A(n20659), .Z(n27427) );
  BUF_X1 U21526 ( .A(n20658), .Z(n27430) );
  BUF_X1 U21527 ( .A(n20657), .Z(n27433) );
  BUF_X1 U21528 ( .A(n20656), .Z(n27436) );
  BUF_X1 U21529 ( .A(n20655), .Z(n27439) );
  BUF_X1 U21530 ( .A(n20654), .Z(n27442) );
  BUF_X1 U21531 ( .A(n20653), .Z(n27445) );
  BUF_X1 U21532 ( .A(n20652), .Z(n27448) );
  BUF_X1 U21533 ( .A(n20651), .Z(n27451) );
  BUF_X1 U21534 ( .A(n20650), .Z(n27454) );
  BUF_X1 U21535 ( .A(n20649), .Z(n27457) );
  BUF_X1 U21536 ( .A(n20648), .Z(n27460) );
  BUF_X1 U21537 ( .A(n20647), .Z(n27463) );
  BUF_X1 U21538 ( .A(n20646), .Z(n27466) );
  BUF_X1 U21539 ( .A(n20645), .Z(n27469) );
  NAND2_X1 U21540 ( .A1(n25153), .A2(n25148), .ZN(n23985) );
  NAND2_X1 U21541 ( .A1(n25153), .A2(n25151), .ZN(n24005) );
  NAND2_X1 U21542 ( .A1(n23954), .A2(n23949), .ZN(n22786) );
  NAND2_X1 U21543 ( .A1(n23954), .A2(n23952), .ZN(n22806) );
  NAND2_X1 U21544 ( .A1(n22716), .A2(n22695), .ZN(n22714) );
  NAND2_X1 U21545 ( .A1(n22707), .A2(n22695), .ZN(n22705) );
  NAND2_X1 U21546 ( .A1(n22713), .A2(n22695), .ZN(n22711) );
  NAND2_X1 U21547 ( .A1(n22710), .A2(n22695), .ZN(n22708) );
  NAND2_X1 U21548 ( .A1(n25144), .A2(n25147), .ZN(n23990) );
  NAND2_X1 U21549 ( .A1(n25144), .A2(n25155), .ZN(n24000) );
  NAND2_X1 U21550 ( .A1(n23945), .A2(n23948), .ZN(n22791) );
  NAND2_X1 U21551 ( .A1(n23945), .A2(n23956), .ZN(n22801) );
  NAND2_X1 U21552 ( .A1(n22720), .A2(n22698), .ZN(n22721) );
  NAND2_X1 U21553 ( .A1(n22754), .A2(n22704), .ZN(n22759) );
  NAND2_X1 U21554 ( .A1(n22754), .A2(n22694), .ZN(n22752) );
  NAND2_X1 U21555 ( .A1(n22720), .A2(n22694), .ZN(n22718) );
  NAND2_X1 U21556 ( .A1(n22720), .A2(n22701), .ZN(n22723) );
  NAND2_X1 U21557 ( .A1(n22737), .A2(n22704), .ZN(n22742) );
  NAND2_X1 U21558 ( .A1(n22754), .A2(n22710), .ZN(n22763) );
  NAND2_X1 U21559 ( .A1(n22754), .A2(n22707), .ZN(n22761) );
  NAND2_X1 U21560 ( .A1(n22720), .A2(n22704), .ZN(n22725) );
  NAND2_X1 U21561 ( .A1(n22737), .A2(n22713), .ZN(n22748) );
  NAND2_X1 U21562 ( .A1(n22737), .A2(n22698), .ZN(n22738) );
  NAND2_X1 U21563 ( .A1(n22737), .A2(n22701), .ZN(n22740) );
  NAND2_X1 U21564 ( .A1(n22754), .A2(n22701), .ZN(n22757) );
  NAND2_X1 U21565 ( .A1(n22737), .A2(n22716), .ZN(n22750) );
  NAND2_X1 U21566 ( .A1(n22737), .A2(n22694), .ZN(n22735) );
  NAND2_X1 U21567 ( .A1(n22754), .A2(n22698), .ZN(n22755) );
  NAND2_X1 U21568 ( .A1(n22720), .A2(n22710), .ZN(n22729) );
  NAND2_X1 U21569 ( .A1(n22720), .A2(n22716), .ZN(n22733) );
  NAND2_X1 U21570 ( .A1(n22737), .A2(n22707), .ZN(n22744) );
  NAND2_X1 U21571 ( .A1(n22737), .A2(n22710), .ZN(n22746) );
  NAND2_X1 U21572 ( .A1(n22754), .A2(n22716), .ZN(n22767) );
  NAND2_X1 U21573 ( .A1(n22754), .A2(n22713), .ZN(n22765) );
  NAND2_X1 U21574 ( .A1(n22720), .A2(n22713), .ZN(n22731) );
  NAND2_X1 U21575 ( .A1(n22720), .A2(n22707), .ZN(n22727) );
  NAND2_X1 U21576 ( .A1(n25146), .A2(n25144), .ZN(n23975) );
  NAND2_X1 U21577 ( .A1(n23947), .A2(n23945), .ZN(n22776) );
  BUF_X1 U21578 ( .A(n24010), .Z(n26493) );
  BUF_X1 U21579 ( .A(n22811), .Z(n26718) );
  BUF_X1 U21580 ( .A(n24015), .Z(n26465) );
  BUF_X1 U21581 ( .A(n24015), .Z(n26466) );
  BUF_X1 U21582 ( .A(n24015), .Z(n26467) );
  BUF_X1 U21583 ( .A(n24015), .Z(n26468) );
  BUF_X1 U21584 ( .A(n24015), .Z(n26469) );
  BUF_X1 U21585 ( .A(n22816), .Z(n26690) );
  BUF_X1 U21586 ( .A(n22816), .Z(n26691) );
  BUF_X1 U21587 ( .A(n22816), .Z(n26692) );
  BUF_X1 U21588 ( .A(n22816), .Z(n26693) );
  BUF_X1 U21589 ( .A(n22816), .Z(n26694) );
  BUF_X1 U21590 ( .A(n24014), .Z(n26475) );
  BUF_X1 U21591 ( .A(n24009), .Z(n26499) );
  BUF_X1 U21592 ( .A(n22815), .Z(n26700) );
  BUF_X1 U21593 ( .A(n22810), .Z(n26724) );
  BUF_X1 U21594 ( .A(n20626), .Z(n27474) );
  BUF_X1 U21595 ( .A(n20626), .Z(n27475) );
  BUF_X1 U21596 ( .A(n20707), .Z(n27284) );
  BUF_X1 U21597 ( .A(n20706), .Z(n27287) );
  BUF_X1 U21598 ( .A(n20705), .Z(n27290) );
  BUF_X1 U21599 ( .A(n20704), .Z(n27293) );
  BUF_X1 U21600 ( .A(n20703), .Z(n27296) );
  BUF_X1 U21601 ( .A(n20702), .Z(n27299) );
  BUF_X1 U21602 ( .A(n20701), .Z(n27302) );
  BUF_X1 U21603 ( .A(n20700), .Z(n27305) );
  BUF_X1 U21604 ( .A(n20699), .Z(n27308) );
  BUF_X1 U21605 ( .A(n20698), .Z(n27311) );
  BUF_X1 U21606 ( .A(n20697), .Z(n27314) );
  BUF_X1 U21607 ( .A(n20696), .Z(n27317) );
  BUF_X1 U21608 ( .A(n20695), .Z(n27320) );
  BUF_X1 U21609 ( .A(n20694), .Z(n27323) );
  BUF_X1 U21610 ( .A(n20693), .Z(n27326) );
  BUF_X1 U21611 ( .A(n20692), .Z(n27329) );
  BUF_X1 U21612 ( .A(n20691), .Z(n27332) );
  BUF_X1 U21613 ( .A(n20690), .Z(n27335) );
  BUF_X1 U21614 ( .A(n20689), .Z(n27338) );
  BUF_X1 U21615 ( .A(n20688), .Z(n27341) );
  BUF_X1 U21616 ( .A(n20687), .Z(n27344) );
  BUF_X1 U21617 ( .A(n20686), .Z(n27347) );
  BUF_X1 U21618 ( .A(n20685), .Z(n27350) );
  BUF_X1 U21619 ( .A(n20684), .Z(n27353) );
  BUF_X1 U21620 ( .A(n20683), .Z(n27356) );
  BUF_X1 U21621 ( .A(n20682), .Z(n27359) );
  BUF_X1 U21622 ( .A(n20681), .Z(n27362) );
  BUF_X1 U21623 ( .A(n20680), .Z(n27365) );
  BUF_X1 U21624 ( .A(n20679), .Z(n27368) );
  BUF_X1 U21625 ( .A(n20678), .Z(n27371) );
  BUF_X1 U21626 ( .A(n20677), .Z(n27374) );
  BUF_X1 U21627 ( .A(n20676), .Z(n27377) );
  BUF_X1 U21628 ( .A(n20675), .Z(n27380) );
  BUF_X1 U21629 ( .A(n20674), .Z(n27383) );
  BUF_X1 U21630 ( .A(n20673), .Z(n27386) );
  BUF_X1 U21631 ( .A(n20672), .Z(n27389) );
  BUF_X1 U21632 ( .A(n20671), .Z(n27392) );
  BUF_X1 U21633 ( .A(n20670), .Z(n27395) );
  BUF_X1 U21634 ( .A(n20669), .Z(n27398) );
  BUF_X1 U21635 ( .A(n20668), .Z(n27401) );
  BUF_X1 U21636 ( .A(n20667), .Z(n27404) );
  BUF_X1 U21637 ( .A(n20666), .Z(n27407) );
  BUF_X1 U21638 ( .A(n20665), .Z(n27410) );
  BUF_X1 U21639 ( .A(n20664), .Z(n27413) );
  BUF_X1 U21640 ( .A(n20663), .Z(n27416) );
  BUF_X1 U21641 ( .A(n20662), .Z(n27419) );
  BUF_X1 U21642 ( .A(n20661), .Z(n27422) );
  BUF_X1 U21643 ( .A(n20660), .Z(n27425) );
  BUF_X1 U21644 ( .A(n20659), .Z(n27428) );
  BUF_X1 U21645 ( .A(n20658), .Z(n27431) );
  BUF_X1 U21646 ( .A(n20657), .Z(n27434) );
  BUF_X1 U21647 ( .A(n20656), .Z(n27437) );
  BUF_X1 U21648 ( .A(n20655), .Z(n27440) );
  BUF_X1 U21649 ( .A(n20654), .Z(n27443) );
  BUF_X1 U21650 ( .A(n20653), .Z(n27446) );
  BUF_X1 U21651 ( .A(n20652), .Z(n27449) );
  BUF_X1 U21652 ( .A(n20651), .Z(n27452) );
  BUF_X1 U21653 ( .A(n20650), .Z(n27455) );
  BUF_X1 U21654 ( .A(n20649), .Z(n27458) );
  BUF_X1 U21655 ( .A(n20648), .Z(n27461) );
  BUF_X1 U21656 ( .A(n20647), .Z(n27464) );
  BUF_X1 U21657 ( .A(n20646), .Z(n27467) );
  BUF_X1 U21658 ( .A(n20645), .Z(n27470) );
  BUF_X1 U21659 ( .A(n20644), .Z(n27473) );
  BUF_X1 U21660 ( .A(n20626), .Z(n27476) );
  NAND2_X1 U21661 ( .A1(n25147), .A2(n25151), .ZN(n23989) );
  NAND2_X1 U21662 ( .A1(n25147), .A2(n25148), .ZN(n23974) );
  NAND2_X1 U21663 ( .A1(n23948), .A2(n23952), .ZN(n22790) );
  NAND2_X1 U21664 ( .A1(n23948), .A2(n23949), .ZN(n22775) );
  NAND2_X1 U21665 ( .A1(n25153), .A2(n25145), .ZN(n23999) );
  NAND2_X1 U21666 ( .A1(n23954), .A2(n23946), .ZN(n22800) );
  NAND2_X1 U21667 ( .A1(n25146), .A2(n25151), .ZN(n23979) );
  NAND2_X1 U21668 ( .A1(n23947), .A2(n23952), .ZN(n22780) );
  NAND2_X1 U21669 ( .A1(n25150), .A2(n25145), .ZN(n23984) );
  NAND2_X1 U21670 ( .A1(n23951), .A2(n23946), .ZN(n22785) );
  NAND2_X1 U21671 ( .A1(n25151), .A2(n25155), .ZN(n24004) );
  NAND2_X1 U21672 ( .A1(n23952), .A2(n23956), .ZN(n22805) );
  NAND2_X1 U21673 ( .A1(n22694), .A2(n22695), .ZN(n22692) );
  AND3_X1 U21674 ( .A1(n20642), .A2(n20641), .A3(n25165), .ZN(n24012) );
  AND3_X1 U21675 ( .A1(n20637), .A2(n20636), .A3(n23966), .ZN(n22813) );
  AND2_X1 U21676 ( .A1(n25147), .A2(n25145), .ZN(n23988) );
  AND2_X1 U21677 ( .A1(n23948), .A2(n23946), .ZN(n22789) );
  AND2_X1 U21678 ( .A1(n25153), .A2(n25144), .ZN(n24002) );
  AND2_X1 U21679 ( .A1(n23954), .A2(n23945), .ZN(n22803) );
  AND2_X1 U21680 ( .A1(n25155), .A2(n25148), .ZN(n23993) );
  AND2_X1 U21681 ( .A1(n23956), .A2(n23949), .ZN(n22794) );
  AND2_X1 U21682 ( .A1(n25146), .A2(n25145), .ZN(n23983) );
  AND2_X1 U21683 ( .A1(n25146), .A2(n25148), .ZN(n24008) );
  AND2_X1 U21684 ( .A1(n23947), .A2(n23946), .ZN(n22784) );
  AND2_X1 U21685 ( .A1(n23947), .A2(n23949), .ZN(n22809) );
  AND2_X1 U21686 ( .A1(n25150), .A2(n25148), .ZN(n23982) );
  AND2_X1 U21687 ( .A1(n23951), .A2(n23949), .ZN(n22783) );
  AND2_X1 U21688 ( .A1(n25143), .A2(n25145), .ZN(n23977) );
  AND2_X1 U21689 ( .A1(n25143), .A2(n25144), .ZN(n23978) );
  AND2_X1 U21690 ( .A1(n25143), .A2(n25148), .ZN(n24007) );
  AND2_X1 U21691 ( .A1(n23944), .A2(n23946), .ZN(n22778) );
  AND2_X1 U21692 ( .A1(n23944), .A2(n23945), .ZN(n22779) );
  AND2_X1 U21693 ( .A1(n23944), .A2(n23949), .ZN(n22808) );
  AND2_X1 U21694 ( .A1(n25145), .A2(n25155), .ZN(n23994) );
  AND2_X1 U21695 ( .A1(n23946), .A2(n23956), .ZN(n22795) );
  AND2_X1 U21696 ( .A1(n25163), .A2(n25148), .ZN(n24017) );
  AND2_X1 U21697 ( .A1(n25163), .A2(n25145), .ZN(n24018) );
  AND2_X1 U21698 ( .A1(n25163), .A2(n25151), .ZN(n24019) );
  AND2_X1 U21699 ( .A1(n25163), .A2(n25144), .ZN(n24013) );
  AND2_X1 U21700 ( .A1(n23964), .A2(n23949), .ZN(n22818) );
  AND2_X1 U21701 ( .A1(n23964), .A2(n23946), .ZN(n22819) );
  AND2_X1 U21702 ( .A1(n23964), .A2(n23952), .ZN(n22820) );
  AND2_X1 U21703 ( .A1(n23964), .A2(n23945), .ZN(n22814) );
  AND2_X1 U21704 ( .A1(n25151), .A2(n25150), .ZN(n23992) );
  AND2_X1 U21705 ( .A1(n25144), .A2(n25150), .ZN(n23987) );
  AND2_X1 U21706 ( .A1(n23952), .A2(n23951), .ZN(n22793) );
  AND2_X1 U21707 ( .A1(n23945), .A2(n23951), .ZN(n22788) );
  BUF_X1 U21708 ( .A(n24003), .Z(n26531) );
  BUF_X1 U21709 ( .A(n24003), .Z(n26532) );
  BUF_X1 U21710 ( .A(n22804), .Z(n26756) );
  BUF_X1 U21711 ( .A(n22804), .Z(n26757) );
  OAI221_X1 U21712 ( .B1(n21347), .B2(n26667), .C1(n21627), .C2(n26661), .A(
        n24926), .ZN(n24925) );
  AOI22_X1 U21713 ( .A1(n26655), .A2(n9402), .B1(n26649), .B2(n19234), .ZN(
        n24926) );
  OAI221_X1 U21714 ( .B1(n20759), .B2(n26565), .C1(n21987), .C2(n26559), .A(
        n24934), .ZN(n24933) );
  AOI22_X1 U21715 ( .A1(n26553), .A2(n19249), .B1(n26549), .B2(n4328), .ZN(
        n24934) );
  OAI221_X1 U21716 ( .B1(n21346), .B2(n26667), .C1(n21626), .C2(n26661), .A(
        n24908), .ZN(n24907) );
  AOI22_X1 U21717 ( .A1(n26655), .A2(n9399), .B1(n26649), .B2(n19217), .ZN(
        n24908) );
  OAI221_X1 U21718 ( .B1(n20758), .B2(n26565), .C1(n21986), .C2(n26559), .A(
        n24916), .ZN(n24915) );
  AOI22_X1 U21719 ( .A1(n26553), .A2(n19232), .B1(n26548), .B2(n4326), .ZN(
        n24916) );
  OAI221_X1 U21720 ( .B1(n21345), .B2(n26667), .C1(n21625), .C2(n26661), .A(
        n24890), .ZN(n24889) );
  AOI22_X1 U21721 ( .A1(n26655), .A2(n9396), .B1(n26649), .B2(n19200), .ZN(
        n24890) );
  OAI221_X1 U21722 ( .B1(n20757), .B2(n26565), .C1(n21985), .C2(n26559), .A(
        n24898), .ZN(n24897) );
  AOI22_X1 U21723 ( .A1(n26553), .A2(n19215), .B1(n26548), .B2(n4324), .ZN(
        n24898) );
  OAI221_X1 U21724 ( .B1(n21344), .B2(n26667), .C1(n21624), .C2(n26661), .A(
        n24872), .ZN(n24871) );
  AOI22_X1 U21725 ( .A1(n26655), .A2(n9393), .B1(n26649), .B2(n19183), .ZN(
        n24872) );
  OAI221_X1 U21726 ( .B1(n20756), .B2(n26565), .C1(n21984), .C2(n26559), .A(
        n24880), .ZN(n24879) );
  AOI22_X1 U21727 ( .A1(n26553), .A2(n19198), .B1(n26548), .B2(n4322), .ZN(
        n24880) );
  OAI221_X1 U21728 ( .B1(n21343), .B2(n26667), .C1(n21623), .C2(n26661), .A(
        n24854), .ZN(n24853) );
  AOI22_X1 U21729 ( .A1(n26655), .A2(n9390), .B1(n26649), .B2(n19166), .ZN(
        n24854) );
  OAI221_X1 U21730 ( .B1(n20755), .B2(n26565), .C1(n21983), .C2(n26559), .A(
        n24862), .ZN(n24861) );
  AOI22_X1 U21731 ( .A1(n26553), .A2(n19181), .B1(n26548), .B2(n4320), .ZN(
        n24862) );
  OAI221_X1 U21732 ( .B1(n21342), .B2(n26667), .C1(n21622), .C2(n26661), .A(
        n24836), .ZN(n24835) );
  AOI22_X1 U21733 ( .A1(n26655), .A2(n9387), .B1(n26649), .B2(n19149), .ZN(
        n24836) );
  OAI221_X1 U21734 ( .B1(n20754), .B2(n26565), .C1(n21982), .C2(n26559), .A(
        n24844), .ZN(n24843) );
  AOI22_X1 U21735 ( .A1(n26553), .A2(n19164), .B1(n26547), .B2(n4318), .ZN(
        n24844) );
  OAI221_X1 U21736 ( .B1(n21341), .B2(n26667), .C1(n21621), .C2(n26661), .A(
        n24818), .ZN(n24817) );
  AOI22_X1 U21737 ( .A1(n26655), .A2(n9384), .B1(n26649), .B2(n19132), .ZN(
        n24818) );
  OAI221_X1 U21738 ( .B1(n20753), .B2(n26565), .C1(n21981), .C2(n26559), .A(
        n24826), .ZN(n24825) );
  AOI22_X1 U21739 ( .A1(n26553), .A2(n19147), .B1(n26547), .B2(n4316), .ZN(
        n24826) );
  OAI221_X1 U21740 ( .B1(n21340), .B2(n26667), .C1(n21620), .C2(n26661), .A(
        n24800), .ZN(n24799) );
  AOI22_X1 U21741 ( .A1(n26655), .A2(n9381), .B1(n26649), .B2(n19115), .ZN(
        n24800) );
  OAI221_X1 U21742 ( .B1(n20752), .B2(n26565), .C1(n21980), .C2(n26559), .A(
        n24808), .ZN(n24807) );
  AOI22_X1 U21743 ( .A1(n26553), .A2(n19130), .B1(n26547), .B2(n4314), .ZN(
        n24808) );
  OAI221_X1 U21744 ( .B1(n21339), .B2(n26667), .C1(n21619), .C2(n26661), .A(
        n24782), .ZN(n24781) );
  AOI22_X1 U21745 ( .A1(n26655), .A2(n9378), .B1(n26649), .B2(n19098), .ZN(
        n24782) );
  OAI221_X1 U21746 ( .B1(n20751), .B2(n26565), .C1(n21979), .C2(n26559), .A(
        n24790), .ZN(n24789) );
  AOI22_X1 U21747 ( .A1(n26553), .A2(n19113), .B1(n26547), .B2(n4312), .ZN(
        n24790) );
  OAI221_X1 U21748 ( .B1(n21338), .B2(n26667), .C1(n21618), .C2(n26661), .A(
        n24764), .ZN(n24763) );
  AOI22_X1 U21749 ( .A1(n26655), .A2(n9375), .B1(n26649), .B2(n19081), .ZN(
        n24764) );
  OAI221_X1 U21750 ( .B1(n20750), .B2(n26565), .C1(n21978), .C2(n26559), .A(
        n24772), .ZN(n24771) );
  AOI22_X1 U21751 ( .A1(n26553), .A2(n19096), .B1(n26546), .B2(n4310), .ZN(
        n24772) );
  OAI221_X1 U21752 ( .B1(n21337), .B2(n26667), .C1(n21617), .C2(n26661), .A(
        n24746), .ZN(n24745) );
  AOI22_X1 U21753 ( .A1(n26655), .A2(n9372), .B1(n26649), .B2(n19064), .ZN(
        n24746) );
  OAI221_X1 U21754 ( .B1(n20749), .B2(n26565), .C1(n21977), .C2(n26559), .A(
        n24754), .ZN(n24753) );
  AOI22_X1 U21755 ( .A1(n26553), .A2(n19079), .B1(n26546), .B2(n4308), .ZN(
        n24754) );
  OAI221_X1 U21756 ( .B1(n21336), .B2(n26667), .C1(n21616), .C2(n26661), .A(
        n24728), .ZN(n24727) );
  AOI22_X1 U21757 ( .A1(n26655), .A2(n9369), .B1(n26649), .B2(n19047), .ZN(
        n24728) );
  OAI221_X1 U21758 ( .B1(n20748), .B2(n26565), .C1(n21976), .C2(n26559), .A(
        n24736), .ZN(n24735) );
  AOI22_X1 U21759 ( .A1(n26553), .A2(n19062), .B1(n26546), .B2(n4306), .ZN(
        n24736) );
  OAI221_X1 U21760 ( .B1(n21335), .B2(n26668), .C1(n21615), .C2(n26662), .A(
        n24710), .ZN(n24709) );
  AOI22_X1 U21761 ( .A1(n26656), .A2(n9366), .B1(n26650), .B2(n19030), .ZN(
        n24710) );
  OAI221_X1 U21762 ( .B1(n20747), .B2(n26566), .C1(n21975), .C2(n26560), .A(
        n24718), .ZN(n24717) );
  AOI22_X1 U21763 ( .A1(n26554), .A2(n19045), .B1(n26546), .B2(n4304), .ZN(
        n24718) );
  OAI221_X1 U21764 ( .B1(n21334), .B2(n26668), .C1(n21614), .C2(n26662), .A(
        n24692), .ZN(n24691) );
  AOI22_X1 U21765 ( .A1(n26656), .A2(n9363), .B1(n26650), .B2(n19013), .ZN(
        n24692) );
  OAI221_X1 U21766 ( .B1(n20746), .B2(n26566), .C1(n21974), .C2(n26560), .A(
        n24700), .ZN(n24699) );
  AOI22_X1 U21767 ( .A1(n26554), .A2(n19028), .B1(n26545), .B2(n4302), .ZN(
        n24700) );
  OAI221_X1 U21768 ( .B1(n21333), .B2(n26668), .C1(n21613), .C2(n26662), .A(
        n24674), .ZN(n24673) );
  AOI22_X1 U21769 ( .A1(n26656), .A2(n9360), .B1(n26650), .B2(n18996), .ZN(
        n24674) );
  OAI221_X1 U21770 ( .B1(n20745), .B2(n26566), .C1(n21973), .C2(n26560), .A(
        n24682), .ZN(n24681) );
  AOI22_X1 U21771 ( .A1(n26554), .A2(n19011), .B1(n26545), .B2(n4300), .ZN(
        n24682) );
  OAI221_X1 U21772 ( .B1(n21332), .B2(n26668), .C1(n21612), .C2(n26662), .A(
        n24656), .ZN(n24655) );
  AOI22_X1 U21773 ( .A1(n26656), .A2(n9357), .B1(n26650), .B2(n18979), .ZN(
        n24656) );
  OAI221_X1 U21774 ( .B1(n20744), .B2(n26566), .C1(n21972), .C2(n26560), .A(
        n24664), .ZN(n24663) );
  AOI22_X1 U21775 ( .A1(n26554), .A2(n18994), .B1(n26545), .B2(n4298), .ZN(
        n24664) );
  OAI221_X1 U21776 ( .B1(n21331), .B2(n26668), .C1(n21611), .C2(n26662), .A(
        n24638), .ZN(n24637) );
  AOI22_X1 U21777 ( .A1(n26656), .A2(n9354), .B1(n26650), .B2(n18962), .ZN(
        n24638) );
  OAI221_X1 U21778 ( .B1(n20743), .B2(n26566), .C1(n21971), .C2(n26560), .A(
        n24646), .ZN(n24645) );
  AOI22_X1 U21779 ( .A1(n26554), .A2(n18977), .B1(n26545), .B2(n4296), .ZN(
        n24646) );
  OAI221_X1 U21780 ( .B1(n21330), .B2(n26668), .C1(n21610), .C2(n26662), .A(
        n24620), .ZN(n24619) );
  AOI22_X1 U21781 ( .A1(n26656), .A2(n9351), .B1(n26650), .B2(n18945), .ZN(
        n24620) );
  OAI221_X1 U21782 ( .B1(n20742), .B2(n26566), .C1(n21970), .C2(n26560), .A(
        n24628), .ZN(n24627) );
  AOI22_X1 U21783 ( .A1(n26554), .A2(n18960), .B1(n26544), .B2(n4294), .ZN(
        n24628) );
  OAI221_X1 U21784 ( .B1(n21329), .B2(n26668), .C1(n21609), .C2(n26662), .A(
        n24602), .ZN(n24601) );
  AOI22_X1 U21785 ( .A1(n26656), .A2(n9348), .B1(n26650), .B2(n18928), .ZN(
        n24602) );
  OAI221_X1 U21786 ( .B1(n20741), .B2(n26566), .C1(n21969), .C2(n26560), .A(
        n24610), .ZN(n24609) );
  AOI22_X1 U21787 ( .A1(n26554), .A2(n18943), .B1(n26544), .B2(n4292), .ZN(
        n24610) );
  OAI221_X1 U21788 ( .B1(n21328), .B2(n26668), .C1(n21608), .C2(n26662), .A(
        n24584), .ZN(n24583) );
  AOI22_X1 U21789 ( .A1(n26656), .A2(n9345), .B1(n26650), .B2(n18911), .ZN(
        n24584) );
  OAI221_X1 U21790 ( .B1(n20740), .B2(n26566), .C1(n21968), .C2(n26560), .A(
        n24592), .ZN(n24591) );
  AOI22_X1 U21791 ( .A1(n26554), .A2(n18926), .B1(n26544), .B2(n4290), .ZN(
        n24592) );
  OAI221_X1 U21792 ( .B1(n21327), .B2(n26668), .C1(n21607), .C2(n26662), .A(
        n24566), .ZN(n24565) );
  AOI22_X1 U21793 ( .A1(n26656), .A2(n9342), .B1(n26650), .B2(n18894), .ZN(
        n24566) );
  OAI221_X1 U21794 ( .B1(n20739), .B2(n26566), .C1(n21967), .C2(n26560), .A(
        n24574), .ZN(n24573) );
  AOI22_X1 U21795 ( .A1(n26554), .A2(n18909), .B1(n26543), .B2(n4288), .ZN(
        n24574) );
  OAI221_X1 U21796 ( .B1(n21326), .B2(n26668), .C1(n21606), .C2(n26662), .A(
        n24548), .ZN(n24547) );
  AOI22_X1 U21797 ( .A1(n26656), .A2(n9339), .B1(n26650), .B2(n18877), .ZN(
        n24548) );
  OAI221_X1 U21798 ( .B1(n20738), .B2(n26566), .C1(n21966), .C2(n26560), .A(
        n24556), .ZN(n24555) );
  AOI22_X1 U21799 ( .A1(n26554), .A2(n18892), .B1(n26543), .B2(n4286), .ZN(
        n24556) );
  OAI221_X1 U21800 ( .B1(n21325), .B2(n26668), .C1(n21605), .C2(n26662), .A(
        n24530), .ZN(n24529) );
  AOI22_X1 U21801 ( .A1(n26656), .A2(n9336), .B1(n26650), .B2(n18860), .ZN(
        n24530) );
  OAI221_X1 U21802 ( .B1(n20737), .B2(n26566), .C1(n21965), .C2(n26560), .A(
        n24538), .ZN(n24537) );
  AOI22_X1 U21803 ( .A1(n26554), .A2(n18875), .B1(n26543), .B2(n4284), .ZN(
        n24538) );
  OAI221_X1 U21804 ( .B1(n21324), .B2(n26668), .C1(n21604), .C2(n26662), .A(
        n24512), .ZN(n24511) );
  AOI22_X1 U21805 ( .A1(n26656), .A2(n9333), .B1(n26650), .B2(n18843), .ZN(
        n24512) );
  OAI221_X1 U21806 ( .B1(n20736), .B2(n26566), .C1(n21964), .C2(n26560), .A(
        n24520), .ZN(n24519) );
  AOI22_X1 U21807 ( .A1(n26554), .A2(n18858), .B1(n26543), .B2(n4282), .ZN(
        n24520) );
  OAI221_X1 U21808 ( .B1(n21323), .B2(n26669), .C1(n21603), .C2(n26663), .A(
        n24494), .ZN(n24493) );
  AOI22_X1 U21809 ( .A1(n26657), .A2(n9330), .B1(n26651), .B2(n18826), .ZN(
        n24494) );
  OAI221_X1 U21810 ( .B1(n20735), .B2(n26567), .C1(n21963), .C2(n26561), .A(
        n24502), .ZN(n24501) );
  AOI22_X1 U21811 ( .A1(n26555), .A2(n18841), .B1(n26542), .B2(n4280), .ZN(
        n24502) );
  OAI221_X1 U21812 ( .B1(n21322), .B2(n26669), .C1(n21602), .C2(n26663), .A(
        n24476), .ZN(n24475) );
  AOI22_X1 U21813 ( .A1(n26657), .A2(n9327), .B1(n26651), .B2(n18809), .ZN(
        n24476) );
  OAI221_X1 U21814 ( .B1(n20734), .B2(n26567), .C1(n21962), .C2(n26561), .A(
        n24484), .ZN(n24483) );
  AOI22_X1 U21815 ( .A1(n26555), .A2(n18824), .B1(n26542), .B2(n4278), .ZN(
        n24484) );
  OAI221_X1 U21816 ( .B1(n21321), .B2(n26669), .C1(n21601), .C2(n26663), .A(
        n24458), .ZN(n24457) );
  AOI22_X1 U21817 ( .A1(n26657), .A2(n9324), .B1(n26651), .B2(n18792), .ZN(
        n24458) );
  OAI221_X1 U21818 ( .B1(n20733), .B2(n26567), .C1(n21961), .C2(n26561), .A(
        n24466), .ZN(n24465) );
  AOI22_X1 U21819 ( .A1(n26555), .A2(n18807), .B1(n26542), .B2(n4276), .ZN(
        n24466) );
  OAI221_X1 U21820 ( .B1(n21320), .B2(n26669), .C1(n21600), .C2(n26663), .A(
        n24440), .ZN(n24439) );
  AOI22_X1 U21821 ( .A1(n26657), .A2(n9321), .B1(n26651), .B2(n18775), .ZN(
        n24440) );
  OAI221_X1 U21822 ( .B1(n20732), .B2(n26567), .C1(n21960), .C2(n26561), .A(
        n24448), .ZN(n24447) );
  AOI22_X1 U21823 ( .A1(n26555), .A2(n18790), .B1(n26542), .B2(n4274), .ZN(
        n24448) );
  OAI221_X1 U21824 ( .B1(n21319), .B2(n26669), .C1(n21599), .C2(n26663), .A(
        n24422), .ZN(n24421) );
  AOI22_X1 U21825 ( .A1(n26657), .A2(n9318), .B1(n26651), .B2(n18758), .ZN(
        n24422) );
  OAI221_X1 U21826 ( .B1(n20731), .B2(n26567), .C1(n21959), .C2(n26561), .A(
        n24430), .ZN(n24429) );
  AOI22_X1 U21827 ( .A1(n26555), .A2(n18773), .B1(n26541), .B2(n4272), .ZN(
        n24430) );
  OAI221_X1 U21828 ( .B1(n21318), .B2(n26669), .C1(n21598), .C2(n26663), .A(
        n24404), .ZN(n24403) );
  AOI22_X1 U21829 ( .A1(n26657), .A2(n9315), .B1(n26651), .B2(n18741), .ZN(
        n24404) );
  OAI221_X1 U21830 ( .B1(n20730), .B2(n26567), .C1(n21958), .C2(n26561), .A(
        n24412), .ZN(n24411) );
  AOI22_X1 U21831 ( .A1(n26555), .A2(n18756), .B1(n26541), .B2(n4270), .ZN(
        n24412) );
  OAI221_X1 U21832 ( .B1(n21317), .B2(n26669), .C1(n21597), .C2(n26663), .A(
        n24386), .ZN(n24385) );
  AOI22_X1 U21833 ( .A1(n26657), .A2(n9312), .B1(n26651), .B2(n18724), .ZN(
        n24386) );
  OAI221_X1 U21834 ( .B1(n20729), .B2(n26567), .C1(n21957), .C2(n26561), .A(
        n24394), .ZN(n24393) );
  AOI22_X1 U21835 ( .A1(n26555), .A2(n18739), .B1(n26541), .B2(n4268), .ZN(
        n24394) );
  OAI221_X1 U21836 ( .B1(n21316), .B2(n26669), .C1(n21596), .C2(n26663), .A(
        n24368), .ZN(n24367) );
  AOI22_X1 U21837 ( .A1(n26657), .A2(n9309), .B1(n26651), .B2(n18707), .ZN(
        n24368) );
  OAI221_X1 U21838 ( .B1(n20728), .B2(n26567), .C1(n21956), .C2(n26561), .A(
        n24376), .ZN(n24375) );
  AOI22_X1 U21839 ( .A1(n26555), .A2(n18722), .B1(n26541), .B2(n4266), .ZN(
        n24376) );
  OAI221_X1 U21840 ( .B1(n21315), .B2(n26669), .C1(n21595), .C2(n26663), .A(
        n24350), .ZN(n24349) );
  AOI22_X1 U21841 ( .A1(n26657), .A2(n9306), .B1(n26651), .B2(n18690), .ZN(
        n24350) );
  OAI221_X1 U21842 ( .B1(n20727), .B2(n26567), .C1(n21955), .C2(n26561), .A(
        n24358), .ZN(n24357) );
  AOI22_X1 U21843 ( .A1(n26555), .A2(n18705), .B1(n26540), .B2(n4264), .ZN(
        n24358) );
  OAI221_X1 U21844 ( .B1(n21314), .B2(n26669), .C1(n21594), .C2(n26663), .A(
        n24332), .ZN(n24331) );
  AOI22_X1 U21845 ( .A1(n26657), .A2(n9303), .B1(n26651), .B2(n18673), .ZN(
        n24332) );
  OAI221_X1 U21846 ( .B1(n20726), .B2(n26567), .C1(n21954), .C2(n26561), .A(
        n24340), .ZN(n24339) );
  AOI22_X1 U21847 ( .A1(n26555), .A2(n18688), .B1(n26540), .B2(n4262), .ZN(
        n24340) );
  OAI221_X1 U21848 ( .B1(n21313), .B2(n26669), .C1(n21593), .C2(n26663), .A(
        n24314), .ZN(n24313) );
  AOI22_X1 U21849 ( .A1(n26657), .A2(n9300), .B1(n26651), .B2(n18656), .ZN(
        n24314) );
  OAI221_X1 U21850 ( .B1(n20725), .B2(n26567), .C1(n21953), .C2(n26561), .A(
        n24322), .ZN(n24321) );
  AOI22_X1 U21851 ( .A1(n26555), .A2(n18671), .B1(n26540), .B2(n4260), .ZN(
        n24322) );
  OAI221_X1 U21852 ( .B1(n21312), .B2(n26669), .C1(n21592), .C2(n26663), .A(
        n24296), .ZN(n24295) );
  AOI22_X1 U21853 ( .A1(n26657), .A2(n9297), .B1(n26651), .B2(n18639), .ZN(
        n24296) );
  OAI221_X1 U21854 ( .B1(n20724), .B2(n26567), .C1(n21952), .C2(n26561), .A(
        n24304), .ZN(n24303) );
  AOI22_X1 U21855 ( .A1(n26555), .A2(n18654), .B1(n26540), .B2(n4258), .ZN(
        n24304) );
  OAI221_X1 U21856 ( .B1(n21311), .B2(n26670), .C1(n21591), .C2(n26664), .A(
        n24278), .ZN(n24277) );
  AOI22_X1 U21857 ( .A1(n26658), .A2(n9294), .B1(n26652), .B2(n18622), .ZN(
        n24278) );
  OAI221_X1 U21858 ( .B1(n20723), .B2(n26568), .C1(n21951), .C2(n26562), .A(
        n24286), .ZN(n24285) );
  AOI22_X1 U21859 ( .A1(n26556), .A2(n18637), .B1(n26539), .B2(n4256), .ZN(
        n24286) );
  OAI221_X1 U21860 ( .B1(n21310), .B2(n26670), .C1(n21590), .C2(n26664), .A(
        n24260), .ZN(n24259) );
  AOI22_X1 U21861 ( .A1(n26658), .A2(n9291), .B1(n26652), .B2(n18605), .ZN(
        n24260) );
  OAI221_X1 U21862 ( .B1(n20722), .B2(n26568), .C1(n21950), .C2(n26562), .A(
        n24268), .ZN(n24267) );
  AOI22_X1 U21863 ( .A1(n26556), .A2(n18620), .B1(n26539), .B2(n4254), .ZN(
        n24268) );
  OAI221_X1 U21864 ( .B1(n21309), .B2(n26670), .C1(n21589), .C2(n26664), .A(
        n24242), .ZN(n24241) );
  AOI22_X1 U21865 ( .A1(n26658), .A2(n9288), .B1(n26652), .B2(n18588), .ZN(
        n24242) );
  OAI221_X1 U21866 ( .B1(n20721), .B2(n26568), .C1(n21949), .C2(n26562), .A(
        n24250), .ZN(n24249) );
  AOI22_X1 U21867 ( .A1(n26556), .A2(n18603), .B1(n26539), .B2(n4252), .ZN(
        n24250) );
  OAI221_X1 U21868 ( .B1(n21308), .B2(n26670), .C1(n21588), .C2(n26664), .A(
        n24224), .ZN(n24223) );
  AOI22_X1 U21869 ( .A1(n26658), .A2(n9285), .B1(n26652), .B2(n18571), .ZN(
        n24224) );
  OAI221_X1 U21870 ( .B1(n20720), .B2(n26568), .C1(n21948), .C2(n26562), .A(
        n24232), .ZN(n24231) );
  AOI22_X1 U21871 ( .A1(n26556), .A2(n18586), .B1(n26539), .B2(n4250), .ZN(
        n24232) );
  OAI221_X1 U21872 ( .B1(n21307), .B2(n26670), .C1(n21587), .C2(n26664), .A(
        n24206), .ZN(n24205) );
  AOI22_X1 U21873 ( .A1(n26658), .A2(n9282), .B1(n26652), .B2(n18554), .ZN(
        n24206) );
  OAI221_X1 U21874 ( .B1(n20719), .B2(n26568), .C1(n21947), .C2(n26562), .A(
        n24214), .ZN(n24213) );
  AOI22_X1 U21875 ( .A1(n26556), .A2(n18569), .B1(n26538), .B2(n4248), .ZN(
        n24214) );
  OAI221_X1 U21876 ( .B1(n21306), .B2(n26670), .C1(n21586), .C2(n26664), .A(
        n24188), .ZN(n24187) );
  AOI22_X1 U21877 ( .A1(n26658), .A2(n9279), .B1(n26652), .B2(n18537), .ZN(
        n24188) );
  OAI221_X1 U21878 ( .B1(n20718), .B2(n26568), .C1(n21946), .C2(n26562), .A(
        n24196), .ZN(n24195) );
  AOI22_X1 U21879 ( .A1(n26556), .A2(n18552), .B1(n26538), .B2(n4246), .ZN(
        n24196) );
  OAI221_X1 U21880 ( .B1(n21305), .B2(n26670), .C1(n21585), .C2(n26664), .A(
        n24170), .ZN(n24169) );
  AOI22_X1 U21881 ( .A1(n26658), .A2(n9276), .B1(n26652), .B2(n18520), .ZN(
        n24170) );
  OAI221_X1 U21882 ( .B1(n20717), .B2(n26568), .C1(n21945), .C2(n26562), .A(
        n24178), .ZN(n24177) );
  AOI22_X1 U21883 ( .A1(n26556), .A2(n18535), .B1(n26538), .B2(n4244), .ZN(
        n24178) );
  OAI221_X1 U21884 ( .B1(n21304), .B2(n26670), .C1(n21584), .C2(n26664), .A(
        n24152), .ZN(n24151) );
  AOI22_X1 U21885 ( .A1(n26658), .A2(n9273), .B1(n26652), .B2(n18503), .ZN(
        n24152) );
  OAI221_X1 U21886 ( .B1(n20716), .B2(n26568), .C1(n21944), .C2(n26562), .A(
        n24160), .ZN(n24159) );
  AOI22_X1 U21887 ( .A1(n26556), .A2(n18518), .B1(n26538), .B2(n4242), .ZN(
        n24160) );
  OAI221_X1 U21888 ( .B1(n21303), .B2(n26670), .C1(n21583), .C2(n26664), .A(
        n24134), .ZN(n24133) );
  AOI22_X1 U21889 ( .A1(n26658), .A2(n9270), .B1(n26652), .B2(n18486), .ZN(
        n24134) );
  OAI221_X1 U21890 ( .B1(n20715), .B2(n26568), .C1(n21943), .C2(n26562), .A(
        n24142), .ZN(n24141) );
  AOI22_X1 U21891 ( .A1(n26556), .A2(n18501), .B1(n26537), .B2(n4240), .ZN(
        n24142) );
  OAI221_X1 U21892 ( .B1(n21302), .B2(n26670), .C1(n21582), .C2(n26664), .A(
        n24116), .ZN(n24115) );
  AOI22_X1 U21893 ( .A1(n26658), .A2(n9267), .B1(n26652), .B2(n18469), .ZN(
        n24116) );
  OAI221_X1 U21894 ( .B1(n20714), .B2(n26568), .C1(n21942), .C2(n26562), .A(
        n24124), .ZN(n24123) );
  AOI22_X1 U21895 ( .A1(n26556), .A2(n18484), .B1(n26537), .B2(n4238), .ZN(
        n24124) );
  OAI221_X1 U21896 ( .B1(n21301), .B2(n26670), .C1(n21581), .C2(n26664), .A(
        n24098), .ZN(n24097) );
  AOI22_X1 U21897 ( .A1(n26658), .A2(n9264), .B1(n26652), .B2(n18452), .ZN(
        n24098) );
  OAI221_X1 U21898 ( .B1(n20713), .B2(n26568), .C1(n21941), .C2(n26562), .A(
        n24106), .ZN(n24105) );
  AOI22_X1 U21899 ( .A1(n26556), .A2(n18467), .B1(n26537), .B2(n4236), .ZN(
        n24106) );
  OAI221_X1 U21900 ( .B1(n21300), .B2(n26670), .C1(n21580), .C2(n26664), .A(
        n24080), .ZN(n24079) );
  AOI22_X1 U21901 ( .A1(n26658), .A2(n9261), .B1(n26652), .B2(n18435), .ZN(
        n24080) );
  OAI221_X1 U21902 ( .B1(n20712), .B2(n26568), .C1(n21940), .C2(n26562), .A(
        n24088), .ZN(n24087) );
  AOI22_X1 U21903 ( .A1(n26556), .A2(n18450), .B1(n26537), .B2(n4234), .ZN(
        n24088) );
  OAI221_X1 U21904 ( .B1(n21347), .B2(n26892), .C1(n21627), .C2(n26886), .A(
        n23727), .ZN(n23726) );
  AOI22_X1 U21905 ( .A1(n26880), .A2(n9402), .B1(n26874), .B2(n19234), .ZN(
        n23727) );
  OAI221_X1 U21906 ( .B1(n20759), .B2(n26790), .C1(n21987), .C2(n26784), .A(
        n23735), .ZN(n23734) );
  AOI22_X1 U21907 ( .A1(n26778), .A2(n19249), .B1(n26774), .B2(n4200), .ZN(
        n23735) );
  OAI221_X1 U21908 ( .B1(n21346), .B2(n26892), .C1(n21626), .C2(n26886), .A(
        n23709), .ZN(n23708) );
  AOI22_X1 U21909 ( .A1(n26880), .A2(n9399), .B1(n26874), .B2(n19217), .ZN(
        n23709) );
  OAI221_X1 U21910 ( .B1(n20758), .B2(n26790), .C1(n21986), .C2(n26784), .A(
        n23717), .ZN(n23716) );
  AOI22_X1 U21911 ( .A1(n26778), .A2(n19232), .B1(n26773), .B2(n4198), .ZN(
        n23717) );
  OAI221_X1 U21912 ( .B1(n21345), .B2(n26892), .C1(n21625), .C2(n26886), .A(
        n23691), .ZN(n23690) );
  AOI22_X1 U21913 ( .A1(n26880), .A2(n9396), .B1(n26874), .B2(n19200), .ZN(
        n23691) );
  OAI221_X1 U21914 ( .B1(n20757), .B2(n26790), .C1(n21985), .C2(n26784), .A(
        n23699), .ZN(n23698) );
  AOI22_X1 U21915 ( .A1(n26778), .A2(n19215), .B1(n26773), .B2(n4196), .ZN(
        n23699) );
  OAI221_X1 U21916 ( .B1(n21344), .B2(n26892), .C1(n21624), .C2(n26886), .A(
        n23673), .ZN(n23672) );
  AOI22_X1 U21917 ( .A1(n26880), .A2(n9393), .B1(n26874), .B2(n19183), .ZN(
        n23673) );
  OAI221_X1 U21918 ( .B1(n20756), .B2(n26790), .C1(n21984), .C2(n26784), .A(
        n23681), .ZN(n23680) );
  AOI22_X1 U21919 ( .A1(n26778), .A2(n19198), .B1(n26773), .B2(n4194), .ZN(
        n23681) );
  OAI221_X1 U21920 ( .B1(n21343), .B2(n26892), .C1(n21623), .C2(n26886), .A(
        n23655), .ZN(n23654) );
  AOI22_X1 U21921 ( .A1(n26880), .A2(n9390), .B1(n26874), .B2(n19166), .ZN(
        n23655) );
  OAI221_X1 U21922 ( .B1(n20755), .B2(n26790), .C1(n21983), .C2(n26784), .A(
        n23663), .ZN(n23662) );
  AOI22_X1 U21923 ( .A1(n26778), .A2(n19181), .B1(n26773), .B2(n4192), .ZN(
        n23663) );
  OAI221_X1 U21924 ( .B1(n21342), .B2(n26892), .C1(n21622), .C2(n26886), .A(
        n23637), .ZN(n23636) );
  AOI22_X1 U21925 ( .A1(n26880), .A2(n9387), .B1(n26874), .B2(n19149), .ZN(
        n23637) );
  OAI221_X1 U21926 ( .B1(n20754), .B2(n26790), .C1(n21982), .C2(n26784), .A(
        n23645), .ZN(n23644) );
  AOI22_X1 U21927 ( .A1(n26778), .A2(n19164), .B1(n26772), .B2(n4190), .ZN(
        n23645) );
  OAI221_X1 U21928 ( .B1(n21341), .B2(n26892), .C1(n21621), .C2(n26886), .A(
        n23619), .ZN(n23618) );
  AOI22_X1 U21929 ( .A1(n26880), .A2(n9384), .B1(n26874), .B2(n19132), .ZN(
        n23619) );
  OAI221_X1 U21930 ( .B1(n20753), .B2(n26790), .C1(n21981), .C2(n26784), .A(
        n23627), .ZN(n23626) );
  AOI22_X1 U21931 ( .A1(n26778), .A2(n19147), .B1(n26772), .B2(n4188), .ZN(
        n23627) );
  OAI221_X1 U21932 ( .B1(n21340), .B2(n26892), .C1(n21620), .C2(n26886), .A(
        n23601), .ZN(n23600) );
  AOI22_X1 U21933 ( .A1(n26880), .A2(n9381), .B1(n26874), .B2(n19115), .ZN(
        n23601) );
  OAI221_X1 U21934 ( .B1(n20752), .B2(n26790), .C1(n21980), .C2(n26784), .A(
        n23609), .ZN(n23608) );
  AOI22_X1 U21935 ( .A1(n26778), .A2(n19130), .B1(n26772), .B2(n4186), .ZN(
        n23609) );
  OAI221_X1 U21936 ( .B1(n21339), .B2(n26892), .C1(n21619), .C2(n26886), .A(
        n23583), .ZN(n23582) );
  AOI22_X1 U21937 ( .A1(n26880), .A2(n9378), .B1(n26874), .B2(n19098), .ZN(
        n23583) );
  OAI221_X1 U21938 ( .B1(n20751), .B2(n26790), .C1(n21979), .C2(n26784), .A(
        n23591), .ZN(n23590) );
  AOI22_X1 U21939 ( .A1(n26778), .A2(n19113), .B1(n26772), .B2(n4184), .ZN(
        n23591) );
  OAI221_X1 U21940 ( .B1(n21338), .B2(n26892), .C1(n21618), .C2(n26886), .A(
        n23565), .ZN(n23564) );
  AOI22_X1 U21941 ( .A1(n26880), .A2(n9375), .B1(n26874), .B2(n19081), .ZN(
        n23565) );
  OAI221_X1 U21942 ( .B1(n20750), .B2(n26790), .C1(n21978), .C2(n26784), .A(
        n23573), .ZN(n23572) );
  AOI22_X1 U21943 ( .A1(n26778), .A2(n19096), .B1(n26771), .B2(n4182), .ZN(
        n23573) );
  OAI221_X1 U21944 ( .B1(n21337), .B2(n26892), .C1(n21617), .C2(n26886), .A(
        n23547), .ZN(n23546) );
  AOI22_X1 U21945 ( .A1(n26880), .A2(n9372), .B1(n26874), .B2(n19064), .ZN(
        n23547) );
  OAI221_X1 U21946 ( .B1(n20749), .B2(n26790), .C1(n21977), .C2(n26784), .A(
        n23555), .ZN(n23554) );
  AOI22_X1 U21947 ( .A1(n26778), .A2(n19079), .B1(n26771), .B2(n4180), .ZN(
        n23555) );
  OAI221_X1 U21948 ( .B1(n21336), .B2(n26892), .C1(n21616), .C2(n26886), .A(
        n23529), .ZN(n23528) );
  AOI22_X1 U21949 ( .A1(n26880), .A2(n9369), .B1(n26874), .B2(n19047), .ZN(
        n23529) );
  OAI221_X1 U21950 ( .B1(n20748), .B2(n26790), .C1(n21976), .C2(n26784), .A(
        n23537), .ZN(n23536) );
  AOI22_X1 U21951 ( .A1(n26778), .A2(n19062), .B1(n26771), .B2(n4178), .ZN(
        n23537) );
  OAI221_X1 U21952 ( .B1(n21335), .B2(n26893), .C1(n21615), .C2(n26887), .A(
        n23511), .ZN(n23510) );
  AOI22_X1 U21953 ( .A1(n26881), .A2(n9366), .B1(n26875), .B2(n19030), .ZN(
        n23511) );
  OAI221_X1 U21954 ( .B1(n20747), .B2(n26791), .C1(n21975), .C2(n26785), .A(
        n23519), .ZN(n23518) );
  AOI22_X1 U21955 ( .A1(n26779), .A2(n19045), .B1(n26771), .B2(n4176), .ZN(
        n23519) );
  OAI221_X1 U21956 ( .B1(n21334), .B2(n26893), .C1(n21614), .C2(n26887), .A(
        n23493), .ZN(n23492) );
  AOI22_X1 U21957 ( .A1(n26881), .A2(n9363), .B1(n26875), .B2(n19013), .ZN(
        n23493) );
  OAI221_X1 U21958 ( .B1(n20746), .B2(n26791), .C1(n21974), .C2(n26785), .A(
        n23501), .ZN(n23500) );
  AOI22_X1 U21959 ( .A1(n26779), .A2(n19028), .B1(n26770), .B2(n4174), .ZN(
        n23501) );
  OAI221_X1 U21960 ( .B1(n21333), .B2(n26893), .C1(n21613), .C2(n26887), .A(
        n23475), .ZN(n23474) );
  AOI22_X1 U21961 ( .A1(n26881), .A2(n9360), .B1(n26875), .B2(n18996), .ZN(
        n23475) );
  OAI221_X1 U21962 ( .B1(n20745), .B2(n26791), .C1(n21973), .C2(n26785), .A(
        n23483), .ZN(n23482) );
  AOI22_X1 U21963 ( .A1(n26779), .A2(n19011), .B1(n26770), .B2(n4172), .ZN(
        n23483) );
  OAI221_X1 U21964 ( .B1(n21332), .B2(n26893), .C1(n21612), .C2(n26887), .A(
        n23457), .ZN(n23456) );
  AOI22_X1 U21965 ( .A1(n26881), .A2(n9357), .B1(n26875), .B2(n18979), .ZN(
        n23457) );
  OAI221_X1 U21966 ( .B1(n20744), .B2(n26791), .C1(n21972), .C2(n26785), .A(
        n23465), .ZN(n23464) );
  AOI22_X1 U21967 ( .A1(n26779), .A2(n18994), .B1(n26770), .B2(n4170), .ZN(
        n23465) );
  OAI221_X1 U21968 ( .B1(n21331), .B2(n26893), .C1(n21611), .C2(n26887), .A(
        n23439), .ZN(n23438) );
  AOI22_X1 U21969 ( .A1(n26881), .A2(n9354), .B1(n26875), .B2(n18962), .ZN(
        n23439) );
  OAI221_X1 U21970 ( .B1(n20743), .B2(n26791), .C1(n21971), .C2(n26785), .A(
        n23447), .ZN(n23446) );
  AOI22_X1 U21971 ( .A1(n26779), .A2(n18977), .B1(n26770), .B2(n4168), .ZN(
        n23447) );
  OAI221_X1 U21972 ( .B1(n21330), .B2(n26893), .C1(n21610), .C2(n26887), .A(
        n23421), .ZN(n23420) );
  AOI22_X1 U21973 ( .A1(n26881), .A2(n9351), .B1(n26875), .B2(n18945), .ZN(
        n23421) );
  OAI221_X1 U21974 ( .B1(n20742), .B2(n26791), .C1(n21970), .C2(n26785), .A(
        n23429), .ZN(n23428) );
  AOI22_X1 U21975 ( .A1(n26779), .A2(n18960), .B1(n26769), .B2(n4166), .ZN(
        n23429) );
  OAI221_X1 U21976 ( .B1(n21329), .B2(n26893), .C1(n21609), .C2(n26887), .A(
        n23403), .ZN(n23402) );
  AOI22_X1 U21977 ( .A1(n26881), .A2(n9348), .B1(n26875), .B2(n18928), .ZN(
        n23403) );
  OAI221_X1 U21978 ( .B1(n20741), .B2(n26791), .C1(n21969), .C2(n26785), .A(
        n23411), .ZN(n23410) );
  AOI22_X1 U21979 ( .A1(n26779), .A2(n18943), .B1(n26769), .B2(n4164), .ZN(
        n23411) );
  OAI221_X1 U21980 ( .B1(n21328), .B2(n26893), .C1(n21608), .C2(n26887), .A(
        n23385), .ZN(n23384) );
  AOI22_X1 U21981 ( .A1(n26881), .A2(n9345), .B1(n26875), .B2(n18911), .ZN(
        n23385) );
  OAI221_X1 U21982 ( .B1(n20740), .B2(n26791), .C1(n21968), .C2(n26785), .A(
        n23393), .ZN(n23392) );
  AOI22_X1 U21983 ( .A1(n26779), .A2(n18926), .B1(n26769), .B2(n4162), .ZN(
        n23393) );
  OAI221_X1 U21984 ( .B1(n21327), .B2(n26893), .C1(n21607), .C2(n26887), .A(
        n23367), .ZN(n23366) );
  AOI22_X1 U21985 ( .A1(n26881), .A2(n9342), .B1(n26875), .B2(n18894), .ZN(
        n23367) );
  OAI221_X1 U21986 ( .B1(n20739), .B2(n26791), .C1(n21967), .C2(n26785), .A(
        n23375), .ZN(n23374) );
  AOI22_X1 U21987 ( .A1(n26779), .A2(n18909), .B1(n26768), .B2(n4160), .ZN(
        n23375) );
  OAI221_X1 U21988 ( .B1(n21326), .B2(n26893), .C1(n21606), .C2(n26887), .A(
        n23349), .ZN(n23348) );
  AOI22_X1 U21989 ( .A1(n26881), .A2(n9339), .B1(n26875), .B2(n18877), .ZN(
        n23349) );
  OAI221_X1 U21990 ( .B1(n20738), .B2(n26791), .C1(n21966), .C2(n26785), .A(
        n23357), .ZN(n23356) );
  AOI22_X1 U21991 ( .A1(n26779), .A2(n18892), .B1(n26768), .B2(n4158), .ZN(
        n23357) );
  OAI221_X1 U21992 ( .B1(n21325), .B2(n26893), .C1(n21605), .C2(n26887), .A(
        n23331), .ZN(n23330) );
  AOI22_X1 U21993 ( .A1(n26881), .A2(n9336), .B1(n26875), .B2(n18860), .ZN(
        n23331) );
  OAI221_X1 U21994 ( .B1(n20737), .B2(n26791), .C1(n21965), .C2(n26785), .A(
        n23339), .ZN(n23338) );
  AOI22_X1 U21995 ( .A1(n26779), .A2(n18875), .B1(n26768), .B2(n4156), .ZN(
        n23339) );
  OAI221_X1 U21996 ( .B1(n21324), .B2(n26893), .C1(n21604), .C2(n26887), .A(
        n23313), .ZN(n23312) );
  AOI22_X1 U21997 ( .A1(n26881), .A2(n9333), .B1(n26875), .B2(n18843), .ZN(
        n23313) );
  OAI221_X1 U21998 ( .B1(n20736), .B2(n26791), .C1(n21964), .C2(n26785), .A(
        n23321), .ZN(n23320) );
  AOI22_X1 U21999 ( .A1(n26779), .A2(n18858), .B1(n26768), .B2(n4154), .ZN(
        n23321) );
  OAI221_X1 U22000 ( .B1(n21323), .B2(n26894), .C1(n21603), .C2(n26888), .A(
        n23295), .ZN(n23294) );
  AOI22_X1 U22001 ( .A1(n26882), .A2(n9330), .B1(n26876), .B2(n18826), .ZN(
        n23295) );
  OAI221_X1 U22002 ( .B1(n20735), .B2(n26792), .C1(n21963), .C2(n26786), .A(
        n23303), .ZN(n23302) );
  AOI22_X1 U22003 ( .A1(n26780), .A2(n18841), .B1(n26767), .B2(n4152), .ZN(
        n23303) );
  OAI221_X1 U22004 ( .B1(n21322), .B2(n26894), .C1(n21602), .C2(n26888), .A(
        n23277), .ZN(n23276) );
  AOI22_X1 U22005 ( .A1(n26882), .A2(n9327), .B1(n26876), .B2(n18809), .ZN(
        n23277) );
  OAI221_X1 U22006 ( .B1(n20734), .B2(n26792), .C1(n21962), .C2(n26786), .A(
        n23285), .ZN(n23284) );
  AOI22_X1 U22007 ( .A1(n26780), .A2(n18824), .B1(n26767), .B2(n4150), .ZN(
        n23285) );
  OAI221_X1 U22008 ( .B1(n21321), .B2(n26894), .C1(n21601), .C2(n26888), .A(
        n23259), .ZN(n23258) );
  AOI22_X1 U22009 ( .A1(n26882), .A2(n9324), .B1(n26876), .B2(n18792), .ZN(
        n23259) );
  OAI221_X1 U22010 ( .B1(n20733), .B2(n26792), .C1(n21961), .C2(n26786), .A(
        n23267), .ZN(n23266) );
  AOI22_X1 U22011 ( .A1(n26780), .A2(n18807), .B1(n26767), .B2(n4148), .ZN(
        n23267) );
  OAI221_X1 U22012 ( .B1(n21320), .B2(n26894), .C1(n21600), .C2(n26888), .A(
        n23241), .ZN(n23240) );
  AOI22_X1 U22013 ( .A1(n26882), .A2(n9321), .B1(n26876), .B2(n18775), .ZN(
        n23241) );
  OAI221_X1 U22014 ( .B1(n20732), .B2(n26792), .C1(n21960), .C2(n26786), .A(
        n23249), .ZN(n23248) );
  AOI22_X1 U22015 ( .A1(n26780), .A2(n18790), .B1(n26767), .B2(n4146), .ZN(
        n23249) );
  OAI221_X1 U22016 ( .B1(n21319), .B2(n26894), .C1(n21599), .C2(n26888), .A(
        n23223), .ZN(n23222) );
  AOI22_X1 U22017 ( .A1(n26882), .A2(n9318), .B1(n26876), .B2(n18758), .ZN(
        n23223) );
  OAI221_X1 U22018 ( .B1(n20731), .B2(n26792), .C1(n21959), .C2(n26786), .A(
        n23231), .ZN(n23230) );
  AOI22_X1 U22019 ( .A1(n26780), .A2(n18773), .B1(n26766), .B2(n4144), .ZN(
        n23231) );
  OAI221_X1 U22020 ( .B1(n21318), .B2(n26894), .C1(n21598), .C2(n26888), .A(
        n23205), .ZN(n23204) );
  AOI22_X1 U22021 ( .A1(n26882), .A2(n9315), .B1(n26876), .B2(n18741), .ZN(
        n23205) );
  OAI221_X1 U22022 ( .B1(n20730), .B2(n26792), .C1(n21958), .C2(n26786), .A(
        n23213), .ZN(n23212) );
  AOI22_X1 U22023 ( .A1(n26780), .A2(n18756), .B1(n26766), .B2(n4142), .ZN(
        n23213) );
  OAI221_X1 U22024 ( .B1(n21317), .B2(n26894), .C1(n21597), .C2(n26888), .A(
        n23187), .ZN(n23186) );
  AOI22_X1 U22025 ( .A1(n26882), .A2(n9312), .B1(n26876), .B2(n18724), .ZN(
        n23187) );
  OAI221_X1 U22026 ( .B1(n20729), .B2(n26792), .C1(n21957), .C2(n26786), .A(
        n23195), .ZN(n23194) );
  AOI22_X1 U22027 ( .A1(n26780), .A2(n18739), .B1(n26766), .B2(n4140), .ZN(
        n23195) );
  OAI221_X1 U22028 ( .B1(n21316), .B2(n26894), .C1(n21596), .C2(n26888), .A(
        n23169), .ZN(n23168) );
  AOI22_X1 U22029 ( .A1(n26882), .A2(n9309), .B1(n26876), .B2(n18707), .ZN(
        n23169) );
  OAI221_X1 U22030 ( .B1(n20728), .B2(n26792), .C1(n21956), .C2(n26786), .A(
        n23177), .ZN(n23176) );
  AOI22_X1 U22031 ( .A1(n26780), .A2(n18722), .B1(n26766), .B2(n4138), .ZN(
        n23177) );
  OAI221_X1 U22032 ( .B1(n21315), .B2(n26894), .C1(n21595), .C2(n26888), .A(
        n23151), .ZN(n23150) );
  AOI22_X1 U22033 ( .A1(n26882), .A2(n9306), .B1(n26876), .B2(n18690), .ZN(
        n23151) );
  OAI221_X1 U22034 ( .B1(n20727), .B2(n26792), .C1(n21955), .C2(n26786), .A(
        n23159), .ZN(n23158) );
  AOI22_X1 U22035 ( .A1(n26780), .A2(n18705), .B1(n26765), .B2(n4136), .ZN(
        n23159) );
  OAI221_X1 U22036 ( .B1(n21314), .B2(n26894), .C1(n21594), .C2(n26888), .A(
        n23133), .ZN(n23132) );
  AOI22_X1 U22037 ( .A1(n26882), .A2(n9303), .B1(n26876), .B2(n18673), .ZN(
        n23133) );
  OAI221_X1 U22038 ( .B1(n20726), .B2(n26792), .C1(n21954), .C2(n26786), .A(
        n23141), .ZN(n23140) );
  AOI22_X1 U22039 ( .A1(n26780), .A2(n18688), .B1(n26765), .B2(n4134), .ZN(
        n23141) );
  OAI221_X1 U22040 ( .B1(n21313), .B2(n26894), .C1(n21593), .C2(n26888), .A(
        n23115), .ZN(n23114) );
  AOI22_X1 U22041 ( .A1(n26882), .A2(n9300), .B1(n26876), .B2(n18656), .ZN(
        n23115) );
  OAI221_X1 U22042 ( .B1(n20725), .B2(n26792), .C1(n21953), .C2(n26786), .A(
        n23123), .ZN(n23122) );
  AOI22_X1 U22043 ( .A1(n26780), .A2(n18671), .B1(n26765), .B2(n4132), .ZN(
        n23123) );
  OAI221_X1 U22044 ( .B1(n21312), .B2(n26894), .C1(n21592), .C2(n26888), .A(
        n23097), .ZN(n23096) );
  AOI22_X1 U22045 ( .A1(n26882), .A2(n9297), .B1(n26876), .B2(n18639), .ZN(
        n23097) );
  OAI221_X1 U22046 ( .B1(n20724), .B2(n26792), .C1(n21952), .C2(n26786), .A(
        n23105), .ZN(n23104) );
  AOI22_X1 U22047 ( .A1(n26780), .A2(n18654), .B1(n26765), .B2(n4130), .ZN(
        n23105) );
  OAI221_X1 U22048 ( .B1(n21311), .B2(n26895), .C1(n21591), .C2(n26889), .A(
        n23079), .ZN(n23078) );
  AOI22_X1 U22049 ( .A1(n26883), .A2(n9294), .B1(n26877), .B2(n18622), .ZN(
        n23079) );
  OAI221_X1 U22050 ( .B1(n20723), .B2(n26793), .C1(n21951), .C2(n26787), .A(
        n23087), .ZN(n23086) );
  AOI22_X1 U22051 ( .A1(n26781), .A2(n18637), .B1(n26764), .B2(n4128), .ZN(
        n23087) );
  OAI221_X1 U22052 ( .B1(n21310), .B2(n26895), .C1(n21590), .C2(n26889), .A(
        n23061), .ZN(n23060) );
  AOI22_X1 U22053 ( .A1(n26883), .A2(n9291), .B1(n26877), .B2(n18605), .ZN(
        n23061) );
  OAI221_X1 U22054 ( .B1(n20722), .B2(n26793), .C1(n21950), .C2(n26787), .A(
        n23069), .ZN(n23068) );
  AOI22_X1 U22055 ( .A1(n26781), .A2(n18620), .B1(n26764), .B2(n4126), .ZN(
        n23069) );
  OAI221_X1 U22056 ( .B1(n21309), .B2(n26895), .C1(n21589), .C2(n26889), .A(
        n23043), .ZN(n23042) );
  AOI22_X1 U22057 ( .A1(n26883), .A2(n9288), .B1(n26877), .B2(n18588), .ZN(
        n23043) );
  OAI221_X1 U22058 ( .B1(n20721), .B2(n26793), .C1(n21949), .C2(n26787), .A(
        n23051), .ZN(n23050) );
  AOI22_X1 U22059 ( .A1(n26781), .A2(n18603), .B1(n26764), .B2(n4124), .ZN(
        n23051) );
  OAI221_X1 U22060 ( .B1(n21308), .B2(n26895), .C1(n21588), .C2(n26889), .A(
        n23025), .ZN(n23024) );
  AOI22_X1 U22061 ( .A1(n26883), .A2(n9285), .B1(n26877), .B2(n18571), .ZN(
        n23025) );
  OAI221_X1 U22062 ( .B1(n20720), .B2(n26793), .C1(n21948), .C2(n26787), .A(
        n23033), .ZN(n23032) );
  AOI22_X1 U22063 ( .A1(n26781), .A2(n18586), .B1(n26764), .B2(n4122), .ZN(
        n23033) );
  OAI221_X1 U22064 ( .B1(n21307), .B2(n26895), .C1(n21587), .C2(n26889), .A(
        n23007), .ZN(n23006) );
  AOI22_X1 U22065 ( .A1(n26883), .A2(n9282), .B1(n26877), .B2(n18554), .ZN(
        n23007) );
  OAI221_X1 U22066 ( .B1(n20719), .B2(n26793), .C1(n21947), .C2(n26787), .A(
        n23015), .ZN(n23014) );
  AOI22_X1 U22067 ( .A1(n26781), .A2(n18569), .B1(n26763), .B2(n4120), .ZN(
        n23015) );
  OAI221_X1 U22068 ( .B1(n21306), .B2(n26895), .C1(n21586), .C2(n26889), .A(
        n22989), .ZN(n22988) );
  AOI22_X1 U22069 ( .A1(n26883), .A2(n9279), .B1(n26877), .B2(n18537), .ZN(
        n22989) );
  OAI221_X1 U22070 ( .B1(n20718), .B2(n26793), .C1(n21946), .C2(n26787), .A(
        n22997), .ZN(n22996) );
  AOI22_X1 U22071 ( .A1(n26781), .A2(n18552), .B1(n26763), .B2(n4118), .ZN(
        n22997) );
  OAI221_X1 U22072 ( .B1(n21305), .B2(n26895), .C1(n21585), .C2(n26889), .A(
        n22971), .ZN(n22970) );
  AOI22_X1 U22073 ( .A1(n26883), .A2(n9276), .B1(n26877), .B2(n18520), .ZN(
        n22971) );
  OAI221_X1 U22074 ( .B1(n20717), .B2(n26793), .C1(n21945), .C2(n26787), .A(
        n22979), .ZN(n22978) );
  AOI22_X1 U22075 ( .A1(n26781), .A2(n18535), .B1(n26763), .B2(n4116), .ZN(
        n22979) );
  OAI221_X1 U22076 ( .B1(n21304), .B2(n26895), .C1(n21584), .C2(n26889), .A(
        n22953), .ZN(n22952) );
  AOI22_X1 U22077 ( .A1(n26883), .A2(n9273), .B1(n26877), .B2(n18503), .ZN(
        n22953) );
  OAI221_X1 U22078 ( .B1(n20716), .B2(n26793), .C1(n21944), .C2(n26787), .A(
        n22961), .ZN(n22960) );
  AOI22_X1 U22079 ( .A1(n26781), .A2(n18518), .B1(n26763), .B2(n4114), .ZN(
        n22961) );
  OAI221_X1 U22080 ( .B1(n21303), .B2(n26895), .C1(n21583), .C2(n26889), .A(
        n22935), .ZN(n22934) );
  AOI22_X1 U22081 ( .A1(n26883), .A2(n9270), .B1(n26877), .B2(n18486), .ZN(
        n22935) );
  OAI221_X1 U22082 ( .B1(n20715), .B2(n26793), .C1(n21943), .C2(n26787), .A(
        n22943), .ZN(n22942) );
  AOI22_X1 U22083 ( .A1(n26781), .A2(n18501), .B1(n26762), .B2(n4112), .ZN(
        n22943) );
  OAI221_X1 U22084 ( .B1(n21302), .B2(n26895), .C1(n21582), .C2(n26889), .A(
        n22917), .ZN(n22916) );
  AOI22_X1 U22085 ( .A1(n26883), .A2(n9267), .B1(n26877), .B2(n18469), .ZN(
        n22917) );
  OAI221_X1 U22086 ( .B1(n20714), .B2(n26793), .C1(n21942), .C2(n26787), .A(
        n22925), .ZN(n22924) );
  AOI22_X1 U22087 ( .A1(n26781), .A2(n18484), .B1(n26762), .B2(n4110), .ZN(
        n22925) );
  OAI221_X1 U22088 ( .B1(n21301), .B2(n26895), .C1(n21581), .C2(n26889), .A(
        n22899), .ZN(n22898) );
  AOI22_X1 U22089 ( .A1(n26883), .A2(n9264), .B1(n26877), .B2(n18452), .ZN(
        n22899) );
  OAI221_X1 U22090 ( .B1(n20713), .B2(n26793), .C1(n21941), .C2(n26787), .A(
        n22907), .ZN(n22906) );
  AOI22_X1 U22091 ( .A1(n26781), .A2(n18467), .B1(n26762), .B2(n4108), .ZN(
        n22907) );
  OAI221_X1 U22092 ( .B1(n21300), .B2(n26895), .C1(n21580), .C2(n26889), .A(
        n22881), .ZN(n22880) );
  AOI22_X1 U22093 ( .A1(n26883), .A2(n9261), .B1(n26877), .B2(n18435), .ZN(
        n22881) );
  OAI221_X1 U22094 ( .B1(n20712), .B2(n26793), .C1(n21940), .C2(n26787), .A(
        n22889), .ZN(n22888) );
  AOI22_X1 U22095 ( .A1(n26781), .A2(n18450), .B1(n26762), .B2(n4106), .ZN(
        n22889) );
  OAI221_X1 U22096 ( .B1(n21164), .B2(n26671), .C1(n21480), .C2(n26665), .A(
        n23976), .ZN(n23973) );
  AOI22_X1 U22097 ( .A1(n26659), .A2(n9249), .B1(n26653), .B2(n18367), .ZN(
        n23976) );
  OAI221_X1 U22098 ( .B1(n20708), .B2(n26569), .C1(n21504), .C2(n26563), .A(
        n24001), .ZN(n23998) );
  AOI22_X1 U22099 ( .A1(n26557), .A2(n18382), .B1(n26544), .B2(n4226), .ZN(
        n24001) );
  OAI221_X1 U22100 ( .B1(n21167), .B2(n26671), .C1(n21483), .C2(n26665), .A(
        n24062), .ZN(n24061) );
  AOI22_X1 U22101 ( .A1(n26659), .A2(n9258), .B1(n26653), .B2(n18418), .ZN(
        n24062) );
  OAI221_X1 U22102 ( .B1(n20711), .B2(n26569), .C1(n21507), .C2(n26563), .A(
        n24070), .ZN(n24069) );
  AOI22_X1 U22103 ( .A1(n26557), .A2(n18433), .B1(n26536), .B2(n4232), .ZN(
        n24070) );
  OAI221_X1 U22104 ( .B1(n21166), .B2(n26671), .C1(n21482), .C2(n26665), .A(
        n24044), .ZN(n24043) );
  AOI22_X1 U22105 ( .A1(n26659), .A2(n9255), .B1(n26653), .B2(n18401), .ZN(
        n24044) );
  OAI221_X1 U22106 ( .B1(n20710), .B2(n26569), .C1(n21506), .C2(n26563), .A(
        n24052), .ZN(n24051) );
  AOI22_X1 U22107 ( .A1(n26557), .A2(n18416), .B1(n26536), .B2(n4230), .ZN(
        n24052) );
  OAI221_X1 U22108 ( .B1(n21165), .B2(n26671), .C1(n21481), .C2(n26665), .A(
        n24026), .ZN(n24025) );
  AOI22_X1 U22109 ( .A1(n26659), .A2(n9252), .B1(n26653), .B2(n18384), .ZN(
        n24026) );
  OAI221_X1 U22110 ( .B1(n20709), .B2(n26569), .C1(n21505), .C2(n26563), .A(
        n24034), .ZN(n24033) );
  AOI22_X1 U22111 ( .A1(n26557), .A2(n18399), .B1(n26536), .B2(n4228), .ZN(
        n24034) );
  OAI221_X1 U22112 ( .B1(n21167), .B2(n26896), .C1(n21483), .C2(n26890), .A(
        n22863), .ZN(n22862) );
  AOI22_X1 U22113 ( .A1(n26884), .A2(n9258), .B1(n26878), .B2(n18418), .ZN(
        n22863) );
  OAI221_X1 U22114 ( .B1(n20711), .B2(n26794), .C1(n21507), .C2(n26788), .A(
        n22871), .ZN(n22870) );
  AOI22_X1 U22115 ( .A1(n26782), .A2(n18433), .B1(n26761), .B2(n4104), .ZN(
        n22871) );
  OAI221_X1 U22116 ( .B1(n21166), .B2(n26896), .C1(n21482), .C2(n26890), .A(
        n22845), .ZN(n22844) );
  AOI22_X1 U22117 ( .A1(n26884), .A2(n9255), .B1(n26878), .B2(n18401), .ZN(
        n22845) );
  OAI221_X1 U22118 ( .B1(n20710), .B2(n26794), .C1(n21506), .C2(n26788), .A(
        n22853), .ZN(n22852) );
  AOI22_X1 U22119 ( .A1(n26782), .A2(n18416), .B1(n26761), .B2(n4102), .ZN(
        n22853) );
  OAI221_X1 U22120 ( .B1(n21165), .B2(n26896), .C1(n21481), .C2(n26890), .A(
        n22827), .ZN(n22826) );
  AOI22_X1 U22121 ( .A1(n26884), .A2(n9252), .B1(n26878), .B2(n18384), .ZN(
        n22827) );
  OAI221_X1 U22122 ( .B1(n20709), .B2(n26794), .C1(n21505), .C2(n26788), .A(
        n22835), .ZN(n22834) );
  AOI22_X1 U22123 ( .A1(n26782), .A2(n18399), .B1(n26761), .B2(n4100), .ZN(
        n22835) );
  OAI221_X1 U22124 ( .B1(n21164), .B2(n26896), .C1(n21480), .C2(n26890), .A(
        n22777), .ZN(n22774) );
  AOI22_X1 U22125 ( .A1(n26884), .A2(n9249), .B1(n26878), .B2(n18367), .ZN(
        n22777) );
  OAI221_X1 U22126 ( .B1(n20708), .B2(n26794), .C1(n21504), .C2(n26788), .A(
        n22802), .ZN(n22799) );
  AOI22_X1 U22127 ( .A1(n26782), .A2(n18382), .B1(n26769), .B2(n4098), .ZN(
        n22802) );
  OAI221_X1 U22128 ( .B1(n21359), .B2(n26666), .C1(n21639), .C2(n26660), .A(
        n25142), .ZN(n25141) );
  AOI22_X1 U22129 ( .A1(n26654), .A2(n9438), .B1(n26648), .B2(n19438), .ZN(
        n25142) );
  OAI221_X1 U22130 ( .B1(n20771), .B2(n26564), .C1(n21999), .C2(n26558), .A(
        n25160), .ZN(n25159) );
  AOI22_X1 U22131 ( .A1(n26552), .A2(n19453), .B1(n26530), .B2(n4352), .ZN(
        n25160) );
  OAI221_X1 U22132 ( .B1(n21358), .B2(n26666), .C1(n21638), .C2(n26660), .A(
        n25124), .ZN(n25123) );
  AOI22_X1 U22133 ( .A1(n26654), .A2(n9435), .B1(n26648), .B2(n19421), .ZN(
        n25124) );
  OAI221_X1 U22134 ( .B1(n20770), .B2(n26564), .C1(n21998), .C2(n26558), .A(
        n25132), .ZN(n25131) );
  AOI22_X1 U22135 ( .A1(n26552), .A2(n19436), .B1(n26551), .B2(n4350), .ZN(
        n25132) );
  OAI221_X1 U22136 ( .B1(n21357), .B2(n26666), .C1(n21637), .C2(n26660), .A(
        n25106), .ZN(n25105) );
  AOI22_X1 U22137 ( .A1(n26654), .A2(n9432), .B1(n26648), .B2(n19404), .ZN(
        n25106) );
  OAI221_X1 U22138 ( .B1(n20769), .B2(n26564), .C1(n21997), .C2(n26558), .A(
        n25114), .ZN(n25113) );
  AOI22_X1 U22139 ( .A1(n26552), .A2(n19419), .B1(n26551), .B2(n4348), .ZN(
        n25114) );
  OAI221_X1 U22140 ( .B1(n21356), .B2(n26666), .C1(n21636), .C2(n26660), .A(
        n25088), .ZN(n25087) );
  AOI22_X1 U22141 ( .A1(n26654), .A2(n9429), .B1(n26648), .B2(n19387), .ZN(
        n25088) );
  OAI221_X1 U22142 ( .B1(n20768), .B2(n26564), .C1(n21996), .C2(n26558), .A(
        n25096), .ZN(n25095) );
  AOI22_X1 U22143 ( .A1(n26552), .A2(n19402), .B1(n26551), .B2(n4346), .ZN(
        n25096) );
  OAI221_X1 U22144 ( .B1(n21355), .B2(n26666), .C1(n21635), .C2(n26660), .A(
        n25070), .ZN(n25069) );
  AOI22_X1 U22145 ( .A1(n26654), .A2(n9426), .B1(n26648), .B2(n19370), .ZN(
        n25070) );
  OAI221_X1 U22146 ( .B1(n20767), .B2(n26564), .C1(n21995), .C2(n26558), .A(
        n25078), .ZN(n25077) );
  AOI22_X1 U22147 ( .A1(n26552), .A2(n19385), .B1(n26551), .B2(n4344), .ZN(
        n25078) );
  OAI221_X1 U22148 ( .B1(n21354), .B2(n26666), .C1(n21634), .C2(n26660), .A(
        n25052), .ZN(n25051) );
  AOI22_X1 U22149 ( .A1(n26654), .A2(n9423), .B1(n26648), .B2(n19353), .ZN(
        n25052) );
  OAI221_X1 U22150 ( .B1(n20766), .B2(n26564), .C1(n21994), .C2(n26558), .A(
        n25060), .ZN(n25059) );
  AOI22_X1 U22151 ( .A1(n26552), .A2(n19368), .B1(n26550), .B2(n4342), .ZN(
        n25060) );
  OAI221_X1 U22152 ( .B1(n21353), .B2(n26666), .C1(n21633), .C2(n26660), .A(
        n25034), .ZN(n25033) );
  AOI22_X1 U22153 ( .A1(n26654), .A2(n9420), .B1(n26648), .B2(n19336), .ZN(
        n25034) );
  OAI221_X1 U22154 ( .B1(n20765), .B2(n26564), .C1(n21993), .C2(n26558), .A(
        n25042), .ZN(n25041) );
  AOI22_X1 U22155 ( .A1(n26552), .A2(n19351), .B1(n26550), .B2(n4340), .ZN(
        n25042) );
  OAI221_X1 U22156 ( .B1(n21352), .B2(n26666), .C1(n21632), .C2(n26660), .A(
        n25016), .ZN(n25015) );
  AOI22_X1 U22157 ( .A1(n26654), .A2(n9417), .B1(n26648), .B2(n19319), .ZN(
        n25016) );
  OAI221_X1 U22158 ( .B1(n20764), .B2(n26564), .C1(n21992), .C2(n26558), .A(
        n25024), .ZN(n25023) );
  AOI22_X1 U22159 ( .A1(n26552), .A2(n19334), .B1(n26550), .B2(n4338), .ZN(
        n25024) );
  OAI221_X1 U22160 ( .B1(n21351), .B2(n26666), .C1(n21631), .C2(n26660), .A(
        n24998), .ZN(n24997) );
  AOI22_X1 U22161 ( .A1(n26654), .A2(n9414), .B1(n26648), .B2(n19302), .ZN(
        n24998) );
  OAI221_X1 U22162 ( .B1(n20763), .B2(n26564), .C1(n21991), .C2(n26558), .A(
        n25006), .ZN(n25005) );
  AOI22_X1 U22163 ( .A1(n26552), .A2(n19317), .B1(n26550), .B2(n4336), .ZN(
        n25006) );
  OAI221_X1 U22164 ( .B1(n21350), .B2(n26666), .C1(n21630), .C2(n26660), .A(
        n24980), .ZN(n24979) );
  AOI22_X1 U22165 ( .A1(n26654), .A2(n9411), .B1(n26648), .B2(n19285), .ZN(
        n24980) );
  OAI221_X1 U22166 ( .B1(n20762), .B2(n26564), .C1(n21990), .C2(n26558), .A(
        n24988), .ZN(n24987) );
  AOI22_X1 U22167 ( .A1(n26552), .A2(n19300), .B1(n26549), .B2(n4334), .ZN(
        n24988) );
  OAI221_X1 U22168 ( .B1(n21349), .B2(n26666), .C1(n21629), .C2(n26660), .A(
        n24962), .ZN(n24961) );
  AOI22_X1 U22169 ( .A1(n26654), .A2(n9408), .B1(n26648), .B2(n19268), .ZN(
        n24962) );
  OAI221_X1 U22170 ( .B1(n20761), .B2(n26564), .C1(n21989), .C2(n26558), .A(
        n24970), .ZN(n24969) );
  AOI22_X1 U22171 ( .A1(n26552), .A2(n19283), .B1(n26549), .B2(n4332), .ZN(
        n24970) );
  OAI221_X1 U22172 ( .B1(n21348), .B2(n26666), .C1(n21628), .C2(n26660), .A(
        n24944), .ZN(n24943) );
  AOI22_X1 U22173 ( .A1(n26654), .A2(n9405), .B1(n26648), .B2(n19251), .ZN(
        n24944) );
  OAI221_X1 U22174 ( .B1(n20760), .B2(n26564), .C1(n21988), .C2(n26558), .A(
        n24952), .ZN(n24951) );
  AOI22_X1 U22175 ( .A1(n26552), .A2(n19266), .B1(n26549), .B2(n4330), .ZN(
        n24952) );
  OAI221_X1 U22176 ( .B1(n21359), .B2(n26891), .C1(n21639), .C2(n26885), .A(
        n23943), .ZN(n23942) );
  AOI22_X1 U22177 ( .A1(n26879), .A2(n9438), .B1(n26873), .B2(n19438), .ZN(
        n23943) );
  OAI221_X1 U22178 ( .B1(n20771), .B2(n26789), .C1(n21999), .C2(n26783), .A(
        n23961), .ZN(n23960) );
  AOI22_X1 U22179 ( .A1(n26777), .A2(n19453), .B1(n26755), .B2(n4224), .ZN(
        n23961) );
  OAI221_X1 U22180 ( .B1(n21358), .B2(n26891), .C1(n21638), .C2(n26885), .A(
        n23925), .ZN(n23924) );
  AOI22_X1 U22181 ( .A1(n26879), .A2(n9435), .B1(n26873), .B2(n19421), .ZN(
        n23925) );
  OAI221_X1 U22182 ( .B1(n20770), .B2(n26789), .C1(n21998), .C2(n26783), .A(
        n23933), .ZN(n23932) );
  AOI22_X1 U22183 ( .A1(n26777), .A2(n19436), .B1(n26776), .B2(n4222), .ZN(
        n23933) );
  OAI221_X1 U22184 ( .B1(n21357), .B2(n26891), .C1(n21637), .C2(n26885), .A(
        n23907), .ZN(n23906) );
  AOI22_X1 U22185 ( .A1(n26879), .A2(n9432), .B1(n26873), .B2(n19404), .ZN(
        n23907) );
  OAI221_X1 U22186 ( .B1(n20769), .B2(n26789), .C1(n21997), .C2(n26783), .A(
        n23915), .ZN(n23914) );
  AOI22_X1 U22187 ( .A1(n26777), .A2(n19419), .B1(n26776), .B2(n4220), .ZN(
        n23915) );
  OAI221_X1 U22188 ( .B1(n21356), .B2(n26891), .C1(n21636), .C2(n26885), .A(
        n23889), .ZN(n23888) );
  AOI22_X1 U22189 ( .A1(n26879), .A2(n9429), .B1(n26873), .B2(n19387), .ZN(
        n23889) );
  OAI221_X1 U22190 ( .B1(n20768), .B2(n26789), .C1(n21996), .C2(n26783), .A(
        n23897), .ZN(n23896) );
  AOI22_X1 U22191 ( .A1(n26777), .A2(n19402), .B1(n26776), .B2(n4218), .ZN(
        n23897) );
  OAI221_X1 U22192 ( .B1(n21355), .B2(n26891), .C1(n21635), .C2(n26885), .A(
        n23871), .ZN(n23870) );
  AOI22_X1 U22193 ( .A1(n26879), .A2(n9426), .B1(n26873), .B2(n19370), .ZN(
        n23871) );
  OAI221_X1 U22194 ( .B1(n20767), .B2(n26789), .C1(n21995), .C2(n26783), .A(
        n23879), .ZN(n23878) );
  AOI22_X1 U22195 ( .A1(n26777), .A2(n19385), .B1(n26776), .B2(n4216), .ZN(
        n23879) );
  OAI221_X1 U22196 ( .B1(n21354), .B2(n26891), .C1(n21634), .C2(n26885), .A(
        n23853), .ZN(n23852) );
  AOI22_X1 U22197 ( .A1(n26879), .A2(n9423), .B1(n26873), .B2(n19353), .ZN(
        n23853) );
  OAI221_X1 U22198 ( .B1(n20766), .B2(n26789), .C1(n21994), .C2(n26783), .A(
        n23861), .ZN(n23860) );
  AOI22_X1 U22199 ( .A1(n26777), .A2(n19368), .B1(n26775), .B2(n4214), .ZN(
        n23861) );
  OAI221_X1 U22200 ( .B1(n21353), .B2(n26891), .C1(n21633), .C2(n26885), .A(
        n23835), .ZN(n23834) );
  AOI22_X1 U22201 ( .A1(n26879), .A2(n9420), .B1(n26873), .B2(n19336), .ZN(
        n23835) );
  OAI221_X1 U22202 ( .B1(n20765), .B2(n26789), .C1(n21993), .C2(n26783), .A(
        n23843), .ZN(n23842) );
  AOI22_X1 U22203 ( .A1(n26777), .A2(n19351), .B1(n26775), .B2(n4212), .ZN(
        n23843) );
  OAI221_X1 U22204 ( .B1(n21352), .B2(n26891), .C1(n21632), .C2(n26885), .A(
        n23817), .ZN(n23816) );
  AOI22_X1 U22205 ( .A1(n26879), .A2(n9417), .B1(n26873), .B2(n19319), .ZN(
        n23817) );
  OAI221_X1 U22206 ( .B1(n20764), .B2(n26789), .C1(n21992), .C2(n26783), .A(
        n23825), .ZN(n23824) );
  AOI22_X1 U22207 ( .A1(n26777), .A2(n19334), .B1(n26775), .B2(n4210), .ZN(
        n23825) );
  OAI221_X1 U22208 ( .B1(n21351), .B2(n26891), .C1(n21631), .C2(n26885), .A(
        n23799), .ZN(n23798) );
  AOI22_X1 U22209 ( .A1(n26879), .A2(n9414), .B1(n26873), .B2(n19302), .ZN(
        n23799) );
  OAI221_X1 U22210 ( .B1(n20763), .B2(n26789), .C1(n21991), .C2(n26783), .A(
        n23807), .ZN(n23806) );
  AOI22_X1 U22211 ( .A1(n26777), .A2(n19317), .B1(n26775), .B2(n4208), .ZN(
        n23807) );
  OAI221_X1 U22212 ( .B1(n21350), .B2(n26891), .C1(n21630), .C2(n26885), .A(
        n23781), .ZN(n23780) );
  AOI22_X1 U22213 ( .A1(n26879), .A2(n9411), .B1(n26873), .B2(n19285), .ZN(
        n23781) );
  OAI221_X1 U22214 ( .B1(n20762), .B2(n26789), .C1(n21990), .C2(n26783), .A(
        n23789), .ZN(n23788) );
  AOI22_X1 U22215 ( .A1(n26777), .A2(n19300), .B1(n26774), .B2(n4206), .ZN(
        n23789) );
  OAI221_X1 U22216 ( .B1(n21349), .B2(n26891), .C1(n21629), .C2(n26885), .A(
        n23763), .ZN(n23762) );
  AOI22_X1 U22217 ( .A1(n26879), .A2(n9408), .B1(n26873), .B2(n19268), .ZN(
        n23763) );
  OAI221_X1 U22218 ( .B1(n20761), .B2(n26789), .C1(n21989), .C2(n26783), .A(
        n23771), .ZN(n23770) );
  AOI22_X1 U22219 ( .A1(n26777), .A2(n19283), .B1(n26774), .B2(n4204), .ZN(
        n23771) );
  OAI221_X1 U22220 ( .B1(n21348), .B2(n26891), .C1(n21628), .C2(n26885), .A(
        n23745), .ZN(n23744) );
  AOI22_X1 U22221 ( .A1(n26879), .A2(n9405), .B1(n26873), .B2(n19251), .ZN(
        n23745) );
  OAI221_X1 U22222 ( .B1(n20760), .B2(n26789), .C1(n21988), .C2(n26783), .A(
        n23753), .ZN(n23752) );
  AOI22_X1 U22223 ( .A1(n26777), .A2(n19266), .B1(n26774), .B2(n4202), .ZN(
        n23753) );
  OAI221_X1 U22224 ( .B1(n22559), .B2(n26643), .C1(n21227), .C2(n26637), .A(
        n24927), .ZN(n24924) );
  AOI22_X1 U22225 ( .A1(n26631), .A2(n25760), .B1(n26625), .B2(n8603), .ZN(
        n24927) );
  OAI221_X1 U22226 ( .B1(n22679), .B2(n26520), .C1(n22487), .C2(n26514), .A(
        n24935), .ZN(n24932) );
  AOI22_X1 U22227 ( .A1(n26508), .A2(n26219), .B1(n26502), .B2(n26339), .ZN(
        n24935) );
  OAI221_X1 U22228 ( .B1(n22558), .B2(n26643), .C1(n21226), .C2(n26637), .A(
        n24909), .ZN(n24906) );
  AOI22_X1 U22229 ( .A1(n26631), .A2(n25765), .B1(n26625), .B2(n8600), .ZN(
        n24909) );
  OAI221_X1 U22230 ( .B1(n22678), .B2(n26520), .C1(n22486), .C2(n26514), .A(
        n24917), .ZN(n24914) );
  AOI22_X1 U22231 ( .A1(n26508), .A2(n26220), .B1(n26502), .B2(n26340), .ZN(
        n24917) );
  OAI221_X1 U22232 ( .B1(n22557), .B2(n26643), .C1(n21225), .C2(n26637), .A(
        n24891), .ZN(n24888) );
  AOI22_X1 U22233 ( .A1(n26631), .A2(n25770), .B1(n26625), .B2(n8597), .ZN(
        n24891) );
  OAI221_X1 U22234 ( .B1(n22677), .B2(n26520), .C1(n22485), .C2(n26514), .A(
        n24899), .ZN(n24896) );
  AOI22_X1 U22235 ( .A1(n26508), .A2(n26221), .B1(n26502), .B2(n26341), .ZN(
        n24899) );
  OAI221_X1 U22236 ( .B1(n22556), .B2(n26643), .C1(n21224), .C2(n26637), .A(
        n24873), .ZN(n24870) );
  AOI22_X1 U22237 ( .A1(n26631), .A2(n25775), .B1(n26625), .B2(n8594), .ZN(
        n24873) );
  OAI221_X1 U22238 ( .B1(n22676), .B2(n26520), .C1(n22484), .C2(n26514), .A(
        n24881), .ZN(n24878) );
  AOI22_X1 U22239 ( .A1(n26508), .A2(n26222), .B1(n26502), .B2(n26342), .ZN(
        n24881) );
  OAI221_X1 U22240 ( .B1(n22555), .B2(n26643), .C1(n21223), .C2(n26637), .A(
        n24855), .ZN(n24852) );
  AOI22_X1 U22241 ( .A1(n26631), .A2(n25780), .B1(n26625), .B2(n8591), .ZN(
        n24855) );
  OAI221_X1 U22242 ( .B1(n22675), .B2(n26520), .C1(n22483), .C2(n26514), .A(
        n24863), .ZN(n24860) );
  AOI22_X1 U22243 ( .A1(n26508), .A2(n26223), .B1(n26502), .B2(n26343), .ZN(
        n24863) );
  OAI221_X1 U22244 ( .B1(n22554), .B2(n26643), .C1(n21222), .C2(n26637), .A(
        n24837), .ZN(n24834) );
  AOI22_X1 U22245 ( .A1(n26631), .A2(n25785), .B1(n26625), .B2(n8588), .ZN(
        n24837) );
  OAI221_X1 U22246 ( .B1(n22674), .B2(n26520), .C1(n22482), .C2(n26514), .A(
        n24845), .ZN(n24842) );
  AOI22_X1 U22247 ( .A1(n26508), .A2(n26224), .B1(n26502), .B2(n26344), .ZN(
        n24845) );
  OAI221_X1 U22248 ( .B1(n22553), .B2(n26643), .C1(n21221), .C2(n26637), .A(
        n24819), .ZN(n24816) );
  AOI22_X1 U22249 ( .A1(n26631), .A2(n25790), .B1(n26625), .B2(n8585), .ZN(
        n24819) );
  OAI221_X1 U22250 ( .B1(n22673), .B2(n26520), .C1(n22481), .C2(n26514), .A(
        n24827), .ZN(n24824) );
  AOI22_X1 U22251 ( .A1(n26508), .A2(n26225), .B1(n26502), .B2(n26345), .ZN(
        n24827) );
  OAI221_X1 U22252 ( .B1(n22552), .B2(n26643), .C1(n21220), .C2(n26637), .A(
        n24801), .ZN(n24798) );
  AOI22_X1 U22253 ( .A1(n26631), .A2(n25795), .B1(n26625), .B2(n8582), .ZN(
        n24801) );
  OAI221_X1 U22254 ( .B1(n22672), .B2(n26520), .C1(n22480), .C2(n26514), .A(
        n24809), .ZN(n24806) );
  AOI22_X1 U22255 ( .A1(n26508), .A2(n26226), .B1(n26502), .B2(n26346), .ZN(
        n24809) );
  OAI221_X1 U22256 ( .B1(n22551), .B2(n26643), .C1(n21219), .C2(n26637), .A(
        n24783), .ZN(n24780) );
  AOI22_X1 U22257 ( .A1(n26631), .A2(n25800), .B1(n26625), .B2(n8579), .ZN(
        n24783) );
  OAI221_X1 U22258 ( .B1(n22671), .B2(n26520), .C1(n22479), .C2(n26514), .A(
        n24791), .ZN(n24788) );
  AOI22_X1 U22259 ( .A1(n26508), .A2(n26227), .B1(n26502), .B2(n26347), .ZN(
        n24791) );
  OAI221_X1 U22260 ( .B1(n22550), .B2(n26643), .C1(n21218), .C2(n26637), .A(
        n24765), .ZN(n24762) );
  AOI22_X1 U22261 ( .A1(n26631), .A2(n25805), .B1(n26625), .B2(n8576), .ZN(
        n24765) );
  OAI221_X1 U22262 ( .B1(n22670), .B2(n26520), .C1(n22478), .C2(n26514), .A(
        n24773), .ZN(n24770) );
  AOI22_X1 U22263 ( .A1(n26508), .A2(n26228), .B1(n26502), .B2(n26348), .ZN(
        n24773) );
  OAI221_X1 U22264 ( .B1(n22549), .B2(n26643), .C1(n21217), .C2(n26637), .A(
        n24747), .ZN(n24744) );
  AOI22_X1 U22265 ( .A1(n26631), .A2(n25810), .B1(n26625), .B2(n8573), .ZN(
        n24747) );
  OAI221_X1 U22266 ( .B1(n22669), .B2(n26520), .C1(n22477), .C2(n26514), .A(
        n24755), .ZN(n24752) );
  AOI22_X1 U22267 ( .A1(n26508), .A2(n26229), .B1(n26502), .B2(n26349), .ZN(
        n24755) );
  OAI221_X1 U22268 ( .B1(n22548), .B2(n26643), .C1(n21216), .C2(n26637), .A(
        n24729), .ZN(n24726) );
  AOI22_X1 U22269 ( .A1(n26631), .A2(n25815), .B1(n26625), .B2(n8570), .ZN(
        n24729) );
  OAI221_X1 U22270 ( .B1(n22668), .B2(n26520), .C1(n22476), .C2(n26514), .A(
        n24737), .ZN(n24734) );
  AOI22_X1 U22271 ( .A1(n26508), .A2(n26230), .B1(n26502), .B2(n26350), .ZN(
        n24737) );
  OAI221_X1 U22272 ( .B1(n22547), .B2(n26644), .C1(n21215), .C2(n26638), .A(
        n24711), .ZN(n24708) );
  AOI22_X1 U22273 ( .A1(n26632), .A2(n25820), .B1(n26626), .B2(n8567), .ZN(
        n24711) );
  OAI221_X1 U22274 ( .B1(n22667), .B2(n26521), .C1(n22475), .C2(n26515), .A(
        n24719), .ZN(n24716) );
  AOI22_X1 U22275 ( .A1(n26509), .A2(n26231), .B1(n26503), .B2(n26351), .ZN(
        n24719) );
  OAI221_X1 U22276 ( .B1(n22546), .B2(n26644), .C1(n21214), .C2(n26638), .A(
        n24693), .ZN(n24690) );
  AOI22_X1 U22277 ( .A1(n26632), .A2(n25825), .B1(n26626), .B2(n8564), .ZN(
        n24693) );
  OAI221_X1 U22278 ( .B1(n22666), .B2(n26521), .C1(n22474), .C2(n26515), .A(
        n24701), .ZN(n24698) );
  AOI22_X1 U22279 ( .A1(n26509), .A2(n26232), .B1(n26503), .B2(n26352), .ZN(
        n24701) );
  OAI221_X1 U22280 ( .B1(n22545), .B2(n26644), .C1(n21213), .C2(n26638), .A(
        n24675), .ZN(n24672) );
  AOI22_X1 U22281 ( .A1(n26632), .A2(n25830), .B1(n26626), .B2(n8561), .ZN(
        n24675) );
  OAI221_X1 U22282 ( .B1(n22665), .B2(n26521), .C1(n22473), .C2(n26515), .A(
        n24683), .ZN(n24680) );
  AOI22_X1 U22283 ( .A1(n26509), .A2(n26233), .B1(n26503), .B2(n26353), .ZN(
        n24683) );
  OAI221_X1 U22284 ( .B1(n22544), .B2(n26644), .C1(n21212), .C2(n26638), .A(
        n24657), .ZN(n24654) );
  AOI22_X1 U22285 ( .A1(n26632), .A2(n25835), .B1(n26626), .B2(n8558), .ZN(
        n24657) );
  OAI221_X1 U22286 ( .B1(n22664), .B2(n26521), .C1(n22472), .C2(n26515), .A(
        n24665), .ZN(n24662) );
  AOI22_X1 U22287 ( .A1(n26509), .A2(n26234), .B1(n26503), .B2(n26354), .ZN(
        n24665) );
  OAI221_X1 U22288 ( .B1(n22543), .B2(n26644), .C1(n21211), .C2(n26638), .A(
        n24639), .ZN(n24636) );
  AOI22_X1 U22289 ( .A1(n26632), .A2(n25840), .B1(n26626), .B2(n8555), .ZN(
        n24639) );
  OAI221_X1 U22290 ( .B1(n22663), .B2(n26521), .C1(n22471), .C2(n26515), .A(
        n24647), .ZN(n24644) );
  AOI22_X1 U22291 ( .A1(n26509), .A2(n26235), .B1(n26503), .B2(n26355), .ZN(
        n24647) );
  OAI221_X1 U22292 ( .B1(n22542), .B2(n26644), .C1(n21210), .C2(n26638), .A(
        n24621), .ZN(n24618) );
  AOI22_X1 U22293 ( .A1(n26632), .A2(n25845), .B1(n26626), .B2(n8552), .ZN(
        n24621) );
  OAI221_X1 U22294 ( .B1(n22662), .B2(n26521), .C1(n22470), .C2(n26515), .A(
        n24629), .ZN(n24626) );
  AOI22_X1 U22295 ( .A1(n26509), .A2(n26236), .B1(n26503), .B2(n26356), .ZN(
        n24629) );
  OAI221_X1 U22296 ( .B1(n22541), .B2(n26644), .C1(n21209), .C2(n26638), .A(
        n24603), .ZN(n24600) );
  AOI22_X1 U22297 ( .A1(n26632), .A2(n25850), .B1(n26626), .B2(n8549), .ZN(
        n24603) );
  OAI221_X1 U22298 ( .B1(n22661), .B2(n26521), .C1(n22469), .C2(n26515), .A(
        n24611), .ZN(n24608) );
  AOI22_X1 U22299 ( .A1(n26509), .A2(n26237), .B1(n26503), .B2(n26357), .ZN(
        n24611) );
  OAI221_X1 U22300 ( .B1(n22540), .B2(n26644), .C1(n21208), .C2(n26638), .A(
        n24585), .ZN(n24582) );
  AOI22_X1 U22301 ( .A1(n26632), .A2(n25855), .B1(n26626), .B2(n8546), .ZN(
        n24585) );
  OAI221_X1 U22302 ( .B1(n22660), .B2(n26521), .C1(n22468), .C2(n26515), .A(
        n24593), .ZN(n24590) );
  AOI22_X1 U22303 ( .A1(n26509), .A2(n26238), .B1(n26503), .B2(n26358), .ZN(
        n24593) );
  OAI221_X1 U22304 ( .B1(n22539), .B2(n26644), .C1(n21207), .C2(n26638), .A(
        n24567), .ZN(n24564) );
  AOI22_X1 U22305 ( .A1(n26632), .A2(n25860), .B1(n26626), .B2(n8543), .ZN(
        n24567) );
  OAI221_X1 U22306 ( .B1(n22659), .B2(n26521), .C1(n22467), .C2(n26515), .A(
        n24575), .ZN(n24572) );
  AOI22_X1 U22307 ( .A1(n26509), .A2(n26239), .B1(n26503), .B2(n26359), .ZN(
        n24575) );
  OAI221_X1 U22308 ( .B1(n22538), .B2(n26644), .C1(n21206), .C2(n26638), .A(
        n24549), .ZN(n24546) );
  AOI22_X1 U22309 ( .A1(n26632), .A2(n25865), .B1(n26626), .B2(n8540), .ZN(
        n24549) );
  OAI221_X1 U22310 ( .B1(n22658), .B2(n26521), .C1(n22466), .C2(n26515), .A(
        n24557), .ZN(n24554) );
  AOI22_X1 U22311 ( .A1(n26509), .A2(n26240), .B1(n26503), .B2(n26360), .ZN(
        n24557) );
  OAI221_X1 U22312 ( .B1(n22537), .B2(n26644), .C1(n21205), .C2(n26638), .A(
        n24531), .ZN(n24528) );
  AOI22_X1 U22313 ( .A1(n26632), .A2(n25870), .B1(n26626), .B2(n8537), .ZN(
        n24531) );
  OAI221_X1 U22314 ( .B1(n22657), .B2(n26521), .C1(n22465), .C2(n26515), .A(
        n24539), .ZN(n24536) );
  AOI22_X1 U22315 ( .A1(n26509), .A2(n26241), .B1(n26503), .B2(n26361), .ZN(
        n24539) );
  OAI221_X1 U22316 ( .B1(n22536), .B2(n26644), .C1(n21204), .C2(n26638), .A(
        n24513), .ZN(n24510) );
  AOI22_X1 U22317 ( .A1(n26632), .A2(n25875), .B1(n26626), .B2(n8534), .ZN(
        n24513) );
  OAI221_X1 U22318 ( .B1(n22656), .B2(n26521), .C1(n22464), .C2(n26515), .A(
        n24521), .ZN(n24518) );
  AOI22_X1 U22319 ( .A1(n26509), .A2(n26242), .B1(n26503), .B2(n26362), .ZN(
        n24521) );
  OAI221_X1 U22320 ( .B1(n22535), .B2(n26645), .C1(n21203), .C2(n26639), .A(
        n24495), .ZN(n24492) );
  AOI22_X1 U22321 ( .A1(n26633), .A2(n25880), .B1(n26627), .B2(n8531), .ZN(
        n24495) );
  OAI221_X1 U22322 ( .B1(n22655), .B2(n26522), .C1(n22463), .C2(n26516), .A(
        n24503), .ZN(n24500) );
  AOI22_X1 U22323 ( .A1(n26510), .A2(n26243), .B1(n26504), .B2(n26363), .ZN(
        n24503) );
  OAI221_X1 U22324 ( .B1(n22534), .B2(n26645), .C1(n21202), .C2(n26639), .A(
        n24477), .ZN(n24474) );
  AOI22_X1 U22325 ( .A1(n26633), .A2(n25885), .B1(n26627), .B2(n8528), .ZN(
        n24477) );
  OAI221_X1 U22326 ( .B1(n22654), .B2(n26522), .C1(n22462), .C2(n26516), .A(
        n24485), .ZN(n24482) );
  AOI22_X1 U22327 ( .A1(n26510), .A2(n26244), .B1(n26504), .B2(n26364), .ZN(
        n24485) );
  OAI221_X1 U22328 ( .B1(n22533), .B2(n26645), .C1(n21201), .C2(n26639), .A(
        n24459), .ZN(n24456) );
  AOI22_X1 U22329 ( .A1(n26633), .A2(n25890), .B1(n26627), .B2(n8525), .ZN(
        n24459) );
  OAI221_X1 U22330 ( .B1(n22653), .B2(n26522), .C1(n22461), .C2(n26516), .A(
        n24467), .ZN(n24464) );
  AOI22_X1 U22331 ( .A1(n26510), .A2(n26245), .B1(n26504), .B2(n26365), .ZN(
        n24467) );
  OAI221_X1 U22332 ( .B1(n22532), .B2(n26645), .C1(n21200), .C2(n26639), .A(
        n24441), .ZN(n24438) );
  AOI22_X1 U22333 ( .A1(n26633), .A2(n25895), .B1(n26627), .B2(n8522), .ZN(
        n24441) );
  OAI221_X1 U22334 ( .B1(n22652), .B2(n26522), .C1(n22460), .C2(n26516), .A(
        n24449), .ZN(n24446) );
  AOI22_X1 U22335 ( .A1(n26510), .A2(n26246), .B1(n26504), .B2(n26366), .ZN(
        n24449) );
  OAI221_X1 U22336 ( .B1(n22531), .B2(n26645), .C1(n21199), .C2(n26639), .A(
        n24423), .ZN(n24420) );
  AOI22_X1 U22337 ( .A1(n26633), .A2(n25900), .B1(n26627), .B2(n8519), .ZN(
        n24423) );
  OAI221_X1 U22338 ( .B1(n22651), .B2(n26522), .C1(n22459), .C2(n26516), .A(
        n24431), .ZN(n24428) );
  AOI22_X1 U22339 ( .A1(n26510), .A2(n26247), .B1(n26504), .B2(n26367), .ZN(
        n24431) );
  OAI221_X1 U22340 ( .B1(n22530), .B2(n26645), .C1(n21198), .C2(n26639), .A(
        n24405), .ZN(n24402) );
  AOI22_X1 U22341 ( .A1(n26633), .A2(n25905), .B1(n26627), .B2(n8516), .ZN(
        n24405) );
  OAI221_X1 U22342 ( .B1(n22650), .B2(n26522), .C1(n22458), .C2(n26516), .A(
        n24413), .ZN(n24410) );
  AOI22_X1 U22343 ( .A1(n26510), .A2(n26248), .B1(n26504), .B2(n26368), .ZN(
        n24413) );
  OAI221_X1 U22344 ( .B1(n22529), .B2(n26645), .C1(n21197), .C2(n26639), .A(
        n24387), .ZN(n24384) );
  AOI22_X1 U22345 ( .A1(n26633), .A2(n25910), .B1(n26627), .B2(n8513), .ZN(
        n24387) );
  OAI221_X1 U22346 ( .B1(n22649), .B2(n26522), .C1(n22457), .C2(n26516), .A(
        n24395), .ZN(n24392) );
  AOI22_X1 U22347 ( .A1(n26510), .A2(n26249), .B1(n26504), .B2(n26369), .ZN(
        n24395) );
  OAI221_X1 U22348 ( .B1(n22528), .B2(n26645), .C1(n21196), .C2(n26639), .A(
        n24369), .ZN(n24366) );
  AOI22_X1 U22349 ( .A1(n26633), .A2(n25915), .B1(n26627), .B2(n8510), .ZN(
        n24369) );
  OAI221_X1 U22350 ( .B1(n22648), .B2(n26522), .C1(n22456), .C2(n26516), .A(
        n24377), .ZN(n24374) );
  AOI22_X1 U22351 ( .A1(n26510), .A2(n26250), .B1(n26504), .B2(n26370), .ZN(
        n24377) );
  OAI221_X1 U22352 ( .B1(n22527), .B2(n26645), .C1(n21195), .C2(n26639), .A(
        n24351), .ZN(n24348) );
  AOI22_X1 U22353 ( .A1(n26633), .A2(n25920), .B1(n26627), .B2(n8507), .ZN(
        n24351) );
  OAI221_X1 U22354 ( .B1(n22647), .B2(n26522), .C1(n22455), .C2(n26516), .A(
        n24359), .ZN(n24356) );
  AOI22_X1 U22355 ( .A1(n26510), .A2(n26251), .B1(n26504), .B2(n26371), .ZN(
        n24359) );
  OAI221_X1 U22356 ( .B1(n22526), .B2(n26645), .C1(n21194), .C2(n26639), .A(
        n24333), .ZN(n24330) );
  AOI22_X1 U22357 ( .A1(n26633), .A2(n25925), .B1(n26627), .B2(n8504), .ZN(
        n24333) );
  OAI221_X1 U22358 ( .B1(n22646), .B2(n26522), .C1(n22454), .C2(n26516), .A(
        n24341), .ZN(n24338) );
  AOI22_X1 U22359 ( .A1(n26510), .A2(n26252), .B1(n26504), .B2(n26372), .ZN(
        n24341) );
  OAI221_X1 U22360 ( .B1(n22525), .B2(n26645), .C1(n21193), .C2(n26639), .A(
        n24315), .ZN(n24312) );
  AOI22_X1 U22361 ( .A1(n26633), .A2(n25930), .B1(n26627), .B2(n8501), .ZN(
        n24315) );
  OAI221_X1 U22362 ( .B1(n22645), .B2(n26522), .C1(n22453), .C2(n26516), .A(
        n24323), .ZN(n24320) );
  AOI22_X1 U22363 ( .A1(n26510), .A2(n26253), .B1(n26504), .B2(n26373), .ZN(
        n24323) );
  OAI221_X1 U22364 ( .B1(n22524), .B2(n26645), .C1(n21192), .C2(n26639), .A(
        n24297), .ZN(n24294) );
  AOI22_X1 U22365 ( .A1(n26633), .A2(n25935), .B1(n26627), .B2(n8498), .ZN(
        n24297) );
  OAI221_X1 U22366 ( .B1(n22644), .B2(n26522), .C1(n22452), .C2(n26516), .A(
        n24305), .ZN(n24302) );
  AOI22_X1 U22367 ( .A1(n26510), .A2(n26254), .B1(n26504), .B2(n26374), .ZN(
        n24305) );
  OAI221_X1 U22368 ( .B1(n22523), .B2(n26646), .C1(n21191), .C2(n26640), .A(
        n24279), .ZN(n24276) );
  AOI22_X1 U22369 ( .A1(n26634), .A2(n25940), .B1(n26628), .B2(n8495), .ZN(
        n24279) );
  OAI221_X1 U22370 ( .B1(n22643), .B2(n26523), .C1(n22451), .C2(n26517), .A(
        n24287), .ZN(n24284) );
  AOI22_X1 U22371 ( .A1(n26511), .A2(n26255), .B1(n26505), .B2(n26375), .ZN(
        n24287) );
  OAI221_X1 U22372 ( .B1(n22522), .B2(n26646), .C1(n21190), .C2(n26640), .A(
        n24261), .ZN(n24258) );
  AOI22_X1 U22373 ( .A1(n26634), .A2(n25945), .B1(n26628), .B2(n8492), .ZN(
        n24261) );
  OAI221_X1 U22374 ( .B1(n22642), .B2(n26523), .C1(n22450), .C2(n26517), .A(
        n24269), .ZN(n24266) );
  AOI22_X1 U22375 ( .A1(n26511), .A2(n26256), .B1(n26505), .B2(n26376), .ZN(
        n24269) );
  OAI221_X1 U22376 ( .B1(n22521), .B2(n26646), .C1(n21189), .C2(n26640), .A(
        n24243), .ZN(n24240) );
  AOI22_X1 U22377 ( .A1(n26634), .A2(n25950), .B1(n26628), .B2(n8489), .ZN(
        n24243) );
  OAI221_X1 U22378 ( .B1(n22641), .B2(n26523), .C1(n22449), .C2(n26517), .A(
        n24251), .ZN(n24248) );
  AOI22_X1 U22379 ( .A1(n26511), .A2(n26257), .B1(n26505), .B2(n26377), .ZN(
        n24251) );
  OAI221_X1 U22380 ( .B1(n22520), .B2(n26646), .C1(n21188), .C2(n26640), .A(
        n24225), .ZN(n24222) );
  AOI22_X1 U22381 ( .A1(n26634), .A2(n25955), .B1(n26628), .B2(n8486), .ZN(
        n24225) );
  OAI221_X1 U22382 ( .B1(n22640), .B2(n26523), .C1(n22448), .C2(n26517), .A(
        n24233), .ZN(n24230) );
  AOI22_X1 U22383 ( .A1(n26511), .A2(n26258), .B1(n26505), .B2(n26378), .ZN(
        n24233) );
  OAI221_X1 U22384 ( .B1(n22519), .B2(n26646), .C1(n21187), .C2(n26640), .A(
        n24207), .ZN(n24204) );
  AOI22_X1 U22385 ( .A1(n26634), .A2(n25960), .B1(n26628), .B2(n8483), .ZN(
        n24207) );
  OAI221_X1 U22386 ( .B1(n22639), .B2(n26523), .C1(n22447), .C2(n26517), .A(
        n24215), .ZN(n24212) );
  AOI22_X1 U22387 ( .A1(n26511), .A2(n26259), .B1(n26505), .B2(n26379), .ZN(
        n24215) );
  OAI221_X1 U22388 ( .B1(n22518), .B2(n26646), .C1(n21186), .C2(n26640), .A(
        n24189), .ZN(n24186) );
  AOI22_X1 U22389 ( .A1(n26634), .A2(n25965), .B1(n26628), .B2(n8480), .ZN(
        n24189) );
  OAI221_X1 U22390 ( .B1(n22638), .B2(n26523), .C1(n22446), .C2(n26517), .A(
        n24197), .ZN(n24194) );
  AOI22_X1 U22391 ( .A1(n26511), .A2(n26260), .B1(n26505), .B2(n26380), .ZN(
        n24197) );
  OAI221_X1 U22392 ( .B1(n22517), .B2(n26646), .C1(n21185), .C2(n26640), .A(
        n24171), .ZN(n24168) );
  AOI22_X1 U22393 ( .A1(n26634), .A2(n25970), .B1(n26628), .B2(n8477), .ZN(
        n24171) );
  OAI221_X1 U22394 ( .B1(n22637), .B2(n26523), .C1(n22445), .C2(n26517), .A(
        n24179), .ZN(n24176) );
  AOI22_X1 U22395 ( .A1(n26511), .A2(n26261), .B1(n26505), .B2(n26381), .ZN(
        n24179) );
  OAI221_X1 U22396 ( .B1(n22516), .B2(n26646), .C1(n21184), .C2(n26640), .A(
        n24153), .ZN(n24150) );
  AOI22_X1 U22397 ( .A1(n26634), .A2(n25975), .B1(n26628), .B2(n8474), .ZN(
        n24153) );
  OAI221_X1 U22398 ( .B1(n22636), .B2(n26523), .C1(n22444), .C2(n26517), .A(
        n24161), .ZN(n24158) );
  AOI22_X1 U22399 ( .A1(n26511), .A2(n26262), .B1(n26505), .B2(n26382), .ZN(
        n24161) );
  OAI221_X1 U22400 ( .B1(n22515), .B2(n26646), .C1(n21183), .C2(n26640), .A(
        n24135), .ZN(n24132) );
  AOI22_X1 U22401 ( .A1(n26634), .A2(n25980), .B1(n26628), .B2(n8471), .ZN(
        n24135) );
  OAI221_X1 U22402 ( .B1(n22635), .B2(n26523), .C1(n22443), .C2(n26517), .A(
        n24143), .ZN(n24140) );
  AOI22_X1 U22403 ( .A1(n26511), .A2(n26263), .B1(n26505), .B2(n26383), .ZN(
        n24143) );
  OAI221_X1 U22404 ( .B1(n22514), .B2(n26646), .C1(n21182), .C2(n26640), .A(
        n24117), .ZN(n24114) );
  AOI22_X1 U22405 ( .A1(n26634), .A2(n25985), .B1(n26628), .B2(n8468), .ZN(
        n24117) );
  OAI221_X1 U22406 ( .B1(n22634), .B2(n26523), .C1(n22442), .C2(n26517), .A(
        n24125), .ZN(n24122) );
  AOI22_X1 U22407 ( .A1(n26511), .A2(n26264), .B1(n26505), .B2(n26384), .ZN(
        n24125) );
  OAI221_X1 U22408 ( .B1(n22513), .B2(n26646), .C1(n21181), .C2(n26640), .A(
        n24099), .ZN(n24096) );
  AOI22_X1 U22409 ( .A1(n26634), .A2(n25990), .B1(n26628), .B2(n8465), .ZN(
        n24099) );
  OAI221_X1 U22410 ( .B1(n22633), .B2(n26523), .C1(n22441), .C2(n26517), .A(
        n24107), .ZN(n24104) );
  AOI22_X1 U22411 ( .A1(n26511), .A2(n26265), .B1(n26505), .B2(n26385), .ZN(
        n24107) );
  OAI221_X1 U22412 ( .B1(n22512), .B2(n26646), .C1(n21180), .C2(n26640), .A(
        n24081), .ZN(n24078) );
  AOI22_X1 U22413 ( .A1(n26634), .A2(n25995), .B1(n26628), .B2(n8462), .ZN(
        n24081) );
  OAI221_X1 U22414 ( .B1(n22632), .B2(n26523), .C1(n22440), .C2(n26517), .A(
        n24089), .ZN(n24086) );
  AOI22_X1 U22415 ( .A1(n26511), .A2(n26266), .B1(n26505), .B2(n26386), .ZN(
        n24089) );
  OAI221_X1 U22416 ( .B1(n22559), .B2(n26868), .C1(n21227), .C2(n26862), .A(
        n23728), .ZN(n23725) );
  AOI22_X1 U22417 ( .A1(n26856), .A2(n25760), .B1(n26850), .B2(n8603), .ZN(
        n23728) );
  OAI221_X1 U22418 ( .B1(n22679), .B2(n26745), .C1(n22487), .C2(n26739), .A(
        n23736), .ZN(n23733) );
  AOI22_X1 U22419 ( .A1(n26733), .A2(n26219), .B1(n26727), .B2(n26339), .ZN(
        n23736) );
  OAI221_X1 U22420 ( .B1(n22558), .B2(n26868), .C1(n21226), .C2(n26862), .A(
        n23710), .ZN(n23707) );
  AOI22_X1 U22421 ( .A1(n26856), .A2(n25765), .B1(n26850), .B2(n8600), .ZN(
        n23710) );
  OAI221_X1 U22422 ( .B1(n22678), .B2(n26745), .C1(n22486), .C2(n26739), .A(
        n23718), .ZN(n23715) );
  AOI22_X1 U22423 ( .A1(n26733), .A2(n26220), .B1(n26727), .B2(n26340), .ZN(
        n23718) );
  OAI221_X1 U22424 ( .B1(n22557), .B2(n26868), .C1(n21225), .C2(n26862), .A(
        n23692), .ZN(n23689) );
  AOI22_X1 U22425 ( .A1(n26856), .A2(n25770), .B1(n26850), .B2(n8597), .ZN(
        n23692) );
  OAI221_X1 U22426 ( .B1(n22677), .B2(n26745), .C1(n22485), .C2(n26739), .A(
        n23700), .ZN(n23697) );
  AOI22_X1 U22427 ( .A1(n26733), .A2(n26221), .B1(n26727), .B2(n26341), .ZN(
        n23700) );
  OAI221_X1 U22428 ( .B1(n22556), .B2(n26868), .C1(n21224), .C2(n26862), .A(
        n23674), .ZN(n23671) );
  AOI22_X1 U22429 ( .A1(n26856), .A2(n25775), .B1(n26850), .B2(n8594), .ZN(
        n23674) );
  OAI221_X1 U22430 ( .B1(n22676), .B2(n26745), .C1(n22484), .C2(n26739), .A(
        n23682), .ZN(n23679) );
  AOI22_X1 U22431 ( .A1(n26733), .A2(n26222), .B1(n26727), .B2(n26342), .ZN(
        n23682) );
  OAI221_X1 U22432 ( .B1(n22555), .B2(n26868), .C1(n21223), .C2(n26862), .A(
        n23656), .ZN(n23653) );
  AOI22_X1 U22433 ( .A1(n26856), .A2(n25780), .B1(n26850), .B2(n8591), .ZN(
        n23656) );
  OAI221_X1 U22434 ( .B1(n22675), .B2(n26745), .C1(n22483), .C2(n26739), .A(
        n23664), .ZN(n23661) );
  AOI22_X1 U22435 ( .A1(n26733), .A2(n26223), .B1(n26727), .B2(n26343), .ZN(
        n23664) );
  OAI221_X1 U22436 ( .B1(n22554), .B2(n26868), .C1(n21222), .C2(n26862), .A(
        n23638), .ZN(n23635) );
  AOI22_X1 U22437 ( .A1(n26856), .A2(n25785), .B1(n26850), .B2(n8588), .ZN(
        n23638) );
  OAI221_X1 U22438 ( .B1(n22674), .B2(n26745), .C1(n22482), .C2(n26739), .A(
        n23646), .ZN(n23643) );
  AOI22_X1 U22439 ( .A1(n26733), .A2(n26224), .B1(n26727), .B2(n26344), .ZN(
        n23646) );
  OAI221_X1 U22440 ( .B1(n22553), .B2(n26868), .C1(n21221), .C2(n26862), .A(
        n23620), .ZN(n23617) );
  AOI22_X1 U22441 ( .A1(n26856), .A2(n25790), .B1(n26850), .B2(n8585), .ZN(
        n23620) );
  OAI221_X1 U22442 ( .B1(n22673), .B2(n26745), .C1(n22481), .C2(n26739), .A(
        n23628), .ZN(n23625) );
  AOI22_X1 U22443 ( .A1(n26733), .A2(n26225), .B1(n26727), .B2(n26345), .ZN(
        n23628) );
  OAI221_X1 U22444 ( .B1(n22552), .B2(n26868), .C1(n21220), .C2(n26862), .A(
        n23602), .ZN(n23599) );
  AOI22_X1 U22445 ( .A1(n26856), .A2(n25795), .B1(n26850), .B2(n8582), .ZN(
        n23602) );
  OAI221_X1 U22446 ( .B1(n22672), .B2(n26745), .C1(n22480), .C2(n26739), .A(
        n23610), .ZN(n23607) );
  AOI22_X1 U22447 ( .A1(n26733), .A2(n26226), .B1(n26727), .B2(n26346), .ZN(
        n23610) );
  OAI221_X1 U22448 ( .B1(n22551), .B2(n26868), .C1(n21219), .C2(n26862), .A(
        n23584), .ZN(n23581) );
  AOI22_X1 U22449 ( .A1(n26856), .A2(n25800), .B1(n26850), .B2(n8579), .ZN(
        n23584) );
  OAI221_X1 U22450 ( .B1(n22671), .B2(n26745), .C1(n22479), .C2(n26739), .A(
        n23592), .ZN(n23589) );
  AOI22_X1 U22451 ( .A1(n26733), .A2(n26227), .B1(n26727), .B2(n26347), .ZN(
        n23592) );
  OAI221_X1 U22452 ( .B1(n22550), .B2(n26868), .C1(n21218), .C2(n26862), .A(
        n23566), .ZN(n23563) );
  AOI22_X1 U22453 ( .A1(n26856), .A2(n25805), .B1(n26850), .B2(n8576), .ZN(
        n23566) );
  OAI221_X1 U22454 ( .B1(n22670), .B2(n26745), .C1(n22478), .C2(n26739), .A(
        n23574), .ZN(n23571) );
  AOI22_X1 U22455 ( .A1(n26733), .A2(n26228), .B1(n26727), .B2(n26348), .ZN(
        n23574) );
  OAI221_X1 U22456 ( .B1(n22549), .B2(n26868), .C1(n21217), .C2(n26862), .A(
        n23548), .ZN(n23545) );
  AOI22_X1 U22457 ( .A1(n26856), .A2(n25810), .B1(n26850), .B2(n8573), .ZN(
        n23548) );
  OAI221_X1 U22458 ( .B1(n22669), .B2(n26745), .C1(n22477), .C2(n26739), .A(
        n23556), .ZN(n23553) );
  AOI22_X1 U22459 ( .A1(n26733), .A2(n26229), .B1(n26727), .B2(n26349), .ZN(
        n23556) );
  OAI221_X1 U22460 ( .B1(n22548), .B2(n26868), .C1(n21216), .C2(n26862), .A(
        n23530), .ZN(n23527) );
  AOI22_X1 U22461 ( .A1(n26856), .A2(n25815), .B1(n26850), .B2(n8570), .ZN(
        n23530) );
  OAI221_X1 U22462 ( .B1(n22668), .B2(n26745), .C1(n22476), .C2(n26739), .A(
        n23538), .ZN(n23535) );
  AOI22_X1 U22463 ( .A1(n26733), .A2(n26230), .B1(n26727), .B2(n26350), .ZN(
        n23538) );
  OAI221_X1 U22464 ( .B1(n22547), .B2(n26869), .C1(n21215), .C2(n26863), .A(
        n23512), .ZN(n23509) );
  AOI22_X1 U22465 ( .A1(n26857), .A2(n25820), .B1(n26851), .B2(n8567), .ZN(
        n23512) );
  OAI221_X1 U22466 ( .B1(n22667), .B2(n26746), .C1(n22475), .C2(n26740), .A(
        n23520), .ZN(n23517) );
  AOI22_X1 U22467 ( .A1(n26734), .A2(n26231), .B1(n26728), .B2(n26351), .ZN(
        n23520) );
  OAI221_X1 U22468 ( .B1(n22546), .B2(n26869), .C1(n21214), .C2(n26863), .A(
        n23494), .ZN(n23491) );
  AOI22_X1 U22469 ( .A1(n26857), .A2(n25825), .B1(n26851), .B2(n8564), .ZN(
        n23494) );
  OAI221_X1 U22470 ( .B1(n22666), .B2(n26746), .C1(n22474), .C2(n26740), .A(
        n23502), .ZN(n23499) );
  AOI22_X1 U22471 ( .A1(n26734), .A2(n26232), .B1(n26728), .B2(n26352), .ZN(
        n23502) );
  OAI221_X1 U22472 ( .B1(n22545), .B2(n26869), .C1(n21213), .C2(n26863), .A(
        n23476), .ZN(n23473) );
  AOI22_X1 U22473 ( .A1(n26857), .A2(n25830), .B1(n26851), .B2(n8561), .ZN(
        n23476) );
  OAI221_X1 U22474 ( .B1(n22665), .B2(n26746), .C1(n22473), .C2(n26740), .A(
        n23484), .ZN(n23481) );
  AOI22_X1 U22475 ( .A1(n26734), .A2(n26233), .B1(n26728), .B2(n26353), .ZN(
        n23484) );
  OAI221_X1 U22476 ( .B1(n22544), .B2(n26869), .C1(n21212), .C2(n26863), .A(
        n23458), .ZN(n23455) );
  AOI22_X1 U22477 ( .A1(n26857), .A2(n25835), .B1(n26851), .B2(n8558), .ZN(
        n23458) );
  OAI221_X1 U22478 ( .B1(n22664), .B2(n26746), .C1(n22472), .C2(n26740), .A(
        n23466), .ZN(n23463) );
  AOI22_X1 U22479 ( .A1(n26734), .A2(n26234), .B1(n26728), .B2(n26354), .ZN(
        n23466) );
  OAI221_X1 U22480 ( .B1(n22543), .B2(n26869), .C1(n21211), .C2(n26863), .A(
        n23440), .ZN(n23437) );
  AOI22_X1 U22481 ( .A1(n26857), .A2(n25840), .B1(n26851), .B2(n8555), .ZN(
        n23440) );
  OAI221_X1 U22482 ( .B1(n22663), .B2(n26746), .C1(n22471), .C2(n26740), .A(
        n23448), .ZN(n23445) );
  AOI22_X1 U22483 ( .A1(n26734), .A2(n26235), .B1(n26728), .B2(n26355), .ZN(
        n23448) );
  OAI221_X1 U22484 ( .B1(n22542), .B2(n26869), .C1(n21210), .C2(n26863), .A(
        n23422), .ZN(n23419) );
  AOI22_X1 U22485 ( .A1(n26857), .A2(n25845), .B1(n26851), .B2(n8552), .ZN(
        n23422) );
  OAI221_X1 U22486 ( .B1(n22662), .B2(n26746), .C1(n22470), .C2(n26740), .A(
        n23430), .ZN(n23427) );
  AOI22_X1 U22487 ( .A1(n26734), .A2(n26236), .B1(n26728), .B2(n26356), .ZN(
        n23430) );
  OAI221_X1 U22488 ( .B1(n22541), .B2(n26869), .C1(n21209), .C2(n26863), .A(
        n23404), .ZN(n23401) );
  AOI22_X1 U22489 ( .A1(n26857), .A2(n25850), .B1(n26851), .B2(n8549), .ZN(
        n23404) );
  OAI221_X1 U22490 ( .B1(n22661), .B2(n26746), .C1(n22469), .C2(n26740), .A(
        n23412), .ZN(n23409) );
  AOI22_X1 U22491 ( .A1(n26734), .A2(n26237), .B1(n26728), .B2(n26357), .ZN(
        n23412) );
  OAI221_X1 U22492 ( .B1(n22540), .B2(n26869), .C1(n21208), .C2(n26863), .A(
        n23386), .ZN(n23383) );
  AOI22_X1 U22493 ( .A1(n26857), .A2(n25855), .B1(n26851), .B2(n8546), .ZN(
        n23386) );
  OAI221_X1 U22494 ( .B1(n22660), .B2(n26746), .C1(n22468), .C2(n26740), .A(
        n23394), .ZN(n23391) );
  AOI22_X1 U22495 ( .A1(n26734), .A2(n26238), .B1(n26728), .B2(n26358), .ZN(
        n23394) );
  OAI221_X1 U22496 ( .B1(n22539), .B2(n26869), .C1(n21207), .C2(n26863), .A(
        n23368), .ZN(n23365) );
  AOI22_X1 U22497 ( .A1(n26857), .A2(n25860), .B1(n26851), .B2(n8543), .ZN(
        n23368) );
  OAI221_X1 U22498 ( .B1(n22659), .B2(n26746), .C1(n22467), .C2(n26740), .A(
        n23376), .ZN(n23373) );
  AOI22_X1 U22499 ( .A1(n26734), .A2(n26239), .B1(n26728), .B2(n26359), .ZN(
        n23376) );
  OAI221_X1 U22500 ( .B1(n22538), .B2(n26869), .C1(n21206), .C2(n26863), .A(
        n23350), .ZN(n23347) );
  AOI22_X1 U22501 ( .A1(n26857), .A2(n25865), .B1(n26851), .B2(n8540), .ZN(
        n23350) );
  OAI221_X1 U22502 ( .B1(n22658), .B2(n26746), .C1(n22466), .C2(n26740), .A(
        n23358), .ZN(n23355) );
  AOI22_X1 U22503 ( .A1(n26734), .A2(n26240), .B1(n26728), .B2(n26360), .ZN(
        n23358) );
  OAI221_X1 U22504 ( .B1(n22537), .B2(n26869), .C1(n21205), .C2(n26863), .A(
        n23332), .ZN(n23329) );
  AOI22_X1 U22505 ( .A1(n26857), .A2(n25870), .B1(n26851), .B2(n8537), .ZN(
        n23332) );
  OAI221_X1 U22506 ( .B1(n22657), .B2(n26746), .C1(n22465), .C2(n26740), .A(
        n23340), .ZN(n23337) );
  AOI22_X1 U22507 ( .A1(n26734), .A2(n26241), .B1(n26728), .B2(n26361), .ZN(
        n23340) );
  OAI221_X1 U22508 ( .B1(n22536), .B2(n26869), .C1(n21204), .C2(n26863), .A(
        n23314), .ZN(n23311) );
  AOI22_X1 U22509 ( .A1(n26857), .A2(n25875), .B1(n26851), .B2(n8534), .ZN(
        n23314) );
  OAI221_X1 U22510 ( .B1(n22656), .B2(n26746), .C1(n22464), .C2(n26740), .A(
        n23322), .ZN(n23319) );
  AOI22_X1 U22511 ( .A1(n26734), .A2(n26242), .B1(n26728), .B2(n26362), .ZN(
        n23322) );
  OAI221_X1 U22512 ( .B1(n22535), .B2(n26870), .C1(n21203), .C2(n26864), .A(
        n23296), .ZN(n23293) );
  AOI22_X1 U22513 ( .A1(n26858), .A2(n25880), .B1(n26852), .B2(n8531), .ZN(
        n23296) );
  OAI221_X1 U22514 ( .B1(n22655), .B2(n26747), .C1(n22463), .C2(n26741), .A(
        n23304), .ZN(n23301) );
  AOI22_X1 U22515 ( .A1(n26735), .A2(n26243), .B1(n26729), .B2(n26363), .ZN(
        n23304) );
  OAI221_X1 U22516 ( .B1(n22534), .B2(n26870), .C1(n21202), .C2(n26864), .A(
        n23278), .ZN(n23275) );
  AOI22_X1 U22517 ( .A1(n26858), .A2(n25885), .B1(n26852), .B2(n8528), .ZN(
        n23278) );
  OAI221_X1 U22518 ( .B1(n22654), .B2(n26747), .C1(n22462), .C2(n26741), .A(
        n23286), .ZN(n23283) );
  AOI22_X1 U22519 ( .A1(n26735), .A2(n26244), .B1(n26729), .B2(n26364), .ZN(
        n23286) );
  OAI221_X1 U22520 ( .B1(n22533), .B2(n26870), .C1(n21201), .C2(n26864), .A(
        n23260), .ZN(n23257) );
  AOI22_X1 U22521 ( .A1(n26858), .A2(n25890), .B1(n26852), .B2(n8525), .ZN(
        n23260) );
  OAI221_X1 U22522 ( .B1(n22653), .B2(n26747), .C1(n22461), .C2(n26741), .A(
        n23268), .ZN(n23265) );
  AOI22_X1 U22523 ( .A1(n26735), .A2(n26245), .B1(n26729), .B2(n26365), .ZN(
        n23268) );
  OAI221_X1 U22524 ( .B1(n22532), .B2(n26870), .C1(n21200), .C2(n26864), .A(
        n23242), .ZN(n23239) );
  AOI22_X1 U22525 ( .A1(n26858), .A2(n25895), .B1(n26852), .B2(n8522), .ZN(
        n23242) );
  OAI221_X1 U22526 ( .B1(n22652), .B2(n26747), .C1(n22460), .C2(n26741), .A(
        n23250), .ZN(n23247) );
  AOI22_X1 U22527 ( .A1(n26735), .A2(n26246), .B1(n26729), .B2(n26366), .ZN(
        n23250) );
  OAI221_X1 U22528 ( .B1(n22531), .B2(n26870), .C1(n21199), .C2(n26864), .A(
        n23224), .ZN(n23221) );
  AOI22_X1 U22529 ( .A1(n26858), .A2(n25900), .B1(n26852), .B2(n8519), .ZN(
        n23224) );
  OAI221_X1 U22530 ( .B1(n22651), .B2(n26747), .C1(n22459), .C2(n26741), .A(
        n23232), .ZN(n23229) );
  AOI22_X1 U22531 ( .A1(n26735), .A2(n26247), .B1(n26729), .B2(n26367), .ZN(
        n23232) );
  OAI221_X1 U22532 ( .B1(n22530), .B2(n26870), .C1(n21198), .C2(n26864), .A(
        n23206), .ZN(n23203) );
  AOI22_X1 U22533 ( .A1(n26858), .A2(n25905), .B1(n26852), .B2(n8516), .ZN(
        n23206) );
  OAI221_X1 U22534 ( .B1(n22650), .B2(n26747), .C1(n22458), .C2(n26741), .A(
        n23214), .ZN(n23211) );
  AOI22_X1 U22535 ( .A1(n26735), .A2(n26248), .B1(n26729), .B2(n26368), .ZN(
        n23214) );
  OAI221_X1 U22536 ( .B1(n22529), .B2(n26870), .C1(n21197), .C2(n26864), .A(
        n23188), .ZN(n23185) );
  AOI22_X1 U22537 ( .A1(n26858), .A2(n25910), .B1(n26852), .B2(n8513), .ZN(
        n23188) );
  OAI221_X1 U22538 ( .B1(n22649), .B2(n26747), .C1(n22457), .C2(n26741), .A(
        n23196), .ZN(n23193) );
  AOI22_X1 U22539 ( .A1(n26735), .A2(n26249), .B1(n26729), .B2(n26369), .ZN(
        n23196) );
  OAI221_X1 U22540 ( .B1(n22528), .B2(n26870), .C1(n21196), .C2(n26864), .A(
        n23170), .ZN(n23167) );
  AOI22_X1 U22541 ( .A1(n26858), .A2(n25915), .B1(n26852), .B2(n8510), .ZN(
        n23170) );
  OAI221_X1 U22542 ( .B1(n22648), .B2(n26747), .C1(n22456), .C2(n26741), .A(
        n23178), .ZN(n23175) );
  AOI22_X1 U22543 ( .A1(n26735), .A2(n26250), .B1(n26729), .B2(n26370), .ZN(
        n23178) );
  OAI221_X1 U22544 ( .B1(n22527), .B2(n26870), .C1(n21195), .C2(n26864), .A(
        n23152), .ZN(n23149) );
  AOI22_X1 U22545 ( .A1(n26858), .A2(n25920), .B1(n26852), .B2(n8507), .ZN(
        n23152) );
  OAI221_X1 U22546 ( .B1(n22647), .B2(n26747), .C1(n22455), .C2(n26741), .A(
        n23160), .ZN(n23157) );
  AOI22_X1 U22547 ( .A1(n26735), .A2(n26251), .B1(n26729), .B2(n26371), .ZN(
        n23160) );
  OAI221_X1 U22548 ( .B1(n22526), .B2(n26870), .C1(n21194), .C2(n26864), .A(
        n23134), .ZN(n23131) );
  AOI22_X1 U22549 ( .A1(n26858), .A2(n25925), .B1(n26852), .B2(n8504), .ZN(
        n23134) );
  OAI221_X1 U22550 ( .B1(n22646), .B2(n26747), .C1(n22454), .C2(n26741), .A(
        n23142), .ZN(n23139) );
  AOI22_X1 U22551 ( .A1(n26735), .A2(n26252), .B1(n26729), .B2(n26372), .ZN(
        n23142) );
  OAI221_X1 U22552 ( .B1(n22525), .B2(n26870), .C1(n21193), .C2(n26864), .A(
        n23116), .ZN(n23113) );
  AOI22_X1 U22553 ( .A1(n26858), .A2(n25930), .B1(n26852), .B2(n8501), .ZN(
        n23116) );
  OAI221_X1 U22554 ( .B1(n22645), .B2(n26747), .C1(n22453), .C2(n26741), .A(
        n23124), .ZN(n23121) );
  AOI22_X1 U22555 ( .A1(n26735), .A2(n26253), .B1(n26729), .B2(n26373), .ZN(
        n23124) );
  OAI221_X1 U22556 ( .B1(n22524), .B2(n26870), .C1(n21192), .C2(n26864), .A(
        n23098), .ZN(n23095) );
  AOI22_X1 U22557 ( .A1(n26858), .A2(n25935), .B1(n26852), .B2(n8498), .ZN(
        n23098) );
  OAI221_X1 U22558 ( .B1(n22644), .B2(n26747), .C1(n22452), .C2(n26741), .A(
        n23106), .ZN(n23103) );
  AOI22_X1 U22559 ( .A1(n26735), .A2(n26254), .B1(n26729), .B2(n26374), .ZN(
        n23106) );
  OAI221_X1 U22560 ( .B1(n22523), .B2(n26871), .C1(n21191), .C2(n26865), .A(
        n23080), .ZN(n23077) );
  AOI22_X1 U22561 ( .A1(n26859), .A2(n25940), .B1(n26853), .B2(n8495), .ZN(
        n23080) );
  OAI221_X1 U22562 ( .B1(n22643), .B2(n26748), .C1(n22451), .C2(n26742), .A(
        n23088), .ZN(n23085) );
  AOI22_X1 U22563 ( .A1(n26736), .A2(n26255), .B1(n26730), .B2(n26375), .ZN(
        n23088) );
  OAI221_X1 U22564 ( .B1(n22522), .B2(n26871), .C1(n21190), .C2(n26865), .A(
        n23062), .ZN(n23059) );
  AOI22_X1 U22565 ( .A1(n26859), .A2(n25945), .B1(n26853), .B2(n8492), .ZN(
        n23062) );
  OAI221_X1 U22566 ( .B1(n22642), .B2(n26748), .C1(n22450), .C2(n26742), .A(
        n23070), .ZN(n23067) );
  AOI22_X1 U22567 ( .A1(n26736), .A2(n26256), .B1(n26730), .B2(n26376), .ZN(
        n23070) );
  OAI221_X1 U22568 ( .B1(n22521), .B2(n26871), .C1(n21189), .C2(n26865), .A(
        n23044), .ZN(n23041) );
  AOI22_X1 U22569 ( .A1(n26859), .A2(n25950), .B1(n26853), .B2(n8489), .ZN(
        n23044) );
  OAI221_X1 U22570 ( .B1(n22641), .B2(n26748), .C1(n22449), .C2(n26742), .A(
        n23052), .ZN(n23049) );
  AOI22_X1 U22571 ( .A1(n26736), .A2(n26257), .B1(n26730), .B2(n26377), .ZN(
        n23052) );
  OAI221_X1 U22572 ( .B1(n22520), .B2(n26871), .C1(n21188), .C2(n26865), .A(
        n23026), .ZN(n23023) );
  AOI22_X1 U22573 ( .A1(n26859), .A2(n25955), .B1(n26853), .B2(n8486), .ZN(
        n23026) );
  OAI221_X1 U22574 ( .B1(n22640), .B2(n26748), .C1(n22448), .C2(n26742), .A(
        n23034), .ZN(n23031) );
  AOI22_X1 U22575 ( .A1(n26736), .A2(n26258), .B1(n26730), .B2(n26378), .ZN(
        n23034) );
  OAI221_X1 U22576 ( .B1(n22519), .B2(n26871), .C1(n21187), .C2(n26865), .A(
        n23008), .ZN(n23005) );
  AOI22_X1 U22577 ( .A1(n26859), .A2(n25960), .B1(n26853), .B2(n8483), .ZN(
        n23008) );
  OAI221_X1 U22578 ( .B1(n22639), .B2(n26748), .C1(n22447), .C2(n26742), .A(
        n23016), .ZN(n23013) );
  AOI22_X1 U22579 ( .A1(n26736), .A2(n26259), .B1(n26730), .B2(n26379), .ZN(
        n23016) );
  OAI221_X1 U22580 ( .B1(n22518), .B2(n26871), .C1(n21186), .C2(n26865), .A(
        n22990), .ZN(n22987) );
  AOI22_X1 U22581 ( .A1(n26859), .A2(n25965), .B1(n26853), .B2(n8480), .ZN(
        n22990) );
  OAI221_X1 U22582 ( .B1(n22638), .B2(n26748), .C1(n22446), .C2(n26742), .A(
        n22998), .ZN(n22995) );
  AOI22_X1 U22583 ( .A1(n26736), .A2(n26260), .B1(n26730), .B2(n26380), .ZN(
        n22998) );
  OAI221_X1 U22584 ( .B1(n22517), .B2(n26871), .C1(n21185), .C2(n26865), .A(
        n22972), .ZN(n22969) );
  AOI22_X1 U22585 ( .A1(n26859), .A2(n25970), .B1(n26853), .B2(n8477), .ZN(
        n22972) );
  OAI221_X1 U22586 ( .B1(n22637), .B2(n26748), .C1(n22445), .C2(n26742), .A(
        n22980), .ZN(n22977) );
  AOI22_X1 U22587 ( .A1(n26736), .A2(n26261), .B1(n26730), .B2(n26381), .ZN(
        n22980) );
  OAI221_X1 U22588 ( .B1(n22516), .B2(n26871), .C1(n21184), .C2(n26865), .A(
        n22954), .ZN(n22951) );
  AOI22_X1 U22589 ( .A1(n26859), .A2(n25975), .B1(n26853), .B2(n8474), .ZN(
        n22954) );
  OAI221_X1 U22590 ( .B1(n22636), .B2(n26748), .C1(n22444), .C2(n26742), .A(
        n22962), .ZN(n22959) );
  AOI22_X1 U22591 ( .A1(n26736), .A2(n26262), .B1(n26730), .B2(n26382), .ZN(
        n22962) );
  OAI221_X1 U22592 ( .B1(n22515), .B2(n26871), .C1(n21183), .C2(n26865), .A(
        n22936), .ZN(n22933) );
  AOI22_X1 U22593 ( .A1(n26859), .A2(n25980), .B1(n26853), .B2(n8471), .ZN(
        n22936) );
  OAI221_X1 U22594 ( .B1(n22635), .B2(n26748), .C1(n22443), .C2(n26742), .A(
        n22944), .ZN(n22941) );
  AOI22_X1 U22595 ( .A1(n26736), .A2(n26263), .B1(n26730), .B2(n26383), .ZN(
        n22944) );
  OAI221_X1 U22596 ( .B1(n22514), .B2(n26871), .C1(n21182), .C2(n26865), .A(
        n22918), .ZN(n22915) );
  AOI22_X1 U22597 ( .A1(n26859), .A2(n25985), .B1(n26853), .B2(n8468), .ZN(
        n22918) );
  OAI221_X1 U22598 ( .B1(n22634), .B2(n26748), .C1(n22442), .C2(n26742), .A(
        n22926), .ZN(n22923) );
  AOI22_X1 U22599 ( .A1(n26736), .A2(n26264), .B1(n26730), .B2(n26384), .ZN(
        n22926) );
  OAI221_X1 U22600 ( .B1(n22513), .B2(n26871), .C1(n21181), .C2(n26865), .A(
        n22900), .ZN(n22897) );
  AOI22_X1 U22601 ( .A1(n26859), .A2(n25990), .B1(n26853), .B2(n8465), .ZN(
        n22900) );
  OAI221_X1 U22602 ( .B1(n22633), .B2(n26748), .C1(n22441), .C2(n26742), .A(
        n22908), .ZN(n22905) );
  AOI22_X1 U22603 ( .A1(n26736), .A2(n26265), .B1(n26730), .B2(n26385), .ZN(
        n22908) );
  OAI221_X1 U22604 ( .B1(n22512), .B2(n26871), .C1(n21180), .C2(n26865), .A(
        n22882), .ZN(n22879) );
  AOI22_X1 U22605 ( .A1(n26859), .A2(n25995), .B1(n26853), .B2(n8462), .ZN(
        n22882) );
  OAI221_X1 U22606 ( .B1(n22632), .B2(n26748), .C1(n22440), .C2(n26742), .A(
        n22890), .ZN(n22887) );
  AOI22_X1 U22607 ( .A1(n26736), .A2(n26266), .B1(n26730), .B2(n26386), .ZN(
        n22890) );
  OAI221_X1 U22608 ( .B1(n22500), .B2(n26647), .C1(n21156), .C2(n26641), .A(
        n23981), .ZN(n23972) );
  AOI22_X1 U22609 ( .A1(n26635), .A2(n25695), .B1(n26629), .B2(n8450), .ZN(
        n23981) );
  OAI221_X1 U22610 ( .B1(n22508), .B2(n26524), .C1(n22256), .C2(n26518), .A(
        n24006), .ZN(n23997) );
  AOI22_X1 U22611 ( .A1(n26512), .A2(n26194), .B1(n26506), .B2(n26198), .ZN(
        n24006) );
  OAI221_X1 U22612 ( .B1(n22503), .B2(n26647), .C1(n21159), .C2(n26641), .A(
        n24063), .ZN(n24060) );
  AOI22_X1 U22613 ( .A1(n26635), .A2(n25680), .B1(n26629), .B2(n8459), .ZN(
        n24063) );
  OAI221_X1 U22614 ( .B1(n22511), .B2(n26524), .C1(n22259), .C2(n26518), .A(
        n24071), .ZN(n24068) );
  AOI22_X1 U22615 ( .A1(n26512), .A2(n26191), .B1(n26506), .B2(n26195), .ZN(
        n24071) );
  OAI221_X1 U22616 ( .B1(n22502), .B2(n26647), .C1(n21158), .C2(n26641), .A(
        n24045), .ZN(n24042) );
  AOI22_X1 U22617 ( .A1(n26635), .A2(n25685), .B1(n26629), .B2(n8456), .ZN(
        n24045) );
  OAI221_X1 U22618 ( .B1(n22510), .B2(n26524), .C1(n22258), .C2(n26518), .A(
        n24053), .ZN(n24050) );
  AOI22_X1 U22619 ( .A1(n26512), .A2(n26192), .B1(n26506), .B2(n26196), .ZN(
        n24053) );
  OAI221_X1 U22620 ( .B1(n22501), .B2(n26647), .C1(n21157), .C2(n26641), .A(
        n24027), .ZN(n24024) );
  AOI22_X1 U22621 ( .A1(n26635), .A2(n25690), .B1(n26629), .B2(n8453), .ZN(
        n24027) );
  OAI221_X1 U22622 ( .B1(n22509), .B2(n26524), .C1(n22257), .C2(n26518), .A(
        n24035), .ZN(n24032) );
  AOI22_X1 U22623 ( .A1(n26512), .A2(n26193), .B1(n26506), .B2(n26197), .ZN(
        n24035) );
  OAI221_X1 U22624 ( .B1(n22503), .B2(n26872), .C1(n21159), .C2(n26866), .A(
        n22864), .ZN(n22861) );
  AOI22_X1 U22625 ( .A1(n26860), .A2(n25680), .B1(n26854), .B2(n8459), .ZN(
        n22864) );
  OAI221_X1 U22626 ( .B1(n22511), .B2(n26749), .C1(n22259), .C2(n26743), .A(
        n22872), .ZN(n22869) );
  AOI22_X1 U22627 ( .A1(n26737), .A2(n26191), .B1(n26731), .B2(n26195), .ZN(
        n22872) );
  OAI221_X1 U22628 ( .B1(n22502), .B2(n26872), .C1(n21158), .C2(n26866), .A(
        n22846), .ZN(n22843) );
  AOI22_X1 U22629 ( .A1(n26860), .A2(n25685), .B1(n26854), .B2(n8456), .ZN(
        n22846) );
  OAI221_X1 U22630 ( .B1(n22510), .B2(n26749), .C1(n22258), .C2(n26743), .A(
        n22854), .ZN(n22851) );
  AOI22_X1 U22631 ( .A1(n26737), .A2(n26192), .B1(n26731), .B2(n26196), .ZN(
        n22854) );
  OAI221_X1 U22632 ( .B1(n22501), .B2(n26872), .C1(n21157), .C2(n26866), .A(
        n22828), .ZN(n22825) );
  AOI22_X1 U22633 ( .A1(n26860), .A2(n25690), .B1(n26854), .B2(n8453), .ZN(
        n22828) );
  OAI221_X1 U22634 ( .B1(n22509), .B2(n26749), .C1(n22257), .C2(n26743), .A(
        n22836), .ZN(n22833) );
  AOI22_X1 U22635 ( .A1(n26737), .A2(n26193), .B1(n26731), .B2(n26197), .ZN(
        n22836) );
  OAI221_X1 U22636 ( .B1(n22500), .B2(n26872), .C1(n21156), .C2(n26866), .A(
        n22782), .ZN(n22773) );
  AOI22_X1 U22637 ( .A1(n26860), .A2(n25695), .B1(n26854), .B2(n8450), .ZN(
        n22782) );
  OAI221_X1 U22638 ( .B1(n22508), .B2(n26749), .C1(n22256), .C2(n26743), .A(
        n22807), .ZN(n22798) );
  AOI22_X1 U22639 ( .A1(n26737), .A2(n26194), .B1(n26731), .B2(n26198), .ZN(
        n22807) );
  OAI221_X1 U22640 ( .B1(n22571), .B2(n26642), .C1(n21239), .C2(n26636), .A(
        n25149), .ZN(n25140) );
  AOI22_X1 U22641 ( .A1(n26630), .A2(n25700), .B1(n26624), .B2(n8639), .ZN(
        n25149) );
  OAI221_X1 U22642 ( .B1(n22691), .B2(n26519), .C1(n22499), .C2(n26513), .A(
        n25161), .ZN(n25158) );
  AOI22_X1 U22643 ( .A1(n26507), .A2(n26207), .B1(n26501), .B2(n26327), .ZN(
        n25161) );
  OAI221_X1 U22644 ( .B1(n22570), .B2(n26642), .C1(n21238), .C2(n26636), .A(
        n25125), .ZN(n25122) );
  AOI22_X1 U22645 ( .A1(n26630), .A2(n25705), .B1(n26624), .B2(n8636), .ZN(
        n25125) );
  OAI221_X1 U22646 ( .B1(n22690), .B2(n26519), .C1(n22498), .C2(n26513), .A(
        n25133), .ZN(n25130) );
  AOI22_X1 U22647 ( .A1(n26507), .A2(n26208), .B1(n26501), .B2(n26328), .ZN(
        n25133) );
  OAI221_X1 U22648 ( .B1(n22569), .B2(n26642), .C1(n21237), .C2(n26636), .A(
        n25107), .ZN(n25104) );
  AOI22_X1 U22649 ( .A1(n26630), .A2(n25710), .B1(n26624), .B2(n8633), .ZN(
        n25107) );
  OAI221_X1 U22650 ( .B1(n22689), .B2(n26519), .C1(n22497), .C2(n26513), .A(
        n25115), .ZN(n25112) );
  AOI22_X1 U22651 ( .A1(n26507), .A2(n26209), .B1(n26501), .B2(n26329), .ZN(
        n25115) );
  OAI221_X1 U22652 ( .B1(n22568), .B2(n26642), .C1(n21236), .C2(n26636), .A(
        n25089), .ZN(n25086) );
  AOI22_X1 U22653 ( .A1(n26630), .A2(n25715), .B1(n26624), .B2(n8630), .ZN(
        n25089) );
  OAI221_X1 U22654 ( .B1(n22688), .B2(n26519), .C1(n22496), .C2(n26513), .A(
        n25097), .ZN(n25094) );
  AOI22_X1 U22655 ( .A1(n26507), .A2(n26210), .B1(n26501), .B2(n26330), .ZN(
        n25097) );
  OAI221_X1 U22656 ( .B1(n22567), .B2(n26642), .C1(n21235), .C2(n26636), .A(
        n25071), .ZN(n25068) );
  AOI22_X1 U22657 ( .A1(n26630), .A2(n25720), .B1(n26624), .B2(n8627), .ZN(
        n25071) );
  OAI221_X1 U22658 ( .B1(n22687), .B2(n26519), .C1(n22495), .C2(n26513), .A(
        n25079), .ZN(n25076) );
  AOI22_X1 U22659 ( .A1(n26507), .A2(n26211), .B1(n26501), .B2(n26331), .ZN(
        n25079) );
  OAI221_X1 U22660 ( .B1(n22566), .B2(n26642), .C1(n21234), .C2(n26636), .A(
        n25053), .ZN(n25050) );
  AOI22_X1 U22661 ( .A1(n26630), .A2(n25725), .B1(n26624), .B2(n8624), .ZN(
        n25053) );
  OAI221_X1 U22662 ( .B1(n22686), .B2(n26519), .C1(n22494), .C2(n26513), .A(
        n25061), .ZN(n25058) );
  AOI22_X1 U22663 ( .A1(n26507), .A2(n26212), .B1(n26501), .B2(n26332), .ZN(
        n25061) );
  OAI221_X1 U22664 ( .B1(n22565), .B2(n26642), .C1(n21233), .C2(n26636), .A(
        n25035), .ZN(n25032) );
  AOI22_X1 U22665 ( .A1(n26630), .A2(n25730), .B1(n26624), .B2(n8621), .ZN(
        n25035) );
  OAI221_X1 U22666 ( .B1(n22685), .B2(n26519), .C1(n22493), .C2(n26513), .A(
        n25043), .ZN(n25040) );
  AOI22_X1 U22667 ( .A1(n26507), .A2(n26213), .B1(n26501), .B2(n26333), .ZN(
        n25043) );
  OAI221_X1 U22668 ( .B1(n22564), .B2(n26642), .C1(n21232), .C2(n26636), .A(
        n25017), .ZN(n25014) );
  AOI22_X1 U22669 ( .A1(n26630), .A2(n25735), .B1(n26624), .B2(n8618), .ZN(
        n25017) );
  OAI221_X1 U22670 ( .B1(n22684), .B2(n26519), .C1(n22492), .C2(n26513), .A(
        n25025), .ZN(n25022) );
  AOI22_X1 U22671 ( .A1(n26507), .A2(n26214), .B1(n26501), .B2(n26334), .ZN(
        n25025) );
  OAI221_X1 U22672 ( .B1(n22563), .B2(n26642), .C1(n21231), .C2(n26636), .A(
        n24999), .ZN(n24996) );
  AOI22_X1 U22673 ( .A1(n26630), .A2(n25740), .B1(n26624), .B2(n8615), .ZN(
        n24999) );
  OAI221_X1 U22674 ( .B1(n22683), .B2(n26519), .C1(n22491), .C2(n26513), .A(
        n25007), .ZN(n25004) );
  AOI22_X1 U22675 ( .A1(n26507), .A2(n26215), .B1(n26501), .B2(n26335), .ZN(
        n25007) );
  OAI221_X1 U22676 ( .B1(n22562), .B2(n26642), .C1(n21230), .C2(n26636), .A(
        n24981), .ZN(n24978) );
  AOI22_X1 U22677 ( .A1(n26630), .A2(n25745), .B1(n26624), .B2(n8612), .ZN(
        n24981) );
  OAI221_X1 U22678 ( .B1(n22682), .B2(n26519), .C1(n22490), .C2(n26513), .A(
        n24989), .ZN(n24986) );
  AOI22_X1 U22679 ( .A1(n26507), .A2(n26216), .B1(n26501), .B2(n26336), .ZN(
        n24989) );
  OAI221_X1 U22680 ( .B1(n22561), .B2(n26642), .C1(n21229), .C2(n26636), .A(
        n24963), .ZN(n24960) );
  AOI22_X1 U22681 ( .A1(n26630), .A2(n25750), .B1(n26624), .B2(n8609), .ZN(
        n24963) );
  OAI221_X1 U22682 ( .B1(n22681), .B2(n26519), .C1(n22489), .C2(n26513), .A(
        n24971), .ZN(n24968) );
  AOI22_X1 U22683 ( .A1(n26507), .A2(n26217), .B1(n26501), .B2(n26337), .ZN(
        n24971) );
  OAI221_X1 U22684 ( .B1(n22560), .B2(n26642), .C1(n21228), .C2(n26636), .A(
        n24945), .ZN(n24942) );
  AOI22_X1 U22685 ( .A1(n26630), .A2(n25755), .B1(n26624), .B2(n8606), .ZN(
        n24945) );
  OAI221_X1 U22686 ( .B1(n22680), .B2(n26519), .C1(n22488), .C2(n26513), .A(
        n24953), .ZN(n24950) );
  AOI22_X1 U22687 ( .A1(n26507), .A2(n26218), .B1(n26501), .B2(n26338), .ZN(
        n24953) );
  OAI221_X1 U22688 ( .B1(n22571), .B2(n26867), .C1(n21239), .C2(n26861), .A(
        n23950), .ZN(n23941) );
  AOI22_X1 U22689 ( .A1(n26855), .A2(n25700), .B1(n26849), .B2(n8639), .ZN(
        n23950) );
  OAI221_X1 U22690 ( .B1(n22691), .B2(n26744), .C1(n22499), .C2(n26738), .A(
        n23962), .ZN(n23959) );
  AOI22_X1 U22691 ( .A1(n26732), .A2(n26207), .B1(n26726), .B2(n26327), .ZN(
        n23962) );
  OAI221_X1 U22692 ( .B1(n22570), .B2(n26867), .C1(n21238), .C2(n26861), .A(
        n23926), .ZN(n23923) );
  AOI22_X1 U22693 ( .A1(n26855), .A2(n25705), .B1(n26849), .B2(n8636), .ZN(
        n23926) );
  OAI221_X1 U22694 ( .B1(n22690), .B2(n26744), .C1(n22498), .C2(n26738), .A(
        n23934), .ZN(n23931) );
  AOI22_X1 U22695 ( .A1(n26732), .A2(n26208), .B1(n26726), .B2(n26328), .ZN(
        n23934) );
  OAI221_X1 U22696 ( .B1(n22569), .B2(n26867), .C1(n21237), .C2(n26861), .A(
        n23908), .ZN(n23905) );
  AOI22_X1 U22697 ( .A1(n26855), .A2(n25710), .B1(n26849), .B2(n8633), .ZN(
        n23908) );
  OAI221_X1 U22698 ( .B1(n22689), .B2(n26744), .C1(n22497), .C2(n26738), .A(
        n23916), .ZN(n23913) );
  AOI22_X1 U22699 ( .A1(n26732), .A2(n26209), .B1(n26726), .B2(n26329), .ZN(
        n23916) );
  OAI221_X1 U22700 ( .B1(n22568), .B2(n26867), .C1(n21236), .C2(n26861), .A(
        n23890), .ZN(n23887) );
  AOI22_X1 U22701 ( .A1(n26855), .A2(n25715), .B1(n26849), .B2(n8630), .ZN(
        n23890) );
  OAI221_X1 U22702 ( .B1(n22688), .B2(n26744), .C1(n22496), .C2(n26738), .A(
        n23898), .ZN(n23895) );
  AOI22_X1 U22703 ( .A1(n26732), .A2(n26210), .B1(n26726), .B2(n26330), .ZN(
        n23898) );
  OAI221_X1 U22704 ( .B1(n22567), .B2(n26867), .C1(n21235), .C2(n26861), .A(
        n23872), .ZN(n23869) );
  AOI22_X1 U22705 ( .A1(n26855), .A2(n25720), .B1(n26849), .B2(n8627), .ZN(
        n23872) );
  OAI221_X1 U22706 ( .B1(n22687), .B2(n26744), .C1(n22495), .C2(n26738), .A(
        n23880), .ZN(n23877) );
  AOI22_X1 U22707 ( .A1(n26732), .A2(n26211), .B1(n26726), .B2(n26331), .ZN(
        n23880) );
  OAI221_X1 U22708 ( .B1(n22566), .B2(n26867), .C1(n21234), .C2(n26861), .A(
        n23854), .ZN(n23851) );
  AOI22_X1 U22709 ( .A1(n26855), .A2(n25725), .B1(n26849), .B2(n8624), .ZN(
        n23854) );
  OAI221_X1 U22710 ( .B1(n22686), .B2(n26744), .C1(n22494), .C2(n26738), .A(
        n23862), .ZN(n23859) );
  AOI22_X1 U22711 ( .A1(n26732), .A2(n26212), .B1(n26726), .B2(n26332), .ZN(
        n23862) );
  OAI221_X1 U22712 ( .B1(n22565), .B2(n26867), .C1(n21233), .C2(n26861), .A(
        n23836), .ZN(n23833) );
  AOI22_X1 U22713 ( .A1(n26855), .A2(n25730), .B1(n26849), .B2(n8621), .ZN(
        n23836) );
  OAI221_X1 U22714 ( .B1(n22685), .B2(n26744), .C1(n22493), .C2(n26738), .A(
        n23844), .ZN(n23841) );
  AOI22_X1 U22715 ( .A1(n26732), .A2(n26213), .B1(n26726), .B2(n26333), .ZN(
        n23844) );
  OAI221_X1 U22716 ( .B1(n22564), .B2(n26867), .C1(n21232), .C2(n26861), .A(
        n23818), .ZN(n23815) );
  AOI22_X1 U22717 ( .A1(n26855), .A2(n25735), .B1(n26849), .B2(n8618), .ZN(
        n23818) );
  OAI221_X1 U22718 ( .B1(n22684), .B2(n26744), .C1(n22492), .C2(n26738), .A(
        n23826), .ZN(n23823) );
  AOI22_X1 U22719 ( .A1(n26732), .A2(n26214), .B1(n26726), .B2(n26334), .ZN(
        n23826) );
  OAI221_X1 U22720 ( .B1(n22563), .B2(n26867), .C1(n21231), .C2(n26861), .A(
        n23800), .ZN(n23797) );
  AOI22_X1 U22721 ( .A1(n26855), .A2(n25740), .B1(n26849), .B2(n8615), .ZN(
        n23800) );
  OAI221_X1 U22722 ( .B1(n22683), .B2(n26744), .C1(n22491), .C2(n26738), .A(
        n23808), .ZN(n23805) );
  AOI22_X1 U22723 ( .A1(n26732), .A2(n26215), .B1(n26726), .B2(n26335), .ZN(
        n23808) );
  OAI221_X1 U22724 ( .B1(n22562), .B2(n26867), .C1(n21230), .C2(n26861), .A(
        n23782), .ZN(n23779) );
  AOI22_X1 U22725 ( .A1(n26855), .A2(n25745), .B1(n26849), .B2(n8612), .ZN(
        n23782) );
  OAI221_X1 U22726 ( .B1(n22682), .B2(n26744), .C1(n22490), .C2(n26738), .A(
        n23790), .ZN(n23787) );
  AOI22_X1 U22727 ( .A1(n26732), .A2(n26216), .B1(n26726), .B2(n26336), .ZN(
        n23790) );
  OAI221_X1 U22728 ( .B1(n22561), .B2(n26867), .C1(n21229), .C2(n26861), .A(
        n23764), .ZN(n23761) );
  AOI22_X1 U22729 ( .A1(n26855), .A2(n25750), .B1(n26849), .B2(n8609), .ZN(
        n23764) );
  OAI221_X1 U22730 ( .B1(n22681), .B2(n26744), .C1(n22489), .C2(n26738), .A(
        n23772), .ZN(n23769) );
  AOI22_X1 U22731 ( .A1(n26732), .A2(n26217), .B1(n26726), .B2(n26337), .ZN(
        n23772) );
  OAI221_X1 U22732 ( .B1(n22560), .B2(n26867), .C1(n21228), .C2(n26861), .A(
        n23746), .ZN(n23743) );
  AOI22_X1 U22733 ( .A1(n26855), .A2(n25755), .B1(n26849), .B2(n8606), .ZN(
        n23746) );
  OAI221_X1 U22734 ( .B1(n22680), .B2(n26744), .C1(n22488), .C2(n26738), .A(
        n23754), .ZN(n23751) );
  AOI22_X1 U22735 ( .A1(n26732), .A2(n26218), .B1(n26726), .B2(n26338), .ZN(
        n23754) );
  OAI221_X1 U22736 ( .B1(n9620), .B2(n26619), .C1(n20822), .C2(n26613), .A(
        n24928), .ZN(n24923) );
  AOI22_X1 U22737 ( .A1(n26607), .A2(n25761), .B1(n26601), .B2(n21022), .ZN(
        n24928) );
  OAI221_X1 U22738 ( .B1(n9619), .B2(n26619), .C1(n20821), .C2(n26613), .A(
        n24910), .ZN(n24905) );
  AOI22_X1 U22739 ( .A1(n26607), .A2(n25766), .B1(n26601), .B2(n21021), .ZN(
        n24910) );
  OAI221_X1 U22740 ( .B1(n9618), .B2(n26619), .C1(n20820), .C2(n26613), .A(
        n24892), .ZN(n24887) );
  AOI22_X1 U22741 ( .A1(n26607), .A2(n25771), .B1(n26601), .B2(n21020), .ZN(
        n24892) );
  OAI221_X1 U22742 ( .B1(n9617), .B2(n26619), .C1(n20819), .C2(n26613), .A(
        n24874), .ZN(n24869) );
  AOI22_X1 U22743 ( .A1(n26607), .A2(n25776), .B1(n26601), .B2(n21019), .ZN(
        n24874) );
  OAI221_X1 U22744 ( .B1(n9616), .B2(n26619), .C1(n20818), .C2(n26613), .A(
        n24856), .ZN(n24851) );
  AOI22_X1 U22745 ( .A1(n26607), .A2(n25781), .B1(n26601), .B2(n21018), .ZN(
        n24856) );
  OAI221_X1 U22746 ( .B1(n9615), .B2(n26619), .C1(n20817), .C2(n26613), .A(
        n24838), .ZN(n24833) );
  AOI22_X1 U22747 ( .A1(n26607), .A2(n25786), .B1(n26601), .B2(n21017), .ZN(
        n24838) );
  OAI221_X1 U22748 ( .B1(n9614), .B2(n26619), .C1(n20816), .C2(n26613), .A(
        n24820), .ZN(n24815) );
  AOI22_X1 U22749 ( .A1(n26607), .A2(n25791), .B1(n26601), .B2(n21016), .ZN(
        n24820) );
  OAI221_X1 U22750 ( .B1(n9613), .B2(n26619), .C1(n20815), .C2(n26613), .A(
        n24802), .ZN(n24797) );
  AOI22_X1 U22751 ( .A1(n26607), .A2(n25796), .B1(n26601), .B2(n21015), .ZN(
        n24802) );
  OAI221_X1 U22752 ( .B1(n9612), .B2(n26619), .C1(n20814), .C2(n26613), .A(
        n24784), .ZN(n24779) );
  AOI22_X1 U22753 ( .A1(n26607), .A2(n25801), .B1(n26601), .B2(n21014), .ZN(
        n24784) );
  OAI221_X1 U22754 ( .B1(n9611), .B2(n26619), .C1(n20813), .C2(n26613), .A(
        n24766), .ZN(n24761) );
  AOI22_X1 U22755 ( .A1(n26607), .A2(n25806), .B1(n26601), .B2(n21013), .ZN(
        n24766) );
  OAI221_X1 U22756 ( .B1(n9610), .B2(n26619), .C1(n20812), .C2(n26613), .A(
        n24748), .ZN(n24743) );
  AOI22_X1 U22757 ( .A1(n26607), .A2(n25811), .B1(n26601), .B2(n21012), .ZN(
        n24748) );
  OAI221_X1 U22758 ( .B1(n9609), .B2(n26619), .C1(n20811), .C2(n26613), .A(
        n24730), .ZN(n24725) );
  AOI22_X1 U22759 ( .A1(n26607), .A2(n25816), .B1(n26601), .B2(n21011), .ZN(
        n24730) );
  OAI221_X1 U22760 ( .B1(n9608), .B2(n26620), .C1(n20810), .C2(n26614), .A(
        n24712), .ZN(n24707) );
  AOI22_X1 U22761 ( .A1(n26608), .A2(n25821), .B1(n26602), .B2(n21010), .ZN(
        n24712) );
  OAI221_X1 U22762 ( .B1(n9607), .B2(n26620), .C1(n20809), .C2(n26614), .A(
        n24694), .ZN(n24689) );
  AOI22_X1 U22763 ( .A1(n26608), .A2(n25826), .B1(n26602), .B2(n21009), .ZN(
        n24694) );
  OAI221_X1 U22764 ( .B1(n9606), .B2(n26620), .C1(n20808), .C2(n26614), .A(
        n24676), .ZN(n24671) );
  AOI22_X1 U22765 ( .A1(n26608), .A2(n25831), .B1(n26602), .B2(n21008), .ZN(
        n24676) );
  OAI221_X1 U22766 ( .B1(n9605), .B2(n26620), .C1(n20807), .C2(n26614), .A(
        n24658), .ZN(n24653) );
  AOI22_X1 U22767 ( .A1(n26608), .A2(n25836), .B1(n26602), .B2(n21007), .ZN(
        n24658) );
  OAI221_X1 U22768 ( .B1(n9604), .B2(n26620), .C1(n20806), .C2(n26614), .A(
        n24640), .ZN(n24635) );
  AOI22_X1 U22769 ( .A1(n26608), .A2(n25841), .B1(n26602), .B2(n21006), .ZN(
        n24640) );
  OAI221_X1 U22770 ( .B1(n9603), .B2(n26620), .C1(n20805), .C2(n26614), .A(
        n24622), .ZN(n24617) );
  AOI22_X1 U22771 ( .A1(n26608), .A2(n25846), .B1(n26602), .B2(n21005), .ZN(
        n24622) );
  OAI221_X1 U22772 ( .B1(n9602), .B2(n26620), .C1(n20804), .C2(n26614), .A(
        n24604), .ZN(n24599) );
  AOI22_X1 U22773 ( .A1(n26608), .A2(n25851), .B1(n26602), .B2(n21004), .ZN(
        n24604) );
  OAI221_X1 U22774 ( .B1(n9601), .B2(n26620), .C1(n20803), .C2(n26614), .A(
        n24586), .ZN(n24581) );
  AOI22_X1 U22775 ( .A1(n26608), .A2(n25856), .B1(n26602), .B2(n21003), .ZN(
        n24586) );
  OAI221_X1 U22776 ( .B1(n9600), .B2(n26620), .C1(n20802), .C2(n26614), .A(
        n24568), .ZN(n24563) );
  AOI22_X1 U22777 ( .A1(n26608), .A2(n25861), .B1(n26602), .B2(n21002), .ZN(
        n24568) );
  OAI221_X1 U22778 ( .B1(n9599), .B2(n26620), .C1(n20801), .C2(n26614), .A(
        n24550), .ZN(n24545) );
  AOI22_X1 U22779 ( .A1(n26608), .A2(n25866), .B1(n26602), .B2(n21001), .ZN(
        n24550) );
  OAI221_X1 U22780 ( .B1(n9598), .B2(n26620), .C1(n20800), .C2(n26614), .A(
        n24532), .ZN(n24527) );
  AOI22_X1 U22781 ( .A1(n26608), .A2(n25871), .B1(n26602), .B2(n21000), .ZN(
        n24532) );
  OAI221_X1 U22782 ( .B1(n9597), .B2(n26620), .C1(n20799), .C2(n26614), .A(
        n24514), .ZN(n24509) );
  AOI22_X1 U22783 ( .A1(n26608), .A2(n25876), .B1(n26602), .B2(n20999), .ZN(
        n24514) );
  OAI221_X1 U22784 ( .B1(n9596), .B2(n26621), .C1(n20798), .C2(n26615), .A(
        n24496), .ZN(n24491) );
  AOI22_X1 U22785 ( .A1(n26609), .A2(n25881), .B1(n26603), .B2(n20998), .ZN(
        n24496) );
  OAI221_X1 U22786 ( .B1(n9595), .B2(n26621), .C1(n20797), .C2(n26615), .A(
        n24478), .ZN(n24473) );
  AOI22_X1 U22787 ( .A1(n26609), .A2(n25886), .B1(n26603), .B2(n20997), .ZN(
        n24478) );
  OAI221_X1 U22788 ( .B1(n9594), .B2(n26621), .C1(n20796), .C2(n26615), .A(
        n24460), .ZN(n24455) );
  AOI22_X1 U22789 ( .A1(n26609), .A2(n25891), .B1(n26603), .B2(n20996), .ZN(
        n24460) );
  OAI221_X1 U22790 ( .B1(n9593), .B2(n26621), .C1(n20795), .C2(n26615), .A(
        n24442), .ZN(n24437) );
  AOI22_X1 U22791 ( .A1(n26609), .A2(n25896), .B1(n26603), .B2(n20995), .ZN(
        n24442) );
  OAI221_X1 U22792 ( .B1(n9592), .B2(n26621), .C1(n20794), .C2(n26615), .A(
        n24424), .ZN(n24419) );
  AOI22_X1 U22793 ( .A1(n26609), .A2(n25901), .B1(n26603), .B2(n20994), .ZN(
        n24424) );
  OAI221_X1 U22794 ( .B1(n9591), .B2(n26621), .C1(n20793), .C2(n26615), .A(
        n24406), .ZN(n24401) );
  AOI22_X1 U22795 ( .A1(n26609), .A2(n25906), .B1(n26603), .B2(n20993), .ZN(
        n24406) );
  OAI221_X1 U22796 ( .B1(n9590), .B2(n26621), .C1(n20792), .C2(n26615), .A(
        n24388), .ZN(n24383) );
  AOI22_X1 U22797 ( .A1(n26609), .A2(n25911), .B1(n26603), .B2(n20992), .ZN(
        n24388) );
  OAI221_X1 U22798 ( .B1(n9589), .B2(n26621), .C1(n20791), .C2(n26615), .A(
        n24370), .ZN(n24365) );
  AOI22_X1 U22799 ( .A1(n26609), .A2(n25916), .B1(n26603), .B2(n20991), .ZN(
        n24370) );
  OAI221_X1 U22800 ( .B1(n9588), .B2(n26621), .C1(n20790), .C2(n26615), .A(
        n24352), .ZN(n24347) );
  AOI22_X1 U22801 ( .A1(n26609), .A2(n25921), .B1(n26603), .B2(n20990), .ZN(
        n24352) );
  OAI221_X1 U22802 ( .B1(n9587), .B2(n26621), .C1(n20789), .C2(n26615), .A(
        n24334), .ZN(n24329) );
  AOI22_X1 U22803 ( .A1(n26609), .A2(n25926), .B1(n26603), .B2(n20989), .ZN(
        n24334) );
  OAI221_X1 U22804 ( .B1(n9586), .B2(n26621), .C1(n20788), .C2(n26615), .A(
        n24316), .ZN(n24311) );
  AOI22_X1 U22805 ( .A1(n26609), .A2(n25931), .B1(n26603), .B2(n20988), .ZN(
        n24316) );
  OAI221_X1 U22806 ( .B1(n9585), .B2(n26621), .C1(n20787), .C2(n26615), .A(
        n24298), .ZN(n24293) );
  AOI22_X1 U22807 ( .A1(n26609), .A2(n25936), .B1(n26603), .B2(n20987), .ZN(
        n24298) );
  OAI221_X1 U22808 ( .B1(n9620), .B2(n26844), .C1(n20822), .C2(n26838), .A(
        n23729), .ZN(n23724) );
  AOI22_X1 U22809 ( .A1(n26832), .A2(n25761), .B1(n26826), .B2(n21022), .ZN(
        n23729) );
  OAI221_X1 U22810 ( .B1(n9619), .B2(n26844), .C1(n20821), .C2(n26838), .A(
        n23711), .ZN(n23706) );
  AOI22_X1 U22811 ( .A1(n26832), .A2(n25766), .B1(n26826), .B2(n21021), .ZN(
        n23711) );
  OAI221_X1 U22812 ( .B1(n9618), .B2(n26844), .C1(n20820), .C2(n26838), .A(
        n23693), .ZN(n23688) );
  AOI22_X1 U22813 ( .A1(n26832), .A2(n25771), .B1(n26826), .B2(n21020), .ZN(
        n23693) );
  OAI221_X1 U22814 ( .B1(n9617), .B2(n26844), .C1(n20819), .C2(n26838), .A(
        n23675), .ZN(n23670) );
  AOI22_X1 U22815 ( .A1(n26832), .A2(n25776), .B1(n26826), .B2(n21019), .ZN(
        n23675) );
  OAI221_X1 U22816 ( .B1(n9616), .B2(n26844), .C1(n20818), .C2(n26838), .A(
        n23657), .ZN(n23652) );
  AOI22_X1 U22817 ( .A1(n26832), .A2(n25781), .B1(n26826), .B2(n21018), .ZN(
        n23657) );
  OAI221_X1 U22818 ( .B1(n9615), .B2(n26844), .C1(n20817), .C2(n26838), .A(
        n23639), .ZN(n23634) );
  AOI22_X1 U22819 ( .A1(n26832), .A2(n25786), .B1(n26826), .B2(n21017), .ZN(
        n23639) );
  OAI221_X1 U22820 ( .B1(n9614), .B2(n26844), .C1(n20816), .C2(n26838), .A(
        n23621), .ZN(n23616) );
  AOI22_X1 U22821 ( .A1(n26832), .A2(n25791), .B1(n26826), .B2(n21016), .ZN(
        n23621) );
  OAI221_X1 U22822 ( .B1(n9613), .B2(n26844), .C1(n20815), .C2(n26838), .A(
        n23603), .ZN(n23598) );
  AOI22_X1 U22823 ( .A1(n26832), .A2(n25796), .B1(n26826), .B2(n21015), .ZN(
        n23603) );
  OAI221_X1 U22824 ( .B1(n9612), .B2(n26844), .C1(n20814), .C2(n26838), .A(
        n23585), .ZN(n23580) );
  AOI22_X1 U22825 ( .A1(n26832), .A2(n25801), .B1(n26826), .B2(n21014), .ZN(
        n23585) );
  OAI221_X1 U22826 ( .B1(n9611), .B2(n26844), .C1(n20813), .C2(n26838), .A(
        n23567), .ZN(n23562) );
  AOI22_X1 U22827 ( .A1(n26832), .A2(n25806), .B1(n26826), .B2(n21013), .ZN(
        n23567) );
  OAI221_X1 U22828 ( .B1(n9610), .B2(n26844), .C1(n20812), .C2(n26838), .A(
        n23549), .ZN(n23544) );
  AOI22_X1 U22829 ( .A1(n26832), .A2(n25811), .B1(n26826), .B2(n21012), .ZN(
        n23549) );
  OAI221_X1 U22830 ( .B1(n9609), .B2(n26844), .C1(n20811), .C2(n26838), .A(
        n23531), .ZN(n23526) );
  AOI22_X1 U22831 ( .A1(n26832), .A2(n25816), .B1(n26826), .B2(n21011), .ZN(
        n23531) );
  OAI221_X1 U22832 ( .B1(n9608), .B2(n26845), .C1(n20810), .C2(n26839), .A(
        n23513), .ZN(n23508) );
  AOI22_X1 U22833 ( .A1(n26833), .A2(n25821), .B1(n26827), .B2(n21010), .ZN(
        n23513) );
  OAI221_X1 U22834 ( .B1(n9607), .B2(n26845), .C1(n20809), .C2(n26839), .A(
        n23495), .ZN(n23490) );
  AOI22_X1 U22835 ( .A1(n26833), .A2(n25826), .B1(n26827), .B2(n21009), .ZN(
        n23495) );
  OAI221_X1 U22836 ( .B1(n9606), .B2(n26845), .C1(n20808), .C2(n26839), .A(
        n23477), .ZN(n23472) );
  AOI22_X1 U22837 ( .A1(n26833), .A2(n25831), .B1(n26827), .B2(n21008), .ZN(
        n23477) );
  OAI221_X1 U22838 ( .B1(n9605), .B2(n26845), .C1(n20807), .C2(n26839), .A(
        n23459), .ZN(n23454) );
  AOI22_X1 U22839 ( .A1(n26833), .A2(n25836), .B1(n26827), .B2(n21007), .ZN(
        n23459) );
  OAI221_X1 U22840 ( .B1(n9604), .B2(n26845), .C1(n20806), .C2(n26839), .A(
        n23441), .ZN(n23436) );
  AOI22_X1 U22841 ( .A1(n26833), .A2(n25841), .B1(n26827), .B2(n21006), .ZN(
        n23441) );
  OAI221_X1 U22842 ( .B1(n9603), .B2(n26845), .C1(n20805), .C2(n26839), .A(
        n23423), .ZN(n23418) );
  AOI22_X1 U22843 ( .A1(n26833), .A2(n25846), .B1(n26827), .B2(n21005), .ZN(
        n23423) );
  OAI221_X1 U22844 ( .B1(n9602), .B2(n26845), .C1(n20804), .C2(n26839), .A(
        n23405), .ZN(n23400) );
  AOI22_X1 U22845 ( .A1(n26833), .A2(n25851), .B1(n26827), .B2(n21004), .ZN(
        n23405) );
  OAI221_X1 U22846 ( .B1(n9601), .B2(n26845), .C1(n20803), .C2(n26839), .A(
        n23387), .ZN(n23382) );
  AOI22_X1 U22847 ( .A1(n26833), .A2(n25856), .B1(n26827), .B2(n21003), .ZN(
        n23387) );
  OAI221_X1 U22848 ( .B1(n9600), .B2(n26845), .C1(n20802), .C2(n26839), .A(
        n23369), .ZN(n23364) );
  AOI22_X1 U22849 ( .A1(n26833), .A2(n25861), .B1(n26827), .B2(n21002), .ZN(
        n23369) );
  OAI221_X1 U22850 ( .B1(n9599), .B2(n26845), .C1(n20801), .C2(n26839), .A(
        n23351), .ZN(n23346) );
  AOI22_X1 U22851 ( .A1(n26833), .A2(n25866), .B1(n26827), .B2(n21001), .ZN(
        n23351) );
  OAI221_X1 U22852 ( .B1(n9598), .B2(n26845), .C1(n20800), .C2(n26839), .A(
        n23333), .ZN(n23328) );
  AOI22_X1 U22853 ( .A1(n26833), .A2(n25871), .B1(n26827), .B2(n21000), .ZN(
        n23333) );
  OAI221_X1 U22854 ( .B1(n9597), .B2(n26845), .C1(n20799), .C2(n26839), .A(
        n23315), .ZN(n23310) );
  AOI22_X1 U22855 ( .A1(n26833), .A2(n25876), .B1(n26827), .B2(n20999), .ZN(
        n23315) );
  OAI221_X1 U22856 ( .B1(n9596), .B2(n26846), .C1(n20798), .C2(n26840), .A(
        n23297), .ZN(n23292) );
  AOI22_X1 U22857 ( .A1(n26834), .A2(n25881), .B1(n26828), .B2(n20998), .ZN(
        n23297) );
  OAI221_X1 U22858 ( .B1(n9595), .B2(n26846), .C1(n20797), .C2(n26840), .A(
        n23279), .ZN(n23274) );
  AOI22_X1 U22859 ( .A1(n26834), .A2(n25886), .B1(n26828), .B2(n20997), .ZN(
        n23279) );
  OAI221_X1 U22860 ( .B1(n9594), .B2(n26846), .C1(n20796), .C2(n26840), .A(
        n23261), .ZN(n23256) );
  AOI22_X1 U22861 ( .A1(n26834), .A2(n25891), .B1(n26828), .B2(n20996), .ZN(
        n23261) );
  OAI221_X1 U22862 ( .B1(n9593), .B2(n26846), .C1(n20795), .C2(n26840), .A(
        n23243), .ZN(n23238) );
  AOI22_X1 U22863 ( .A1(n26834), .A2(n25896), .B1(n26828), .B2(n20995), .ZN(
        n23243) );
  OAI221_X1 U22864 ( .B1(n9592), .B2(n26846), .C1(n20794), .C2(n26840), .A(
        n23225), .ZN(n23220) );
  AOI22_X1 U22865 ( .A1(n26834), .A2(n25901), .B1(n26828), .B2(n20994), .ZN(
        n23225) );
  OAI221_X1 U22866 ( .B1(n9591), .B2(n26846), .C1(n20793), .C2(n26840), .A(
        n23207), .ZN(n23202) );
  AOI22_X1 U22867 ( .A1(n26834), .A2(n25906), .B1(n26828), .B2(n20993), .ZN(
        n23207) );
  OAI221_X1 U22868 ( .B1(n9590), .B2(n26846), .C1(n20792), .C2(n26840), .A(
        n23189), .ZN(n23184) );
  AOI22_X1 U22869 ( .A1(n26834), .A2(n25911), .B1(n26828), .B2(n20992), .ZN(
        n23189) );
  OAI221_X1 U22870 ( .B1(n9589), .B2(n26846), .C1(n20791), .C2(n26840), .A(
        n23171), .ZN(n23166) );
  AOI22_X1 U22871 ( .A1(n26834), .A2(n25916), .B1(n26828), .B2(n20991), .ZN(
        n23171) );
  OAI221_X1 U22872 ( .B1(n9588), .B2(n26846), .C1(n20790), .C2(n26840), .A(
        n23153), .ZN(n23148) );
  AOI22_X1 U22873 ( .A1(n26834), .A2(n25921), .B1(n26828), .B2(n20990), .ZN(
        n23153) );
  OAI221_X1 U22874 ( .B1(n9587), .B2(n26846), .C1(n20789), .C2(n26840), .A(
        n23135), .ZN(n23130) );
  AOI22_X1 U22875 ( .A1(n26834), .A2(n25926), .B1(n26828), .B2(n20989), .ZN(
        n23135) );
  OAI221_X1 U22876 ( .B1(n9586), .B2(n26846), .C1(n20788), .C2(n26840), .A(
        n23117), .ZN(n23112) );
  AOI22_X1 U22877 ( .A1(n26834), .A2(n25931), .B1(n26828), .B2(n20988), .ZN(
        n23117) );
  OAI221_X1 U22878 ( .B1(n9585), .B2(n26846), .C1(n20787), .C2(n26840), .A(
        n23099), .ZN(n23094) );
  AOI22_X1 U22879 ( .A1(n26834), .A2(n25936), .B1(n26828), .B2(n20987), .ZN(
        n23099) );
  OAI221_X1 U22880 ( .B1(n9569), .B2(n26623), .C1(n21155), .C2(n26617), .A(
        n23986), .ZN(n23971) );
  AOI22_X1 U22881 ( .A1(n26611), .A2(n25696), .B1(n26605), .B2(n20963), .ZN(
        n23986) );
  OAI221_X1 U22882 ( .B1(n9572), .B2(n26623), .C1(n20774), .C2(n26617), .A(
        n24064), .ZN(n24059) );
  AOI22_X1 U22883 ( .A1(n26611), .A2(n25681), .B1(n26605), .B2(n20966), .ZN(
        n24064) );
  OAI221_X1 U22884 ( .B1(n9571), .B2(n26623), .C1(n20773), .C2(n26617), .A(
        n24046), .ZN(n24041) );
  AOI22_X1 U22885 ( .A1(n26611), .A2(n25686), .B1(n26605), .B2(n20965), .ZN(
        n24046) );
  OAI221_X1 U22886 ( .B1(n9570), .B2(n26623), .C1(n20772), .C2(n26617), .A(
        n24028), .ZN(n24023) );
  AOI22_X1 U22887 ( .A1(n26611), .A2(n25691), .B1(n26605), .B2(n20964), .ZN(
        n24028) );
  OAI221_X1 U22888 ( .B1(n9572), .B2(n26848), .C1(n20774), .C2(n26842), .A(
        n22865), .ZN(n22860) );
  AOI22_X1 U22889 ( .A1(n26836), .A2(n25681), .B1(n26830), .B2(n20966), .ZN(
        n22865) );
  OAI221_X1 U22890 ( .B1(n9571), .B2(n26848), .C1(n20773), .C2(n26842), .A(
        n22847), .ZN(n22842) );
  AOI22_X1 U22891 ( .A1(n26836), .A2(n25686), .B1(n26830), .B2(n20965), .ZN(
        n22847) );
  OAI221_X1 U22892 ( .B1(n9570), .B2(n26848), .C1(n20772), .C2(n26842), .A(
        n22829), .ZN(n22824) );
  AOI22_X1 U22893 ( .A1(n26836), .A2(n25691), .B1(n26830), .B2(n20964), .ZN(
        n22829) );
  OAI221_X1 U22894 ( .B1(n9569), .B2(n26848), .C1(n21155), .C2(n26842), .A(
        n22787), .ZN(n22772) );
  AOI22_X1 U22895 ( .A1(n26836), .A2(n25696), .B1(n26830), .B2(n20963), .ZN(
        n22787) );
  OAI221_X1 U22896 ( .B1(n21747), .B2(n26595), .C1(n22367), .C2(n26589), .A(
        n24929), .ZN(n24922) );
  AOI222_X1 U22897 ( .A1(n26583), .A2(n25762), .B1(n26577), .B2(n21082), .C1(
        n26571), .C2(n21142), .ZN(n24929) );
  OAI221_X1 U22898 ( .B1(n21746), .B2(n26595), .C1(n22366), .C2(n26589), .A(
        n24911), .ZN(n24904) );
  AOI222_X1 U22899 ( .A1(n26583), .A2(n25767), .B1(n26577), .B2(n21081), .C1(
        n26571), .C2(n21141), .ZN(n24911) );
  OAI221_X1 U22900 ( .B1(n21745), .B2(n26595), .C1(n22365), .C2(n26589), .A(
        n24893), .ZN(n24886) );
  AOI222_X1 U22901 ( .A1(n26583), .A2(n25772), .B1(n26577), .B2(n21080), .C1(
        n26571), .C2(n21140), .ZN(n24893) );
  OAI221_X1 U22902 ( .B1(n21744), .B2(n26595), .C1(n22364), .C2(n26589), .A(
        n24875), .ZN(n24868) );
  AOI222_X1 U22903 ( .A1(n26583), .A2(n25777), .B1(n26577), .B2(n21079), .C1(
        n26571), .C2(n21139), .ZN(n24875) );
  OAI221_X1 U22904 ( .B1(n21743), .B2(n26595), .C1(n22363), .C2(n26589), .A(
        n24857), .ZN(n24850) );
  AOI222_X1 U22905 ( .A1(n26583), .A2(n25782), .B1(n26577), .B2(n21078), .C1(
        n26571), .C2(n21138), .ZN(n24857) );
  OAI221_X1 U22906 ( .B1(n21742), .B2(n26595), .C1(n22362), .C2(n26589), .A(
        n24839), .ZN(n24832) );
  AOI222_X1 U22907 ( .A1(n26583), .A2(n25787), .B1(n26577), .B2(n21077), .C1(
        n26571), .C2(n21137), .ZN(n24839) );
  OAI221_X1 U22908 ( .B1(n21741), .B2(n26595), .C1(n22361), .C2(n26589), .A(
        n24821), .ZN(n24814) );
  AOI222_X1 U22909 ( .A1(n26583), .A2(n25792), .B1(n26577), .B2(n21076), .C1(
        n26571), .C2(n21136), .ZN(n24821) );
  OAI221_X1 U22910 ( .B1(n21740), .B2(n26595), .C1(n22360), .C2(n26589), .A(
        n24803), .ZN(n24796) );
  AOI222_X1 U22911 ( .A1(n26583), .A2(n25797), .B1(n26577), .B2(n21075), .C1(
        n26571), .C2(n21135), .ZN(n24803) );
  OAI221_X1 U22912 ( .B1(n21739), .B2(n26595), .C1(n22359), .C2(n26589), .A(
        n24785), .ZN(n24778) );
  AOI222_X1 U22913 ( .A1(n26583), .A2(n25802), .B1(n26577), .B2(n21074), .C1(
        n26571), .C2(n21134), .ZN(n24785) );
  OAI221_X1 U22914 ( .B1(n21738), .B2(n26595), .C1(n22358), .C2(n26589), .A(
        n24767), .ZN(n24760) );
  AOI222_X1 U22915 ( .A1(n26583), .A2(n25807), .B1(n26577), .B2(n21073), .C1(
        n26571), .C2(n21133), .ZN(n24767) );
  OAI221_X1 U22916 ( .B1(n21737), .B2(n26595), .C1(n22357), .C2(n26589), .A(
        n24749), .ZN(n24742) );
  AOI222_X1 U22917 ( .A1(n26583), .A2(n25812), .B1(n26577), .B2(n21072), .C1(
        n26571), .C2(n21132), .ZN(n24749) );
  OAI221_X1 U22918 ( .B1(n21736), .B2(n26595), .C1(n22356), .C2(n26589), .A(
        n24731), .ZN(n24724) );
  AOI222_X1 U22919 ( .A1(n26583), .A2(n25817), .B1(n26577), .B2(n21071), .C1(
        n26571), .C2(n21131), .ZN(n24731) );
  OAI221_X1 U22920 ( .B1(n21735), .B2(n26596), .C1(n22355), .C2(n26590), .A(
        n24713), .ZN(n24706) );
  AOI222_X1 U22921 ( .A1(n26584), .A2(n25822), .B1(n26578), .B2(n21070), .C1(
        n26572), .C2(n21130), .ZN(n24713) );
  OAI221_X1 U22922 ( .B1(n21734), .B2(n26596), .C1(n22354), .C2(n26590), .A(
        n24695), .ZN(n24688) );
  AOI222_X1 U22923 ( .A1(n26584), .A2(n25827), .B1(n26578), .B2(n21069), .C1(
        n26572), .C2(n21129), .ZN(n24695) );
  OAI221_X1 U22924 ( .B1(n21733), .B2(n26596), .C1(n22353), .C2(n26590), .A(
        n24677), .ZN(n24670) );
  AOI222_X1 U22925 ( .A1(n26584), .A2(n25832), .B1(n26578), .B2(n21068), .C1(
        n26572), .C2(n21128), .ZN(n24677) );
  OAI221_X1 U22926 ( .B1(n21732), .B2(n26596), .C1(n22352), .C2(n26590), .A(
        n24659), .ZN(n24652) );
  AOI222_X1 U22927 ( .A1(n26584), .A2(n25837), .B1(n26578), .B2(n21067), .C1(
        n26572), .C2(n21127), .ZN(n24659) );
  OAI221_X1 U22928 ( .B1(n21731), .B2(n26596), .C1(n22351), .C2(n26590), .A(
        n24641), .ZN(n24634) );
  AOI222_X1 U22929 ( .A1(n26584), .A2(n25842), .B1(n26578), .B2(n21066), .C1(
        n26572), .C2(n21126), .ZN(n24641) );
  OAI221_X1 U22930 ( .B1(n21730), .B2(n26596), .C1(n22350), .C2(n26590), .A(
        n24623), .ZN(n24616) );
  AOI222_X1 U22931 ( .A1(n26584), .A2(n25847), .B1(n26578), .B2(n21065), .C1(
        n26572), .C2(n21125), .ZN(n24623) );
  OAI221_X1 U22932 ( .B1(n21729), .B2(n26596), .C1(n22349), .C2(n26590), .A(
        n24605), .ZN(n24598) );
  AOI222_X1 U22933 ( .A1(n26584), .A2(n25852), .B1(n26578), .B2(n21064), .C1(
        n26572), .C2(n21124), .ZN(n24605) );
  OAI221_X1 U22934 ( .B1(n21728), .B2(n26596), .C1(n22348), .C2(n26590), .A(
        n24587), .ZN(n24580) );
  AOI222_X1 U22935 ( .A1(n26584), .A2(n25857), .B1(n26578), .B2(n21063), .C1(
        n26572), .C2(n21123), .ZN(n24587) );
  OAI221_X1 U22936 ( .B1(n21727), .B2(n26596), .C1(n22347), .C2(n26590), .A(
        n24569), .ZN(n24562) );
  AOI222_X1 U22937 ( .A1(n26584), .A2(n25862), .B1(n26578), .B2(n21062), .C1(
        n26572), .C2(n21122), .ZN(n24569) );
  OAI221_X1 U22938 ( .B1(n21726), .B2(n26596), .C1(n22346), .C2(n26590), .A(
        n24551), .ZN(n24544) );
  AOI222_X1 U22939 ( .A1(n26584), .A2(n25867), .B1(n26578), .B2(n21061), .C1(
        n26572), .C2(n21121), .ZN(n24551) );
  OAI221_X1 U22940 ( .B1(n21725), .B2(n26596), .C1(n22345), .C2(n26590), .A(
        n24533), .ZN(n24526) );
  AOI222_X1 U22941 ( .A1(n26584), .A2(n25872), .B1(n26578), .B2(n21060), .C1(
        n26572), .C2(n21120), .ZN(n24533) );
  OAI221_X1 U22942 ( .B1(n21724), .B2(n26596), .C1(n22344), .C2(n26590), .A(
        n24515), .ZN(n24508) );
  AOI222_X1 U22943 ( .A1(n26584), .A2(n25877), .B1(n26578), .B2(n21059), .C1(
        n26572), .C2(n21119), .ZN(n24515) );
  OAI221_X1 U22944 ( .B1(n21723), .B2(n26597), .C1(n22343), .C2(n26591), .A(
        n24497), .ZN(n24490) );
  AOI222_X1 U22945 ( .A1(n26585), .A2(n25882), .B1(n26579), .B2(n21058), .C1(
        n26573), .C2(n21118), .ZN(n24497) );
  OAI221_X1 U22946 ( .B1(n21722), .B2(n26597), .C1(n22342), .C2(n26591), .A(
        n24479), .ZN(n24472) );
  AOI222_X1 U22947 ( .A1(n26585), .A2(n25887), .B1(n26579), .B2(n21057), .C1(
        n26573), .C2(n21117), .ZN(n24479) );
  OAI221_X1 U22948 ( .B1(n21721), .B2(n26597), .C1(n22341), .C2(n26591), .A(
        n24461), .ZN(n24454) );
  AOI222_X1 U22949 ( .A1(n26585), .A2(n25892), .B1(n26579), .B2(n21056), .C1(
        n26573), .C2(n21116), .ZN(n24461) );
  OAI221_X1 U22950 ( .B1(n21720), .B2(n26597), .C1(n22340), .C2(n26591), .A(
        n24443), .ZN(n24436) );
  AOI222_X1 U22951 ( .A1(n26585), .A2(n25897), .B1(n26579), .B2(n21055), .C1(
        n26573), .C2(n21115), .ZN(n24443) );
  OAI221_X1 U22952 ( .B1(n21719), .B2(n26597), .C1(n22339), .C2(n26591), .A(
        n24425), .ZN(n24418) );
  AOI222_X1 U22953 ( .A1(n26585), .A2(n25902), .B1(n26579), .B2(n21054), .C1(
        n26573), .C2(n21114), .ZN(n24425) );
  OAI221_X1 U22954 ( .B1(n21718), .B2(n26597), .C1(n22338), .C2(n26591), .A(
        n24407), .ZN(n24400) );
  AOI222_X1 U22955 ( .A1(n26585), .A2(n25907), .B1(n26579), .B2(n21053), .C1(
        n26573), .C2(n21113), .ZN(n24407) );
  OAI221_X1 U22956 ( .B1(n21717), .B2(n26597), .C1(n22337), .C2(n26591), .A(
        n24389), .ZN(n24382) );
  AOI222_X1 U22957 ( .A1(n26585), .A2(n25912), .B1(n26579), .B2(n21052), .C1(
        n26573), .C2(n21112), .ZN(n24389) );
  OAI221_X1 U22958 ( .B1(n21716), .B2(n26597), .C1(n22336), .C2(n26591), .A(
        n24371), .ZN(n24364) );
  AOI222_X1 U22959 ( .A1(n26585), .A2(n25917), .B1(n26579), .B2(n21051), .C1(
        n26573), .C2(n21111), .ZN(n24371) );
  OAI221_X1 U22960 ( .B1(n21715), .B2(n26597), .C1(n22335), .C2(n26591), .A(
        n24353), .ZN(n24346) );
  AOI222_X1 U22961 ( .A1(n26585), .A2(n25922), .B1(n26579), .B2(n21050), .C1(
        n26573), .C2(n21110), .ZN(n24353) );
  OAI221_X1 U22962 ( .B1(n21714), .B2(n26597), .C1(n22334), .C2(n26591), .A(
        n24335), .ZN(n24328) );
  AOI222_X1 U22963 ( .A1(n26585), .A2(n25927), .B1(n26579), .B2(n21049), .C1(
        n26573), .C2(n21109), .ZN(n24335) );
  OAI221_X1 U22964 ( .B1(n21713), .B2(n26597), .C1(n22333), .C2(n26591), .A(
        n24317), .ZN(n24310) );
  AOI222_X1 U22965 ( .A1(n26585), .A2(n25932), .B1(n26579), .B2(n21048), .C1(
        n26573), .C2(n21108), .ZN(n24317) );
  OAI221_X1 U22966 ( .B1(n21712), .B2(n26597), .C1(n22332), .C2(n26591), .A(
        n24299), .ZN(n24292) );
  AOI222_X1 U22967 ( .A1(n26585), .A2(n25937), .B1(n26579), .B2(n21047), .C1(
        n26573), .C2(n21107), .ZN(n24299) );
  OAI221_X1 U22968 ( .B1(n21711), .B2(n26598), .C1(n22331), .C2(n26592), .A(
        n24281), .ZN(n24274) );
  AOI222_X1 U22969 ( .A1(n26586), .A2(n25942), .B1(n26580), .B2(n21046), .C1(
        n26574), .C2(n21106), .ZN(n24281) );
  OAI221_X1 U22970 ( .B1(n21710), .B2(n26598), .C1(n22330), .C2(n26592), .A(
        n24263), .ZN(n24256) );
  AOI222_X1 U22971 ( .A1(n26586), .A2(n25947), .B1(n26580), .B2(n21045), .C1(
        n26574), .C2(n21105), .ZN(n24263) );
  OAI221_X1 U22972 ( .B1(n21709), .B2(n26598), .C1(n22329), .C2(n26592), .A(
        n24245), .ZN(n24238) );
  AOI222_X1 U22973 ( .A1(n26586), .A2(n25952), .B1(n26580), .B2(n21044), .C1(
        n26574), .C2(n21104), .ZN(n24245) );
  OAI221_X1 U22974 ( .B1(n21708), .B2(n26598), .C1(n22328), .C2(n26592), .A(
        n24227), .ZN(n24220) );
  AOI222_X1 U22975 ( .A1(n26586), .A2(n25957), .B1(n26580), .B2(n21043), .C1(
        n26574), .C2(n21103), .ZN(n24227) );
  OAI221_X1 U22976 ( .B1(n21707), .B2(n26598), .C1(n22327), .C2(n26592), .A(
        n24209), .ZN(n24202) );
  AOI222_X1 U22977 ( .A1(n26586), .A2(n25962), .B1(n26580), .B2(n21042), .C1(
        n26574), .C2(n21102), .ZN(n24209) );
  OAI221_X1 U22978 ( .B1(n21706), .B2(n26598), .C1(n22326), .C2(n26592), .A(
        n24191), .ZN(n24184) );
  AOI222_X1 U22979 ( .A1(n26586), .A2(n25967), .B1(n26580), .B2(n21041), .C1(
        n26574), .C2(n21101), .ZN(n24191) );
  OAI221_X1 U22980 ( .B1(n21705), .B2(n26598), .C1(n22325), .C2(n26592), .A(
        n24173), .ZN(n24166) );
  AOI222_X1 U22981 ( .A1(n26586), .A2(n25972), .B1(n26580), .B2(n21040), .C1(
        n26574), .C2(n21100), .ZN(n24173) );
  OAI221_X1 U22982 ( .B1(n21704), .B2(n26598), .C1(n22324), .C2(n26592), .A(
        n24155), .ZN(n24148) );
  AOI222_X1 U22983 ( .A1(n26586), .A2(n25977), .B1(n26580), .B2(n21039), .C1(
        n26574), .C2(n21099), .ZN(n24155) );
  OAI221_X1 U22984 ( .B1(n21703), .B2(n26598), .C1(n22323), .C2(n26592), .A(
        n24137), .ZN(n24130) );
  AOI222_X1 U22985 ( .A1(n26586), .A2(n25982), .B1(n26580), .B2(n21038), .C1(
        n26574), .C2(n21098), .ZN(n24137) );
  OAI221_X1 U22986 ( .B1(n21702), .B2(n26598), .C1(n22322), .C2(n26592), .A(
        n24119), .ZN(n24112) );
  AOI222_X1 U22987 ( .A1(n26586), .A2(n25987), .B1(n26580), .B2(n21037), .C1(
        n26574), .C2(n21097), .ZN(n24119) );
  OAI221_X1 U22988 ( .B1(n21701), .B2(n26598), .C1(n22321), .C2(n26592), .A(
        n24101), .ZN(n24094) );
  AOI222_X1 U22989 ( .A1(n26586), .A2(n25992), .B1(n26580), .B2(n21036), .C1(
        n26574), .C2(n21096), .ZN(n24101) );
  OAI221_X1 U22990 ( .B1(n21700), .B2(n26598), .C1(n22320), .C2(n26592), .A(
        n24083), .ZN(n24076) );
  AOI222_X1 U22991 ( .A1(n26586), .A2(n25997), .B1(n26580), .B2(n21035), .C1(
        n26574), .C2(n21095), .ZN(n24083) );
  OAI221_X1 U22992 ( .B1(n21747), .B2(n26820), .C1(n22367), .C2(n26814), .A(
        n23730), .ZN(n23723) );
  AOI222_X1 U22993 ( .A1(n26808), .A2(n25762), .B1(n26802), .B2(n21082), .C1(
        n26796), .C2(n21142), .ZN(n23730) );
  OAI221_X1 U22994 ( .B1(n21746), .B2(n26820), .C1(n22366), .C2(n26814), .A(
        n23712), .ZN(n23705) );
  AOI222_X1 U22995 ( .A1(n26808), .A2(n25767), .B1(n26802), .B2(n21081), .C1(
        n26796), .C2(n21141), .ZN(n23712) );
  OAI221_X1 U22996 ( .B1(n21745), .B2(n26820), .C1(n22365), .C2(n26814), .A(
        n23694), .ZN(n23687) );
  AOI222_X1 U22997 ( .A1(n26808), .A2(n25772), .B1(n26802), .B2(n21080), .C1(
        n26796), .C2(n21140), .ZN(n23694) );
  OAI221_X1 U22998 ( .B1(n21744), .B2(n26820), .C1(n22364), .C2(n26814), .A(
        n23676), .ZN(n23669) );
  AOI222_X1 U22999 ( .A1(n26808), .A2(n25777), .B1(n26802), .B2(n21079), .C1(
        n26796), .C2(n21139), .ZN(n23676) );
  OAI221_X1 U23000 ( .B1(n21743), .B2(n26820), .C1(n22363), .C2(n26814), .A(
        n23658), .ZN(n23651) );
  AOI222_X1 U23001 ( .A1(n26808), .A2(n25782), .B1(n26802), .B2(n21078), .C1(
        n26796), .C2(n21138), .ZN(n23658) );
  OAI221_X1 U23002 ( .B1(n21742), .B2(n26820), .C1(n22362), .C2(n26814), .A(
        n23640), .ZN(n23633) );
  AOI222_X1 U23003 ( .A1(n26808), .A2(n25787), .B1(n26802), .B2(n21077), .C1(
        n26796), .C2(n21137), .ZN(n23640) );
  OAI221_X1 U23004 ( .B1(n21741), .B2(n26820), .C1(n22361), .C2(n26814), .A(
        n23622), .ZN(n23615) );
  AOI222_X1 U23005 ( .A1(n26808), .A2(n25792), .B1(n26802), .B2(n21076), .C1(
        n26796), .C2(n21136), .ZN(n23622) );
  OAI221_X1 U23006 ( .B1(n21740), .B2(n26820), .C1(n22360), .C2(n26814), .A(
        n23604), .ZN(n23597) );
  AOI222_X1 U23007 ( .A1(n26808), .A2(n25797), .B1(n26802), .B2(n21075), .C1(
        n26796), .C2(n21135), .ZN(n23604) );
  OAI221_X1 U23008 ( .B1(n21739), .B2(n26820), .C1(n22359), .C2(n26814), .A(
        n23586), .ZN(n23579) );
  AOI222_X1 U23009 ( .A1(n26808), .A2(n25802), .B1(n26802), .B2(n21074), .C1(
        n26796), .C2(n21134), .ZN(n23586) );
  OAI221_X1 U23010 ( .B1(n21738), .B2(n26820), .C1(n22358), .C2(n26814), .A(
        n23568), .ZN(n23561) );
  AOI222_X1 U23011 ( .A1(n26808), .A2(n25807), .B1(n26802), .B2(n21073), .C1(
        n26796), .C2(n21133), .ZN(n23568) );
  OAI221_X1 U23012 ( .B1(n21737), .B2(n26820), .C1(n22357), .C2(n26814), .A(
        n23550), .ZN(n23543) );
  AOI222_X1 U23013 ( .A1(n26808), .A2(n25812), .B1(n26802), .B2(n21072), .C1(
        n26796), .C2(n21132), .ZN(n23550) );
  OAI221_X1 U23014 ( .B1(n21736), .B2(n26820), .C1(n22356), .C2(n26814), .A(
        n23532), .ZN(n23525) );
  AOI222_X1 U23015 ( .A1(n26808), .A2(n25817), .B1(n26802), .B2(n21071), .C1(
        n26796), .C2(n21131), .ZN(n23532) );
  OAI221_X1 U23016 ( .B1(n21735), .B2(n26821), .C1(n22355), .C2(n26815), .A(
        n23514), .ZN(n23507) );
  AOI222_X1 U23017 ( .A1(n26809), .A2(n25822), .B1(n26803), .B2(n21070), .C1(
        n26797), .C2(n21130), .ZN(n23514) );
  OAI221_X1 U23018 ( .B1(n21734), .B2(n26821), .C1(n22354), .C2(n26815), .A(
        n23496), .ZN(n23489) );
  AOI222_X1 U23019 ( .A1(n26809), .A2(n25827), .B1(n26803), .B2(n21069), .C1(
        n26797), .C2(n21129), .ZN(n23496) );
  OAI221_X1 U23020 ( .B1(n21733), .B2(n26821), .C1(n22353), .C2(n26815), .A(
        n23478), .ZN(n23471) );
  AOI222_X1 U23021 ( .A1(n26809), .A2(n25832), .B1(n26803), .B2(n21068), .C1(
        n26797), .C2(n21128), .ZN(n23478) );
  OAI221_X1 U23022 ( .B1(n21732), .B2(n26821), .C1(n22352), .C2(n26815), .A(
        n23460), .ZN(n23453) );
  AOI222_X1 U23023 ( .A1(n26809), .A2(n25837), .B1(n26803), .B2(n21067), .C1(
        n26797), .C2(n21127), .ZN(n23460) );
  OAI221_X1 U23024 ( .B1(n21731), .B2(n26821), .C1(n22351), .C2(n26815), .A(
        n23442), .ZN(n23435) );
  AOI222_X1 U23025 ( .A1(n26809), .A2(n25842), .B1(n26803), .B2(n21066), .C1(
        n26797), .C2(n21126), .ZN(n23442) );
  OAI221_X1 U23026 ( .B1(n21730), .B2(n26821), .C1(n22350), .C2(n26815), .A(
        n23424), .ZN(n23417) );
  AOI222_X1 U23027 ( .A1(n26809), .A2(n25847), .B1(n26803), .B2(n21065), .C1(
        n26797), .C2(n21125), .ZN(n23424) );
  OAI221_X1 U23028 ( .B1(n21729), .B2(n26821), .C1(n22349), .C2(n26815), .A(
        n23406), .ZN(n23399) );
  AOI222_X1 U23029 ( .A1(n26809), .A2(n25852), .B1(n26803), .B2(n21064), .C1(
        n26797), .C2(n21124), .ZN(n23406) );
  OAI221_X1 U23030 ( .B1(n21728), .B2(n26821), .C1(n22348), .C2(n26815), .A(
        n23388), .ZN(n23381) );
  AOI222_X1 U23031 ( .A1(n26809), .A2(n25857), .B1(n26803), .B2(n21063), .C1(
        n26797), .C2(n21123), .ZN(n23388) );
  OAI221_X1 U23032 ( .B1(n21727), .B2(n26821), .C1(n22347), .C2(n26815), .A(
        n23370), .ZN(n23363) );
  AOI222_X1 U23033 ( .A1(n26809), .A2(n25862), .B1(n26803), .B2(n21062), .C1(
        n26797), .C2(n21122), .ZN(n23370) );
  OAI221_X1 U23034 ( .B1(n21726), .B2(n26821), .C1(n22346), .C2(n26815), .A(
        n23352), .ZN(n23345) );
  AOI222_X1 U23035 ( .A1(n26809), .A2(n25867), .B1(n26803), .B2(n21061), .C1(
        n26797), .C2(n21121), .ZN(n23352) );
  OAI221_X1 U23036 ( .B1(n21725), .B2(n26821), .C1(n22345), .C2(n26815), .A(
        n23334), .ZN(n23327) );
  AOI222_X1 U23037 ( .A1(n26809), .A2(n25872), .B1(n26803), .B2(n21060), .C1(
        n26797), .C2(n21120), .ZN(n23334) );
  OAI221_X1 U23038 ( .B1(n21724), .B2(n26821), .C1(n22344), .C2(n26815), .A(
        n23316), .ZN(n23309) );
  AOI222_X1 U23039 ( .A1(n26809), .A2(n25877), .B1(n26803), .B2(n21059), .C1(
        n26797), .C2(n21119), .ZN(n23316) );
  OAI221_X1 U23040 ( .B1(n21723), .B2(n26822), .C1(n22343), .C2(n26816), .A(
        n23298), .ZN(n23291) );
  AOI222_X1 U23041 ( .A1(n26810), .A2(n25882), .B1(n26804), .B2(n21058), .C1(
        n26798), .C2(n21118), .ZN(n23298) );
  OAI221_X1 U23042 ( .B1(n21722), .B2(n26822), .C1(n22342), .C2(n26816), .A(
        n23280), .ZN(n23273) );
  AOI222_X1 U23043 ( .A1(n26810), .A2(n25887), .B1(n26804), .B2(n21057), .C1(
        n26798), .C2(n21117), .ZN(n23280) );
  OAI221_X1 U23044 ( .B1(n21721), .B2(n26822), .C1(n22341), .C2(n26816), .A(
        n23262), .ZN(n23255) );
  AOI222_X1 U23045 ( .A1(n26810), .A2(n25892), .B1(n26804), .B2(n21056), .C1(
        n26798), .C2(n21116), .ZN(n23262) );
  OAI221_X1 U23046 ( .B1(n21720), .B2(n26822), .C1(n22340), .C2(n26816), .A(
        n23244), .ZN(n23237) );
  AOI222_X1 U23047 ( .A1(n26810), .A2(n25897), .B1(n26804), .B2(n21055), .C1(
        n26798), .C2(n21115), .ZN(n23244) );
  OAI221_X1 U23048 ( .B1(n21719), .B2(n26822), .C1(n22339), .C2(n26816), .A(
        n23226), .ZN(n23219) );
  AOI222_X1 U23049 ( .A1(n26810), .A2(n25902), .B1(n26804), .B2(n21054), .C1(
        n26798), .C2(n21114), .ZN(n23226) );
  OAI221_X1 U23050 ( .B1(n21718), .B2(n26822), .C1(n22338), .C2(n26816), .A(
        n23208), .ZN(n23201) );
  AOI222_X1 U23051 ( .A1(n26810), .A2(n25907), .B1(n26804), .B2(n21053), .C1(
        n26798), .C2(n21113), .ZN(n23208) );
  OAI221_X1 U23052 ( .B1(n21717), .B2(n26822), .C1(n22337), .C2(n26816), .A(
        n23190), .ZN(n23183) );
  AOI222_X1 U23053 ( .A1(n26810), .A2(n25912), .B1(n26804), .B2(n21052), .C1(
        n26798), .C2(n21112), .ZN(n23190) );
  OAI221_X1 U23054 ( .B1(n21716), .B2(n26822), .C1(n22336), .C2(n26816), .A(
        n23172), .ZN(n23165) );
  AOI222_X1 U23055 ( .A1(n26810), .A2(n25917), .B1(n26804), .B2(n21051), .C1(
        n26798), .C2(n21111), .ZN(n23172) );
  OAI221_X1 U23056 ( .B1(n21715), .B2(n26822), .C1(n22335), .C2(n26816), .A(
        n23154), .ZN(n23147) );
  AOI222_X1 U23057 ( .A1(n26810), .A2(n25922), .B1(n26804), .B2(n21050), .C1(
        n26798), .C2(n21110), .ZN(n23154) );
  OAI221_X1 U23058 ( .B1(n21714), .B2(n26822), .C1(n22334), .C2(n26816), .A(
        n23136), .ZN(n23129) );
  AOI222_X1 U23059 ( .A1(n26810), .A2(n25927), .B1(n26804), .B2(n21049), .C1(
        n26798), .C2(n21109), .ZN(n23136) );
  OAI221_X1 U23060 ( .B1(n21713), .B2(n26822), .C1(n22333), .C2(n26816), .A(
        n23118), .ZN(n23111) );
  AOI222_X1 U23061 ( .A1(n26810), .A2(n25932), .B1(n26804), .B2(n21048), .C1(
        n26798), .C2(n21108), .ZN(n23118) );
  OAI221_X1 U23062 ( .B1(n21712), .B2(n26822), .C1(n22332), .C2(n26816), .A(
        n23100), .ZN(n23093) );
  AOI222_X1 U23063 ( .A1(n26810), .A2(n25937), .B1(n26804), .B2(n21047), .C1(
        n26798), .C2(n21107), .ZN(n23100) );
  OAI221_X1 U23064 ( .B1(n21711), .B2(n26823), .C1(n22331), .C2(n26817), .A(
        n23082), .ZN(n23075) );
  AOI222_X1 U23065 ( .A1(n26811), .A2(n25942), .B1(n26805), .B2(n21046), .C1(
        n26799), .C2(n21106), .ZN(n23082) );
  OAI221_X1 U23066 ( .B1(n21710), .B2(n26823), .C1(n22330), .C2(n26817), .A(
        n23064), .ZN(n23057) );
  AOI222_X1 U23067 ( .A1(n26811), .A2(n25947), .B1(n26805), .B2(n21045), .C1(
        n26799), .C2(n21105), .ZN(n23064) );
  OAI221_X1 U23068 ( .B1(n21709), .B2(n26823), .C1(n22329), .C2(n26817), .A(
        n23046), .ZN(n23039) );
  AOI222_X1 U23069 ( .A1(n26811), .A2(n25952), .B1(n26805), .B2(n21044), .C1(
        n26799), .C2(n21104), .ZN(n23046) );
  OAI221_X1 U23070 ( .B1(n21708), .B2(n26823), .C1(n22328), .C2(n26817), .A(
        n23028), .ZN(n23021) );
  AOI222_X1 U23071 ( .A1(n26811), .A2(n25957), .B1(n26805), .B2(n21043), .C1(
        n26799), .C2(n21103), .ZN(n23028) );
  OAI221_X1 U23072 ( .B1(n21707), .B2(n26823), .C1(n22327), .C2(n26817), .A(
        n23010), .ZN(n23003) );
  AOI222_X1 U23073 ( .A1(n26811), .A2(n25962), .B1(n26805), .B2(n21042), .C1(
        n26799), .C2(n21102), .ZN(n23010) );
  OAI221_X1 U23074 ( .B1(n21706), .B2(n26823), .C1(n22326), .C2(n26817), .A(
        n22992), .ZN(n22985) );
  AOI222_X1 U23075 ( .A1(n26811), .A2(n25967), .B1(n26805), .B2(n21041), .C1(
        n26799), .C2(n21101), .ZN(n22992) );
  OAI221_X1 U23076 ( .B1(n21705), .B2(n26823), .C1(n22325), .C2(n26817), .A(
        n22974), .ZN(n22967) );
  AOI222_X1 U23077 ( .A1(n26811), .A2(n25972), .B1(n26805), .B2(n21040), .C1(
        n26799), .C2(n21100), .ZN(n22974) );
  OAI221_X1 U23078 ( .B1(n21704), .B2(n26823), .C1(n22324), .C2(n26817), .A(
        n22956), .ZN(n22949) );
  AOI222_X1 U23079 ( .A1(n26811), .A2(n25977), .B1(n26805), .B2(n21039), .C1(
        n26799), .C2(n21099), .ZN(n22956) );
  OAI221_X1 U23080 ( .B1(n21703), .B2(n26823), .C1(n22323), .C2(n26817), .A(
        n22938), .ZN(n22931) );
  AOI222_X1 U23081 ( .A1(n26811), .A2(n25982), .B1(n26805), .B2(n21038), .C1(
        n26799), .C2(n21098), .ZN(n22938) );
  OAI221_X1 U23082 ( .B1(n21702), .B2(n26823), .C1(n22322), .C2(n26817), .A(
        n22920), .ZN(n22913) );
  AOI222_X1 U23083 ( .A1(n26811), .A2(n25987), .B1(n26805), .B2(n21037), .C1(
        n26799), .C2(n21097), .ZN(n22920) );
  OAI221_X1 U23084 ( .B1(n21701), .B2(n26823), .C1(n22321), .C2(n26817), .A(
        n22902), .ZN(n22895) );
  AOI222_X1 U23085 ( .A1(n26811), .A2(n25992), .B1(n26805), .B2(n21036), .C1(
        n26799), .C2(n21096), .ZN(n22902) );
  OAI221_X1 U23086 ( .B1(n21700), .B2(n26823), .C1(n22320), .C2(n26817), .A(
        n22884), .ZN(n22877) );
  AOI222_X1 U23087 ( .A1(n26811), .A2(n25997), .B1(n26805), .B2(n21035), .C1(
        n26799), .C2(n21095), .ZN(n22884) );
  OAI221_X1 U23088 ( .B1(n21508), .B2(n26476), .C1(n27473), .C2(n26470), .A(
        n24016), .ZN(n23995) );
  AOI222_X1 U23089 ( .A1(n26464), .A2(n25558), .B1(n26458), .B2(n25574), .C1(
        n26452), .C2(n25582), .ZN(n24016) );
  OAI221_X1 U23090 ( .B1(n21511), .B2(n26476), .C1(n27464), .C2(n26470), .A(
        n24073), .ZN(n24066) );
  AOI222_X1 U23091 ( .A1(n26464), .A2(n25555), .B1(n26458), .B2(n25571), .C1(
        n26452), .C2(n25579), .ZN(n24073) );
  OAI221_X1 U23092 ( .B1(n21510), .B2(n26476), .C1(n27467), .C2(n26470), .A(
        n24055), .ZN(n24048) );
  AOI222_X1 U23093 ( .A1(n26464), .A2(n25556), .B1(n26458), .B2(n25572), .C1(
        n26452), .C2(n25580), .ZN(n24055) );
  OAI221_X1 U23094 ( .B1(n21509), .B2(n26476), .C1(n27470), .C2(n26470), .A(
        n24037), .ZN(n24030) );
  AOI222_X1 U23095 ( .A1(n26464), .A2(n25557), .B1(n26458), .B2(n25573), .C1(
        n26452), .C2(n25581), .ZN(n24037) );
  OAI221_X1 U23096 ( .B1(n21511), .B2(n26701), .C1(n27464), .C2(n26695), .A(
        n22874), .ZN(n22867) );
  AOI222_X1 U23097 ( .A1(n26689), .A2(n25555), .B1(n26683), .B2(n25571), .C1(
        n26677), .C2(n25579), .ZN(n22874) );
  OAI221_X1 U23098 ( .B1(n21510), .B2(n26701), .C1(n27467), .C2(n26695), .A(
        n22856), .ZN(n22849) );
  AOI222_X1 U23099 ( .A1(n26689), .A2(n25556), .B1(n26683), .B2(n25572), .C1(
        n26677), .C2(n25580), .ZN(n22856) );
  OAI221_X1 U23100 ( .B1(n21509), .B2(n26701), .C1(n27470), .C2(n26695), .A(
        n22838), .ZN(n22831) );
  AOI222_X1 U23101 ( .A1(n26689), .A2(n25557), .B1(n26683), .B2(n25573), .C1(
        n26677), .C2(n25581), .ZN(n22838) );
  OAI221_X1 U23102 ( .B1(n21508), .B2(n26701), .C1(n27473), .C2(n26695), .A(
        n22817), .ZN(n22796) );
  AOI222_X1 U23103 ( .A1(n26689), .A2(n25558), .B1(n26683), .B2(n25574), .C1(
        n26677), .C2(n25582), .ZN(n22817) );
  OAI221_X1 U23104 ( .B1(n21488), .B2(n26599), .C1(n22248), .C2(n26593), .A(
        n23991), .ZN(n23970) );
  AOI222_X1 U23105 ( .A1(n26587), .A2(n25697), .B1(n26581), .B2(n20967), .C1(
        n26575), .C2(n20971), .ZN(n23991) );
  OAI221_X1 U23106 ( .B1(n21491), .B2(n26599), .C1(n22251), .C2(n26593), .A(
        n24065), .ZN(n24058) );
  AOI222_X1 U23107 ( .A1(n26587), .A2(n25682), .B1(n26581), .B2(n20970), .C1(
        n26575), .C2(n20974), .ZN(n24065) );
  OAI221_X1 U23108 ( .B1(n21490), .B2(n26599), .C1(n22250), .C2(n26593), .A(
        n24047), .ZN(n24040) );
  AOI222_X1 U23109 ( .A1(n26587), .A2(n25687), .B1(n26581), .B2(n20969), .C1(
        n26575), .C2(n20973), .ZN(n24047) );
  OAI221_X1 U23110 ( .B1(n21489), .B2(n26599), .C1(n22249), .C2(n26593), .A(
        n24029), .ZN(n24022) );
  AOI222_X1 U23111 ( .A1(n26587), .A2(n25692), .B1(n26581), .B2(n20968), .C1(
        n26575), .C2(n20972), .ZN(n24029) );
  OAI221_X1 U23112 ( .B1(n21491), .B2(n26824), .C1(n22251), .C2(n26818), .A(
        n22866), .ZN(n22859) );
  AOI222_X1 U23113 ( .A1(n26812), .A2(n25682), .B1(n26806), .B2(n20970), .C1(
        n26800), .C2(n20974), .ZN(n22866) );
  OAI221_X1 U23114 ( .B1(n21490), .B2(n26824), .C1(n22250), .C2(n26818), .A(
        n22848), .ZN(n22841) );
  AOI222_X1 U23115 ( .A1(n26812), .A2(n25687), .B1(n26806), .B2(n20969), .C1(
        n26800), .C2(n20973), .ZN(n22848) );
  OAI221_X1 U23116 ( .B1(n21489), .B2(n26824), .C1(n22249), .C2(n26818), .A(
        n22830), .ZN(n22823) );
  AOI222_X1 U23117 ( .A1(n26812), .A2(n25692), .B1(n26806), .B2(n20968), .C1(
        n26800), .C2(n20972), .ZN(n22830) );
  OAI221_X1 U23118 ( .B1(n21488), .B2(n26824), .C1(n22248), .C2(n26818), .A(
        n22792), .ZN(n22771) );
  AOI222_X1 U23119 ( .A1(n26812), .A2(n25697), .B1(n26806), .B2(n20967), .C1(
        n26800), .C2(n20971), .ZN(n22792) );
  OAI221_X1 U23120 ( .B1(n9632), .B2(n26618), .C1(n20834), .C2(n26612), .A(
        n25152), .ZN(n25139) );
  AOI22_X1 U23121 ( .A1(n26606), .A2(n25701), .B1(n26600), .B2(n21034), .ZN(
        n25152) );
  OAI221_X1 U23122 ( .B1(n9631), .B2(n26618), .C1(n20833), .C2(n26612), .A(
        n25126), .ZN(n25121) );
  AOI22_X1 U23123 ( .A1(n26606), .A2(n25706), .B1(n26600), .B2(n21033), .ZN(
        n25126) );
  OAI221_X1 U23124 ( .B1(n9630), .B2(n26618), .C1(n20832), .C2(n26612), .A(
        n25108), .ZN(n25103) );
  AOI22_X1 U23125 ( .A1(n26606), .A2(n25711), .B1(n26600), .B2(n21032), .ZN(
        n25108) );
  OAI221_X1 U23126 ( .B1(n9629), .B2(n26618), .C1(n20831), .C2(n26612), .A(
        n25090), .ZN(n25085) );
  AOI22_X1 U23127 ( .A1(n26606), .A2(n25716), .B1(n26600), .B2(n21031), .ZN(
        n25090) );
  OAI221_X1 U23128 ( .B1(n9628), .B2(n26618), .C1(n20830), .C2(n26612), .A(
        n25072), .ZN(n25067) );
  AOI22_X1 U23129 ( .A1(n26606), .A2(n25721), .B1(n26600), .B2(n21030), .ZN(
        n25072) );
  OAI221_X1 U23130 ( .B1(n9627), .B2(n26618), .C1(n20829), .C2(n26612), .A(
        n25054), .ZN(n25049) );
  AOI22_X1 U23131 ( .A1(n26606), .A2(n25726), .B1(n26600), .B2(n21029), .ZN(
        n25054) );
  OAI221_X1 U23132 ( .B1(n9626), .B2(n26618), .C1(n20828), .C2(n26612), .A(
        n25036), .ZN(n25031) );
  AOI22_X1 U23133 ( .A1(n26606), .A2(n25731), .B1(n26600), .B2(n21028), .ZN(
        n25036) );
  OAI221_X1 U23134 ( .B1(n9625), .B2(n26618), .C1(n20827), .C2(n26612), .A(
        n25018), .ZN(n25013) );
  AOI22_X1 U23135 ( .A1(n26606), .A2(n25736), .B1(n26600), .B2(n21027), .ZN(
        n25018) );
  OAI221_X1 U23136 ( .B1(n9624), .B2(n26618), .C1(n20826), .C2(n26612), .A(
        n25000), .ZN(n24995) );
  AOI22_X1 U23137 ( .A1(n26606), .A2(n25741), .B1(n26600), .B2(n21026), .ZN(
        n25000) );
  OAI221_X1 U23138 ( .B1(n9623), .B2(n26618), .C1(n20825), .C2(n26612), .A(
        n24982), .ZN(n24977) );
  AOI22_X1 U23139 ( .A1(n26606), .A2(n25746), .B1(n26600), .B2(n21025), .ZN(
        n24982) );
  OAI221_X1 U23140 ( .B1(n9622), .B2(n26618), .C1(n20824), .C2(n26612), .A(
        n24964), .ZN(n24959) );
  AOI22_X1 U23141 ( .A1(n26606), .A2(n25751), .B1(n26600), .B2(n21024), .ZN(
        n24964) );
  OAI221_X1 U23142 ( .B1(n9621), .B2(n26618), .C1(n20823), .C2(n26612), .A(
        n24946), .ZN(n24941) );
  AOI22_X1 U23143 ( .A1(n26606), .A2(n25756), .B1(n26600), .B2(n21023), .ZN(
        n24946) );
  OAI221_X1 U23144 ( .B1(n9632), .B2(n26843), .C1(n20834), .C2(n26837), .A(
        n23953), .ZN(n23940) );
  AOI22_X1 U23145 ( .A1(n26831), .A2(n25701), .B1(n26825), .B2(n21034), .ZN(
        n23953) );
  OAI221_X1 U23146 ( .B1(n9631), .B2(n26843), .C1(n20833), .C2(n26837), .A(
        n23927), .ZN(n23922) );
  AOI22_X1 U23147 ( .A1(n26831), .A2(n25706), .B1(n26825), .B2(n21033), .ZN(
        n23927) );
  OAI221_X1 U23148 ( .B1(n9630), .B2(n26843), .C1(n20832), .C2(n26837), .A(
        n23909), .ZN(n23904) );
  AOI22_X1 U23149 ( .A1(n26831), .A2(n25711), .B1(n26825), .B2(n21032), .ZN(
        n23909) );
  OAI221_X1 U23150 ( .B1(n9629), .B2(n26843), .C1(n20831), .C2(n26837), .A(
        n23891), .ZN(n23886) );
  AOI22_X1 U23151 ( .A1(n26831), .A2(n25716), .B1(n26825), .B2(n21031), .ZN(
        n23891) );
  OAI221_X1 U23152 ( .B1(n9628), .B2(n26843), .C1(n20830), .C2(n26837), .A(
        n23873), .ZN(n23868) );
  AOI22_X1 U23153 ( .A1(n26831), .A2(n25721), .B1(n26825), .B2(n21030), .ZN(
        n23873) );
  OAI221_X1 U23154 ( .B1(n9627), .B2(n26843), .C1(n20829), .C2(n26837), .A(
        n23855), .ZN(n23850) );
  AOI22_X1 U23155 ( .A1(n26831), .A2(n25726), .B1(n26825), .B2(n21029), .ZN(
        n23855) );
  OAI221_X1 U23156 ( .B1(n9626), .B2(n26843), .C1(n20828), .C2(n26837), .A(
        n23837), .ZN(n23832) );
  AOI22_X1 U23157 ( .A1(n26831), .A2(n25731), .B1(n26825), .B2(n21028), .ZN(
        n23837) );
  OAI221_X1 U23158 ( .B1(n9625), .B2(n26843), .C1(n20827), .C2(n26837), .A(
        n23819), .ZN(n23814) );
  AOI22_X1 U23159 ( .A1(n26831), .A2(n25736), .B1(n26825), .B2(n21027), .ZN(
        n23819) );
  OAI221_X1 U23160 ( .B1(n9624), .B2(n26843), .C1(n20826), .C2(n26837), .A(
        n23801), .ZN(n23796) );
  AOI22_X1 U23161 ( .A1(n26831), .A2(n25741), .B1(n26825), .B2(n21026), .ZN(
        n23801) );
  OAI221_X1 U23162 ( .B1(n9623), .B2(n26843), .C1(n20825), .C2(n26837), .A(
        n23783), .ZN(n23778) );
  AOI22_X1 U23163 ( .A1(n26831), .A2(n25746), .B1(n26825), .B2(n21025), .ZN(
        n23783) );
  OAI221_X1 U23164 ( .B1(n9622), .B2(n26843), .C1(n20824), .C2(n26837), .A(
        n23765), .ZN(n23760) );
  AOI22_X1 U23165 ( .A1(n26831), .A2(n25751), .B1(n26825), .B2(n21024), .ZN(
        n23765) );
  OAI221_X1 U23166 ( .B1(n9621), .B2(n26843), .C1(n20823), .C2(n26837), .A(
        n23747), .ZN(n23742) );
  AOI22_X1 U23167 ( .A1(n26831), .A2(n25756), .B1(n26825), .B2(n21023), .ZN(
        n23747) );
  OAI221_X1 U23168 ( .B1(n22059), .B2(n26471), .C1(n27284), .C2(n26465), .A(
        n25166), .ZN(n25156) );
  AOI222_X1 U23169 ( .A1(n26459), .A2(n25595), .B1(n26453), .B2(n25619), .C1(
        n26447), .C2(n25667), .ZN(n25166) );
  OAI221_X1 U23170 ( .B1(n22058), .B2(n26471), .C1(n27287), .C2(n26465), .A(
        n25135), .ZN(n25128) );
  AOI222_X1 U23171 ( .A1(n26459), .A2(n25596), .B1(n26453), .B2(n25620), .C1(
        n26447), .C2(n25668), .ZN(n25135) );
  OAI221_X1 U23172 ( .B1(n22057), .B2(n26471), .C1(n27290), .C2(n26465), .A(
        n25117), .ZN(n25110) );
  AOI222_X1 U23173 ( .A1(n26459), .A2(n25597), .B1(n26453), .B2(n25621), .C1(
        n26447), .C2(n25669), .ZN(n25117) );
  OAI221_X1 U23174 ( .B1(n22056), .B2(n26471), .C1(n27293), .C2(n26465), .A(
        n25099), .ZN(n25092) );
  AOI222_X1 U23175 ( .A1(n26459), .A2(n25598), .B1(n26453), .B2(n25622), .C1(
        n26447), .C2(n25670), .ZN(n25099) );
  OAI221_X1 U23176 ( .B1(n22055), .B2(n26471), .C1(n27296), .C2(n26465), .A(
        n25081), .ZN(n25074) );
  AOI222_X1 U23177 ( .A1(n26459), .A2(n25599), .B1(n26453), .B2(n25623), .C1(
        n26447), .C2(n25671), .ZN(n25081) );
  OAI221_X1 U23178 ( .B1(n22054), .B2(n26471), .C1(n27299), .C2(n26465), .A(
        n25063), .ZN(n25056) );
  AOI222_X1 U23179 ( .A1(n26459), .A2(n25600), .B1(n26453), .B2(n25624), .C1(
        n26447), .C2(n25672), .ZN(n25063) );
  OAI221_X1 U23180 ( .B1(n22053), .B2(n26471), .C1(n27302), .C2(n26465), .A(
        n25045), .ZN(n25038) );
  AOI222_X1 U23181 ( .A1(n26459), .A2(n25601), .B1(n26453), .B2(n25625), .C1(
        n26447), .C2(n25673), .ZN(n25045) );
  OAI221_X1 U23182 ( .B1(n22052), .B2(n26471), .C1(n27305), .C2(n26465), .A(
        n25027), .ZN(n25020) );
  AOI222_X1 U23183 ( .A1(n26459), .A2(n25602), .B1(n26453), .B2(n25626), .C1(
        n26447), .C2(n25674), .ZN(n25027) );
  OAI221_X1 U23184 ( .B1(n22051), .B2(n26471), .C1(n27308), .C2(n26465), .A(
        n25009), .ZN(n25002) );
  AOI222_X1 U23185 ( .A1(n26459), .A2(n25603), .B1(n26453), .B2(n25627), .C1(
        n26447), .C2(n25675), .ZN(n25009) );
  OAI221_X1 U23186 ( .B1(n22050), .B2(n26471), .C1(n27311), .C2(n26465), .A(
        n24991), .ZN(n24984) );
  AOI222_X1 U23187 ( .A1(n26459), .A2(n25604), .B1(n26453), .B2(n25628), .C1(
        n26447), .C2(n25676), .ZN(n24991) );
  OAI221_X1 U23188 ( .B1(n22049), .B2(n26471), .C1(n27314), .C2(n26465), .A(
        n24973), .ZN(n24966) );
  AOI222_X1 U23189 ( .A1(n26459), .A2(n25605), .B1(n26453), .B2(n25629), .C1(
        n26447), .C2(n25677), .ZN(n24973) );
  OAI221_X1 U23190 ( .B1(n22048), .B2(n26471), .C1(n27317), .C2(n26465), .A(
        n24955), .ZN(n24948) );
  AOI222_X1 U23191 ( .A1(n26459), .A2(n25606), .B1(n26453), .B2(n25630), .C1(
        n26447), .C2(n25678), .ZN(n24955) );
  OAI221_X1 U23192 ( .B1(n22047), .B2(n26472), .C1(n27320), .C2(n26466), .A(
        n24937), .ZN(n24930) );
  AOI222_X1 U23193 ( .A1(n26460), .A2(n25215), .B1(n26454), .B2(n25407), .C1(
        n26448), .C2(n25503), .ZN(n24937) );
  OAI221_X1 U23194 ( .B1(n22046), .B2(n26472), .C1(n27323), .C2(n26466), .A(
        n24919), .ZN(n24912) );
  AOI222_X1 U23195 ( .A1(n26460), .A2(n25216), .B1(n26454), .B2(n25408), .C1(
        n26448), .C2(n25504), .ZN(n24919) );
  OAI221_X1 U23196 ( .B1(n22045), .B2(n26472), .C1(n27326), .C2(n26466), .A(
        n24901), .ZN(n24894) );
  AOI222_X1 U23197 ( .A1(n26460), .A2(n25217), .B1(n26454), .B2(n25409), .C1(
        n26448), .C2(n25505), .ZN(n24901) );
  OAI221_X1 U23198 ( .B1(n22044), .B2(n26472), .C1(n27329), .C2(n26466), .A(
        n24883), .ZN(n24876) );
  AOI222_X1 U23199 ( .A1(n26460), .A2(n25218), .B1(n26454), .B2(n25410), .C1(
        n26448), .C2(n25506), .ZN(n24883) );
  OAI221_X1 U23200 ( .B1(n22043), .B2(n26472), .C1(n27332), .C2(n26466), .A(
        n24865), .ZN(n24858) );
  AOI222_X1 U23201 ( .A1(n26460), .A2(n25219), .B1(n26454), .B2(n25411), .C1(
        n26448), .C2(n25507), .ZN(n24865) );
  OAI221_X1 U23202 ( .B1(n22042), .B2(n26472), .C1(n27335), .C2(n26466), .A(
        n24847), .ZN(n24840) );
  AOI222_X1 U23203 ( .A1(n26460), .A2(n25220), .B1(n26454), .B2(n25412), .C1(
        n26448), .C2(n25508), .ZN(n24847) );
  OAI221_X1 U23204 ( .B1(n22041), .B2(n26472), .C1(n27338), .C2(n26466), .A(
        n24829), .ZN(n24822) );
  AOI222_X1 U23205 ( .A1(n26460), .A2(n25221), .B1(n26454), .B2(n25413), .C1(
        n26448), .C2(n25509), .ZN(n24829) );
  OAI221_X1 U23206 ( .B1(n22040), .B2(n26472), .C1(n27341), .C2(n26466), .A(
        n24811), .ZN(n24804) );
  AOI222_X1 U23207 ( .A1(n26460), .A2(n25222), .B1(n26454), .B2(n25414), .C1(
        n26448), .C2(n25510), .ZN(n24811) );
  OAI221_X1 U23208 ( .B1(n22039), .B2(n26472), .C1(n27344), .C2(n26466), .A(
        n24793), .ZN(n24786) );
  AOI222_X1 U23209 ( .A1(n26460), .A2(n25223), .B1(n26454), .B2(n25415), .C1(
        n26448), .C2(n25511), .ZN(n24793) );
  OAI221_X1 U23210 ( .B1(n22038), .B2(n26472), .C1(n27347), .C2(n26466), .A(
        n24775), .ZN(n24768) );
  AOI222_X1 U23211 ( .A1(n26460), .A2(n25224), .B1(n26454), .B2(n25416), .C1(
        n26448), .C2(n25512), .ZN(n24775) );
  OAI221_X1 U23212 ( .B1(n22037), .B2(n26472), .C1(n27350), .C2(n26466), .A(
        n24757), .ZN(n24750) );
  AOI222_X1 U23213 ( .A1(n26460), .A2(n25225), .B1(n26454), .B2(n25417), .C1(
        n26448), .C2(n25513), .ZN(n24757) );
  OAI221_X1 U23214 ( .B1(n22036), .B2(n26472), .C1(n27353), .C2(n26466), .A(
        n24739), .ZN(n24732) );
  AOI222_X1 U23215 ( .A1(n26460), .A2(n25226), .B1(n26454), .B2(n25418), .C1(
        n26448), .C2(n25514), .ZN(n24739) );
  OAI221_X1 U23216 ( .B1(n22035), .B2(n26473), .C1(n27356), .C2(n26467), .A(
        n24721), .ZN(n24714) );
  AOI222_X1 U23217 ( .A1(n26461), .A2(n25227), .B1(n26455), .B2(n25419), .C1(
        n26449), .C2(n25515), .ZN(n24721) );
  OAI221_X1 U23218 ( .B1(n22034), .B2(n26473), .C1(n27359), .C2(n26467), .A(
        n24703), .ZN(n24696) );
  AOI222_X1 U23219 ( .A1(n26461), .A2(n25228), .B1(n26455), .B2(n25420), .C1(
        n26449), .C2(n25516), .ZN(n24703) );
  OAI221_X1 U23220 ( .B1(n22033), .B2(n26473), .C1(n27362), .C2(n26467), .A(
        n24685), .ZN(n24678) );
  AOI222_X1 U23221 ( .A1(n26461), .A2(n25229), .B1(n26455), .B2(n25421), .C1(
        n26449), .C2(n25517), .ZN(n24685) );
  OAI221_X1 U23222 ( .B1(n22032), .B2(n26473), .C1(n27365), .C2(n26467), .A(
        n24667), .ZN(n24660) );
  AOI222_X1 U23223 ( .A1(n26461), .A2(n25230), .B1(n26455), .B2(n25422), .C1(
        n26449), .C2(n25518), .ZN(n24667) );
  OAI221_X1 U23224 ( .B1(n22031), .B2(n26473), .C1(n27368), .C2(n26467), .A(
        n24649), .ZN(n24642) );
  AOI222_X1 U23225 ( .A1(n26461), .A2(n25231), .B1(n26455), .B2(n25423), .C1(
        n26449), .C2(n25519), .ZN(n24649) );
  OAI221_X1 U23226 ( .B1(n22030), .B2(n26473), .C1(n27371), .C2(n26467), .A(
        n24631), .ZN(n24624) );
  AOI222_X1 U23227 ( .A1(n26461), .A2(n25232), .B1(n26455), .B2(n25424), .C1(
        n26449), .C2(n25520), .ZN(n24631) );
  OAI221_X1 U23228 ( .B1(n22029), .B2(n26473), .C1(n27374), .C2(n26467), .A(
        n24613), .ZN(n24606) );
  AOI222_X1 U23229 ( .A1(n26461), .A2(n25233), .B1(n26455), .B2(n25425), .C1(
        n26449), .C2(n25521), .ZN(n24613) );
  OAI221_X1 U23230 ( .B1(n22028), .B2(n26473), .C1(n27377), .C2(n26467), .A(
        n24595), .ZN(n24588) );
  AOI222_X1 U23231 ( .A1(n26461), .A2(n25234), .B1(n26455), .B2(n25426), .C1(
        n26449), .C2(n25522), .ZN(n24595) );
  OAI221_X1 U23232 ( .B1(n22027), .B2(n26473), .C1(n27380), .C2(n26467), .A(
        n24577), .ZN(n24570) );
  AOI222_X1 U23233 ( .A1(n26461), .A2(n25235), .B1(n26455), .B2(n25427), .C1(
        n26449), .C2(n25523), .ZN(n24577) );
  OAI221_X1 U23234 ( .B1(n22026), .B2(n26473), .C1(n27383), .C2(n26467), .A(
        n24559), .ZN(n24552) );
  AOI222_X1 U23235 ( .A1(n26461), .A2(n25236), .B1(n26455), .B2(n25428), .C1(
        n26449), .C2(n25524), .ZN(n24559) );
  OAI221_X1 U23236 ( .B1(n22025), .B2(n26473), .C1(n27386), .C2(n26467), .A(
        n24541), .ZN(n24534) );
  AOI222_X1 U23237 ( .A1(n26461), .A2(n25237), .B1(n26455), .B2(n25429), .C1(
        n26449), .C2(n25525), .ZN(n24541) );
  OAI221_X1 U23238 ( .B1(n22024), .B2(n26473), .C1(n27389), .C2(n26467), .A(
        n24523), .ZN(n24516) );
  AOI222_X1 U23239 ( .A1(n26461), .A2(n25238), .B1(n26455), .B2(n25430), .C1(
        n26449), .C2(n25526), .ZN(n24523) );
  OAI221_X1 U23240 ( .B1(n22023), .B2(n26474), .C1(n27392), .C2(n26468), .A(
        n24505), .ZN(n24498) );
  AOI222_X1 U23241 ( .A1(n26462), .A2(n25239), .B1(n26456), .B2(n25431), .C1(
        n26450), .C2(n25527), .ZN(n24505) );
  OAI221_X1 U23242 ( .B1(n22022), .B2(n26474), .C1(n27395), .C2(n26468), .A(
        n24487), .ZN(n24480) );
  AOI222_X1 U23243 ( .A1(n26462), .A2(n25240), .B1(n26456), .B2(n25432), .C1(
        n26450), .C2(n25528), .ZN(n24487) );
  OAI221_X1 U23244 ( .B1(n22021), .B2(n26474), .C1(n27398), .C2(n26468), .A(
        n24469), .ZN(n24462) );
  AOI222_X1 U23245 ( .A1(n26462), .A2(n25241), .B1(n26456), .B2(n25433), .C1(
        n26450), .C2(n25529), .ZN(n24469) );
  OAI221_X1 U23246 ( .B1(n22020), .B2(n26474), .C1(n27401), .C2(n26468), .A(
        n24451), .ZN(n24444) );
  AOI222_X1 U23247 ( .A1(n26462), .A2(n25242), .B1(n26456), .B2(n25434), .C1(
        n26450), .C2(n25530), .ZN(n24451) );
  OAI221_X1 U23248 ( .B1(n22019), .B2(n26474), .C1(n27404), .C2(n26468), .A(
        n24433), .ZN(n24426) );
  AOI222_X1 U23249 ( .A1(n26462), .A2(n25243), .B1(n26456), .B2(n25435), .C1(
        n26450), .C2(n25531), .ZN(n24433) );
  OAI221_X1 U23250 ( .B1(n22018), .B2(n26474), .C1(n27407), .C2(n26468), .A(
        n24415), .ZN(n24408) );
  AOI222_X1 U23251 ( .A1(n26462), .A2(n25244), .B1(n26456), .B2(n25436), .C1(
        n26450), .C2(n25532), .ZN(n24415) );
  OAI221_X1 U23252 ( .B1(n22017), .B2(n26474), .C1(n27410), .C2(n26468), .A(
        n24397), .ZN(n24390) );
  AOI222_X1 U23253 ( .A1(n26462), .A2(n25245), .B1(n26456), .B2(n25437), .C1(
        n26450), .C2(n25533), .ZN(n24397) );
  OAI221_X1 U23254 ( .B1(n22016), .B2(n26474), .C1(n27413), .C2(n26468), .A(
        n24379), .ZN(n24372) );
  AOI222_X1 U23255 ( .A1(n26462), .A2(n25246), .B1(n26456), .B2(n25438), .C1(
        n26450), .C2(n25534), .ZN(n24379) );
  OAI221_X1 U23256 ( .B1(n22015), .B2(n26474), .C1(n27416), .C2(n26468), .A(
        n24361), .ZN(n24354) );
  AOI222_X1 U23257 ( .A1(n26462), .A2(n25247), .B1(n26456), .B2(n25439), .C1(
        n26450), .C2(n25535), .ZN(n24361) );
  OAI221_X1 U23258 ( .B1(n22014), .B2(n26474), .C1(n27419), .C2(n26468), .A(
        n24343), .ZN(n24336) );
  AOI222_X1 U23259 ( .A1(n26462), .A2(n25248), .B1(n26456), .B2(n25440), .C1(
        n26450), .C2(n25536), .ZN(n24343) );
  OAI221_X1 U23260 ( .B1(n22013), .B2(n26474), .C1(n27422), .C2(n26468), .A(
        n24325), .ZN(n24318) );
  AOI222_X1 U23261 ( .A1(n26462), .A2(n25249), .B1(n26456), .B2(n25441), .C1(
        n26450), .C2(n25537), .ZN(n24325) );
  OAI221_X1 U23262 ( .B1(n22012), .B2(n26474), .C1(n27425), .C2(n26468), .A(
        n24307), .ZN(n24300) );
  AOI222_X1 U23263 ( .A1(n26462), .A2(n25250), .B1(n26456), .B2(n25442), .C1(
        n26450), .C2(n25538), .ZN(n24307) );
  OAI221_X1 U23264 ( .B1(n22059), .B2(n26696), .C1(n27284), .C2(n26690), .A(
        n23967), .ZN(n23957) );
  AOI222_X1 U23265 ( .A1(n26684), .A2(n25595), .B1(n26678), .B2(n25619), .C1(
        n26672), .C2(n25667), .ZN(n23967) );
  OAI221_X1 U23266 ( .B1(n22058), .B2(n26696), .C1(n27287), .C2(n26690), .A(
        n23936), .ZN(n23929) );
  AOI222_X1 U23267 ( .A1(n26684), .A2(n25596), .B1(n26678), .B2(n25620), .C1(
        n26672), .C2(n25668), .ZN(n23936) );
  OAI221_X1 U23268 ( .B1(n22057), .B2(n26696), .C1(n27290), .C2(n26690), .A(
        n23918), .ZN(n23911) );
  AOI222_X1 U23269 ( .A1(n26684), .A2(n25597), .B1(n26678), .B2(n25621), .C1(
        n26672), .C2(n25669), .ZN(n23918) );
  OAI221_X1 U23270 ( .B1(n22056), .B2(n26696), .C1(n27293), .C2(n26690), .A(
        n23900), .ZN(n23893) );
  AOI222_X1 U23271 ( .A1(n26684), .A2(n25598), .B1(n26678), .B2(n25622), .C1(
        n26672), .C2(n25670), .ZN(n23900) );
  OAI221_X1 U23272 ( .B1(n22055), .B2(n26696), .C1(n27296), .C2(n26690), .A(
        n23882), .ZN(n23875) );
  AOI222_X1 U23273 ( .A1(n26684), .A2(n25599), .B1(n26678), .B2(n25623), .C1(
        n26672), .C2(n25671), .ZN(n23882) );
  OAI221_X1 U23274 ( .B1(n22054), .B2(n26696), .C1(n27299), .C2(n26690), .A(
        n23864), .ZN(n23857) );
  AOI222_X1 U23275 ( .A1(n26684), .A2(n25600), .B1(n26678), .B2(n25624), .C1(
        n26672), .C2(n25672), .ZN(n23864) );
  OAI221_X1 U23276 ( .B1(n22053), .B2(n26696), .C1(n27302), .C2(n26690), .A(
        n23846), .ZN(n23839) );
  AOI222_X1 U23277 ( .A1(n26684), .A2(n25601), .B1(n26678), .B2(n25625), .C1(
        n26672), .C2(n25673), .ZN(n23846) );
  OAI221_X1 U23278 ( .B1(n22052), .B2(n26696), .C1(n27305), .C2(n26690), .A(
        n23828), .ZN(n23821) );
  AOI222_X1 U23279 ( .A1(n26684), .A2(n25602), .B1(n26678), .B2(n25626), .C1(
        n26672), .C2(n25674), .ZN(n23828) );
  OAI221_X1 U23280 ( .B1(n22051), .B2(n26696), .C1(n27308), .C2(n26690), .A(
        n23810), .ZN(n23803) );
  AOI222_X1 U23281 ( .A1(n26684), .A2(n25603), .B1(n26678), .B2(n25627), .C1(
        n26672), .C2(n25675), .ZN(n23810) );
  OAI221_X1 U23282 ( .B1(n22050), .B2(n26696), .C1(n27311), .C2(n26690), .A(
        n23792), .ZN(n23785) );
  AOI222_X1 U23283 ( .A1(n26684), .A2(n25604), .B1(n26678), .B2(n25628), .C1(
        n26672), .C2(n25676), .ZN(n23792) );
  OAI221_X1 U23284 ( .B1(n22049), .B2(n26696), .C1(n27314), .C2(n26690), .A(
        n23774), .ZN(n23767) );
  AOI222_X1 U23285 ( .A1(n26684), .A2(n25605), .B1(n26678), .B2(n25629), .C1(
        n26672), .C2(n25677), .ZN(n23774) );
  OAI221_X1 U23286 ( .B1(n22048), .B2(n26696), .C1(n27317), .C2(n26690), .A(
        n23756), .ZN(n23749) );
  AOI222_X1 U23287 ( .A1(n26684), .A2(n25606), .B1(n26678), .B2(n25630), .C1(
        n26672), .C2(n25678), .ZN(n23756) );
  OAI221_X1 U23288 ( .B1(n22047), .B2(n26697), .C1(n27320), .C2(n26691), .A(
        n23738), .ZN(n23731) );
  AOI222_X1 U23289 ( .A1(n26685), .A2(n25215), .B1(n26679), .B2(n25407), .C1(
        n26673), .C2(n25503), .ZN(n23738) );
  OAI221_X1 U23290 ( .B1(n22046), .B2(n26697), .C1(n27323), .C2(n26691), .A(
        n23720), .ZN(n23713) );
  AOI222_X1 U23291 ( .A1(n26685), .A2(n25216), .B1(n26679), .B2(n25408), .C1(
        n26673), .C2(n25504), .ZN(n23720) );
  OAI221_X1 U23292 ( .B1(n22045), .B2(n26697), .C1(n27326), .C2(n26691), .A(
        n23702), .ZN(n23695) );
  AOI222_X1 U23293 ( .A1(n26685), .A2(n25217), .B1(n26679), .B2(n25409), .C1(
        n26673), .C2(n25505), .ZN(n23702) );
  OAI221_X1 U23294 ( .B1(n22044), .B2(n26697), .C1(n27329), .C2(n26691), .A(
        n23684), .ZN(n23677) );
  AOI222_X1 U23295 ( .A1(n26685), .A2(n25218), .B1(n26679), .B2(n25410), .C1(
        n26673), .C2(n25506), .ZN(n23684) );
  OAI221_X1 U23296 ( .B1(n22043), .B2(n26697), .C1(n27332), .C2(n26691), .A(
        n23666), .ZN(n23659) );
  AOI222_X1 U23297 ( .A1(n26685), .A2(n25219), .B1(n26679), .B2(n25411), .C1(
        n26673), .C2(n25507), .ZN(n23666) );
  OAI221_X1 U23298 ( .B1(n22042), .B2(n26697), .C1(n27335), .C2(n26691), .A(
        n23648), .ZN(n23641) );
  AOI222_X1 U23299 ( .A1(n26685), .A2(n25220), .B1(n26679), .B2(n25412), .C1(
        n26673), .C2(n25508), .ZN(n23648) );
  OAI221_X1 U23300 ( .B1(n22041), .B2(n26697), .C1(n27338), .C2(n26691), .A(
        n23630), .ZN(n23623) );
  AOI222_X1 U23301 ( .A1(n26685), .A2(n25221), .B1(n26679), .B2(n25413), .C1(
        n26673), .C2(n25509), .ZN(n23630) );
  OAI221_X1 U23302 ( .B1(n22040), .B2(n26697), .C1(n27341), .C2(n26691), .A(
        n23612), .ZN(n23605) );
  AOI222_X1 U23303 ( .A1(n26685), .A2(n25222), .B1(n26679), .B2(n25414), .C1(
        n26673), .C2(n25510), .ZN(n23612) );
  OAI221_X1 U23304 ( .B1(n22039), .B2(n26697), .C1(n27344), .C2(n26691), .A(
        n23594), .ZN(n23587) );
  AOI222_X1 U23305 ( .A1(n26685), .A2(n25223), .B1(n26679), .B2(n25415), .C1(
        n26673), .C2(n25511), .ZN(n23594) );
  OAI221_X1 U23306 ( .B1(n22038), .B2(n26697), .C1(n27347), .C2(n26691), .A(
        n23576), .ZN(n23569) );
  AOI222_X1 U23307 ( .A1(n26685), .A2(n25224), .B1(n26679), .B2(n25416), .C1(
        n26673), .C2(n25512), .ZN(n23576) );
  OAI221_X1 U23308 ( .B1(n22037), .B2(n26697), .C1(n27350), .C2(n26691), .A(
        n23558), .ZN(n23551) );
  AOI222_X1 U23309 ( .A1(n26685), .A2(n25225), .B1(n26679), .B2(n25417), .C1(
        n26673), .C2(n25513), .ZN(n23558) );
  OAI221_X1 U23310 ( .B1(n22036), .B2(n26697), .C1(n27353), .C2(n26691), .A(
        n23540), .ZN(n23533) );
  AOI222_X1 U23311 ( .A1(n26685), .A2(n25226), .B1(n26679), .B2(n25418), .C1(
        n26673), .C2(n25514), .ZN(n23540) );
  OAI221_X1 U23312 ( .B1(n22035), .B2(n26698), .C1(n27356), .C2(n26692), .A(
        n23522), .ZN(n23515) );
  AOI222_X1 U23313 ( .A1(n26686), .A2(n25227), .B1(n26680), .B2(n25419), .C1(
        n26674), .C2(n25515), .ZN(n23522) );
  OAI221_X1 U23314 ( .B1(n22034), .B2(n26698), .C1(n27359), .C2(n26692), .A(
        n23504), .ZN(n23497) );
  AOI222_X1 U23315 ( .A1(n26686), .A2(n25228), .B1(n26680), .B2(n25420), .C1(
        n26674), .C2(n25516), .ZN(n23504) );
  OAI221_X1 U23316 ( .B1(n22033), .B2(n26698), .C1(n27362), .C2(n26692), .A(
        n23486), .ZN(n23479) );
  AOI222_X1 U23317 ( .A1(n26686), .A2(n25229), .B1(n26680), .B2(n25421), .C1(
        n26674), .C2(n25517), .ZN(n23486) );
  OAI221_X1 U23318 ( .B1(n22032), .B2(n26698), .C1(n27365), .C2(n26692), .A(
        n23468), .ZN(n23461) );
  AOI222_X1 U23319 ( .A1(n26686), .A2(n25230), .B1(n26680), .B2(n25422), .C1(
        n26674), .C2(n25518), .ZN(n23468) );
  OAI221_X1 U23320 ( .B1(n22031), .B2(n26698), .C1(n27368), .C2(n26692), .A(
        n23450), .ZN(n23443) );
  AOI222_X1 U23321 ( .A1(n26686), .A2(n25231), .B1(n26680), .B2(n25423), .C1(
        n26674), .C2(n25519), .ZN(n23450) );
  OAI221_X1 U23322 ( .B1(n22030), .B2(n26698), .C1(n27371), .C2(n26692), .A(
        n23432), .ZN(n23425) );
  AOI222_X1 U23323 ( .A1(n26686), .A2(n25232), .B1(n26680), .B2(n25424), .C1(
        n26674), .C2(n25520), .ZN(n23432) );
  OAI221_X1 U23324 ( .B1(n22029), .B2(n26698), .C1(n27374), .C2(n26692), .A(
        n23414), .ZN(n23407) );
  AOI222_X1 U23325 ( .A1(n26686), .A2(n25233), .B1(n26680), .B2(n25425), .C1(
        n26674), .C2(n25521), .ZN(n23414) );
  OAI221_X1 U23326 ( .B1(n22028), .B2(n26698), .C1(n27377), .C2(n26692), .A(
        n23396), .ZN(n23389) );
  AOI222_X1 U23327 ( .A1(n26686), .A2(n25234), .B1(n26680), .B2(n25426), .C1(
        n26674), .C2(n25522), .ZN(n23396) );
  OAI221_X1 U23328 ( .B1(n22027), .B2(n26698), .C1(n27380), .C2(n26692), .A(
        n23378), .ZN(n23371) );
  AOI222_X1 U23329 ( .A1(n26686), .A2(n25235), .B1(n26680), .B2(n25427), .C1(
        n26674), .C2(n25523), .ZN(n23378) );
  OAI221_X1 U23330 ( .B1(n22026), .B2(n26698), .C1(n27383), .C2(n26692), .A(
        n23360), .ZN(n23353) );
  AOI222_X1 U23331 ( .A1(n26686), .A2(n25236), .B1(n26680), .B2(n25428), .C1(
        n26674), .C2(n25524), .ZN(n23360) );
  OAI221_X1 U23332 ( .B1(n22025), .B2(n26698), .C1(n27386), .C2(n26692), .A(
        n23342), .ZN(n23335) );
  AOI222_X1 U23333 ( .A1(n26686), .A2(n25237), .B1(n26680), .B2(n25429), .C1(
        n26674), .C2(n25525), .ZN(n23342) );
  OAI221_X1 U23334 ( .B1(n22024), .B2(n26698), .C1(n27389), .C2(n26692), .A(
        n23324), .ZN(n23317) );
  AOI222_X1 U23335 ( .A1(n26686), .A2(n25238), .B1(n26680), .B2(n25430), .C1(
        n26674), .C2(n25526), .ZN(n23324) );
  OAI221_X1 U23336 ( .B1(n22023), .B2(n26699), .C1(n27392), .C2(n26693), .A(
        n23306), .ZN(n23299) );
  AOI222_X1 U23337 ( .A1(n26687), .A2(n25239), .B1(n26681), .B2(n25431), .C1(
        n26675), .C2(n25527), .ZN(n23306) );
  OAI221_X1 U23338 ( .B1(n22022), .B2(n26699), .C1(n27395), .C2(n26693), .A(
        n23288), .ZN(n23281) );
  AOI222_X1 U23339 ( .A1(n26687), .A2(n25240), .B1(n26681), .B2(n25432), .C1(
        n26675), .C2(n25528), .ZN(n23288) );
  OAI221_X1 U23340 ( .B1(n22021), .B2(n26699), .C1(n27398), .C2(n26693), .A(
        n23270), .ZN(n23263) );
  AOI222_X1 U23341 ( .A1(n26687), .A2(n25241), .B1(n26681), .B2(n25433), .C1(
        n26675), .C2(n25529), .ZN(n23270) );
  OAI221_X1 U23342 ( .B1(n22020), .B2(n26699), .C1(n27401), .C2(n26693), .A(
        n23252), .ZN(n23245) );
  AOI222_X1 U23343 ( .A1(n26687), .A2(n25242), .B1(n26681), .B2(n25434), .C1(
        n26675), .C2(n25530), .ZN(n23252) );
  OAI221_X1 U23344 ( .B1(n22019), .B2(n26699), .C1(n27404), .C2(n26693), .A(
        n23234), .ZN(n23227) );
  AOI222_X1 U23345 ( .A1(n26687), .A2(n25243), .B1(n26681), .B2(n25435), .C1(
        n26675), .C2(n25531), .ZN(n23234) );
  OAI221_X1 U23346 ( .B1(n22018), .B2(n26699), .C1(n27407), .C2(n26693), .A(
        n23216), .ZN(n23209) );
  AOI222_X1 U23347 ( .A1(n26687), .A2(n25244), .B1(n26681), .B2(n25436), .C1(
        n26675), .C2(n25532), .ZN(n23216) );
  OAI221_X1 U23348 ( .B1(n22017), .B2(n26699), .C1(n27410), .C2(n26693), .A(
        n23198), .ZN(n23191) );
  AOI222_X1 U23349 ( .A1(n26687), .A2(n25245), .B1(n26681), .B2(n25437), .C1(
        n26675), .C2(n25533), .ZN(n23198) );
  OAI221_X1 U23350 ( .B1(n22016), .B2(n26699), .C1(n27413), .C2(n26693), .A(
        n23180), .ZN(n23173) );
  AOI222_X1 U23351 ( .A1(n26687), .A2(n25246), .B1(n26681), .B2(n25438), .C1(
        n26675), .C2(n25534), .ZN(n23180) );
  OAI221_X1 U23352 ( .B1(n22015), .B2(n26699), .C1(n27416), .C2(n26693), .A(
        n23162), .ZN(n23155) );
  AOI222_X1 U23353 ( .A1(n26687), .A2(n25247), .B1(n26681), .B2(n25439), .C1(
        n26675), .C2(n25535), .ZN(n23162) );
  OAI221_X1 U23354 ( .B1(n22014), .B2(n26699), .C1(n27419), .C2(n26693), .A(
        n23144), .ZN(n23137) );
  AOI222_X1 U23355 ( .A1(n26687), .A2(n25248), .B1(n26681), .B2(n25440), .C1(
        n26675), .C2(n25536), .ZN(n23144) );
  OAI221_X1 U23356 ( .B1(n22013), .B2(n26699), .C1(n27422), .C2(n26693), .A(
        n23126), .ZN(n23119) );
  AOI222_X1 U23357 ( .A1(n26687), .A2(n25249), .B1(n26681), .B2(n25441), .C1(
        n26675), .C2(n25537), .ZN(n23126) );
  OAI221_X1 U23358 ( .B1(n22012), .B2(n26699), .C1(n27425), .C2(n26693), .A(
        n23108), .ZN(n23101) );
  AOI222_X1 U23359 ( .A1(n26687), .A2(n25250), .B1(n26681), .B2(n25442), .C1(
        n26675), .C2(n25538), .ZN(n23108) );
  OAI221_X1 U23360 ( .B1(n21759), .B2(n26594), .C1(n22379), .C2(n26588), .A(
        n25154), .ZN(n25138) );
  AOI222_X1 U23361 ( .A1(n26582), .A2(n25702), .B1(n26576), .B2(n21094), .C1(
        n26570), .C2(n21154), .ZN(n25154) );
  OAI221_X1 U23362 ( .B1(n21758), .B2(n26594), .C1(n22378), .C2(n26588), .A(
        n25127), .ZN(n25120) );
  AOI222_X1 U23363 ( .A1(n26582), .A2(n25707), .B1(n26576), .B2(n21093), .C1(
        n26570), .C2(n21153), .ZN(n25127) );
  OAI221_X1 U23364 ( .B1(n21757), .B2(n26594), .C1(n22377), .C2(n26588), .A(
        n25109), .ZN(n25102) );
  AOI222_X1 U23365 ( .A1(n26582), .A2(n25712), .B1(n26576), .B2(n21092), .C1(
        n26570), .C2(n21152), .ZN(n25109) );
  OAI221_X1 U23366 ( .B1(n21756), .B2(n26594), .C1(n22376), .C2(n26588), .A(
        n25091), .ZN(n25084) );
  AOI222_X1 U23367 ( .A1(n26582), .A2(n25717), .B1(n26576), .B2(n21091), .C1(
        n26570), .C2(n21151), .ZN(n25091) );
  OAI221_X1 U23368 ( .B1(n21755), .B2(n26594), .C1(n22375), .C2(n26588), .A(
        n25073), .ZN(n25066) );
  AOI222_X1 U23369 ( .A1(n26582), .A2(n25722), .B1(n26576), .B2(n21090), .C1(
        n26570), .C2(n21150), .ZN(n25073) );
  OAI221_X1 U23370 ( .B1(n21754), .B2(n26594), .C1(n22374), .C2(n26588), .A(
        n25055), .ZN(n25048) );
  AOI222_X1 U23371 ( .A1(n26582), .A2(n25727), .B1(n26576), .B2(n21089), .C1(
        n26570), .C2(n21149), .ZN(n25055) );
  OAI221_X1 U23372 ( .B1(n21753), .B2(n26594), .C1(n22373), .C2(n26588), .A(
        n25037), .ZN(n25030) );
  AOI222_X1 U23373 ( .A1(n26582), .A2(n25732), .B1(n26576), .B2(n21088), .C1(
        n26570), .C2(n21148), .ZN(n25037) );
  OAI221_X1 U23374 ( .B1(n21752), .B2(n26594), .C1(n22372), .C2(n26588), .A(
        n25019), .ZN(n25012) );
  AOI222_X1 U23375 ( .A1(n26582), .A2(n25737), .B1(n26576), .B2(n21087), .C1(
        n26570), .C2(n21147), .ZN(n25019) );
  OAI221_X1 U23376 ( .B1(n21751), .B2(n26594), .C1(n22371), .C2(n26588), .A(
        n25001), .ZN(n24994) );
  AOI222_X1 U23377 ( .A1(n26582), .A2(n25742), .B1(n26576), .B2(n21086), .C1(
        n26570), .C2(n21146), .ZN(n25001) );
  OAI221_X1 U23378 ( .B1(n21750), .B2(n26594), .C1(n22370), .C2(n26588), .A(
        n24983), .ZN(n24976) );
  AOI222_X1 U23379 ( .A1(n26582), .A2(n25747), .B1(n26576), .B2(n21085), .C1(
        n26570), .C2(n21145), .ZN(n24983) );
  OAI221_X1 U23380 ( .B1(n21749), .B2(n26594), .C1(n22369), .C2(n26588), .A(
        n24965), .ZN(n24958) );
  AOI222_X1 U23381 ( .A1(n26582), .A2(n25752), .B1(n26576), .B2(n21084), .C1(
        n26570), .C2(n21144), .ZN(n24965) );
  OAI221_X1 U23382 ( .B1(n21748), .B2(n26594), .C1(n22368), .C2(n26588), .A(
        n24947), .ZN(n24940) );
  AOI222_X1 U23383 ( .A1(n26582), .A2(n25757), .B1(n26576), .B2(n21083), .C1(
        n26570), .C2(n21143), .ZN(n24947) );
  OAI221_X1 U23384 ( .B1(n22011), .B2(n26475), .C1(n27428), .C2(n26469), .A(
        n24289), .ZN(n24282) );
  AOI222_X1 U23385 ( .A1(n26463), .A2(n25251), .B1(n26457), .B2(n25443), .C1(
        n26451), .C2(n25539), .ZN(n24289) );
  OAI221_X1 U23386 ( .B1(n22010), .B2(n26475), .C1(n27431), .C2(n26469), .A(
        n24271), .ZN(n24264) );
  AOI222_X1 U23387 ( .A1(n26463), .A2(n25252), .B1(n26457), .B2(n25444), .C1(
        n26451), .C2(n25540), .ZN(n24271) );
  OAI221_X1 U23388 ( .B1(n22009), .B2(n26475), .C1(n27434), .C2(n26469), .A(
        n24253), .ZN(n24246) );
  AOI222_X1 U23389 ( .A1(n26463), .A2(n25253), .B1(n26457), .B2(n25445), .C1(
        n26451), .C2(n25541), .ZN(n24253) );
  OAI221_X1 U23390 ( .B1(n22008), .B2(n26475), .C1(n27437), .C2(n26469), .A(
        n24235), .ZN(n24228) );
  AOI222_X1 U23391 ( .A1(n26463), .A2(n25254), .B1(n26457), .B2(n25446), .C1(
        n26451), .C2(n25542), .ZN(n24235) );
  OAI221_X1 U23392 ( .B1(n22007), .B2(n26475), .C1(n27440), .C2(n26469), .A(
        n24217), .ZN(n24210) );
  AOI222_X1 U23393 ( .A1(n26463), .A2(n25255), .B1(n26457), .B2(n25447), .C1(
        n26451), .C2(n25543), .ZN(n24217) );
  OAI221_X1 U23394 ( .B1(n22006), .B2(n26475), .C1(n27443), .C2(n26469), .A(
        n24199), .ZN(n24192) );
  AOI222_X1 U23395 ( .A1(n26463), .A2(n25256), .B1(n26457), .B2(n25448), .C1(
        n26451), .C2(n25544), .ZN(n24199) );
  OAI221_X1 U23396 ( .B1(n22005), .B2(n26475), .C1(n27446), .C2(n26469), .A(
        n24181), .ZN(n24174) );
  AOI222_X1 U23397 ( .A1(n26463), .A2(n25257), .B1(n26457), .B2(n25449), .C1(
        n26451), .C2(n25545), .ZN(n24181) );
  OAI221_X1 U23398 ( .B1(n22004), .B2(n26475), .C1(n27449), .C2(n26469), .A(
        n24163), .ZN(n24156) );
  AOI222_X1 U23399 ( .A1(n26463), .A2(n25258), .B1(n26457), .B2(n25450), .C1(
        n26451), .C2(n25546), .ZN(n24163) );
  OAI221_X1 U23400 ( .B1(n22003), .B2(n26475), .C1(n27452), .C2(n26469), .A(
        n24145), .ZN(n24138) );
  AOI222_X1 U23401 ( .A1(n26463), .A2(n25259), .B1(n26457), .B2(n25451), .C1(
        n26451), .C2(n25547), .ZN(n24145) );
  OAI221_X1 U23402 ( .B1(n22002), .B2(n26475), .C1(n27455), .C2(n26469), .A(
        n24127), .ZN(n24120) );
  AOI222_X1 U23403 ( .A1(n26463), .A2(n25260), .B1(n26457), .B2(n25452), .C1(
        n26451), .C2(n25548), .ZN(n24127) );
  OAI221_X1 U23404 ( .B1(n22001), .B2(n26475), .C1(n27458), .C2(n26469), .A(
        n24109), .ZN(n24102) );
  AOI222_X1 U23405 ( .A1(n26463), .A2(n25261), .B1(n26457), .B2(n25453), .C1(
        n26451), .C2(n25549), .ZN(n24109) );
  OAI221_X1 U23406 ( .B1(n22000), .B2(n26475), .C1(n27461), .C2(n26469), .A(
        n24091), .ZN(n24084) );
  AOI222_X1 U23407 ( .A1(n26463), .A2(n25262), .B1(n26457), .B2(n25454), .C1(
        n26451), .C2(n25550), .ZN(n24091) );
  OAI221_X1 U23408 ( .B1(n21759), .B2(n26819), .C1(n22379), .C2(n26813), .A(
        n23955), .ZN(n23939) );
  AOI222_X1 U23409 ( .A1(n26807), .A2(n25702), .B1(n26801), .B2(n21094), .C1(
        n26795), .C2(n21154), .ZN(n23955) );
  OAI221_X1 U23410 ( .B1(n21758), .B2(n26819), .C1(n22378), .C2(n26813), .A(
        n23928), .ZN(n23921) );
  AOI222_X1 U23411 ( .A1(n26807), .A2(n25707), .B1(n26801), .B2(n21093), .C1(
        n26795), .C2(n21153), .ZN(n23928) );
  OAI221_X1 U23412 ( .B1(n21757), .B2(n26819), .C1(n22377), .C2(n26813), .A(
        n23910), .ZN(n23903) );
  AOI222_X1 U23413 ( .A1(n26807), .A2(n25712), .B1(n26801), .B2(n21092), .C1(
        n26795), .C2(n21152), .ZN(n23910) );
  OAI221_X1 U23414 ( .B1(n21756), .B2(n26819), .C1(n22376), .C2(n26813), .A(
        n23892), .ZN(n23885) );
  AOI222_X1 U23415 ( .A1(n26807), .A2(n25717), .B1(n26801), .B2(n21091), .C1(
        n26795), .C2(n21151), .ZN(n23892) );
  OAI221_X1 U23416 ( .B1(n21755), .B2(n26819), .C1(n22375), .C2(n26813), .A(
        n23874), .ZN(n23867) );
  AOI222_X1 U23417 ( .A1(n26807), .A2(n25722), .B1(n26801), .B2(n21090), .C1(
        n26795), .C2(n21150), .ZN(n23874) );
  OAI221_X1 U23418 ( .B1(n21754), .B2(n26819), .C1(n22374), .C2(n26813), .A(
        n23856), .ZN(n23849) );
  AOI222_X1 U23419 ( .A1(n26807), .A2(n25727), .B1(n26801), .B2(n21089), .C1(
        n26795), .C2(n21149), .ZN(n23856) );
  OAI221_X1 U23420 ( .B1(n21753), .B2(n26819), .C1(n22373), .C2(n26813), .A(
        n23838), .ZN(n23831) );
  AOI222_X1 U23421 ( .A1(n26807), .A2(n25732), .B1(n26801), .B2(n21088), .C1(
        n26795), .C2(n21148), .ZN(n23838) );
  OAI221_X1 U23422 ( .B1(n21752), .B2(n26819), .C1(n22372), .C2(n26813), .A(
        n23820), .ZN(n23813) );
  AOI222_X1 U23423 ( .A1(n26807), .A2(n25737), .B1(n26801), .B2(n21087), .C1(
        n26795), .C2(n21147), .ZN(n23820) );
  OAI221_X1 U23424 ( .B1(n21751), .B2(n26819), .C1(n22371), .C2(n26813), .A(
        n23802), .ZN(n23795) );
  AOI222_X1 U23425 ( .A1(n26807), .A2(n25742), .B1(n26801), .B2(n21086), .C1(
        n26795), .C2(n21146), .ZN(n23802) );
  OAI221_X1 U23426 ( .B1(n21750), .B2(n26819), .C1(n22370), .C2(n26813), .A(
        n23784), .ZN(n23777) );
  AOI222_X1 U23427 ( .A1(n26807), .A2(n25747), .B1(n26801), .B2(n21085), .C1(
        n26795), .C2(n21145), .ZN(n23784) );
  OAI221_X1 U23428 ( .B1(n21749), .B2(n26819), .C1(n22369), .C2(n26813), .A(
        n23766), .ZN(n23759) );
  AOI222_X1 U23429 ( .A1(n26807), .A2(n25752), .B1(n26801), .B2(n21084), .C1(
        n26795), .C2(n21144), .ZN(n23766) );
  OAI221_X1 U23430 ( .B1(n21748), .B2(n26819), .C1(n22368), .C2(n26813), .A(
        n23748), .ZN(n23741) );
  AOI222_X1 U23431 ( .A1(n26807), .A2(n25757), .B1(n26801), .B2(n21083), .C1(
        n26795), .C2(n21143), .ZN(n23748) );
  OAI221_X1 U23432 ( .B1(n22011), .B2(n26700), .C1(n27428), .C2(n26694), .A(
        n23090), .ZN(n23083) );
  AOI222_X1 U23433 ( .A1(n26688), .A2(n25251), .B1(n26682), .B2(n25443), .C1(
        n26676), .C2(n25539), .ZN(n23090) );
  OAI221_X1 U23434 ( .B1(n22010), .B2(n26700), .C1(n27431), .C2(n26694), .A(
        n23072), .ZN(n23065) );
  AOI222_X1 U23435 ( .A1(n26688), .A2(n25252), .B1(n26682), .B2(n25444), .C1(
        n26676), .C2(n25540), .ZN(n23072) );
  OAI221_X1 U23436 ( .B1(n22009), .B2(n26700), .C1(n27434), .C2(n26694), .A(
        n23054), .ZN(n23047) );
  AOI222_X1 U23437 ( .A1(n26688), .A2(n25253), .B1(n26682), .B2(n25445), .C1(
        n26676), .C2(n25541), .ZN(n23054) );
  OAI221_X1 U23438 ( .B1(n22008), .B2(n26700), .C1(n27437), .C2(n26694), .A(
        n23036), .ZN(n23029) );
  AOI222_X1 U23439 ( .A1(n26688), .A2(n25254), .B1(n26682), .B2(n25446), .C1(
        n26676), .C2(n25542), .ZN(n23036) );
  OAI221_X1 U23440 ( .B1(n22007), .B2(n26700), .C1(n27440), .C2(n26694), .A(
        n23018), .ZN(n23011) );
  AOI222_X1 U23441 ( .A1(n26688), .A2(n25255), .B1(n26682), .B2(n25447), .C1(
        n26676), .C2(n25543), .ZN(n23018) );
  OAI221_X1 U23442 ( .B1(n22006), .B2(n26700), .C1(n27443), .C2(n26694), .A(
        n23000), .ZN(n22993) );
  AOI222_X1 U23443 ( .A1(n26688), .A2(n25256), .B1(n26682), .B2(n25448), .C1(
        n26676), .C2(n25544), .ZN(n23000) );
  OAI221_X1 U23444 ( .B1(n22005), .B2(n26700), .C1(n27446), .C2(n26694), .A(
        n22982), .ZN(n22975) );
  AOI222_X1 U23445 ( .A1(n26688), .A2(n25257), .B1(n26682), .B2(n25449), .C1(
        n26676), .C2(n25545), .ZN(n22982) );
  OAI221_X1 U23446 ( .B1(n22004), .B2(n26700), .C1(n27449), .C2(n26694), .A(
        n22964), .ZN(n22957) );
  AOI222_X1 U23447 ( .A1(n26688), .A2(n25258), .B1(n26682), .B2(n25450), .C1(
        n26676), .C2(n25546), .ZN(n22964) );
  OAI221_X1 U23448 ( .B1(n22003), .B2(n26700), .C1(n27452), .C2(n26694), .A(
        n22946), .ZN(n22939) );
  AOI222_X1 U23449 ( .A1(n26688), .A2(n25259), .B1(n26682), .B2(n25451), .C1(
        n26676), .C2(n25547), .ZN(n22946) );
  OAI221_X1 U23450 ( .B1(n22002), .B2(n26700), .C1(n27455), .C2(n26694), .A(
        n22928), .ZN(n22921) );
  AOI222_X1 U23451 ( .A1(n26688), .A2(n25260), .B1(n26682), .B2(n25452), .C1(
        n26676), .C2(n25548), .ZN(n22928) );
  OAI221_X1 U23452 ( .B1(n22001), .B2(n26700), .C1(n27458), .C2(n26694), .A(
        n22910), .ZN(n22903) );
  AOI222_X1 U23453 ( .A1(n26688), .A2(n25261), .B1(n26682), .B2(n25453), .C1(
        n26676), .C2(n25549), .ZN(n22910) );
  OAI221_X1 U23454 ( .B1(n22000), .B2(n26700), .C1(n27461), .C2(n26694), .A(
        n22892), .ZN(n22885) );
  AOI222_X1 U23455 ( .A1(n26688), .A2(n25262), .B1(n26682), .B2(n25454), .C1(
        n26676), .C2(n25550), .ZN(n22892) );
  OAI22_X1 U23456 ( .A1(n27320), .A2(n26952), .B1(n26946), .B2(n22619), .ZN(
        n6286) );
  OAI22_X1 U23457 ( .A1(n27323), .A2(n26952), .B1(n26946), .B2(n22618), .ZN(
        n6287) );
  OAI22_X1 U23458 ( .A1(n27326), .A2(n26952), .B1(n26946), .B2(n22617), .ZN(
        n6288) );
  OAI22_X1 U23459 ( .A1(n27329), .A2(n26952), .B1(n26946), .B2(n22616), .ZN(
        n6289) );
  OAI22_X1 U23460 ( .A1(n27332), .A2(n26952), .B1(n26946), .B2(n22615), .ZN(
        n6290) );
  OAI22_X1 U23461 ( .A1(n27335), .A2(n26952), .B1(n26946), .B2(n22614), .ZN(
        n6291) );
  OAI22_X1 U23462 ( .A1(n27338), .A2(n26952), .B1(n26946), .B2(n22613), .ZN(
        n6292) );
  OAI22_X1 U23463 ( .A1(n27341), .A2(n26952), .B1(n26946), .B2(n22612), .ZN(
        n6293) );
  OAI22_X1 U23464 ( .A1(n27344), .A2(n26952), .B1(n26946), .B2(n22611), .ZN(
        n6294) );
  OAI22_X1 U23465 ( .A1(n27347), .A2(n26952), .B1(n26946), .B2(n22610), .ZN(
        n6295) );
  OAI22_X1 U23466 ( .A1(n27350), .A2(n26952), .B1(n26946), .B2(n22609), .ZN(
        n6296) );
  OAI22_X1 U23467 ( .A1(n27353), .A2(n26953), .B1(n26946), .B2(n22608), .ZN(
        n6297) );
  OAI22_X1 U23468 ( .A1(n27356), .A2(n26953), .B1(n26947), .B2(n22607), .ZN(
        n6298) );
  OAI22_X1 U23469 ( .A1(n27359), .A2(n26953), .B1(n26947), .B2(n22606), .ZN(
        n6299) );
  OAI22_X1 U23470 ( .A1(n27362), .A2(n26953), .B1(n26947), .B2(n22605), .ZN(
        n6300) );
  OAI22_X1 U23471 ( .A1(n27365), .A2(n26953), .B1(n26947), .B2(n22604), .ZN(
        n6301) );
  OAI22_X1 U23472 ( .A1(n27368), .A2(n26953), .B1(n26947), .B2(n22603), .ZN(
        n6302) );
  OAI22_X1 U23473 ( .A1(n27371), .A2(n26953), .B1(n26947), .B2(n22602), .ZN(
        n6303) );
  OAI22_X1 U23474 ( .A1(n27374), .A2(n26953), .B1(n26947), .B2(n22601), .ZN(
        n6304) );
  OAI22_X1 U23475 ( .A1(n27377), .A2(n26953), .B1(n26947), .B2(n22600), .ZN(
        n6305) );
  OAI22_X1 U23476 ( .A1(n27380), .A2(n26953), .B1(n26947), .B2(n22599), .ZN(
        n6306) );
  OAI22_X1 U23477 ( .A1(n27383), .A2(n26953), .B1(n26947), .B2(n22598), .ZN(
        n6307) );
  OAI22_X1 U23478 ( .A1(n27386), .A2(n26953), .B1(n26947), .B2(n22597), .ZN(
        n6308) );
  OAI22_X1 U23479 ( .A1(n27389), .A2(n26954), .B1(n26947), .B2(n22596), .ZN(
        n6309) );
  OAI22_X1 U23480 ( .A1(n27392), .A2(n26954), .B1(n26948), .B2(n22595), .ZN(
        n6310) );
  OAI22_X1 U23481 ( .A1(n27395), .A2(n26954), .B1(n26948), .B2(n22594), .ZN(
        n6311) );
  OAI22_X1 U23482 ( .A1(n27398), .A2(n26954), .B1(n26948), .B2(n22593), .ZN(
        n6312) );
  OAI22_X1 U23483 ( .A1(n27401), .A2(n26954), .B1(n26948), .B2(n22592), .ZN(
        n6313) );
  OAI22_X1 U23484 ( .A1(n27404), .A2(n26954), .B1(n26948), .B2(n22591), .ZN(
        n6314) );
  OAI22_X1 U23485 ( .A1(n27407), .A2(n26954), .B1(n26948), .B2(n22590), .ZN(
        n6315) );
  OAI22_X1 U23486 ( .A1(n27410), .A2(n26954), .B1(n26948), .B2(n22589), .ZN(
        n6316) );
  OAI22_X1 U23487 ( .A1(n27413), .A2(n26954), .B1(n26948), .B2(n22588), .ZN(
        n6317) );
  OAI22_X1 U23488 ( .A1(n27416), .A2(n26954), .B1(n26948), .B2(n22587), .ZN(
        n6318) );
  OAI22_X1 U23489 ( .A1(n27419), .A2(n26954), .B1(n26948), .B2(n22586), .ZN(
        n6319) );
  OAI22_X1 U23490 ( .A1(n27422), .A2(n26954), .B1(n26948), .B2(n22585), .ZN(
        n6320) );
  OAI22_X1 U23491 ( .A1(n27425), .A2(n26955), .B1(n26948), .B2(n22584), .ZN(
        n6321) );
  OAI22_X1 U23492 ( .A1(n27428), .A2(n26955), .B1(n26949), .B2(n22583), .ZN(
        n6322) );
  OAI22_X1 U23493 ( .A1(n27431), .A2(n26955), .B1(n26949), .B2(n22582), .ZN(
        n6323) );
  OAI22_X1 U23494 ( .A1(n27434), .A2(n26955), .B1(n26949), .B2(n22581), .ZN(
        n6324) );
  OAI22_X1 U23495 ( .A1(n27437), .A2(n26955), .B1(n26949), .B2(n22580), .ZN(
        n6325) );
  OAI22_X1 U23496 ( .A1(n27440), .A2(n26955), .B1(n26949), .B2(n22579), .ZN(
        n6326) );
  OAI22_X1 U23497 ( .A1(n27443), .A2(n26955), .B1(n26949), .B2(n22578), .ZN(
        n6327) );
  OAI22_X1 U23498 ( .A1(n27446), .A2(n26955), .B1(n26949), .B2(n22577), .ZN(
        n6328) );
  OAI22_X1 U23499 ( .A1(n27449), .A2(n26955), .B1(n26949), .B2(n22576), .ZN(
        n6329) );
  OAI22_X1 U23500 ( .A1(n27452), .A2(n26955), .B1(n26949), .B2(n22575), .ZN(
        n6330) );
  OAI22_X1 U23501 ( .A1(n27455), .A2(n26955), .B1(n26949), .B2(n22574), .ZN(
        n6331) );
  OAI22_X1 U23502 ( .A1(n27458), .A2(n26955), .B1(n26949), .B2(n22573), .ZN(
        n6332) );
  OAI22_X1 U23503 ( .A1(n27461), .A2(n26956), .B1(n26949), .B2(n22572), .ZN(
        n6333) );
  OAI22_X1 U23504 ( .A1(n27318), .A2(n27156), .B1(n27150), .B2(n22427), .ZN(
        n7374) );
  OAI22_X1 U23505 ( .A1(n27321), .A2(n27156), .B1(n27150), .B2(n22426), .ZN(
        n7375) );
  OAI22_X1 U23506 ( .A1(n27324), .A2(n27156), .B1(n27150), .B2(n22425), .ZN(
        n7376) );
  OAI22_X1 U23507 ( .A1(n27327), .A2(n27156), .B1(n27150), .B2(n22424), .ZN(
        n7377) );
  OAI22_X1 U23508 ( .A1(n27330), .A2(n27156), .B1(n27150), .B2(n22423), .ZN(
        n7378) );
  OAI22_X1 U23509 ( .A1(n27333), .A2(n27156), .B1(n27150), .B2(n22422), .ZN(
        n7379) );
  OAI22_X1 U23510 ( .A1(n27336), .A2(n27156), .B1(n27150), .B2(n22421), .ZN(
        n7380) );
  OAI22_X1 U23511 ( .A1(n27339), .A2(n27156), .B1(n27150), .B2(n22420), .ZN(
        n7381) );
  OAI22_X1 U23512 ( .A1(n27342), .A2(n27156), .B1(n27150), .B2(n22419), .ZN(
        n7382) );
  OAI22_X1 U23513 ( .A1(n27345), .A2(n27156), .B1(n27150), .B2(n22418), .ZN(
        n7383) );
  OAI22_X1 U23514 ( .A1(n27348), .A2(n27156), .B1(n27150), .B2(n22417), .ZN(
        n7384) );
  OAI22_X1 U23515 ( .A1(n27351), .A2(n27157), .B1(n27150), .B2(n22416), .ZN(
        n7385) );
  OAI22_X1 U23516 ( .A1(n27354), .A2(n27157), .B1(n27151), .B2(n22415), .ZN(
        n7386) );
  OAI22_X1 U23517 ( .A1(n27357), .A2(n27157), .B1(n27151), .B2(n22414), .ZN(
        n7387) );
  OAI22_X1 U23518 ( .A1(n27360), .A2(n27157), .B1(n27151), .B2(n22413), .ZN(
        n7388) );
  OAI22_X1 U23519 ( .A1(n27363), .A2(n27157), .B1(n27151), .B2(n22412), .ZN(
        n7389) );
  OAI22_X1 U23520 ( .A1(n27366), .A2(n27157), .B1(n27151), .B2(n22411), .ZN(
        n7390) );
  OAI22_X1 U23521 ( .A1(n27369), .A2(n27157), .B1(n27151), .B2(n22410), .ZN(
        n7391) );
  OAI22_X1 U23522 ( .A1(n27372), .A2(n27157), .B1(n27151), .B2(n22409), .ZN(
        n7392) );
  OAI22_X1 U23523 ( .A1(n27375), .A2(n27157), .B1(n27151), .B2(n22408), .ZN(
        n7393) );
  OAI22_X1 U23524 ( .A1(n27378), .A2(n27157), .B1(n27151), .B2(n22407), .ZN(
        n7394) );
  OAI22_X1 U23525 ( .A1(n27381), .A2(n27157), .B1(n27151), .B2(n22406), .ZN(
        n7395) );
  OAI22_X1 U23526 ( .A1(n27384), .A2(n27157), .B1(n27151), .B2(n22405), .ZN(
        n7396) );
  OAI22_X1 U23527 ( .A1(n27387), .A2(n27158), .B1(n27151), .B2(n22404), .ZN(
        n7397) );
  OAI22_X1 U23528 ( .A1(n27390), .A2(n27158), .B1(n27152), .B2(n22403), .ZN(
        n7398) );
  OAI22_X1 U23529 ( .A1(n27393), .A2(n27158), .B1(n27152), .B2(n22402), .ZN(
        n7399) );
  OAI22_X1 U23530 ( .A1(n27396), .A2(n27158), .B1(n27152), .B2(n22401), .ZN(
        n7400) );
  OAI22_X1 U23531 ( .A1(n27399), .A2(n27158), .B1(n27152), .B2(n22400), .ZN(
        n7401) );
  OAI22_X1 U23532 ( .A1(n27402), .A2(n27158), .B1(n27152), .B2(n22399), .ZN(
        n7402) );
  OAI22_X1 U23533 ( .A1(n27405), .A2(n27158), .B1(n27152), .B2(n22398), .ZN(
        n7403) );
  OAI22_X1 U23534 ( .A1(n27408), .A2(n27158), .B1(n27152), .B2(n22397), .ZN(
        n7404) );
  OAI22_X1 U23535 ( .A1(n27411), .A2(n27158), .B1(n27152), .B2(n22396), .ZN(
        n7405) );
  OAI22_X1 U23536 ( .A1(n27414), .A2(n27158), .B1(n27152), .B2(n22395), .ZN(
        n7406) );
  OAI22_X1 U23537 ( .A1(n27417), .A2(n27158), .B1(n27152), .B2(n22394), .ZN(
        n7407) );
  OAI22_X1 U23538 ( .A1(n27420), .A2(n27158), .B1(n27152), .B2(n22393), .ZN(
        n7408) );
  OAI22_X1 U23539 ( .A1(n27423), .A2(n27159), .B1(n27152), .B2(n22392), .ZN(
        n7409) );
  OAI22_X1 U23540 ( .A1(n27426), .A2(n27159), .B1(n27153), .B2(n22391), .ZN(
        n7410) );
  OAI22_X1 U23541 ( .A1(n27429), .A2(n27159), .B1(n27153), .B2(n22390), .ZN(
        n7411) );
  OAI22_X1 U23542 ( .A1(n27432), .A2(n27159), .B1(n27153), .B2(n22389), .ZN(
        n7412) );
  OAI22_X1 U23543 ( .A1(n27435), .A2(n27159), .B1(n27153), .B2(n22388), .ZN(
        n7413) );
  OAI22_X1 U23544 ( .A1(n27438), .A2(n27159), .B1(n27153), .B2(n22387), .ZN(
        n7414) );
  OAI22_X1 U23545 ( .A1(n27441), .A2(n27159), .B1(n27153), .B2(n22386), .ZN(
        n7415) );
  OAI22_X1 U23546 ( .A1(n27444), .A2(n27159), .B1(n27153), .B2(n22385), .ZN(
        n7416) );
  OAI22_X1 U23547 ( .A1(n27447), .A2(n27159), .B1(n27153), .B2(n22384), .ZN(
        n7417) );
  OAI22_X1 U23548 ( .A1(n27450), .A2(n27159), .B1(n27153), .B2(n22383), .ZN(
        n7418) );
  OAI22_X1 U23549 ( .A1(n27453), .A2(n27159), .B1(n27153), .B2(n22382), .ZN(
        n7419) );
  OAI22_X1 U23550 ( .A1(n27456), .A2(n27159), .B1(n27153), .B2(n22381), .ZN(
        n7420) );
  OAI22_X1 U23551 ( .A1(n27459), .A2(n27160), .B1(n27153), .B2(n22380), .ZN(
        n7421) );
  OAI22_X1 U23552 ( .A1(n27320), .A2(n26928), .B1(n26922), .B2(n22307), .ZN(
        n6158) );
  OAI22_X1 U23553 ( .A1(n27323), .A2(n26928), .B1(n26922), .B2(n22306), .ZN(
        n6159) );
  OAI22_X1 U23554 ( .A1(n27326), .A2(n26928), .B1(n26922), .B2(n22305), .ZN(
        n6160) );
  OAI22_X1 U23555 ( .A1(n27329), .A2(n26928), .B1(n26922), .B2(n22304), .ZN(
        n6161) );
  OAI22_X1 U23556 ( .A1(n27332), .A2(n26928), .B1(n26922), .B2(n22303), .ZN(
        n6162) );
  OAI22_X1 U23557 ( .A1(n27335), .A2(n26928), .B1(n26922), .B2(n22302), .ZN(
        n6163) );
  OAI22_X1 U23558 ( .A1(n27338), .A2(n26928), .B1(n26922), .B2(n22301), .ZN(
        n6164) );
  OAI22_X1 U23559 ( .A1(n27341), .A2(n26928), .B1(n26922), .B2(n22300), .ZN(
        n6165) );
  OAI22_X1 U23560 ( .A1(n27344), .A2(n26928), .B1(n26922), .B2(n22299), .ZN(
        n6166) );
  OAI22_X1 U23561 ( .A1(n27347), .A2(n26928), .B1(n26922), .B2(n22298), .ZN(
        n6167) );
  OAI22_X1 U23562 ( .A1(n27350), .A2(n26928), .B1(n26922), .B2(n22297), .ZN(
        n6168) );
  OAI22_X1 U23563 ( .A1(n27353), .A2(n26929), .B1(n26922), .B2(n22296), .ZN(
        n6169) );
  OAI22_X1 U23564 ( .A1(n27356), .A2(n26929), .B1(n26923), .B2(n22295), .ZN(
        n6170) );
  OAI22_X1 U23565 ( .A1(n27359), .A2(n26929), .B1(n26923), .B2(n22294), .ZN(
        n6171) );
  OAI22_X1 U23566 ( .A1(n27362), .A2(n26929), .B1(n26923), .B2(n22293), .ZN(
        n6172) );
  OAI22_X1 U23567 ( .A1(n27365), .A2(n26929), .B1(n26923), .B2(n22292), .ZN(
        n6173) );
  OAI22_X1 U23568 ( .A1(n27368), .A2(n26929), .B1(n26923), .B2(n22291), .ZN(
        n6174) );
  OAI22_X1 U23569 ( .A1(n27371), .A2(n26929), .B1(n26923), .B2(n22290), .ZN(
        n6175) );
  OAI22_X1 U23570 ( .A1(n27374), .A2(n26929), .B1(n26923), .B2(n22289), .ZN(
        n6176) );
  OAI22_X1 U23571 ( .A1(n27377), .A2(n26929), .B1(n26923), .B2(n22288), .ZN(
        n6177) );
  OAI22_X1 U23572 ( .A1(n27380), .A2(n26929), .B1(n26923), .B2(n22287), .ZN(
        n6178) );
  OAI22_X1 U23573 ( .A1(n27383), .A2(n26929), .B1(n26923), .B2(n22286), .ZN(
        n6179) );
  OAI22_X1 U23574 ( .A1(n27386), .A2(n26929), .B1(n26923), .B2(n22285), .ZN(
        n6180) );
  OAI22_X1 U23575 ( .A1(n27389), .A2(n26930), .B1(n26923), .B2(n22284), .ZN(
        n6181) );
  OAI22_X1 U23576 ( .A1(n27392), .A2(n26930), .B1(n26924), .B2(n22283), .ZN(
        n6182) );
  OAI22_X1 U23577 ( .A1(n27395), .A2(n26930), .B1(n26924), .B2(n22282), .ZN(
        n6183) );
  OAI22_X1 U23578 ( .A1(n27398), .A2(n26930), .B1(n26924), .B2(n22281), .ZN(
        n6184) );
  OAI22_X1 U23579 ( .A1(n27401), .A2(n26930), .B1(n26924), .B2(n22280), .ZN(
        n6185) );
  OAI22_X1 U23580 ( .A1(n27404), .A2(n26930), .B1(n26924), .B2(n22279), .ZN(
        n6186) );
  OAI22_X1 U23581 ( .A1(n27407), .A2(n26930), .B1(n26924), .B2(n22278), .ZN(
        n6187) );
  OAI22_X1 U23582 ( .A1(n27410), .A2(n26930), .B1(n26924), .B2(n22277), .ZN(
        n6188) );
  OAI22_X1 U23583 ( .A1(n27413), .A2(n26930), .B1(n26924), .B2(n22276), .ZN(
        n6189) );
  OAI22_X1 U23584 ( .A1(n27416), .A2(n26930), .B1(n26924), .B2(n22275), .ZN(
        n6190) );
  OAI22_X1 U23585 ( .A1(n27419), .A2(n26930), .B1(n26924), .B2(n22274), .ZN(
        n6191) );
  OAI22_X1 U23586 ( .A1(n27422), .A2(n26930), .B1(n26924), .B2(n22273), .ZN(
        n6192) );
  OAI22_X1 U23587 ( .A1(n27425), .A2(n26931), .B1(n26924), .B2(n22272), .ZN(
        n6193) );
  OAI22_X1 U23588 ( .A1(n27428), .A2(n26931), .B1(n26925), .B2(n22271), .ZN(
        n6194) );
  OAI22_X1 U23589 ( .A1(n27431), .A2(n26931), .B1(n26925), .B2(n22270), .ZN(
        n6195) );
  OAI22_X1 U23590 ( .A1(n27434), .A2(n26931), .B1(n26925), .B2(n22269), .ZN(
        n6196) );
  OAI22_X1 U23591 ( .A1(n27437), .A2(n26931), .B1(n26925), .B2(n22268), .ZN(
        n6197) );
  OAI22_X1 U23592 ( .A1(n27440), .A2(n26931), .B1(n26925), .B2(n22267), .ZN(
        n6198) );
  OAI22_X1 U23593 ( .A1(n27443), .A2(n26931), .B1(n26925), .B2(n22266), .ZN(
        n6199) );
  OAI22_X1 U23594 ( .A1(n27446), .A2(n26931), .B1(n26925), .B2(n22265), .ZN(
        n6200) );
  OAI22_X1 U23595 ( .A1(n27449), .A2(n26931), .B1(n26925), .B2(n22264), .ZN(
        n6201) );
  OAI22_X1 U23596 ( .A1(n27452), .A2(n26931), .B1(n26925), .B2(n22263), .ZN(
        n6202) );
  OAI22_X1 U23597 ( .A1(n27455), .A2(n26931), .B1(n26925), .B2(n22262), .ZN(
        n6203) );
  OAI22_X1 U23598 ( .A1(n27458), .A2(n26931), .B1(n26925), .B2(n22261), .ZN(
        n6204) );
  OAI22_X1 U23599 ( .A1(n27461), .A2(n26932), .B1(n26925), .B2(n22260), .ZN(
        n6205) );
  OAI22_X1 U23600 ( .A1(n27320), .A2(n26940), .B1(n26934), .B2(n22231), .ZN(
        n6222) );
  OAI22_X1 U23601 ( .A1(n27323), .A2(n26940), .B1(n26934), .B2(n22230), .ZN(
        n6223) );
  OAI22_X1 U23602 ( .A1(n27326), .A2(n26940), .B1(n26934), .B2(n22229), .ZN(
        n6224) );
  OAI22_X1 U23603 ( .A1(n27329), .A2(n26940), .B1(n26934), .B2(n22228), .ZN(
        n6225) );
  OAI22_X1 U23604 ( .A1(n27332), .A2(n26940), .B1(n26934), .B2(n22227), .ZN(
        n6226) );
  OAI22_X1 U23605 ( .A1(n27335), .A2(n26940), .B1(n26934), .B2(n22226), .ZN(
        n6227) );
  OAI22_X1 U23606 ( .A1(n27338), .A2(n26940), .B1(n26934), .B2(n22225), .ZN(
        n6228) );
  OAI22_X1 U23607 ( .A1(n27341), .A2(n26940), .B1(n26934), .B2(n22224), .ZN(
        n6229) );
  OAI22_X1 U23608 ( .A1(n27344), .A2(n26940), .B1(n26934), .B2(n22223), .ZN(
        n6230) );
  OAI22_X1 U23609 ( .A1(n27347), .A2(n26940), .B1(n26934), .B2(n22222), .ZN(
        n6231) );
  OAI22_X1 U23610 ( .A1(n27350), .A2(n26940), .B1(n26934), .B2(n22221), .ZN(
        n6232) );
  OAI22_X1 U23611 ( .A1(n27353), .A2(n26941), .B1(n26934), .B2(n22220), .ZN(
        n6233) );
  OAI22_X1 U23612 ( .A1(n27356), .A2(n26941), .B1(n26935), .B2(n22219), .ZN(
        n6234) );
  OAI22_X1 U23613 ( .A1(n27359), .A2(n26941), .B1(n26935), .B2(n22218), .ZN(
        n6235) );
  OAI22_X1 U23614 ( .A1(n27362), .A2(n26941), .B1(n26935), .B2(n22217), .ZN(
        n6236) );
  OAI22_X1 U23615 ( .A1(n27365), .A2(n26941), .B1(n26935), .B2(n22216), .ZN(
        n6237) );
  OAI22_X1 U23616 ( .A1(n27368), .A2(n26941), .B1(n26935), .B2(n22215), .ZN(
        n6238) );
  OAI22_X1 U23617 ( .A1(n27371), .A2(n26941), .B1(n26935), .B2(n22214), .ZN(
        n6239) );
  OAI22_X1 U23618 ( .A1(n27374), .A2(n26941), .B1(n26935), .B2(n22213), .ZN(
        n6240) );
  OAI22_X1 U23619 ( .A1(n27377), .A2(n26941), .B1(n26935), .B2(n22212), .ZN(
        n6241) );
  OAI22_X1 U23620 ( .A1(n27380), .A2(n26941), .B1(n26935), .B2(n22211), .ZN(
        n6242) );
  OAI22_X1 U23621 ( .A1(n27383), .A2(n26941), .B1(n26935), .B2(n22210), .ZN(
        n6243) );
  OAI22_X1 U23622 ( .A1(n27386), .A2(n26941), .B1(n26935), .B2(n22209), .ZN(
        n6244) );
  OAI22_X1 U23623 ( .A1(n27389), .A2(n26942), .B1(n26935), .B2(n22208), .ZN(
        n6245) );
  OAI22_X1 U23624 ( .A1(n27392), .A2(n26942), .B1(n26936), .B2(n22207), .ZN(
        n6246) );
  OAI22_X1 U23625 ( .A1(n27395), .A2(n26942), .B1(n26936), .B2(n22206), .ZN(
        n6247) );
  OAI22_X1 U23626 ( .A1(n27398), .A2(n26942), .B1(n26936), .B2(n22205), .ZN(
        n6248) );
  OAI22_X1 U23627 ( .A1(n27401), .A2(n26942), .B1(n26936), .B2(n22204), .ZN(
        n6249) );
  OAI22_X1 U23628 ( .A1(n27404), .A2(n26942), .B1(n26936), .B2(n22203), .ZN(
        n6250) );
  OAI22_X1 U23629 ( .A1(n27407), .A2(n26942), .B1(n26936), .B2(n22202), .ZN(
        n6251) );
  OAI22_X1 U23630 ( .A1(n27410), .A2(n26942), .B1(n26936), .B2(n22201), .ZN(
        n6252) );
  OAI22_X1 U23631 ( .A1(n27413), .A2(n26942), .B1(n26936), .B2(n22200), .ZN(
        n6253) );
  OAI22_X1 U23632 ( .A1(n27416), .A2(n26942), .B1(n26936), .B2(n22199), .ZN(
        n6254) );
  OAI22_X1 U23633 ( .A1(n27419), .A2(n26942), .B1(n26936), .B2(n22198), .ZN(
        n6255) );
  OAI22_X1 U23634 ( .A1(n27422), .A2(n26942), .B1(n26936), .B2(n22197), .ZN(
        n6256) );
  OAI22_X1 U23635 ( .A1(n27425), .A2(n26943), .B1(n26936), .B2(n22196), .ZN(
        n6257) );
  OAI22_X1 U23636 ( .A1(n27428), .A2(n26943), .B1(n26937), .B2(n22195), .ZN(
        n6258) );
  OAI22_X1 U23637 ( .A1(n27431), .A2(n26943), .B1(n26937), .B2(n22194), .ZN(
        n6259) );
  OAI22_X1 U23638 ( .A1(n27434), .A2(n26943), .B1(n26937), .B2(n22193), .ZN(
        n6260) );
  OAI22_X1 U23639 ( .A1(n27437), .A2(n26943), .B1(n26937), .B2(n22192), .ZN(
        n6261) );
  OAI22_X1 U23640 ( .A1(n27440), .A2(n26943), .B1(n26937), .B2(n22191), .ZN(
        n6262) );
  OAI22_X1 U23641 ( .A1(n27443), .A2(n26943), .B1(n26937), .B2(n22190), .ZN(
        n6263) );
  OAI22_X1 U23642 ( .A1(n27446), .A2(n26943), .B1(n26937), .B2(n22189), .ZN(
        n6264) );
  OAI22_X1 U23643 ( .A1(n27449), .A2(n26943), .B1(n26937), .B2(n22188), .ZN(
        n6265) );
  OAI22_X1 U23644 ( .A1(n27452), .A2(n26943), .B1(n26937), .B2(n22187), .ZN(
        n6266) );
  OAI22_X1 U23645 ( .A1(n27455), .A2(n26943), .B1(n26937), .B2(n22186), .ZN(
        n6267) );
  OAI22_X1 U23646 ( .A1(n27458), .A2(n26943), .B1(n26937), .B2(n22185), .ZN(
        n6268) );
  OAI22_X1 U23647 ( .A1(n27461), .A2(n26944), .B1(n26937), .B2(n22184), .ZN(
        n6269) );
  OAI22_X1 U23648 ( .A1(n27278), .A2(n27318), .B1(n27270), .B2(n22167), .ZN(
        n8014) );
  OAI22_X1 U23649 ( .A1(n27278), .A2(n27321), .B1(n27270), .B2(n22166), .ZN(
        n8015) );
  OAI22_X1 U23650 ( .A1(n27278), .A2(n27324), .B1(n27270), .B2(n22165), .ZN(
        n8016) );
  OAI22_X1 U23651 ( .A1(n27278), .A2(n27327), .B1(n27270), .B2(n22164), .ZN(
        n8017) );
  OAI22_X1 U23652 ( .A1(n27278), .A2(n27330), .B1(n27270), .B2(n22163), .ZN(
        n8018) );
  OAI22_X1 U23653 ( .A1(n27278), .A2(n27333), .B1(n27270), .B2(n22162), .ZN(
        n8019) );
  OAI22_X1 U23654 ( .A1(n27278), .A2(n27336), .B1(n27270), .B2(n22161), .ZN(
        n8020) );
  OAI22_X1 U23655 ( .A1(n27278), .A2(n27339), .B1(n27270), .B2(n22160), .ZN(
        n8021) );
  OAI22_X1 U23656 ( .A1(n27278), .A2(n27342), .B1(n27270), .B2(n22159), .ZN(
        n8022) );
  OAI22_X1 U23657 ( .A1(n27278), .A2(n27345), .B1(n27270), .B2(n22158), .ZN(
        n8023) );
  OAI22_X1 U23658 ( .A1(n27278), .A2(n27348), .B1(n27270), .B2(n22157), .ZN(
        n8024) );
  OAI22_X1 U23659 ( .A1(n27278), .A2(n27351), .B1(n27270), .B2(n22156), .ZN(
        n8025) );
  OAI22_X1 U23660 ( .A1(n27278), .A2(n27354), .B1(n27271), .B2(n22155), .ZN(
        n8026) );
  OAI22_X1 U23661 ( .A1(n27279), .A2(n27357), .B1(n27271), .B2(n22154), .ZN(
        n8027) );
  OAI22_X1 U23662 ( .A1(n27279), .A2(n27360), .B1(n27271), .B2(n22153), .ZN(
        n8028) );
  OAI22_X1 U23663 ( .A1(n27279), .A2(n27363), .B1(n27271), .B2(n22152), .ZN(
        n8029) );
  OAI22_X1 U23664 ( .A1(n27279), .A2(n27366), .B1(n27271), .B2(n22151), .ZN(
        n8030) );
  OAI22_X1 U23665 ( .A1(n27279), .A2(n27369), .B1(n27271), .B2(n22150), .ZN(
        n8031) );
  OAI22_X1 U23666 ( .A1(n27279), .A2(n27372), .B1(n27271), .B2(n22149), .ZN(
        n8032) );
  OAI22_X1 U23667 ( .A1(n27279), .A2(n27375), .B1(n27271), .B2(n22148), .ZN(
        n8033) );
  OAI22_X1 U23668 ( .A1(n27279), .A2(n27378), .B1(n27271), .B2(n22147), .ZN(
        n8034) );
  OAI22_X1 U23669 ( .A1(n27279), .A2(n27381), .B1(n27271), .B2(n22146), .ZN(
        n8035) );
  OAI22_X1 U23670 ( .A1(n27279), .A2(n27384), .B1(n27271), .B2(n22145), .ZN(
        n8036) );
  OAI22_X1 U23671 ( .A1(n27279), .A2(n27387), .B1(n27271), .B2(n22144), .ZN(
        n8037) );
  OAI22_X1 U23672 ( .A1(n27279), .A2(n27390), .B1(n27272), .B2(n22143), .ZN(
        n8038) );
  OAI22_X1 U23673 ( .A1(n27279), .A2(n27393), .B1(n27272), .B2(n22142), .ZN(
        n8039) );
  OAI22_X1 U23674 ( .A1(n27280), .A2(n27396), .B1(n27272), .B2(n22141), .ZN(
        n8040) );
  OAI22_X1 U23675 ( .A1(n27280), .A2(n27399), .B1(n27272), .B2(n22140), .ZN(
        n8041) );
  OAI22_X1 U23676 ( .A1(n27280), .A2(n27402), .B1(n27272), .B2(n22139), .ZN(
        n8042) );
  OAI22_X1 U23677 ( .A1(n27280), .A2(n27405), .B1(n27272), .B2(n22138), .ZN(
        n8043) );
  OAI22_X1 U23678 ( .A1(n27280), .A2(n27408), .B1(n27272), .B2(n22137), .ZN(
        n8044) );
  OAI22_X1 U23679 ( .A1(n27280), .A2(n27411), .B1(n27272), .B2(n22136), .ZN(
        n8045) );
  OAI22_X1 U23680 ( .A1(n27280), .A2(n27414), .B1(n27272), .B2(n22135), .ZN(
        n8046) );
  OAI22_X1 U23681 ( .A1(n27280), .A2(n27417), .B1(n27272), .B2(n22134), .ZN(
        n8047) );
  OAI22_X1 U23682 ( .A1(n27280), .A2(n27420), .B1(n27272), .B2(n22133), .ZN(
        n8048) );
  OAI22_X1 U23683 ( .A1(n27280), .A2(n27423), .B1(n27272), .B2(n22132), .ZN(
        n8049) );
  OAI22_X1 U23684 ( .A1(n27280), .A2(n27426), .B1(n27273), .B2(n22131), .ZN(
        n8050) );
  OAI22_X1 U23685 ( .A1(n27280), .A2(n27429), .B1(n27273), .B2(n22130), .ZN(
        n8051) );
  OAI22_X1 U23686 ( .A1(n27280), .A2(n27432), .B1(n27273), .B2(n22129), .ZN(
        n8052) );
  OAI22_X1 U23687 ( .A1(n27281), .A2(n27435), .B1(n27273), .B2(n22128), .ZN(
        n8053) );
  OAI22_X1 U23688 ( .A1(n27281), .A2(n27438), .B1(n27273), .B2(n22127), .ZN(
        n8054) );
  OAI22_X1 U23689 ( .A1(n27281), .A2(n27441), .B1(n27273), .B2(n22126), .ZN(
        n8055) );
  OAI22_X1 U23690 ( .A1(n27281), .A2(n27444), .B1(n27273), .B2(n22125), .ZN(
        n8056) );
  OAI22_X1 U23691 ( .A1(n27281), .A2(n27447), .B1(n27273), .B2(n22124), .ZN(
        n8057) );
  OAI22_X1 U23692 ( .A1(n27281), .A2(n27450), .B1(n27273), .B2(n22123), .ZN(
        n8058) );
  OAI22_X1 U23693 ( .A1(n27281), .A2(n27453), .B1(n27273), .B2(n22122), .ZN(
        n8059) );
  OAI22_X1 U23694 ( .A1(n27281), .A2(n27456), .B1(n27273), .B2(n22121), .ZN(
        n8060) );
  OAI22_X1 U23695 ( .A1(n27281), .A2(n27459), .B1(n27273), .B2(n22120), .ZN(
        n8061) );
  OAI22_X1 U23696 ( .A1(n27318), .A2(n27264), .B1(n27258), .B2(n22107), .ZN(
        n7950) );
  OAI22_X1 U23697 ( .A1(n27321), .A2(n27264), .B1(n27258), .B2(n22106), .ZN(
        n7951) );
  OAI22_X1 U23698 ( .A1(n27324), .A2(n27264), .B1(n27258), .B2(n22105), .ZN(
        n7952) );
  OAI22_X1 U23699 ( .A1(n27327), .A2(n27264), .B1(n27258), .B2(n22104), .ZN(
        n7953) );
  OAI22_X1 U23700 ( .A1(n27330), .A2(n27264), .B1(n27258), .B2(n22103), .ZN(
        n7954) );
  OAI22_X1 U23701 ( .A1(n27333), .A2(n27264), .B1(n27258), .B2(n22102), .ZN(
        n7955) );
  OAI22_X1 U23702 ( .A1(n27336), .A2(n27264), .B1(n27258), .B2(n22101), .ZN(
        n7956) );
  OAI22_X1 U23703 ( .A1(n27339), .A2(n27264), .B1(n27258), .B2(n22100), .ZN(
        n7957) );
  OAI22_X1 U23704 ( .A1(n27342), .A2(n27264), .B1(n27258), .B2(n22099), .ZN(
        n7958) );
  OAI22_X1 U23705 ( .A1(n27345), .A2(n27264), .B1(n27258), .B2(n22098), .ZN(
        n7959) );
  OAI22_X1 U23706 ( .A1(n27348), .A2(n27264), .B1(n27258), .B2(n22097), .ZN(
        n7960) );
  OAI22_X1 U23707 ( .A1(n27351), .A2(n27265), .B1(n27258), .B2(n22096), .ZN(
        n7961) );
  OAI22_X1 U23708 ( .A1(n27354), .A2(n27265), .B1(n27259), .B2(n22095), .ZN(
        n7962) );
  OAI22_X1 U23709 ( .A1(n27357), .A2(n27265), .B1(n27259), .B2(n22094), .ZN(
        n7963) );
  OAI22_X1 U23710 ( .A1(n27360), .A2(n27265), .B1(n27259), .B2(n22093), .ZN(
        n7964) );
  OAI22_X1 U23711 ( .A1(n27363), .A2(n27265), .B1(n27259), .B2(n22092), .ZN(
        n7965) );
  OAI22_X1 U23712 ( .A1(n27366), .A2(n27265), .B1(n27259), .B2(n22091), .ZN(
        n7966) );
  OAI22_X1 U23713 ( .A1(n27369), .A2(n27265), .B1(n27259), .B2(n22090), .ZN(
        n7967) );
  OAI22_X1 U23714 ( .A1(n27372), .A2(n27265), .B1(n27259), .B2(n22089), .ZN(
        n7968) );
  OAI22_X1 U23715 ( .A1(n27375), .A2(n27265), .B1(n27259), .B2(n22088), .ZN(
        n7969) );
  OAI22_X1 U23716 ( .A1(n27378), .A2(n27265), .B1(n27259), .B2(n22087), .ZN(
        n7970) );
  OAI22_X1 U23717 ( .A1(n27381), .A2(n27265), .B1(n27259), .B2(n22086), .ZN(
        n7971) );
  OAI22_X1 U23718 ( .A1(n27384), .A2(n27265), .B1(n27259), .B2(n22085), .ZN(
        n7972) );
  OAI22_X1 U23719 ( .A1(n27387), .A2(n27266), .B1(n27259), .B2(n22084), .ZN(
        n7973) );
  OAI22_X1 U23720 ( .A1(n27390), .A2(n27266), .B1(n27260), .B2(n22083), .ZN(
        n7974) );
  OAI22_X1 U23721 ( .A1(n27393), .A2(n27266), .B1(n27260), .B2(n22082), .ZN(
        n7975) );
  OAI22_X1 U23722 ( .A1(n27396), .A2(n27266), .B1(n27260), .B2(n22081), .ZN(
        n7976) );
  OAI22_X1 U23723 ( .A1(n27399), .A2(n27266), .B1(n27260), .B2(n22080), .ZN(
        n7977) );
  OAI22_X1 U23724 ( .A1(n27402), .A2(n27266), .B1(n27260), .B2(n22079), .ZN(
        n7978) );
  OAI22_X1 U23725 ( .A1(n27405), .A2(n27266), .B1(n27260), .B2(n22078), .ZN(
        n7979) );
  OAI22_X1 U23726 ( .A1(n27408), .A2(n27266), .B1(n27260), .B2(n22077), .ZN(
        n7980) );
  OAI22_X1 U23727 ( .A1(n27411), .A2(n27266), .B1(n27260), .B2(n22076), .ZN(
        n7981) );
  OAI22_X1 U23728 ( .A1(n27414), .A2(n27266), .B1(n27260), .B2(n22075), .ZN(
        n7982) );
  OAI22_X1 U23729 ( .A1(n27417), .A2(n27266), .B1(n27260), .B2(n22074), .ZN(
        n7983) );
  OAI22_X1 U23730 ( .A1(n27420), .A2(n27266), .B1(n27260), .B2(n22073), .ZN(
        n7984) );
  OAI22_X1 U23731 ( .A1(n27423), .A2(n27267), .B1(n27260), .B2(n22072), .ZN(
        n7985) );
  OAI22_X1 U23732 ( .A1(n27426), .A2(n27267), .B1(n27261), .B2(n22071), .ZN(
        n7986) );
  OAI22_X1 U23733 ( .A1(n27429), .A2(n27267), .B1(n27261), .B2(n22070), .ZN(
        n7987) );
  OAI22_X1 U23734 ( .A1(n27432), .A2(n27267), .B1(n27261), .B2(n22069), .ZN(
        n7988) );
  OAI22_X1 U23735 ( .A1(n27435), .A2(n27267), .B1(n27261), .B2(n22068), .ZN(
        n7989) );
  OAI22_X1 U23736 ( .A1(n27438), .A2(n27267), .B1(n27261), .B2(n22067), .ZN(
        n7990) );
  OAI22_X1 U23737 ( .A1(n27441), .A2(n27267), .B1(n27261), .B2(n22066), .ZN(
        n7991) );
  OAI22_X1 U23738 ( .A1(n27444), .A2(n27267), .B1(n27261), .B2(n22065), .ZN(
        n7992) );
  OAI22_X1 U23739 ( .A1(n27447), .A2(n27267), .B1(n27261), .B2(n22064), .ZN(
        n7993) );
  OAI22_X1 U23740 ( .A1(n27450), .A2(n27267), .B1(n27261), .B2(n22063), .ZN(
        n7994) );
  OAI22_X1 U23741 ( .A1(n27453), .A2(n27267), .B1(n27261), .B2(n22062), .ZN(
        n7995) );
  OAI22_X1 U23742 ( .A1(n27456), .A2(n27267), .B1(n27261), .B2(n22061), .ZN(
        n7996) );
  OAI22_X1 U23743 ( .A1(n27459), .A2(n27268), .B1(n27261), .B2(n22060), .ZN(
        n7997) );
  OAI22_X1 U23744 ( .A1(n27318), .A2(n27228), .B1(n27222), .B2(n21927), .ZN(
        n7758) );
  OAI22_X1 U23745 ( .A1(n27321), .A2(n27228), .B1(n27222), .B2(n21926), .ZN(
        n7759) );
  OAI22_X1 U23746 ( .A1(n27324), .A2(n27228), .B1(n27222), .B2(n21925), .ZN(
        n7760) );
  OAI22_X1 U23747 ( .A1(n27327), .A2(n27228), .B1(n27222), .B2(n21924), .ZN(
        n7761) );
  OAI22_X1 U23748 ( .A1(n27330), .A2(n27228), .B1(n27222), .B2(n21923), .ZN(
        n7762) );
  OAI22_X1 U23749 ( .A1(n27333), .A2(n27228), .B1(n27222), .B2(n21922), .ZN(
        n7763) );
  OAI22_X1 U23750 ( .A1(n27336), .A2(n27228), .B1(n27222), .B2(n21921), .ZN(
        n7764) );
  OAI22_X1 U23751 ( .A1(n27339), .A2(n27228), .B1(n27222), .B2(n21920), .ZN(
        n7765) );
  OAI22_X1 U23752 ( .A1(n27342), .A2(n27228), .B1(n27222), .B2(n21919), .ZN(
        n7766) );
  OAI22_X1 U23753 ( .A1(n27345), .A2(n27228), .B1(n27222), .B2(n21918), .ZN(
        n7767) );
  OAI22_X1 U23754 ( .A1(n27348), .A2(n27228), .B1(n27222), .B2(n21917), .ZN(
        n7768) );
  OAI22_X1 U23755 ( .A1(n27351), .A2(n27229), .B1(n27222), .B2(n21916), .ZN(
        n7769) );
  OAI22_X1 U23756 ( .A1(n27354), .A2(n27229), .B1(n27223), .B2(n21915), .ZN(
        n7770) );
  OAI22_X1 U23757 ( .A1(n27357), .A2(n27229), .B1(n27223), .B2(n21914), .ZN(
        n7771) );
  OAI22_X1 U23758 ( .A1(n27360), .A2(n27229), .B1(n27223), .B2(n21913), .ZN(
        n7772) );
  OAI22_X1 U23759 ( .A1(n27363), .A2(n27229), .B1(n27223), .B2(n21912), .ZN(
        n7773) );
  OAI22_X1 U23760 ( .A1(n27366), .A2(n27229), .B1(n27223), .B2(n21911), .ZN(
        n7774) );
  OAI22_X1 U23761 ( .A1(n27369), .A2(n27229), .B1(n27223), .B2(n21910), .ZN(
        n7775) );
  OAI22_X1 U23762 ( .A1(n27372), .A2(n27229), .B1(n27223), .B2(n21909), .ZN(
        n7776) );
  OAI22_X1 U23763 ( .A1(n27375), .A2(n27229), .B1(n27223), .B2(n21908), .ZN(
        n7777) );
  OAI22_X1 U23764 ( .A1(n27378), .A2(n27229), .B1(n27223), .B2(n21907), .ZN(
        n7778) );
  OAI22_X1 U23765 ( .A1(n27381), .A2(n27229), .B1(n27223), .B2(n21906), .ZN(
        n7779) );
  OAI22_X1 U23766 ( .A1(n27384), .A2(n27229), .B1(n27223), .B2(n21905), .ZN(
        n7780) );
  OAI22_X1 U23767 ( .A1(n27387), .A2(n27230), .B1(n27223), .B2(n21904), .ZN(
        n7781) );
  OAI22_X1 U23768 ( .A1(n27390), .A2(n27230), .B1(n27224), .B2(n21903), .ZN(
        n7782) );
  OAI22_X1 U23769 ( .A1(n27393), .A2(n27230), .B1(n27224), .B2(n21902), .ZN(
        n7783) );
  OAI22_X1 U23770 ( .A1(n27396), .A2(n27230), .B1(n27224), .B2(n21901), .ZN(
        n7784) );
  OAI22_X1 U23771 ( .A1(n27399), .A2(n27230), .B1(n27224), .B2(n21900), .ZN(
        n7785) );
  OAI22_X1 U23772 ( .A1(n27402), .A2(n27230), .B1(n27224), .B2(n21899), .ZN(
        n7786) );
  OAI22_X1 U23773 ( .A1(n27405), .A2(n27230), .B1(n27224), .B2(n21898), .ZN(
        n7787) );
  OAI22_X1 U23774 ( .A1(n27408), .A2(n27230), .B1(n27224), .B2(n21897), .ZN(
        n7788) );
  OAI22_X1 U23775 ( .A1(n27411), .A2(n27230), .B1(n27224), .B2(n21896), .ZN(
        n7789) );
  OAI22_X1 U23776 ( .A1(n27414), .A2(n27230), .B1(n27224), .B2(n21895), .ZN(
        n7790) );
  OAI22_X1 U23777 ( .A1(n27417), .A2(n27230), .B1(n27224), .B2(n21894), .ZN(
        n7791) );
  OAI22_X1 U23778 ( .A1(n27420), .A2(n27230), .B1(n27224), .B2(n21893), .ZN(
        n7792) );
  OAI22_X1 U23779 ( .A1(n27423), .A2(n27231), .B1(n27224), .B2(n21892), .ZN(
        n7793) );
  OAI22_X1 U23780 ( .A1(n27426), .A2(n27231), .B1(n27225), .B2(n21891), .ZN(
        n7794) );
  OAI22_X1 U23781 ( .A1(n27429), .A2(n27231), .B1(n27225), .B2(n21890), .ZN(
        n7795) );
  OAI22_X1 U23782 ( .A1(n27432), .A2(n27231), .B1(n27225), .B2(n21889), .ZN(
        n7796) );
  OAI22_X1 U23783 ( .A1(n27435), .A2(n27231), .B1(n27225), .B2(n21888), .ZN(
        n7797) );
  OAI22_X1 U23784 ( .A1(n27438), .A2(n27231), .B1(n27225), .B2(n21887), .ZN(
        n7798) );
  OAI22_X1 U23785 ( .A1(n27441), .A2(n27231), .B1(n27225), .B2(n21886), .ZN(
        n7799) );
  OAI22_X1 U23786 ( .A1(n27444), .A2(n27231), .B1(n27225), .B2(n21885), .ZN(
        n7800) );
  OAI22_X1 U23787 ( .A1(n27447), .A2(n27231), .B1(n27225), .B2(n21884), .ZN(
        n7801) );
  OAI22_X1 U23788 ( .A1(n27450), .A2(n27231), .B1(n27225), .B2(n21883), .ZN(
        n7802) );
  OAI22_X1 U23789 ( .A1(n27453), .A2(n27231), .B1(n27225), .B2(n21882), .ZN(
        n7803) );
  OAI22_X1 U23790 ( .A1(n27456), .A2(n27231), .B1(n27225), .B2(n21881), .ZN(
        n7804) );
  OAI22_X1 U23791 ( .A1(n27459), .A2(n27232), .B1(n27225), .B2(n21880), .ZN(
        n7805) );
  OAI22_X1 U23792 ( .A1(n27318), .A2(n27204), .B1(n27198), .B2(n21867), .ZN(
        n7630) );
  OAI22_X1 U23793 ( .A1(n27321), .A2(n27204), .B1(n27198), .B2(n21866), .ZN(
        n7631) );
  OAI22_X1 U23794 ( .A1(n27324), .A2(n27204), .B1(n27198), .B2(n21865), .ZN(
        n7632) );
  OAI22_X1 U23795 ( .A1(n27327), .A2(n27204), .B1(n27198), .B2(n21864), .ZN(
        n7633) );
  OAI22_X1 U23796 ( .A1(n27330), .A2(n27204), .B1(n27198), .B2(n21863), .ZN(
        n7634) );
  OAI22_X1 U23797 ( .A1(n27333), .A2(n27204), .B1(n27198), .B2(n21862), .ZN(
        n7635) );
  OAI22_X1 U23798 ( .A1(n27336), .A2(n27204), .B1(n27198), .B2(n21861), .ZN(
        n7636) );
  OAI22_X1 U23799 ( .A1(n27339), .A2(n27204), .B1(n27198), .B2(n21860), .ZN(
        n7637) );
  OAI22_X1 U23800 ( .A1(n27342), .A2(n27204), .B1(n27198), .B2(n21859), .ZN(
        n7638) );
  OAI22_X1 U23801 ( .A1(n27345), .A2(n27204), .B1(n27198), .B2(n21858), .ZN(
        n7639) );
  OAI22_X1 U23802 ( .A1(n27348), .A2(n27204), .B1(n27198), .B2(n21857), .ZN(
        n7640) );
  OAI22_X1 U23803 ( .A1(n27351), .A2(n27205), .B1(n27198), .B2(n21856), .ZN(
        n7641) );
  OAI22_X1 U23804 ( .A1(n27354), .A2(n27205), .B1(n27199), .B2(n21855), .ZN(
        n7642) );
  OAI22_X1 U23805 ( .A1(n27357), .A2(n27205), .B1(n27199), .B2(n21854), .ZN(
        n7643) );
  OAI22_X1 U23806 ( .A1(n27360), .A2(n27205), .B1(n27199), .B2(n21853), .ZN(
        n7644) );
  OAI22_X1 U23807 ( .A1(n27363), .A2(n27205), .B1(n27199), .B2(n21852), .ZN(
        n7645) );
  OAI22_X1 U23808 ( .A1(n27366), .A2(n27205), .B1(n27199), .B2(n21851), .ZN(
        n7646) );
  OAI22_X1 U23809 ( .A1(n27369), .A2(n27205), .B1(n27199), .B2(n21850), .ZN(
        n7647) );
  OAI22_X1 U23810 ( .A1(n27372), .A2(n27205), .B1(n27199), .B2(n21849), .ZN(
        n7648) );
  OAI22_X1 U23811 ( .A1(n27375), .A2(n27205), .B1(n27199), .B2(n21848), .ZN(
        n7649) );
  OAI22_X1 U23812 ( .A1(n27378), .A2(n27205), .B1(n27199), .B2(n21847), .ZN(
        n7650) );
  OAI22_X1 U23813 ( .A1(n27381), .A2(n27205), .B1(n27199), .B2(n21846), .ZN(
        n7651) );
  OAI22_X1 U23814 ( .A1(n27384), .A2(n27205), .B1(n27199), .B2(n21845), .ZN(
        n7652) );
  OAI22_X1 U23815 ( .A1(n27387), .A2(n27206), .B1(n27199), .B2(n21844), .ZN(
        n7653) );
  OAI22_X1 U23816 ( .A1(n27390), .A2(n27206), .B1(n27200), .B2(n21843), .ZN(
        n7654) );
  OAI22_X1 U23817 ( .A1(n27393), .A2(n27206), .B1(n27200), .B2(n21842), .ZN(
        n7655) );
  OAI22_X1 U23818 ( .A1(n27396), .A2(n27206), .B1(n27200), .B2(n21841), .ZN(
        n7656) );
  OAI22_X1 U23819 ( .A1(n27399), .A2(n27206), .B1(n27200), .B2(n21840), .ZN(
        n7657) );
  OAI22_X1 U23820 ( .A1(n27402), .A2(n27206), .B1(n27200), .B2(n21839), .ZN(
        n7658) );
  OAI22_X1 U23821 ( .A1(n27405), .A2(n27206), .B1(n27200), .B2(n21838), .ZN(
        n7659) );
  OAI22_X1 U23822 ( .A1(n27408), .A2(n27206), .B1(n27200), .B2(n21837), .ZN(
        n7660) );
  OAI22_X1 U23823 ( .A1(n27411), .A2(n27206), .B1(n27200), .B2(n21836), .ZN(
        n7661) );
  OAI22_X1 U23824 ( .A1(n27414), .A2(n27206), .B1(n27200), .B2(n21835), .ZN(
        n7662) );
  OAI22_X1 U23825 ( .A1(n27417), .A2(n27206), .B1(n27200), .B2(n21834), .ZN(
        n7663) );
  OAI22_X1 U23826 ( .A1(n27420), .A2(n27206), .B1(n27200), .B2(n21833), .ZN(
        n7664) );
  OAI22_X1 U23827 ( .A1(n27423), .A2(n27207), .B1(n27200), .B2(n21832), .ZN(
        n7665) );
  OAI22_X1 U23828 ( .A1(n27426), .A2(n27207), .B1(n27201), .B2(n21831), .ZN(
        n7666) );
  OAI22_X1 U23829 ( .A1(n27429), .A2(n27207), .B1(n27201), .B2(n21830), .ZN(
        n7667) );
  OAI22_X1 U23830 ( .A1(n27432), .A2(n27207), .B1(n27201), .B2(n21829), .ZN(
        n7668) );
  OAI22_X1 U23831 ( .A1(n27435), .A2(n27207), .B1(n27201), .B2(n21828), .ZN(
        n7669) );
  OAI22_X1 U23832 ( .A1(n27438), .A2(n27207), .B1(n27201), .B2(n21827), .ZN(
        n7670) );
  OAI22_X1 U23833 ( .A1(n27441), .A2(n27207), .B1(n27201), .B2(n21826), .ZN(
        n7671) );
  OAI22_X1 U23834 ( .A1(n27444), .A2(n27207), .B1(n27201), .B2(n21825), .ZN(
        n7672) );
  OAI22_X1 U23835 ( .A1(n27447), .A2(n27207), .B1(n27201), .B2(n21824), .ZN(
        n7673) );
  OAI22_X1 U23836 ( .A1(n27450), .A2(n27207), .B1(n27201), .B2(n21823), .ZN(
        n7674) );
  OAI22_X1 U23837 ( .A1(n27453), .A2(n27207), .B1(n27201), .B2(n21822), .ZN(
        n7675) );
  OAI22_X1 U23838 ( .A1(n27456), .A2(n27207), .B1(n27201), .B2(n21821), .ZN(
        n7676) );
  OAI22_X1 U23839 ( .A1(n27459), .A2(n27208), .B1(n27201), .B2(n21820), .ZN(
        n7677) );
  OAI22_X1 U23840 ( .A1(n27319), .A2(n27012), .B1(n27006), .B2(n21807), .ZN(
        n6606) );
  OAI22_X1 U23841 ( .A1(n27322), .A2(n27012), .B1(n27006), .B2(n21806), .ZN(
        n6607) );
  OAI22_X1 U23842 ( .A1(n27325), .A2(n27012), .B1(n27006), .B2(n21805), .ZN(
        n6608) );
  OAI22_X1 U23843 ( .A1(n27328), .A2(n27012), .B1(n27006), .B2(n21804), .ZN(
        n6609) );
  OAI22_X1 U23844 ( .A1(n27331), .A2(n27012), .B1(n27006), .B2(n21803), .ZN(
        n6610) );
  OAI22_X1 U23845 ( .A1(n27334), .A2(n27012), .B1(n27006), .B2(n21802), .ZN(
        n6611) );
  OAI22_X1 U23846 ( .A1(n27337), .A2(n27012), .B1(n27006), .B2(n21801), .ZN(
        n6612) );
  OAI22_X1 U23847 ( .A1(n27340), .A2(n27012), .B1(n27006), .B2(n21800), .ZN(
        n6613) );
  OAI22_X1 U23848 ( .A1(n27343), .A2(n27012), .B1(n27006), .B2(n21799), .ZN(
        n6614) );
  OAI22_X1 U23849 ( .A1(n27346), .A2(n27012), .B1(n27006), .B2(n21798), .ZN(
        n6615) );
  OAI22_X1 U23850 ( .A1(n27349), .A2(n27012), .B1(n27006), .B2(n21797), .ZN(
        n6616) );
  OAI22_X1 U23851 ( .A1(n27352), .A2(n27013), .B1(n27006), .B2(n21796), .ZN(
        n6617) );
  OAI22_X1 U23852 ( .A1(n27355), .A2(n27013), .B1(n27007), .B2(n21795), .ZN(
        n6618) );
  OAI22_X1 U23853 ( .A1(n27358), .A2(n27013), .B1(n27007), .B2(n21794), .ZN(
        n6619) );
  OAI22_X1 U23854 ( .A1(n27361), .A2(n27013), .B1(n27007), .B2(n21793), .ZN(
        n6620) );
  OAI22_X1 U23855 ( .A1(n27364), .A2(n27013), .B1(n27007), .B2(n21792), .ZN(
        n6621) );
  OAI22_X1 U23856 ( .A1(n27367), .A2(n27013), .B1(n27007), .B2(n21791), .ZN(
        n6622) );
  OAI22_X1 U23857 ( .A1(n27370), .A2(n27013), .B1(n27007), .B2(n21790), .ZN(
        n6623) );
  OAI22_X1 U23858 ( .A1(n27373), .A2(n27013), .B1(n27007), .B2(n21789), .ZN(
        n6624) );
  OAI22_X1 U23859 ( .A1(n27376), .A2(n27013), .B1(n27007), .B2(n21788), .ZN(
        n6625) );
  OAI22_X1 U23860 ( .A1(n27379), .A2(n27013), .B1(n27007), .B2(n21787), .ZN(
        n6626) );
  OAI22_X1 U23861 ( .A1(n27382), .A2(n27013), .B1(n27007), .B2(n21786), .ZN(
        n6627) );
  OAI22_X1 U23862 ( .A1(n27385), .A2(n27013), .B1(n27007), .B2(n21785), .ZN(
        n6628) );
  OAI22_X1 U23863 ( .A1(n27388), .A2(n27014), .B1(n27007), .B2(n21784), .ZN(
        n6629) );
  OAI22_X1 U23864 ( .A1(n27391), .A2(n27014), .B1(n27008), .B2(n21783), .ZN(
        n6630) );
  OAI22_X1 U23865 ( .A1(n27394), .A2(n27014), .B1(n27008), .B2(n21782), .ZN(
        n6631) );
  OAI22_X1 U23866 ( .A1(n27397), .A2(n27014), .B1(n27008), .B2(n21781), .ZN(
        n6632) );
  OAI22_X1 U23867 ( .A1(n27400), .A2(n27014), .B1(n27008), .B2(n21780), .ZN(
        n6633) );
  OAI22_X1 U23868 ( .A1(n27403), .A2(n27014), .B1(n27008), .B2(n21779), .ZN(
        n6634) );
  OAI22_X1 U23869 ( .A1(n27406), .A2(n27014), .B1(n27008), .B2(n21778), .ZN(
        n6635) );
  OAI22_X1 U23870 ( .A1(n27409), .A2(n27014), .B1(n27008), .B2(n21777), .ZN(
        n6636) );
  OAI22_X1 U23871 ( .A1(n27412), .A2(n27014), .B1(n27008), .B2(n21776), .ZN(
        n6637) );
  OAI22_X1 U23872 ( .A1(n27415), .A2(n27014), .B1(n27008), .B2(n21775), .ZN(
        n6638) );
  OAI22_X1 U23873 ( .A1(n27418), .A2(n27014), .B1(n27008), .B2(n21774), .ZN(
        n6639) );
  OAI22_X1 U23874 ( .A1(n27421), .A2(n27014), .B1(n27008), .B2(n21773), .ZN(
        n6640) );
  OAI22_X1 U23875 ( .A1(n27424), .A2(n27015), .B1(n27008), .B2(n21772), .ZN(
        n6641) );
  OAI22_X1 U23876 ( .A1(n27427), .A2(n27015), .B1(n27009), .B2(n21771), .ZN(
        n6642) );
  OAI22_X1 U23877 ( .A1(n27430), .A2(n27015), .B1(n27009), .B2(n21770), .ZN(
        n6643) );
  OAI22_X1 U23878 ( .A1(n27433), .A2(n27015), .B1(n27009), .B2(n21769), .ZN(
        n6644) );
  OAI22_X1 U23879 ( .A1(n27436), .A2(n27015), .B1(n27009), .B2(n21768), .ZN(
        n6645) );
  OAI22_X1 U23880 ( .A1(n27439), .A2(n27015), .B1(n27009), .B2(n21767), .ZN(
        n6646) );
  OAI22_X1 U23881 ( .A1(n27442), .A2(n27015), .B1(n27009), .B2(n21766), .ZN(
        n6647) );
  OAI22_X1 U23882 ( .A1(n27445), .A2(n27015), .B1(n27009), .B2(n21765), .ZN(
        n6648) );
  OAI22_X1 U23883 ( .A1(n27448), .A2(n27015), .B1(n27009), .B2(n21764), .ZN(
        n6649) );
  OAI22_X1 U23884 ( .A1(n27451), .A2(n27015), .B1(n27009), .B2(n21763), .ZN(
        n6650) );
  OAI22_X1 U23885 ( .A1(n27454), .A2(n27015), .B1(n27009), .B2(n21762), .ZN(
        n6651) );
  OAI22_X1 U23886 ( .A1(n27457), .A2(n27015), .B1(n27009), .B2(n21761), .ZN(
        n6652) );
  OAI22_X1 U23887 ( .A1(n27460), .A2(n27016), .B1(n27009), .B2(n21760), .ZN(
        n6653) );
  OAI22_X1 U23888 ( .A1(n27319), .A2(n27060), .B1(n27054), .B2(n21687), .ZN(
        n6862) );
  OAI22_X1 U23889 ( .A1(n27322), .A2(n27060), .B1(n27054), .B2(n21686), .ZN(
        n6863) );
  OAI22_X1 U23890 ( .A1(n27325), .A2(n27060), .B1(n27054), .B2(n21685), .ZN(
        n6864) );
  OAI22_X1 U23891 ( .A1(n27328), .A2(n27060), .B1(n27054), .B2(n21684), .ZN(
        n6865) );
  OAI22_X1 U23892 ( .A1(n27331), .A2(n27060), .B1(n27054), .B2(n21683), .ZN(
        n6866) );
  OAI22_X1 U23893 ( .A1(n27334), .A2(n27060), .B1(n27054), .B2(n21682), .ZN(
        n6867) );
  OAI22_X1 U23894 ( .A1(n27337), .A2(n27060), .B1(n27054), .B2(n21681), .ZN(
        n6868) );
  OAI22_X1 U23895 ( .A1(n27340), .A2(n27060), .B1(n27054), .B2(n21680), .ZN(
        n6869) );
  OAI22_X1 U23896 ( .A1(n27343), .A2(n27060), .B1(n27054), .B2(n21679), .ZN(
        n6870) );
  OAI22_X1 U23897 ( .A1(n27346), .A2(n27060), .B1(n27054), .B2(n21678), .ZN(
        n6871) );
  OAI22_X1 U23898 ( .A1(n27349), .A2(n27060), .B1(n27054), .B2(n21677), .ZN(
        n6872) );
  OAI22_X1 U23899 ( .A1(n27352), .A2(n27061), .B1(n27054), .B2(n21676), .ZN(
        n6873) );
  OAI22_X1 U23900 ( .A1(n27355), .A2(n27061), .B1(n27055), .B2(n21675), .ZN(
        n6874) );
  OAI22_X1 U23901 ( .A1(n27358), .A2(n27061), .B1(n27055), .B2(n21674), .ZN(
        n6875) );
  OAI22_X1 U23902 ( .A1(n27361), .A2(n27061), .B1(n27055), .B2(n21673), .ZN(
        n6876) );
  OAI22_X1 U23903 ( .A1(n27364), .A2(n27061), .B1(n27055), .B2(n21672), .ZN(
        n6877) );
  OAI22_X1 U23904 ( .A1(n27367), .A2(n27061), .B1(n27055), .B2(n21671), .ZN(
        n6878) );
  OAI22_X1 U23905 ( .A1(n27370), .A2(n27061), .B1(n27055), .B2(n21670), .ZN(
        n6879) );
  OAI22_X1 U23906 ( .A1(n27373), .A2(n27061), .B1(n27055), .B2(n21669), .ZN(
        n6880) );
  OAI22_X1 U23907 ( .A1(n27376), .A2(n27061), .B1(n27055), .B2(n21668), .ZN(
        n6881) );
  OAI22_X1 U23908 ( .A1(n27379), .A2(n27061), .B1(n27055), .B2(n21667), .ZN(
        n6882) );
  OAI22_X1 U23909 ( .A1(n27382), .A2(n27061), .B1(n27055), .B2(n21666), .ZN(
        n6883) );
  OAI22_X1 U23910 ( .A1(n27385), .A2(n27061), .B1(n27055), .B2(n21665), .ZN(
        n6884) );
  OAI22_X1 U23911 ( .A1(n27388), .A2(n27062), .B1(n27055), .B2(n21664), .ZN(
        n6885) );
  OAI22_X1 U23912 ( .A1(n27391), .A2(n27062), .B1(n27056), .B2(n21663), .ZN(
        n6886) );
  OAI22_X1 U23913 ( .A1(n27394), .A2(n27062), .B1(n27056), .B2(n21662), .ZN(
        n6887) );
  OAI22_X1 U23914 ( .A1(n27397), .A2(n27062), .B1(n27056), .B2(n21661), .ZN(
        n6888) );
  OAI22_X1 U23915 ( .A1(n27400), .A2(n27062), .B1(n27056), .B2(n21660), .ZN(
        n6889) );
  OAI22_X1 U23916 ( .A1(n27403), .A2(n27062), .B1(n27056), .B2(n21659), .ZN(
        n6890) );
  OAI22_X1 U23917 ( .A1(n27406), .A2(n27062), .B1(n27056), .B2(n21658), .ZN(
        n6891) );
  OAI22_X1 U23918 ( .A1(n27409), .A2(n27062), .B1(n27056), .B2(n21657), .ZN(
        n6892) );
  OAI22_X1 U23919 ( .A1(n27412), .A2(n27062), .B1(n27056), .B2(n21656), .ZN(
        n6893) );
  OAI22_X1 U23920 ( .A1(n27415), .A2(n27062), .B1(n27056), .B2(n21655), .ZN(
        n6894) );
  OAI22_X1 U23921 ( .A1(n27418), .A2(n27062), .B1(n27056), .B2(n21654), .ZN(
        n6895) );
  OAI22_X1 U23922 ( .A1(n27421), .A2(n27062), .B1(n27056), .B2(n21653), .ZN(
        n6896) );
  OAI22_X1 U23923 ( .A1(n27424), .A2(n27063), .B1(n27056), .B2(n21652), .ZN(
        n6897) );
  OAI22_X1 U23924 ( .A1(n27427), .A2(n27063), .B1(n27057), .B2(n21651), .ZN(
        n6898) );
  OAI22_X1 U23925 ( .A1(n27430), .A2(n27063), .B1(n27057), .B2(n21650), .ZN(
        n6899) );
  OAI22_X1 U23926 ( .A1(n27433), .A2(n27063), .B1(n27057), .B2(n21649), .ZN(
        n6900) );
  OAI22_X1 U23927 ( .A1(n27436), .A2(n27063), .B1(n27057), .B2(n21648), .ZN(
        n6901) );
  OAI22_X1 U23928 ( .A1(n27439), .A2(n27063), .B1(n27057), .B2(n21647), .ZN(
        n6902) );
  OAI22_X1 U23929 ( .A1(n27442), .A2(n27063), .B1(n27057), .B2(n21646), .ZN(
        n6903) );
  OAI22_X1 U23930 ( .A1(n27445), .A2(n27063), .B1(n27057), .B2(n21645), .ZN(
        n6904) );
  OAI22_X1 U23931 ( .A1(n27448), .A2(n27063), .B1(n27057), .B2(n21644), .ZN(
        n6905) );
  OAI22_X1 U23932 ( .A1(n27451), .A2(n27063), .B1(n27057), .B2(n21643), .ZN(
        n6906) );
  OAI22_X1 U23933 ( .A1(n27454), .A2(n27063), .B1(n27057), .B2(n21642), .ZN(
        n6907) );
  OAI22_X1 U23934 ( .A1(n27457), .A2(n27063), .B1(n27057), .B2(n21641), .ZN(
        n6908) );
  OAI22_X1 U23935 ( .A1(n27460), .A2(n27064), .B1(n27057), .B2(n21640), .ZN(
        n6909) );
  OAI22_X1 U23936 ( .A1(n27318), .A2(n27252), .B1(n27246), .B2(n21467), .ZN(
        n7886) );
  OAI22_X1 U23937 ( .A1(n27321), .A2(n27252), .B1(n27246), .B2(n21466), .ZN(
        n7887) );
  OAI22_X1 U23938 ( .A1(n27324), .A2(n27252), .B1(n27246), .B2(n21465), .ZN(
        n7888) );
  OAI22_X1 U23939 ( .A1(n27327), .A2(n27252), .B1(n27246), .B2(n21464), .ZN(
        n7889) );
  OAI22_X1 U23940 ( .A1(n27330), .A2(n27252), .B1(n27246), .B2(n21463), .ZN(
        n7890) );
  OAI22_X1 U23941 ( .A1(n27333), .A2(n27252), .B1(n27246), .B2(n21462), .ZN(
        n7891) );
  OAI22_X1 U23942 ( .A1(n27336), .A2(n27252), .B1(n27246), .B2(n21461), .ZN(
        n7892) );
  OAI22_X1 U23943 ( .A1(n27339), .A2(n27252), .B1(n27246), .B2(n21460), .ZN(
        n7893) );
  OAI22_X1 U23944 ( .A1(n27342), .A2(n27252), .B1(n27246), .B2(n21459), .ZN(
        n7894) );
  OAI22_X1 U23945 ( .A1(n27345), .A2(n27252), .B1(n27246), .B2(n21458), .ZN(
        n7895) );
  OAI22_X1 U23946 ( .A1(n27348), .A2(n27252), .B1(n27246), .B2(n21457), .ZN(
        n7896) );
  OAI22_X1 U23947 ( .A1(n27351), .A2(n27253), .B1(n27246), .B2(n21456), .ZN(
        n7897) );
  OAI22_X1 U23948 ( .A1(n27354), .A2(n27253), .B1(n27247), .B2(n21455), .ZN(
        n7898) );
  OAI22_X1 U23949 ( .A1(n27357), .A2(n27253), .B1(n27247), .B2(n21454), .ZN(
        n7899) );
  OAI22_X1 U23950 ( .A1(n27360), .A2(n27253), .B1(n27247), .B2(n21453), .ZN(
        n7900) );
  OAI22_X1 U23951 ( .A1(n27363), .A2(n27253), .B1(n27247), .B2(n21452), .ZN(
        n7901) );
  OAI22_X1 U23952 ( .A1(n27366), .A2(n27253), .B1(n27247), .B2(n21451), .ZN(
        n7902) );
  OAI22_X1 U23953 ( .A1(n27369), .A2(n27253), .B1(n27247), .B2(n21450), .ZN(
        n7903) );
  OAI22_X1 U23954 ( .A1(n27372), .A2(n27253), .B1(n27247), .B2(n21449), .ZN(
        n7904) );
  OAI22_X1 U23955 ( .A1(n27375), .A2(n27253), .B1(n27247), .B2(n21448), .ZN(
        n7905) );
  OAI22_X1 U23956 ( .A1(n27378), .A2(n27253), .B1(n27247), .B2(n21447), .ZN(
        n7906) );
  OAI22_X1 U23957 ( .A1(n27381), .A2(n27253), .B1(n27247), .B2(n21446), .ZN(
        n7907) );
  OAI22_X1 U23958 ( .A1(n27384), .A2(n27253), .B1(n27247), .B2(n21445), .ZN(
        n7908) );
  OAI22_X1 U23959 ( .A1(n27387), .A2(n27254), .B1(n27247), .B2(n21444), .ZN(
        n7909) );
  OAI22_X1 U23960 ( .A1(n27390), .A2(n27254), .B1(n27248), .B2(n21443), .ZN(
        n7910) );
  OAI22_X1 U23961 ( .A1(n27393), .A2(n27254), .B1(n27248), .B2(n21442), .ZN(
        n7911) );
  OAI22_X1 U23962 ( .A1(n27396), .A2(n27254), .B1(n27248), .B2(n21441), .ZN(
        n7912) );
  OAI22_X1 U23963 ( .A1(n27399), .A2(n27254), .B1(n27248), .B2(n21440), .ZN(
        n7913) );
  OAI22_X1 U23964 ( .A1(n27402), .A2(n27254), .B1(n27248), .B2(n21439), .ZN(
        n7914) );
  OAI22_X1 U23965 ( .A1(n27405), .A2(n27254), .B1(n27248), .B2(n21438), .ZN(
        n7915) );
  OAI22_X1 U23966 ( .A1(n27408), .A2(n27254), .B1(n27248), .B2(n21437), .ZN(
        n7916) );
  OAI22_X1 U23967 ( .A1(n27411), .A2(n27254), .B1(n27248), .B2(n21436), .ZN(
        n7917) );
  OAI22_X1 U23968 ( .A1(n27414), .A2(n27254), .B1(n27248), .B2(n21435), .ZN(
        n7918) );
  OAI22_X1 U23969 ( .A1(n27417), .A2(n27254), .B1(n27248), .B2(n21434), .ZN(
        n7919) );
  OAI22_X1 U23970 ( .A1(n27420), .A2(n27254), .B1(n27248), .B2(n21433), .ZN(
        n7920) );
  OAI22_X1 U23971 ( .A1(n27423), .A2(n27255), .B1(n27248), .B2(n21432), .ZN(
        n7921) );
  OAI22_X1 U23972 ( .A1(n27426), .A2(n27255), .B1(n27249), .B2(n21431), .ZN(
        n7922) );
  OAI22_X1 U23973 ( .A1(n27429), .A2(n27255), .B1(n27249), .B2(n21430), .ZN(
        n7923) );
  OAI22_X1 U23974 ( .A1(n27432), .A2(n27255), .B1(n27249), .B2(n21429), .ZN(
        n7924) );
  OAI22_X1 U23975 ( .A1(n27435), .A2(n27255), .B1(n27249), .B2(n21428), .ZN(
        n7925) );
  OAI22_X1 U23976 ( .A1(n27438), .A2(n27255), .B1(n27249), .B2(n21427), .ZN(
        n7926) );
  OAI22_X1 U23977 ( .A1(n27441), .A2(n27255), .B1(n27249), .B2(n21426), .ZN(
        n7927) );
  OAI22_X1 U23978 ( .A1(n27444), .A2(n27255), .B1(n27249), .B2(n21425), .ZN(
        n7928) );
  OAI22_X1 U23979 ( .A1(n27447), .A2(n27255), .B1(n27249), .B2(n21424), .ZN(
        n7929) );
  OAI22_X1 U23980 ( .A1(n27450), .A2(n27255), .B1(n27249), .B2(n21423), .ZN(
        n7930) );
  OAI22_X1 U23981 ( .A1(n27453), .A2(n27255), .B1(n27249), .B2(n21422), .ZN(
        n7931) );
  OAI22_X1 U23982 ( .A1(n27456), .A2(n27255), .B1(n27249), .B2(n21421), .ZN(
        n7932) );
  OAI22_X1 U23983 ( .A1(n27459), .A2(n27256), .B1(n27249), .B2(n21420), .ZN(
        n7933) );
  OAI22_X1 U23984 ( .A1(n27319), .A2(n27084), .B1(n27078), .B2(n21287), .ZN(
        n6990) );
  OAI22_X1 U23985 ( .A1(n27322), .A2(n27084), .B1(n27078), .B2(n21286), .ZN(
        n6991) );
  OAI22_X1 U23986 ( .A1(n27325), .A2(n27084), .B1(n27078), .B2(n21285), .ZN(
        n6992) );
  OAI22_X1 U23987 ( .A1(n27328), .A2(n27084), .B1(n27078), .B2(n21284), .ZN(
        n6993) );
  OAI22_X1 U23988 ( .A1(n27331), .A2(n27084), .B1(n27078), .B2(n21283), .ZN(
        n6994) );
  OAI22_X1 U23989 ( .A1(n27334), .A2(n27084), .B1(n27078), .B2(n21282), .ZN(
        n6995) );
  OAI22_X1 U23990 ( .A1(n27337), .A2(n27084), .B1(n27078), .B2(n21281), .ZN(
        n6996) );
  OAI22_X1 U23991 ( .A1(n27340), .A2(n27084), .B1(n27078), .B2(n21280), .ZN(
        n6997) );
  OAI22_X1 U23992 ( .A1(n27343), .A2(n27084), .B1(n27078), .B2(n21279), .ZN(
        n6998) );
  OAI22_X1 U23993 ( .A1(n27346), .A2(n27084), .B1(n27078), .B2(n21278), .ZN(
        n6999) );
  OAI22_X1 U23994 ( .A1(n27349), .A2(n27084), .B1(n27078), .B2(n21277), .ZN(
        n7000) );
  OAI22_X1 U23995 ( .A1(n27352), .A2(n27085), .B1(n27078), .B2(n21276), .ZN(
        n7001) );
  OAI22_X1 U23996 ( .A1(n27355), .A2(n27085), .B1(n27079), .B2(n21275), .ZN(
        n7002) );
  OAI22_X1 U23997 ( .A1(n27358), .A2(n27085), .B1(n27079), .B2(n21274), .ZN(
        n7003) );
  OAI22_X1 U23998 ( .A1(n27361), .A2(n27085), .B1(n27079), .B2(n21273), .ZN(
        n7004) );
  OAI22_X1 U23999 ( .A1(n27364), .A2(n27085), .B1(n27079), .B2(n21272), .ZN(
        n7005) );
  OAI22_X1 U24000 ( .A1(n27367), .A2(n27085), .B1(n27079), .B2(n21271), .ZN(
        n7006) );
  OAI22_X1 U24001 ( .A1(n27370), .A2(n27085), .B1(n27079), .B2(n21270), .ZN(
        n7007) );
  OAI22_X1 U24002 ( .A1(n27373), .A2(n27085), .B1(n27079), .B2(n21269), .ZN(
        n7008) );
  OAI22_X1 U24003 ( .A1(n27376), .A2(n27085), .B1(n27079), .B2(n21268), .ZN(
        n7009) );
  OAI22_X1 U24004 ( .A1(n27379), .A2(n27085), .B1(n27079), .B2(n21267), .ZN(
        n7010) );
  OAI22_X1 U24005 ( .A1(n27382), .A2(n27085), .B1(n27079), .B2(n21266), .ZN(
        n7011) );
  OAI22_X1 U24006 ( .A1(n27385), .A2(n27085), .B1(n27079), .B2(n21265), .ZN(
        n7012) );
  OAI22_X1 U24007 ( .A1(n27388), .A2(n27086), .B1(n27079), .B2(n21264), .ZN(
        n7013) );
  OAI22_X1 U24008 ( .A1(n27391), .A2(n27086), .B1(n27080), .B2(n21263), .ZN(
        n7014) );
  OAI22_X1 U24009 ( .A1(n27394), .A2(n27086), .B1(n27080), .B2(n21262), .ZN(
        n7015) );
  OAI22_X1 U24010 ( .A1(n27397), .A2(n27086), .B1(n27080), .B2(n21261), .ZN(
        n7016) );
  OAI22_X1 U24011 ( .A1(n27400), .A2(n27086), .B1(n27080), .B2(n21260), .ZN(
        n7017) );
  OAI22_X1 U24012 ( .A1(n27403), .A2(n27086), .B1(n27080), .B2(n21259), .ZN(
        n7018) );
  OAI22_X1 U24013 ( .A1(n27406), .A2(n27086), .B1(n27080), .B2(n21258), .ZN(
        n7019) );
  OAI22_X1 U24014 ( .A1(n27409), .A2(n27086), .B1(n27080), .B2(n21257), .ZN(
        n7020) );
  OAI22_X1 U24015 ( .A1(n27412), .A2(n27086), .B1(n27080), .B2(n21256), .ZN(
        n7021) );
  OAI22_X1 U24016 ( .A1(n27415), .A2(n27086), .B1(n27080), .B2(n21255), .ZN(
        n7022) );
  OAI22_X1 U24017 ( .A1(n27418), .A2(n27086), .B1(n27080), .B2(n21254), .ZN(
        n7023) );
  OAI22_X1 U24018 ( .A1(n27421), .A2(n27086), .B1(n27080), .B2(n21253), .ZN(
        n7024) );
  OAI22_X1 U24019 ( .A1(n27424), .A2(n27087), .B1(n27080), .B2(n21252), .ZN(
        n7025) );
  OAI22_X1 U24020 ( .A1(n27427), .A2(n27087), .B1(n27081), .B2(n21251), .ZN(
        n7026) );
  OAI22_X1 U24021 ( .A1(n27430), .A2(n27087), .B1(n27081), .B2(n21250), .ZN(
        n7027) );
  OAI22_X1 U24022 ( .A1(n27433), .A2(n27087), .B1(n27081), .B2(n21249), .ZN(
        n7028) );
  OAI22_X1 U24023 ( .A1(n27436), .A2(n27087), .B1(n27081), .B2(n21248), .ZN(
        n7029) );
  OAI22_X1 U24024 ( .A1(n27439), .A2(n27087), .B1(n27081), .B2(n21247), .ZN(
        n7030) );
  OAI22_X1 U24025 ( .A1(n27442), .A2(n27087), .B1(n27081), .B2(n21246), .ZN(
        n7031) );
  OAI22_X1 U24026 ( .A1(n27445), .A2(n27087), .B1(n27081), .B2(n21245), .ZN(
        n7032) );
  OAI22_X1 U24027 ( .A1(n27448), .A2(n27087), .B1(n27081), .B2(n21244), .ZN(
        n7033) );
  OAI22_X1 U24028 ( .A1(n27451), .A2(n27087), .B1(n27081), .B2(n21243), .ZN(
        n7034) );
  OAI22_X1 U24029 ( .A1(n27454), .A2(n27087), .B1(n27081), .B2(n21242), .ZN(
        n7035) );
  OAI22_X1 U24030 ( .A1(n27457), .A2(n27087), .B1(n27081), .B2(n21241), .ZN(
        n7036) );
  OAI22_X1 U24031 ( .A1(n27460), .A2(n27088), .B1(n27081), .B2(n21240), .ZN(
        n7037) );
  OAI22_X1 U24032 ( .A1(n27320), .A2(n26904), .B1(n26898), .B2(n20950), .ZN(
        n6030) );
  OAI22_X1 U24033 ( .A1(n27323), .A2(n26904), .B1(n26898), .B2(n20949), .ZN(
        n6031) );
  OAI22_X1 U24034 ( .A1(n27326), .A2(n26904), .B1(n26898), .B2(n20948), .ZN(
        n6032) );
  OAI22_X1 U24035 ( .A1(n27329), .A2(n26904), .B1(n26898), .B2(n20947), .ZN(
        n6033) );
  OAI22_X1 U24036 ( .A1(n27332), .A2(n26904), .B1(n26898), .B2(n20946), .ZN(
        n6034) );
  OAI22_X1 U24037 ( .A1(n27335), .A2(n26904), .B1(n26898), .B2(n20945), .ZN(
        n6035) );
  OAI22_X1 U24038 ( .A1(n27338), .A2(n26904), .B1(n26898), .B2(n20944), .ZN(
        n6036) );
  OAI22_X1 U24039 ( .A1(n27341), .A2(n26904), .B1(n26898), .B2(n20943), .ZN(
        n6037) );
  OAI22_X1 U24040 ( .A1(n27344), .A2(n26904), .B1(n26898), .B2(n20942), .ZN(
        n6038) );
  OAI22_X1 U24041 ( .A1(n27347), .A2(n26904), .B1(n26898), .B2(n20941), .ZN(
        n6039) );
  OAI22_X1 U24042 ( .A1(n27350), .A2(n26904), .B1(n26898), .B2(n20940), .ZN(
        n6040) );
  OAI22_X1 U24043 ( .A1(n27353), .A2(n26905), .B1(n26898), .B2(n20939), .ZN(
        n6041) );
  OAI22_X1 U24044 ( .A1(n27356), .A2(n26905), .B1(n26899), .B2(n20938), .ZN(
        n6042) );
  OAI22_X1 U24045 ( .A1(n27359), .A2(n26905), .B1(n26899), .B2(n20937), .ZN(
        n6043) );
  OAI22_X1 U24046 ( .A1(n27362), .A2(n26905), .B1(n26899), .B2(n20936), .ZN(
        n6044) );
  OAI22_X1 U24047 ( .A1(n27365), .A2(n26905), .B1(n26899), .B2(n20935), .ZN(
        n6045) );
  OAI22_X1 U24048 ( .A1(n27368), .A2(n26905), .B1(n26899), .B2(n20934), .ZN(
        n6046) );
  OAI22_X1 U24049 ( .A1(n27371), .A2(n26905), .B1(n26899), .B2(n20933), .ZN(
        n6047) );
  OAI22_X1 U24050 ( .A1(n27374), .A2(n26905), .B1(n26899), .B2(n20932), .ZN(
        n6048) );
  OAI22_X1 U24051 ( .A1(n27377), .A2(n26905), .B1(n26899), .B2(n20931), .ZN(
        n6049) );
  OAI22_X1 U24052 ( .A1(n27380), .A2(n26905), .B1(n26899), .B2(n20930), .ZN(
        n6050) );
  OAI22_X1 U24053 ( .A1(n27383), .A2(n26905), .B1(n26899), .B2(n20929), .ZN(
        n6051) );
  OAI22_X1 U24054 ( .A1(n27386), .A2(n26905), .B1(n26899), .B2(n20928), .ZN(
        n6052) );
  OAI22_X1 U24055 ( .A1(n27389), .A2(n26906), .B1(n26899), .B2(n20927), .ZN(
        n6053) );
  OAI22_X1 U24056 ( .A1(n27392), .A2(n26906), .B1(n26900), .B2(n20926), .ZN(
        n6054) );
  OAI22_X1 U24057 ( .A1(n27395), .A2(n26906), .B1(n26900), .B2(n20925), .ZN(
        n6055) );
  OAI22_X1 U24058 ( .A1(n27398), .A2(n26906), .B1(n26900), .B2(n20924), .ZN(
        n6056) );
  OAI22_X1 U24059 ( .A1(n27401), .A2(n26906), .B1(n26900), .B2(n20923), .ZN(
        n6057) );
  OAI22_X1 U24060 ( .A1(n27404), .A2(n26906), .B1(n26900), .B2(n20922), .ZN(
        n6058) );
  OAI22_X1 U24061 ( .A1(n27407), .A2(n26906), .B1(n26900), .B2(n20921), .ZN(
        n6059) );
  OAI22_X1 U24062 ( .A1(n27410), .A2(n26906), .B1(n26900), .B2(n20920), .ZN(
        n6060) );
  OAI22_X1 U24063 ( .A1(n27413), .A2(n26906), .B1(n26900), .B2(n20919), .ZN(
        n6061) );
  OAI22_X1 U24064 ( .A1(n27416), .A2(n26906), .B1(n26900), .B2(n20918), .ZN(
        n6062) );
  OAI22_X1 U24065 ( .A1(n27419), .A2(n26906), .B1(n26900), .B2(n20917), .ZN(
        n6063) );
  OAI22_X1 U24066 ( .A1(n27422), .A2(n26906), .B1(n26900), .B2(n20916), .ZN(
        n6064) );
  OAI22_X1 U24067 ( .A1(n27425), .A2(n26907), .B1(n26900), .B2(n20915), .ZN(
        n6065) );
  OAI22_X1 U24068 ( .A1(n27428), .A2(n26907), .B1(n26901), .B2(n20914), .ZN(
        n6066) );
  OAI22_X1 U24069 ( .A1(n27431), .A2(n26907), .B1(n26901), .B2(n20913), .ZN(
        n6067) );
  OAI22_X1 U24070 ( .A1(n27434), .A2(n26907), .B1(n26901), .B2(n20912), .ZN(
        n6068) );
  OAI22_X1 U24071 ( .A1(n27437), .A2(n26907), .B1(n26901), .B2(n20911), .ZN(
        n6069) );
  OAI22_X1 U24072 ( .A1(n27440), .A2(n26907), .B1(n26901), .B2(n20910), .ZN(
        n6070) );
  OAI22_X1 U24073 ( .A1(n27443), .A2(n26907), .B1(n26901), .B2(n20909), .ZN(
        n6071) );
  OAI22_X1 U24074 ( .A1(n27446), .A2(n26907), .B1(n26901), .B2(n20908), .ZN(
        n6072) );
  OAI22_X1 U24075 ( .A1(n27449), .A2(n26907), .B1(n26901), .B2(n20907), .ZN(
        n6073) );
  OAI22_X1 U24076 ( .A1(n27452), .A2(n26907), .B1(n26901), .B2(n20906), .ZN(
        n6074) );
  OAI22_X1 U24077 ( .A1(n27455), .A2(n26907), .B1(n26901), .B2(n20905), .ZN(
        n6075) );
  OAI22_X1 U24078 ( .A1(n27458), .A2(n26907), .B1(n26901), .B2(n20904), .ZN(
        n6076) );
  OAI22_X1 U24079 ( .A1(n27461), .A2(n26908), .B1(n26901), .B2(n20903), .ZN(
        n6077) );
  OAI22_X1 U24080 ( .A1(n27320), .A2(n26916), .B1(n26910), .B2(n20886), .ZN(
        n6094) );
  OAI22_X1 U24081 ( .A1(n27323), .A2(n26916), .B1(n26910), .B2(n20885), .ZN(
        n6095) );
  OAI22_X1 U24082 ( .A1(n27326), .A2(n26916), .B1(n26910), .B2(n20884), .ZN(
        n6096) );
  OAI22_X1 U24083 ( .A1(n27329), .A2(n26916), .B1(n26910), .B2(n20883), .ZN(
        n6097) );
  OAI22_X1 U24084 ( .A1(n27332), .A2(n26916), .B1(n26910), .B2(n20882), .ZN(
        n6098) );
  OAI22_X1 U24085 ( .A1(n27335), .A2(n26916), .B1(n26910), .B2(n20881), .ZN(
        n6099) );
  OAI22_X1 U24086 ( .A1(n27338), .A2(n26916), .B1(n26910), .B2(n20880), .ZN(
        n6100) );
  OAI22_X1 U24087 ( .A1(n27341), .A2(n26916), .B1(n26910), .B2(n20879), .ZN(
        n6101) );
  OAI22_X1 U24088 ( .A1(n27344), .A2(n26916), .B1(n26910), .B2(n20878), .ZN(
        n6102) );
  OAI22_X1 U24089 ( .A1(n27347), .A2(n26916), .B1(n26910), .B2(n20877), .ZN(
        n6103) );
  OAI22_X1 U24090 ( .A1(n27350), .A2(n26916), .B1(n26910), .B2(n20876), .ZN(
        n6104) );
  OAI22_X1 U24091 ( .A1(n27353), .A2(n26917), .B1(n26910), .B2(n20875), .ZN(
        n6105) );
  OAI22_X1 U24092 ( .A1(n27356), .A2(n26917), .B1(n26911), .B2(n20874), .ZN(
        n6106) );
  OAI22_X1 U24093 ( .A1(n27359), .A2(n26917), .B1(n26911), .B2(n20873), .ZN(
        n6107) );
  OAI22_X1 U24094 ( .A1(n27362), .A2(n26917), .B1(n26911), .B2(n20872), .ZN(
        n6108) );
  OAI22_X1 U24095 ( .A1(n27365), .A2(n26917), .B1(n26911), .B2(n20871), .ZN(
        n6109) );
  OAI22_X1 U24096 ( .A1(n27368), .A2(n26917), .B1(n26911), .B2(n20870), .ZN(
        n6110) );
  OAI22_X1 U24097 ( .A1(n27371), .A2(n26917), .B1(n26911), .B2(n20869), .ZN(
        n6111) );
  OAI22_X1 U24098 ( .A1(n27374), .A2(n26917), .B1(n26911), .B2(n20868), .ZN(
        n6112) );
  OAI22_X1 U24099 ( .A1(n27377), .A2(n26917), .B1(n26911), .B2(n20867), .ZN(
        n6113) );
  OAI22_X1 U24100 ( .A1(n27380), .A2(n26917), .B1(n26911), .B2(n20866), .ZN(
        n6114) );
  OAI22_X1 U24101 ( .A1(n27383), .A2(n26917), .B1(n26911), .B2(n20865), .ZN(
        n6115) );
  OAI22_X1 U24102 ( .A1(n27386), .A2(n26917), .B1(n26911), .B2(n20864), .ZN(
        n6116) );
  OAI22_X1 U24103 ( .A1(n27389), .A2(n26918), .B1(n26911), .B2(n20863), .ZN(
        n6117) );
  OAI22_X1 U24104 ( .A1(n27392), .A2(n26918), .B1(n26912), .B2(n20862), .ZN(
        n6118) );
  OAI22_X1 U24105 ( .A1(n27395), .A2(n26918), .B1(n26912), .B2(n20861), .ZN(
        n6119) );
  OAI22_X1 U24106 ( .A1(n27398), .A2(n26918), .B1(n26912), .B2(n20860), .ZN(
        n6120) );
  OAI22_X1 U24107 ( .A1(n27401), .A2(n26918), .B1(n26912), .B2(n20859), .ZN(
        n6121) );
  OAI22_X1 U24108 ( .A1(n27404), .A2(n26918), .B1(n26912), .B2(n20858), .ZN(
        n6122) );
  OAI22_X1 U24109 ( .A1(n27407), .A2(n26918), .B1(n26912), .B2(n20857), .ZN(
        n6123) );
  OAI22_X1 U24110 ( .A1(n27410), .A2(n26918), .B1(n26912), .B2(n20856), .ZN(
        n6124) );
  OAI22_X1 U24111 ( .A1(n27413), .A2(n26918), .B1(n26912), .B2(n20855), .ZN(
        n6125) );
  OAI22_X1 U24112 ( .A1(n27416), .A2(n26918), .B1(n26912), .B2(n20854), .ZN(
        n6126) );
  OAI22_X1 U24113 ( .A1(n27419), .A2(n26918), .B1(n26912), .B2(n20853), .ZN(
        n6127) );
  OAI22_X1 U24114 ( .A1(n27422), .A2(n26918), .B1(n26912), .B2(n20852), .ZN(
        n6128) );
  OAI22_X1 U24115 ( .A1(n27425), .A2(n26919), .B1(n26912), .B2(n20851), .ZN(
        n6129) );
  OAI22_X1 U24116 ( .A1(n27428), .A2(n26919), .B1(n26913), .B2(n20850), .ZN(
        n6130) );
  OAI22_X1 U24117 ( .A1(n27431), .A2(n26919), .B1(n26913), .B2(n20849), .ZN(
        n6131) );
  OAI22_X1 U24118 ( .A1(n27434), .A2(n26919), .B1(n26913), .B2(n20848), .ZN(
        n6132) );
  OAI22_X1 U24119 ( .A1(n27437), .A2(n26919), .B1(n26913), .B2(n20847), .ZN(
        n6133) );
  OAI22_X1 U24120 ( .A1(n27440), .A2(n26919), .B1(n26913), .B2(n20846), .ZN(
        n6134) );
  OAI22_X1 U24121 ( .A1(n27443), .A2(n26919), .B1(n26913), .B2(n20845), .ZN(
        n6135) );
  OAI22_X1 U24122 ( .A1(n27446), .A2(n26919), .B1(n26913), .B2(n20844), .ZN(
        n6136) );
  OAI22_X1 U24123 ( .A1(n27449), .A2(n26919), .B1(n26913), .B2(n20843), .ZN(
        n6137) );
  OAI22_X1 U24124 ( .A1(n27452), .A2(n26919), .B1(n26913), .B2(n20842), .ZN(
        n6138) );
  OAI22_X1 U24125 ( .A1(n27455), .A2(n26919), .B1(n26913), .B2(n20841), .ZN(
        n6139) );
  OAI22_X1 U24126 ( .A1(n27458), .A2(n26919), .B1(n26913), .B2(n20840), .ZN(
        n6140) );
  OAI22_X1 U24127 ( .A1(n27461), .A2(n26920), .B1(n26913), .B2(n20839), .ZN(
        n6141) );
  OAI22_X1 U24128 ( .A1(n27464), .A2(n26956), .B1(n26950), .B2(n22507), .ZN(
        n6334) );
  OAI22_X1 U24129 ( .A1(n27467), .A2(n26956), .B1(n26950), .B2(n22506), .ZN(
        n6335) );
  OAI22_X1 U24130 ( .A1(n27470), .A2(n26956), .B1(n26950), .B2(n22505), .ZN(
        n6336) );
  OAI22_X1 U24131 ( .A1(n27473), .A2(n26956), .B1(n26950), .B2(n22504), .ZN(
        n6337) );
  OAI22_X1 U24132 ( .A1(n27462), .A2(n27160), .B1(n27154), .B2(n22255), .ZN(
        n7422) );
  OAI22_X1 U24133 ( .A1(n27465), .A2(n27160), .B1(n27154), .B2(n22254), .ZN(
        n7423) );
  OAI22_X1 U24134 ( .A1(n27468), .A2(n27160), .B1(n27154), .B2(n22253), .ZN(
        n7424) );
  OAI22_X1 U24135 ( .A1(n27471), .A2(n27160), .B1(n27154), .B2(n22252), .ZN(
        n7425) );
  OAI22_X1 U24136 ( .A1(n27464), .A2(n26932), .B1(n26926), .B2(n22247), .ZN(
        n6206) );
  OAI22_X1 U24137 ( .A1(n27467), .A2(n26932), .B1(n26926), .B2(n22246), .ZN(
        n6207) );
  OAI22_X1 U24138 ( .A1(n27470), .A2(n26932), .B1(n26926), .B2(n22245), .ZN(
        n6208) );
  OAI22_X1 U24139 ( .A1(n27473), .A2(n26932), .B1(n26926), .B2(n22244), .ZN(
        n6209) );
  OAI22_X1 U24140 ( .A1(n27464), .A2(n26944), .B1(n26938), .B2(n22183), .ZN(
        n6270) );
  OAI22_X1 U24141 ( .A1(n27467), .A2(n26944), .B1(n26938), .B2(n22182), .ZN(
        n6271) );
  OAI22_X1 U24142 ( .A1(n27470), .A2(n26944), .B1(n26938), .B2(n22181), .ZN(
        n6272) );
  OAI22_X1 U24143 ( .A1(n27473), .A2(n26944), .B1(n26938), .B2(n22180), .ZN(
        n6273) );
  OAI22_X1 U24144 ( .A1(n27281), .A2(n27462), .B1(n27274), .B2(n21519), .ZN(
        n8062) );
  OAI22_X1 U24145 ( .A1(n27281), .A2(n27465), .B1(n27274), .B2(n21518), .ZN(
        n8063) );
  OAI22_X1 U24146 ( .A1(n27281), .A2(n27468), .B1(n27274), .B2(n21517), .ZN(
        n8064) );
  OAI22_X1 U24147 ( .A1(n27281), .A2(n27471), .B1(n27274), .B2(n21516), .ZN(
        n8065) );
  OAI22_X1 U24148 ( .A1(n27462), .A2(n27268), .B1(n27262), .B2(n21515), .ZN(
        n7998) );
  OAI22_X1 U24149 ( .A1(n27465), .A2(n27268), .B1(n27262), .B2(n21514), .ZN(
        n7999) );
  OAI22_X1 U24150 ( .A1(n27468), .A2(n27268), .B1(n27262), .B2(n21513), .ZN(
        n8000) );
  OAI22_X1 U24151 ( .A1(n27471), .A2(n27268), .B1(n27262), .B2(n21512), .ZN(
        n8001) );
  OAI22_X1 U24152 ( .A1(n27462), .A2(n27232), .B1(n27226), .B2(n21503), .ZN(
        n7806) );
  OAI22_X1 U24153 ( .A1(n27465), .A2(n27232), .B1(n27226), .B2(n21502), .ZN(
        n7807) );
  OAI22_X1 U24154 ( .A1(n27468), .A2(n27232), .B1(n27226), .B2(n21501), .ZN(
        n7808) );
  OAI22_X1 U24155 ( .A1(n27471), .A2(n27232), .B1(n27226), .B2(n21500), .ZN(
        n7809) );
  OAI22_X1 U24156 ( .A1(n27462), .A2(n27208), .B1(n27202), .B2(n21499), .ZN(
        n7678) );
  OAI22_X1 U24157 ( .A1(n27465), .A2(n27208), .B1(n27202), .B2(n21498), .ZN(
        n7679) );
  OAI22_X1 U24158 ( .A1(n27468), .A2(n27208), .B1(n27202), .B2(n21497), .ZN(
        n7680) );
  OAI22_X1 U24159 ( .A1(n27471), .A2(n27208), .B1(n27202), .B2(n21496), .ZN(
        n7681) );
  OAI22_X1 U24160 ( .A1(n27463), .A2(n27016), .B1(n27010), .B2(n21495), .ZN(
        n6654) );
  OAI22_X1 U24161 ( .A1(n27466), .A2(n27016), .B1(n27010), .B2(n21494), .ZN(
        n6655) );
  OAI22_X1 U24162 ( .A1(n27469), .A2(n27016), .B1(n27010), .B2(n21493), .ZN(
        n6656) );
  OAI22_X1 U24163 ( .A1(n27472), .A2(n27016), .B1(n27010), .B2(n21492), .ZN(
        n6657) );
  OAI22_X1 U24164 ( .A1(n27463), .A2(n27064), .B1(n27058), .B2(n21487), .ZN(
        n6910) );
  OAI22_X1 U24165 ( .A1(n27466), .A2(n27064), .B1(n27058), .B2(n21486), .ZN(
        n6911) );
  OAI22_X1 U24166 ( .A1(n27469), .A2(n27064), .B1(n27058), .B2(n21485), .ZN(
        n6912) );
  OAI22_X1 U24167 ( .A1(n27472), .A2(n27064), .B1(n27058), .B2(n21484), .ZN(
        n6913) );
  OAI22_X1 U24168 ( .A1(n27462), .A2(n27256), .B1(n27250), .B2(n21175), .ZN(
        n7934) );
  OAI22_X1 U24169 ( .A1(n27465), .A2(n27256), .B1(n27250), .B2(n21174), .ZN(
        n7935) );
  OAI22_X1 U24170 ( .A1(n27468), .A2(n27256), .B1(n27250), .B2(n21173), .ZN(
        n7936) );
  OAI22_X1 U24171 ( .A1(n27471), .A2(n27256), .B1(n27250), .B2(n21172), .ZN(
        n7937) );
  OAI22_X1 U24172 ( .A1(n27463), .A2(n27088), .B1(n27082), .B2(n21163), .ZN(
        n7038) );
  OAI22_X1 U24173 ( .A1(n27466), .A2(n27088), .B1(n27082), .B2(n21162), .ZN(
        n7039) );
  OAI22_X1 U24174 ( .A1(n27469), .A2(n27088), .B1(n27082), .B2(n21161), .ZN(
        n7040) );
  OAI22_X1 U24175 ( .A1(n27472), .A2(n27088), .B1(n27082), .B2(n21160), .ZN(
        n7041) );
  OAI22_X1 U24176 ( .A1(n27464), .A2(n26908), .B1(n26902), .B2(n20902), .ZN(
        n6078) );
  OAI22_X1 U24177 ( .A1(n27467), .A2(n26908), .B1(n26902), .B2(n20901), .ZN(
        n6079) );
  OAI22_X1 U24178 ( .A1(n27470), .A2(n26908), .B1(n26902), .B2(n20900), .ZN(
        n6080) );
  OAI22_X1 U24179 ( .A1(n27473), .A2(n26908), .B1(n26902), .B2(n20899), .ZN(
        n6081) );
  OAI22_X1 U24180 ( .A1(n27464), .A2(n26920), .B1(n26914), .B2(n20838), .ZN(
        n6142) );
  OAI22_X1 U24181 ( .A1(n27467), .A2(n26920), .B1(n26914), .B2(n20837), .ZN(
        n6143) );
  OAI22_X1 U24182 ( .A1(n27470), .A2(n26920), .B1(n26914), .B2(n20836), .ZN(
        n6144) );
  OAI22_X1 U24183 ( .A1(n27473), .A2(n26920), .B1(n26914), .B2(n20835), .ZN(
        n6145) );
  OAI22_X1 U24184 ( .A1(n27463), .A2(n27124), .B1(n9700), .B2(n27118), .ZN(
        n7230) );
  OAI22_X1 U24185 ( .A1(n27466), .A2(n27124), .B1(n9699), .B2(n27118), .ZN(
        n7231) );
  OAI22_X1 U24186 ( .A1(n27469), .A2(n27124), .B1(n9698), .B2(n27118), .ZN(
        n7232) );
  OAI22_X1 U24187 ( .A1(n27472), .A2(n27124), .B1(n9697), .B2(n27118), .ZN(
        n7233) );
  OAI22_X1 U24188 ( .A1(n27463), .A2(n27100), .B1(n9508), .B2(n27094), .ZN(
        n7102) );
  OAI22_X1 U24189 ( .A1(n27466), .A2(n27100), .B1(n9507), .B2(n27094), .ZN(
        n7103) );
  OAI22_X1 U24190 ( .A1(n27469), .A2(n27100), .B1(n9506), .B2(n27094), .ZN(
        n7104) );
  OAI22_X1 U24191 ( .A1(n27472), .A2(n27100), .B1(n9505), .B2(n27094), .ZN(
        n7105) );
  OAI22_X1 U24192 ( .A1(n27463), .A2(n27040), .B1(n9572), .B2(n27034), .ZN(
        n6782) );
  OAI22_X1 U24193 ( .A1(n27466), .A2(n27040), .B1(n9571), .B2(n27034), .ZN(
        n6783) );
  OAI22_X1 U24194 ( .A1(n27469), .A2(n27040), .B1(n9570), .B2(n27034), .ZN(
        n6784) );
  OAI22_X1 U24195 ( .A1(n27472), .A2(n27040), .B1(n9569), .B2(n27034), .ZN(
        n6785) );
  OAI22_X1 U24196 ( .A1(n27463), .A2(n27028), .B1(n9636), .B2(n27022), .ZN(
        n6718) );
  OAI22_X1 U24197 ( .A1(n27466), .A2(n27028), .B1(n9635), .B2(n27022), .ZN(
        n6719) );
  OAI22_X1 U24198 ( .A1(n27469), .A2(n27028), .B1(n9634), .B2(n27022), .ZN(
        n6720) );
  OAI22_X1 U24199 ( .A1(n27472), .A2(n27028), .B1(n9633), .B2(n27022), .ZN(
        n6721) );
  AOI22_X1 U24200 ( .A1(n26488), .A2(n25578), .B1(n26482), .B2(n25566), .ZN(
        n24011) );
  AOI22_X1 U24201 ( .A1(n26483), .A2(n25655), .B1(n26477), .B2(n25643), .ZN(
        n25162) );
  AOI22_X1 U24202 ( .A1(n26483), .A2(n25656), .B1(n26477), .B2(n25644), .ZN(
        n25134) );
  AOI22_X1 U24203 ( .A1(n26483), .A2(n25657), .B1(n26477), .B2(n25645), .ZN(
        n25116) );
  AOI22_X1 U24204 ( .A1(n26483), .A2(n25658), .B1(n26477), .B2(n25646), .ZN(
        n25098) );
  AOI22_X1 U24205 ( .A1(n26483), .A2(n25659), .B1(n26477), .B2(n25647), .ZN(
        n25080) );
  AOI22_X1 U24206 ( .A1(n26483), .A2(n25660), .B1(n26477), .B2(n25648), .ZN(
        n25062) );
  AOI22_X1 U24207 ( .A1(n26483), .A2(n25661), .B1(n26477), .B2(n25649), .ZN(
        n25044) );
  AOI22_X1 U24208 ( .A1(n26483), .A2(n25662), .B1(n26477), .B2(n25650), .ZN(
        n25026) );
  AOI22_X1 U24209 ( .A1(n26483), .A2(n25663), .B1(n26477), .B2(n25651), .ZN(
        n25008) );
  AOI22_X1 U24210 ( .A1(n26483), .A2(n25664), .B1(n26477), .B2(n25652), .ZN(
        n24990) );
  AOI22_X1 U24211 ( .A1(n26483), .A2(n25665), .B1(n26477), .B2(n25653), .ZN(
        n24972) );
  AOI22_X1 U24212 ( .A1(n26483), .A2(n25666), .B1(n26477), .B2(n25654), .ZN(
        n24954) );
  AOI22_X1 U24213 ( .A1(n26484), .A2(n25455), .B1(n26478), .B2(n25311), .ZN(
        n24936) );
  AOI22_X1 U24214 ( .A1(n26484), .A2(n25456), .B1(n26478), .B2(n25312), .ZN(
        n24918) );
  AOI22_X1 U24215 ( .A1(n26484), .A2(n25457), .B1(n26478), .B2(n25313), .ZN(
        n24900) );
  AOI22_X1 U24216 ( .A1(n26484), .A2(n25458), .B1(n26478), .B2(n25314), .ZN(
        n24882) );
  AOI22_X1 U24217 ( .A1(n26484), .A2(n25459), .B1(n26478), .B2(n25315), .ZN(
        n24864) );
  AOI22_X1 U24218 ( .A1(n26484), .A2(n25460), .B1(n26478), .B2(n25316), .ZN(
        n24846) );
  AOI22_X1 U24219 ( .A1(n26484), .A2(n25461), .B1(n26478), .B2(n25317), .ZN(
        n24828) );
  AOI22_X1 U24220 ( .A1(n26484), .A2(n25462), .B1(n26478), .B2(n25318), .ZN(
        n24810) );
  AOI22_X1 U24221 ( .A1(n26484), .A2(n25463), .B1(n26478), .B2(n25319), .ZN(
        n24792) );
  AOI22_X1 U24222 ( .A1(n26484), .A2(n25464), .B1(n26478), .B2(n25320), .ZN(
        n24774) );
  AOI22_X1 U24223 ( .A1(n26484), .A2(n25465), .B1(n26478), .B2(n25321), .ZN(
        n24756) );
  AOI22_X1 U24224 ( .A1(n26484), .A2(n25466), .B1(n26478), .B2(n25322), .ZN(
        n24738) );
  AOI22_X1 U24225 ( .A1(n26485), .A2(n25467), .B1(n26479), .B2(n25323), .ZN(
        n24720) );
  AOI22_X1 U24226 ( .A1(n26485), .A2(n25468), .B1(n26479), .B2(n25324), .ZN(
        n24702) );
  AOI22_X1 U24227 ( .A1(n26485), .A2(n25469), .B1(n26479), .B2(n25325), .ZN(
        n24684) );
  AOI22_X1 U24228 ( .A1(n26485), .A2(n25470), .B1(n26479), .B2(n25326), .ZN(
        n24666) );
  AOI22_X1 U24229 ( .A1(n26485), .A2(n25471), .B1(n26479), .B2(n25327), .ZN(
        n24648) );
  AOI22_X1 U24230 ( .A1(n26485), .A2(n25472), .B1(n26479), .B2(n25328), .ZN(
        n24630) );
  AOI22_X1 U24231 ( .A1(n26485), .A2(n25473), .B1(n26479), .B2(n25329), .ZN(
        n24612) );
  AOI22_X1 U24232 ( .A1(n26485), .A2(n25474), .B1(n26479), .B2(n25330), .ZN(
        n24594) );
  AOI22_X1 U24233 ( .A1(n26485), .A2(n25475), .B1(n26479), .B2(n25331), .ZN(
        n24576) );
  AOI22_X1 U24234 ( .A1(n26485), .A2(n25476), .B1(n26479), .B2(n25332), .ZN(
        n24558) );
  AOI22_X1 U24235 ( .A1(n26485), .A2(n25477), .B1(n26479), .B2(n25333), .ZN(
        n24540) );
  AOI22_X1 U24236 ( .A1(n26485), .A2(n25478), .B1(n26479), .B2(n25334), .ZN(
        n24522) );
  AOI22_X1 U24237 ( .A1(n26486), .A2(n25479), .B1(n26480), .B2(n25335), .ZN(
        n24504) );
  AOI22_X1 U24238 ( .A1(n26486), .A2(n25480), .B1(n26480), .B2(n25336), .ZN(
        n24486) );
  AOI22_X1 U24239 ( .A1(n26486), .A2(n25481), .B1(n26480), .B2(n25337), .ZN(
        n24468) );
  AOI22_X1 U24240 ( .A1(n26486), .A2(n25482), .B1(n26480), .B2(n25338), .ZN(
        n24450) );
  AOI22_X1 U24241 ( .A1(n26486), .A2(n25483), .B1(n26480), .B2(n25339), .ZN(
        n24432) );
  AOI22_X1 U24242 ( .A1(n26486), .A2(n25484), .B1(n26480), .B2(n25340), .ZN(
        n24414) );
  AOI22_X1 U24243 ( .A1(n26486), .A2(n25485), .B1(n26480), .B2(n25341), .ZN(
        n24396) );
  AOI22_X1 U24244 ( .A1(n26486), .A2(n25486), .B1(n26480), .B2(n25342), .ZN(
        n24378) );
  AOI22_X1 U24245 ( .A1(n26486), .A2(n25487), .B1(n26480), .B2(n25343), .ZN(
        n24360) );
  AOI22_X1 U24246 ( .A1(n26486), .A2(n25488), .B1(n26480), .B2(n25344), .ZN(
        n24342) );
  AOI22_X1 U24247 ( .A1(n26486), .A2(n25489), .B1(n26480), .B2(n25345), .ZN(
        n24324) );
  AOI22_X1 U24248 ( .A1(n26486), .A2(n25490), .B1(n26480), .B2(n25346), .ZN(
        n24306) );
  AOI22_X1 U24249 ( .A1(n26487), .A2(n25491), .B1(n26481), .B2(n25347), .ZN(
        n24288) );
  AOI22_X1 U24250 ( .A1(n26487), .A2(n25492), .B1(n26481), .B2(n25348), .ZN(
        n24270) );
  AOI22_X1 U24251 ( .A1(n26487), .A2(n25493), .B1(n26481), .B2(n25349), .ZN(
        n24252) );
  AOI22_X1 U24252 ( .A1(n26487), .A2(n25494), .B1(n26481), .B2(n25350), .ZN(
        n24234) );
  AOI22_X1 U24253 ( .A1(n26487), .A2(n25495), .B1(n26481), .B2(n25351), .ZN(
        n24216) );
  AOI22_X1 U24254 ( .A1(n26487), .A2(n25496), .B1(n26481), .B2(n25352), .ZN(
        n24198) );
  AOI22_X1 U24255 ( .A1(n26487), .A2(n25497), .B1(n26481), .B2(n25353), .ZN(
        n24180) );
  AOI22_X1 U24256 ( .A1(n26487), .A2(n25498), .B1(n26481), .B2(n25354), .ZN(
        n24162) );
  AOI22_X1 U24257 ( .A1(n26487), .A2(n25499), .B1(n26481), .B2(n25355), .ZN(
        n24144) );
  AOI22_X1 U24258 ( .A1(n26487), .A2(n25500), .B1(n26481), .B2(n25356), .ZN(
        n24126) );
  AOI22_X1 U24259 ( .A1(n26487), .A2(n25501), .B1(n26481), .B2(n25357), .ZN(
        n24108) );
  AOI22_X1 U24260 ( .A1(n26487), .A2(n25502), .B1(n26481), .B2(n25358), .ZN(
        n24090) );
  AOI22_X1 U24261 ( .A1(n26488), .A2(n25575), .B1(n26482), .B2(n25563), .ZN(
        n24072) );
  AOI22_X1 U24262 ( .A1(n26488), .A2(n25576), .B1(n26482), .B2(n25564), .ZN(
        n24054) );
  AOI22_X1 U24263 ( .A1(n26488), .A2(n25577), .B1(n26482), .B2(n25565), .ZN(
        n24036) );
  AOI22_X1 U24264 ( .A1(n26708), .A2(n25655), .B1(n26702), .B2(n25643), .ZN(
        n23963) );
  AOI22_X1 U24265 ( .A1(n26708), .A2(n25656), .B1(n26702), .B2(n25644), .ZN(
        n23935) );
  AOI22_X1 U24266 ( .A1(n26708), .A2(n25657), .B1(n26702), .B2(n25645), .ZN(
        n23917) );
  AOI22_X1 U24267 ( .A1(n26708), .A2(n25658), .B1(n26702), .B2(n25646), .ZN(
        n23899) );
  AOI22_X1 U24268 ( .A1(n26708), .A2(n25659), .B1(n26702), .B2(n25647), .ZN(
        n23881) );
  AOI22_X1 U24269 ( .A1(n26708), .A2(n25660), .B1(n26702), .B2(n25648), .ZN(
        n23863) );
  AOI22_X1 U24270 ( .A1(n26708), .A2(n25661), .B1(n26702), .B2(n25649), .ZN(
        n23845) );
  AOI22_X1 U24271 ( .A1(n26708), .A2(n25662), .B1(n26702), .B2(n25650), .ZN(
        n23827) );
  AOI22_X1 U24272 ( .A1(n26708), .A2(n25663), .B1(n26702), .B2(n25651), .ZN(
        n23809) );
  AOI22_X1 U24273 ( .A1(n26708), .A2(n25664), .B1(n26702), .B2(n25652), .ZN(
        n23791) );
  AOI22_X1 U24274 ( .A1(n26708), .A2(n25665), .B1(n26702), .B2(n25653), .ZN(
        n23773) );
  AOI22_X1 U24275 ( .A1(n26708), .A2(n25666), .B1(n26702), .B2(n25654), .ZN(
        n23755) );
  AOI22_X1 U24276 ( .A1(n26709), .A2(n25455), .B1(n26703), .B2(n25311), .ZN(
        n23737) );
  AOI22_X1 U24277 ( .A1(n26709), .A2(n25456), .B1(n26703), .B2(n25312), .ZN(
        n23719) );
  AOI22_X1 U24278 ( .A1(n26709), .A2(n25457), .B1(n26703), .B2(n25313), .ZN(
        n23701) );
  AOI22_X1 U24279 ( .A1(n26709), .A2(n25458), .B1(n26703), .B2(n25314), .ZN(
        n23683) );
  AOI22_X1 U24280 ( .A1(n26709), .A2(n25459), .B1(n26703), .B2(n25315), .ZN(
        n23665) );
  AOI22_X1 U24281 ( .A1(n26709), .A2(n25460), .B1(n26703), .B2(n25316), .ZN(
        n23647) );
  AOI22_X1 U24282 ( .A1(n26709), .A2(n25461), .B1(n26703), .B2(n25317), .ZN(
        n23629) );
  AOI22_X1 U24283 ( .A1(n26709), .A2(n25462), .B1(n26703), .B2(n25318), .ZN(
        n23611) );
  AOI22_X1 U24284 ( .A1(n26709), .A2(n25463), .B1(n26703), .B2(n25319), .ZN(
        n23593) );
  AOI22_X1 U24285 ( .A1(n26709), .A2(n25464), .B1(n26703), .B2(n25320), .ZN(
        n23575) );
  AOI22_X1 U24286 ( .A1(n26709), .A2(n25465), .B1(n26703), .B2(n25321), .ZN(
        n23557) );
  AOI22_X1 U24287 ( .A1(n26709), .A2(n25466), .B1(n26703), .B2(n25322), .ZN(
        n23539) );
  AOI22_X1 U24288 ( .A1(n26710), .A2(n25467), .B1(n26704), .B2(n25323), .ZN(
        n23521) );
  AOI22_X1 U24289 ( .A1(n26710), .A2(n25468), .B1(n26704), .B2(n25324), .ZN(
        n23503) );
  AOI22_X1 U24290 ( .A1(n26710), .A2(n25469), .B1(n26704), .B2(n25325), .ZN(
        n23485) );
  AOI22_X1 U24291 ( .A1(n26710), .A2(n25470), .B1(n26704), .B2(n25326), .ZN(
        n23467) );
  AOI22_X1 U24292 ( .A1(n26710), .A2(n25471), .B1(n26704), .B2(n25327), .ZN(
        n23449) );
  AOI22_X1 U24293 ( .A1(n26710), .A2(n25472), .B1(n26704), .B2(n25328), .ZN(
        n23431) );
  AOI22_X1 U24294 ( .A1(n26710), .A2(n25473), .B1(n26704), .B2(n25329), .ZN(
        n23413) );
  AOI22_X1 U24295 ( .A1(n26710), .A2(n25474), .B1(n26704), .B2(n25330), .ZN(
        n23395) );
  AOI22_X1 U24296 ( .A1(n26710), .A2(n25475), .B1(n26704), .B2(n25331), .ZN(
        n23377) );
  AOI22_X1 U24297 ( .A1(n26710), .A2(n25476), .B1(n26704), .B2(n25332), .ZN(
        n23359) );
  AOI22_X1 U24298 ( .A1(n26710), .A2(n25477), .B1(n26704), .B2(n25333), .ZN(
        n23341) );
  AOI22_X1 U24299 ( .A1(n26710), .A2(n25478), .B1(n26704), .B2(n25334), .ZN(
        n23323) );
  AOI22_X1 U24300 ( .A1(n26711), .A2(n25479), .B1(n26705), .B2(n25335), .ZN(
        n23305) );
  AOI22_X1 U24301 ( .A1(n26711), .A2(n25480), .B1(n26705), .B2(n25336), .ZN(
        n23287) );
  AOI22_X1 U24302 ( .A1(n26711), .A2(n25481), .B1(n26705), .B2(n25337), .ZN(
        n23269) );
  AOI22_X1 U24303 ( .A1(n26711), .A2(n25482), .B1(n26705), .B2(n25338), .ZN(
        n23251) );
  AOI22_X1 U24304 ( .A1(n26711), .A2(n25483), .B1(n26705), .B2(n25339), .ZN(
        n23233) );
  AOI22_X1 U24305 ( .A1(n26711), .A2(n25484), .B1(n26705), .B2(n25340), .ZN(
        n23215) );
  AOI22_X1 U24306 ( .A1(n26711), .A2(n25485), .B1(n26705), .B2(n25341), .ZN(
        n23197) );
  AOI22_X1 U24307 ( .A1(n26711), .A2(n25486), .B1(n26705), .B2(n25342), .ZN(
        n23179) );
  AOI22_X1 U24308 ( .A1(n26711), .A2(n25487), .B1(n26705), .B2(n25343), .ZN(
        n23161) );
  AOI22_X1 U24309 ( .A1(n26711), .A2(n25488), .B1(n26705), .B2(n25344), .ZN(
        n23143) );
  AOI22_X1 U24310 ( .A1(n26711), .A2(n25489), .B1(n26705), .B2(n25345), .ZN(
        n23125) );
  AOI22_X1 U24311 ( .A1(n26711), .A2(n25490), .B1(n26705), .B2(n25346), .ZN(
        n23107) );
  AOI22_X1 U24312 ( .A1(n26712), .A2(n25491), .B1(n26706), .B2(n25347), .ZN(
        n23089) );
  AOI22_X1 U24313 ( .A1(n26712), .A2(n25492), .B1(n26706), .B2(n25348), .ZN(
        n23071) );
  AOI22_X1 U24314 ( .A1(n26712), .A2(n25493), .B1(n26706), .B2(n25349), .ZN(
        n23053) );
  AOI22_X1 U24315 ( .A1(n26712), .A2(n25494), .B1(n26706), .B2(n25350), .ZN(
        n23035) );
  AOI22_X1 U24316 ( .A1(n26712), .A2(n25495), .B1(n26706), .B2(n25351), .ZN(
        n23017) );
  AOI22_X1 U24317 ( .A1(n26712), .A2(n25496), .B1(n26706), .B2(n25352), .ZN(
        n22999) );
  AOI22_X1 U24318 ( .A1(n26712), .A2(n25497), .B1(n26706), .B2(n25353), .ZN(
        n22981) );
  AOI22_X1 U24319 ( .A1(n26712), .A2(n25498), .B1(n26706), .B2(n25354), .ZN(
        n22963) );
  AOI22_X1 U24320 ( .A1(n26712), .A2(n25499), .B1(n26706), .B2(n25355), .ZN(
        n22945) );
  AOI22_X1 U24321 ( .A1(n26712), .A2(n25500), .B1(n26706), .B2(n25356), .ZN(
        n22927) );
  AOI22_X1 U24322 ( .A1(n26712), .A2(n25501), .B1(n26706), .B2(n25357), .ZN(
        n22909) );
  AOI22_X1 U24323 ( .A1(n26712), .A2(n25502), .B1(n26706), .B2(n25358), .ZN(
        n22891) );
  AOI22_X1 U24324 ( .A1(n26713), .A2(n25575), .B1(n26707), .B2(n25563), .ZN(
        n22873) );
  AOI22_X1 U24325 ( .A1(n26713), .A2(n25576), .B1(n26707), .B2(n25564), .ZN(
        n22855) );
  AOI22_X1 U24326 ( .A1(n26713), .A2(n25577), .B1(n26707), .B2(n25565), .ZN(
        n22837) );
  AOI22_X1 U24327 ( .A1(n26713), .A2(n25578), .B1(n26707), .B2(n25566), .ZN(
        n22812) );
  OAI221_X1 U24328 ( .B1(n9584), .B2(n26622), .C1(n20786), .C2(n26616), .A(
        n24280), .ZN(n24275) );
  AOI22_X1 U24329 ( .A1(n26610), .A2(n25941), .B1(n26604), .B2(n20986), .ZN(
        n24280) );
  OAI221_X1 U24330 ( .B1(n9583), .B2(n26622), .C1(n20785), .C2(n26616), .A(
        n24262), .ZN(n24257) );
  AOI22_X1 U24331 ( .A1(n26610), .A2(n25946), .B1(n26604), .B2(n20985), .ZN(
        n24262) );
  OAI221_X1 U24332 ( .B1(n9582), .B2(n26622), .C1(n20784), .C2(n26616), .A(
        n24244), .ZN(n24239) );
  AOI22_X1 U24333 ( .A1(n26610), .A2(n25951), .B1(n26604), .B2(n20984), .ZN(
        n24244) );
  OAI221_X1 U24334 ( .B1(n9581), .B2(n26622), .C1(n20783), .C2(n26616), .A(
        n24226), .ZN(n24221) );
  AOI22_X1 U24335 ( .A1(n26610), .A2(n25956), .B1(n26604), .B2(n20983), .ZN(
        n24226) );
  OAI221_X1 U24336 ( .B1(n9580), .B2(n26622), .C1(n20782), .C2(n26616), .A(
        n24208), .ZN(n24203) );
  AOI22_X1 U24337 ( .A1(n26610), .A2(n25961), .B1(n26604), .B2(n20982), .ZN(
        n24208) );
  OAI221_X1 U24338 ( .B1(n9579), .B2(n26622), .C1(n20781), .C2(n26616), .A(
        n24190), .ZN(n24185) );
  AOI22_X1 U24339 ( .A1(n26610), .A2(n25966), .B1(n26604), .B2(n20981), .ZN(
        n24190) );
  OAI221_X1 U24340 ( .B1(n9578), .B2(n26622), .C1(n20780), .C2(n26616), .A(
        n24172), .ZN(n24167) );
  AOI22_X1 U24341 ( .A1(n26610), .A2(n25971), .B1(n26604), .B2(n20980), .ZN(
        n24172) );
  OAI221_X1 U24342 ( .B1(n9577), .B2(n26622), .C1(n20779), .C2(n26616), .A(
        n24154), .ZN(n24149) );
  AOI22_X1 U24343 ( .A1(n26610), .A2(n25976), .B1(n26604), .B2(n20979), .ZN(
        n24154) );
  OAI221_X1 U24344 ( .B1(n9576), .B2(n26622), .C1(n20778), .C2(n26616), .A(
        n24136), .ZN(n24131) );
  AOI22_X1 U24345 ( .A1(n26610), .A2(n25981), .B1(n26604), .B2(n20978), .ZN(
        n24136) );
  OAI221_X1 U24346 ( .B1(n9575), .B2(n26622), .C1(n20777), .C2(n26616), .A(
        n24118), .ZN(n24113) );
  AOI22_X1 U24347 ( .A1(n26610), .A2(n25986), .B1(n26604), .B2(n20977), .ZN(
        n24118) );
  OAI221_X1 U24348 ( .B1(n9574), .B2(n26622), .C1(n20776), .C2(n26616), .A(
        n24100), .ZN(n24095) );
  AOI22_X1 U24349 ( .A1(n26610), .A2(n25991), .B1(n26604), .B2(n20976), .ZN(
        n24100) );
  OAI221_X1 U24350 ( .B1(n9573), .B2(n26622), .C1(n20775), .C2(n26616), .A(
        n24082), .ZN(n24077) );
  AOI22_X1 U24351 ( .A1(n26610), .A2(n25996), .B1(n26604), .B2(n20975), .ZN(
        n24082) );
  OAI221_X1 U24352 ( .B1(n9584), .B2(n26847), .C1(n20786), .C2(n26841), .A(
        n23081), .ZN(n23076) );
  AOI22_X1 U24353 ( .A1(n26835), .A2(n25941), .B1(n26829), .B2(n20986), .ZN(
        n23081) );
  OAI221_X1 U24354 ( .B1(n9583), .B2(n26847), .C1(n20785), .C2(n26841), .A(
        n23063), .ZN(n23058) );
  AOI22_X1 U24355 ( .A1(n26835), .A2(n25946), .B1(n26829), .B2(n20985), .ZN(
        n23063) );
  OAI221_X1 U24356 ( .B1(n9582), .B2(n26847), .C1(n20784), .C2(n26841), .A(
        n23045), .ZN(n23040) );
  AOI22_X1 U24357 ( .A1(n26835), .A2(n25951), .B1(n26829), .B2(n20984), .ZN(
        n23045) );
  OAI221_X1 U24358 ( .B1(n9581), .B2(n26847), .C1(n20783), .C2(n26841), .A(
        n23027), .ZN(n23022) );
  AOI22_X1 U24359 ( .A1(n26835), .A2(n25956), .B1(n26829), .B2(n20983), .ZN(
        n23027) );
  OAI221_X1 U24360 ( .B1(n9580), .B2(n26847), .C1(n20782), .C2(n26841), .A(
        n23009), .ZN(n23004) );
  AOI22_X1 U24361 ( .A1(n26835), .A2(n25961), .B1(n26829), .B2(n20982), .ZN(
        n23009) );
  OAI221_X1 U24362 ( .B1(n9579), .B2(n26847), .C1(n20781), .C2(n26841), .A(
        n22991), .ZN(n22986) );
  AOI22_X1 U24363 ( .A1(n26835), .A2(n25966), .B1(n26829), .B2(n20981), .ZN(
        n22991) );
  OAI221_X1 U24364 ( .B1(n9578), .B2(n26847), .C1(n20780), .C2(n26841), .A(
        n22973), .ZN(n22968) );
  AOI22_X1 U24365 ( .A1(n26835), .A2(n25971), .B1(n26829), .B2(n20980), .ZN(
        n22973) );
  OAI221_X1 U24366 ( .B1(n9577), .B2(n26847), .C1(n20779), .C2(n26841), .A(
        n22955), .ZN(n22950) );
  AOI22_X1 U24367 ( .A1(n26835), .A2(n25976), .B1(n26829), .B2(n20979), .ZN(
        n22955) );
  OAI221_X1 U24368 ( .B1(n9576), .B2(n26847), .C1(n20778), .C2(n26841), .A(
        n22937), .ZN(n22932) );
  AOI22_X1 U24369 ( .A1(n26835), .A2(n25981), .B1(n26829), .B2(n20978), .ZN(
        n22937) );
  OAI221_X1 U24370 ( .B1(n9575), .B2(n26847), .C1(n20777), .C2(n26841), .A(
        n22919), .ZN(n22914) );
  AOI22_X1 U24371 ( .A1(n26835), .A2(n25986), .B1(n26829), .B2(n20977), .ZN(
        n22919) );
  OAI221_X1 U24372 ( .B1(n9574), .B2(n26847), .C1(n20776), .C2(n26841), .A(
        n22901), .ZN(n22896) );
  AOI22_X1 U24373 ( .A1(n26835), .A2(n25991), .B1(n26829), .B2(n20976), .ZN(
        n22901) );
  OAI221_X1 U24374 ( .B1(n9573), .B2(n26847), .C1(n20775), .C2(n26841), .A(
        n22883), .ZN(n22878) );
  AOI22_X1 U24375 ( .A1(n26835), .A2(n25996), .B1(n26829), .B2(n20975), .ZN(
        n22883) );
  OAI22_X1 U24376 ( .A1(n27283), .A2(n27035), .B1(n9632), .B2(n27029), .ZN(
        n6722) );
  OAI22_X1 U24377 ( .A1(n27286), .A2(n27035), .B1(n9631), .B2(n27029), .ZN(
        n6723) );
  OAI22_X1 U24378 ( .A1(n27289), .A2(n27035), .B1(n9630), .B2(n27029), .ZN(
        n6724) );
  OAI22_X1 U24379 ( .A1(n27292), .A2(n27035), .B1(n9629), .B2(n27029), .ZN(
        n6725) );
  OAI22_X1 U24380 ( .A1(n27295), .A2(n27035), .B1(n9628), .B2(n27029), .ZN(
        n6726) );
  OAI22_X1 U24381 ( .A1(n27298), .A2(n27035), .B1(n9627), .B2(n27029), .ZN(
        n6727) );
  OAI22_X1 U24382 ( .A1(n27301), .A2(n27035), .B1(n9626), .B2(n27029), .ZN(
        n6728) );
  OAI22_X1 U24383 ( .A1(n27304), .A2(n27035), .B1(n9625), .B2(n27029), .ZN(
        n6729) );
  OAI22_X1 U24384 ( .A1(n27307), .A2(n27035), .B1(n9624), .B2(n27029), .ZN(
        n6730) );
  OAI22_X1 U24385 ( .A1(n27310), .A2(n27035), .B1(n9623), .B2(n27029), .ZN(
        n6731) );
  OAI22_X1 U24386 ( .A1(n27313), .A2(n27035), .B1(n9622), .B2(n27029), .ZN(
        n6732) );
  OAI22_X1 U24387 ( .A1(n27316), .A2(n27036), .B1(n9621), .B2(n27029), .ZN(
        n6733) );
  OAI22_X1 U24388 ( .A1(n27319), .A2(n27036), .B1(n9620), .B2(n27030), .ZN(
        n6734) );
  OAI22_X1 U24389 ( .A1(n27322), .A2(n27036), .B1(n9619), .B2(n27030), .ZN(
        n6735) );
  OAI22_X1 U24390 ( .A1(n27325), .A2(n27036), .B1(n9618), .B2(n27030), .ZN(
        n6736) );
  OAI22_X1 U24391 ( .A1(n27328), .A2(n27036), .B1(n9617), .B2(n27030), .ZN(
        n6737) );
  OAI22_X1 U24392 ( .A1(n27331), .A2(n27036), .B1(n9616), .B2(n27030), .ZN(
        n6738) );
  OAI22_X1 U24393 ( .A1(n27334), .A2(n27036), .B1(n9615), .B2(n27030), .ZN(
        n6739) );
  OAI22_X1 U24394 ( .A1(n27337), .A2(n27036), .B1(n9614), .B2(n27030), .ZN(
        n6740) );
  OAI22_X1 U24395 ( .A1(n27340), .A2(n27036), .B1(n9613), .B2(n27030), .ZN(
        n6741) );
  OAI22_X1 U24396 ( .A1(n27343), .A2(n27036), .B1(n9612), .B2(n27030), .ZN(
        n6742) );
  OAI22_X1 U24397 ( .A1(n27346), .A2(n27036), .B1(n9611), .B2(n27030), .ZN(
        n6743) );
  OAI22_X1 U24398 ( .A1(n27349), .A2(n27036), .B1(n9610), .B2(n27030), .ZN(
        n6744) );
  OAI22_X1 U24399 ( .A1(n27352), .A2(n27037), .B1(n9609), .B2(n27030), .ZN(
        n6745) );
  OAI22_X1 U24400 ( .A1(n27355), .A2(n27037), .B1(n9608), .B2(n27031), .ZN(
        n6746) );
  OAI22_X1 U24401 ( .A1(n27358), .A2(n27037), .B1(n9607), .B2(n27031), .ZN(
        n6747) );
  OAI22_X1 U24402 ( .A1(n27361), .A2(n27037), .B1(n9606), .B2(n27031), .ZN(
        n6748) );
  OAI22_X1 U24403 ( .A1(n27364), .A2(n27037), .B1(n9605), .B2(n27031), .ZN(
        n6749) );
  OAI22_X1 U24404 ( .A1(n27367), .A2(n27037), .B1(n9604), .B2(n27031), .ZN(
        n6750) );
  OAI22_X1 U24405 ( .A1(n27370), .A2(n27037), .B1(n9603), .B2(n27031), .ZN(
        n6751) );
  OAI22_X1 U24406 ( .A1(n27373), .A2(n27037), .B1(n9602), .B2(n27031), .ZN(
        n6752) );
  OAI22_X1 U24407 ( .A1(n27376), .A2(n27037), .B1(n9601), .B2(n27031), .ZN(
        n6753) );
  OAI22_X1 U24408 ( .A1(n27379), .A2(n27037), .B1(n9600), .B2(n27031), .ZN(
        n6754) );
  OAI22_X1 U24409 ( .A1(n27382), .A2(n27037), .B1(n9599), .B2(n27031), .ZN(
        n6755) );
  OAI22_X1 U24410 ( .A1(n27385), .A2(n27037), .B1(n9598), .B2(n27031), .ZN(
        n6756) );
  OAI22_X1 U24411 ( .A1(n27388), .A2(n27038), .B1(n9597), .B2(n27031), .ZN(
        n6757) );
  OAI22_X1 U24412 ( .A1(n27391), .A2(n27038), .B1(n9596), .B2(n27032), .ZN(
        n6758) );
  OAI22_X1 U24413 ( .A1(n27394), .A2(n27038), .B1(n9595), .B2(n27032), .ZN(
        n6759) );
  OAI22_X1 U24414 ( .A1(n27397), .A2(n27038), .B1(n9594), .B2(n27032), .ZN(
        n6760) );
  OAI22_X1 U24415 ( .A1(n27400), .A2(n27038), .B1(n9593), .B2(n27032), .ZN(
        n6761) );
  OAI22_X1 U24416 ( .A1(n27403), .A2(n27038), .B1(n9592), .B2(n27032), .ZN(
        n6762) );
  OAI22_X1 U24417 ( .A1(n27406), .A2(n27038), .B1(n9591), .B2(n27032), .ZN(
        n6763) );
  OAI22_X1 U24418 ( .A1(n27409), .A2(n27038), .B1(n9590), .B2(n27032), .ZN(
        n6764) );
  OAI22_X1 U24419 ( .A1(n27412), .A2(n27038), .B1(n9589), .B2(n27032), .ZN(
        n6765) );
  OAI22_X1 U24420 ( .A1(n27415), .A2(n27038), .B1(n9588), .B2(n27032), .ZN(
        n6766) );
  OAI22_X1 U24421 ( .A1(n27418), .A2(n27038), .B1(n9587), .B2(n27032), .ZN(
        n6767) );
  OAI22_X1 U24422 ( .A1(n27421), .A2(n27038), .B1(n9586), .B2(n27032), .ZN(
        n6768) );
  OAI22_X1 U24423 ( .A1(n27424), .A2(n27039), .B1(n9585), .B2(n27032), .ZN(
        n6769) );
  OAI22_X1 U24424 ( .A1(n27427), .A2(n27039), .B1(n9584), .B2(n27033), .ZN(
        n6770) );
  OAI22_X1 U24425 ( .A1(n27430), .A2(n27039), .B1(n9583), .B2(n27033), .ZN(
        n6771) );
  OAI22_X1 U24426 ( .A1(n27433), .A2(n27039), .B1(n9582), .B2(n27033), .ZN(
        n6772) );
  OAI22_X1 U24427 ( .A1(n27436), .A2(n27039), .B1(n9581), .B2(n27033), .ZN(
        n6773) );
  OAI22_X1 U24428 ( .A1(n27439), .A2(n27039), .B1(n9580), .B2(n27033), .ZN(
        n6774) );
  OAI22_X1 U24429 ( .A1(n27442), .A2(n27039), .B1(n9579), .B2(n27033), .ZN(
        n6775) );
  OAI22_X1 U24430 ( .A1(n27445), .A2(n27039), .B1(n9578), .B2(n27033), .ZN(
        n6776) );
  OAI22_X1 U24431 ( .A1(n27448), .A2(n27039), .B1(n9577), .B2(n27033), .ZN(
        n6777) );
  OAI22_X1 U24432 ( .A1(n27451), .A2(n27039), .B1(n9576), .B2(n27033), .ZN(
        n6778) );
  OAI22_X1 U24433 ( .A1(n27454), .A2(n27039), .B1(n9575), .B2(n27033), .ZN(
        n6779) );
  OAI22_X1 U24434 ( .A1(n27457), .A2(n27039), .B1(n9574), .B2(n27033), .ZN(
        n6780) );
  OAI22_X1 U24435 ( .A1(n27460), .A2(n27040), .B1(n9573), .B2(n27033), .ZN(
        n6781) );
  OAI22_X1 U24436 ( .A1(n27283), .A2(n27119), .B1(n9760), .B2(n27113), .ZN(
        n7170) );
  OAI22_X1 U24437 ( .A1(n27286), .A2(n27119), .B1(n9759), .B2(n27113), .ZN(
        n7171) );
  OAI22_X1 U24438 ( .A1(n27289), .A2(n27119), .B1(n9758), .B2(n27113), .ZN(
        n7172) );
  OAI22_X1 U24439 ( .A1(n27292), .A2(n27119), .B1(n9757), .B2(n27113), .ZN(
        n7173) );
  OAI22_X1 U24440 ( .A1(n27295), .A2(n27119), .B1(n9756), .B2(n27113), .ZN(
        n7174) );
  OAI22_X1 U24441 ( .A1(n27298), .A2(n27119), .B1(n9755), .B2(n27113), .ZN(
        n7175) );
  OAI22_X1 U24442 ( .A1(n27301), .A2(n27119), .B1(n9754), .B2(n27113), .ZN(
        n7176) );
  OAI22_X1 U24443 ( .A1(n27304), .A2(n27119), .B1(n9753), .B2(n27113), .ZN(
        n7177) );
  OAI22_X1 U24444 ( .A1(n27307), .A2(n27119), .B1(n9752), .B2(n27113), .ZN(
        n7178) );
  OAI22_X1 U24445 ( .A1(n27310), .A2(n27119), .B1(n9751), .B2(n27113), .ZN(
        n7179) );
  OAI22_X1 U24446 ( .A1(n27313), .A2(n27119), .B1(n9750), .B2(n27113), .ZN(
        n7180) );
  OAI22_X1 U24447 ( .A1(n27316), .A2(n27120), .B1(n9749), .B2(n27113), .ZN(
        n7181) );
  OAI22_X1 U24448 ( .A1(n27319), .A2(n27120), .B1(n9748), .B2(n27114), .ZN(
        n7182) );
  OAI22_X1 U24449 ( .A1(n27322), .A2(n27120), .B1(n9747), .B2(n27114), .ZN(
        n7183) );
  OAI22_X1 U24450 ( .A1(n27325), .A2(n27120), .B1(n9746), .B2(n27114), .ZN(
        n7184) );
  OAI22_X1 U24451 ( .A1(n27328), .A2(n27120), .B1(n9745), .B2(n27114), .ZN(
        n7185) );
  OAI22_X1 U24452 ( .A1(n27331), .A2(n27120), .B1(n9744), .B2(n27114), .ZN(
        n7186) );
  OAI22_X1 U24453 ( .A1(n27334), .A2(n27120), .B1(n9743), .B2(n27114), .ZN(
        n7187) );
  OAI22_X1 U24454 ( .A1(n27337), .A2(n27120), .B1(n9742), .B2(n27114), .ZN(
        n7188) );
  OAI22_X1 U24455 ( .A1(n27340), .A2(n27120), .B1(n9741), .B2(n27114), .ZN(
        n7189) );
  OAI22_X1 U24456 ( .A1(n27343), .A2(n27120), .B1(n9740), .B2(n27114), .ZN(
        n7190) );
  OAI22_X1 U24457 ( .A1(n27346), .A2(n27120), .B1(n9739), .B2(n27114), .ZN(
        n7191) );
  OAI22_X1 U24458 ( .A1(n27349), .A2(n27120), .B1(n9738), .B2(n27114), .ZN(
        n7192) );
  OAI22_X1 U24459 ( .A1(n27352), .A2(n27121), .B1(n9737), .B2(n27114), .ZN(
        n7193) );
  OAI22_X1 U24460 ( .A1(n27355), .A2(n27121), .B1(n9736), .B2(n27115), .ZN(
        n7194) );
  OAI22_X1 U24461 ( .A1(n27358), .A2(n27121), .B1(n9735), .B2(n27115), .ZN(
        n7195) );
  OAI22_X1 U24462 ( .A1(n27361), .A2(n27121), .B1(n9734), .B2(n27115), .ZN(
        n7196) );
  OAI22_X1 U24463 ( .A1(n27364), .A2(n27121), .B1(n9733), .B2(n27115), .ZN(
        n7197) );
  OAI22_X1 U24464 ( .A1(n27367), .A2(n27121), .B1(n9732), .B2(n27115), .ZN(
        n7198) );
  OAI22_X1 U24465 ( .A1(n27370), .A2(n27121), .B1(n9731), .B2(n27115), .ZN(
        n7199) );
  OAI22_X1 U24466 ( .A1(n27373), .A2(n27121), .B1(n9730), .B2(n27115), .ZN(
        n7200) );
  OAI22_X1 U24467 ( .A1(n27376), .A2(n27121), .B1(n9729), .B2(n27115), .ZN(
        n7201) );
  OAI22_X1 U24468 ( .A1(n27379), .A2(n27121), .B1(n9728), .B2(n27115), .ZN(
        n7202) );
  OAI22_X1 U24469 ( .A1(n27382), .A2(n27121), .B1(n9727), .B2(n27115), .ZN(
        n7203) );
  OAI22_X1 U24470 ( .A1(n27385), .A2(n27121), .B1(n9726), .B2(n27115), .ZN(
        n7204) );
  OAI22_X1 U24471 ( .A1(n27388), .A2(n27122), .B1(n9725), .B2(n27115), .ZN(
        n7205) );
  OAI22_X1 U24472 ( .A1(n27391), .A2(n27122), .B1(n9724), .B2(n27116), .ZN(
        n7206) );
  OAI22_X1 U24473 ( .A1(n27394), .A2(n27122), .B1(n9723), .B2(n27116), .ZN(
        n7207) );
  OAI22_X1 U24474 ( .A1(n27397), .A2(n27122), .B1(n9722), .B2(n27116), .ZN(
        n7208) );
  OAI22_X1 U24475 ( .A1(n27400), .A2(n27122), .B1(n9721), .B2(n27116), .ZN(
        n7209) );
  OAI22_X1 U24476 ( .A1(n27403), .A2(n27122), .B1(n9720), .B2(n27116), .ZN(
        n7210) );
  OAI22_X1 U24477 ( .A1(n27406), .A2(n27122), .B1(n9719), .B2(n27116), .ZN(
        n7211) );
  OAI22_X1 U24478 ( .A1(n27409), .A2(n27122), .B1(n9718), .B2(n27116), .ZN(
        n7212) );
  OAI22_X1 U24479 ( .A1(n27412), .A2(n27122), .B1(n9717), .B2(n27116), .ZN(
        n7213) );
  OAI22_X1 U24480 ( .A1(n27415), .A2(n27122), .B1(n9716), .B2(n27116), .ZN(
        n7214) );
  OAI22_X1 U24481 ( .A1(n27418), .A2(n27122), .B1(n9715), .B2(n27116), .ZN(
        n7215) );
  OAI22_X1 U24482 ( .A1(n27421), .A2(n27122), .B1(n9714), .B2(n27116), .ZN(
        n7216) );
  OAI22_X1 U24483 ( .A1(n27424), .A2(n27123), .B1(n9713), .B2(n27116), .ZN(
        n7217) );
  OAI22_X1 U24484 ( .A1(n27427), .A2(n27123), .B1(n9712), .B2(n27117), .ZN(
        n7218) );
  OAI22_X1 U24485 ( .A1(n27430), .A2(n27123), .B1(n9711), .B2(n27117), .ZN(
        n7219) );
  OAI22_X1 U24486 ( .A1(n27433), .A2(n27123), .B1(n9710), .B2(n27117), .ZN(
        n7220) );
  OAI22_X1 U24487 ( .A1(n27436), .A2(n27123), .B1(n9709), .B2(n27117), .ZN(
        n7221) );
  OAI22_X1 U24488 ( .A1(n27439), .A2(n27123), .B1(n9708), .B2(n27117), .ZN(
        n7222) );
  OAI22_X1 U24489 ( .A1(n27442), .A2(n27123), .B1(n9707), .B2(n27117), .ZN(
        n7223) );
  OAI22_X1 U24490 ( .A1(n27445), .A2(n27123), .B1(n9706), .B2(n27117), .ZN(
        n7224) );
  OAI22_X1 U24491 ( .A1(n27448), .A2(n27123), .B1(n9705), .B2(n27117), .ZN(
        n7225) );
  OAI22_X1 U24492 ( .A1(n27451), .A2(n27123), .B1(n9704), .B2(n27117), .ZN(
        n7226) );
  OAI22_X1 U24493 ( .A1(n27454), .A2(n27123), .B1(n9703), .B2(n27117), .ZN(
        n7227) );
  OAI22_X1 U24494 ( .A1(n27457), .A2(n27123), .B1(n9702), .B2(n27117), .ZN(
        n7228) );
  OAI22_X1 U24495 ( .A1(n27460), .A2(n27124), .B1(n9701), .B2(n27117), .ZN(
        n7229) );
  OAI22_X1 U24496 ( .A1(n27283), .A2(n27095), .B1(n9568), .B2(n27089), .ZN(
        n7042) );
  OAI22_X1 U24497 ( .A1(n27286), .A2(n27095), .B1(n9567), .B2(n27089), .ZN(
        n7043) );
  OAI22_X1 U24498 ( .A1(n27289), .A2(n27095), .B1(n9566), .B2(n27089), .ZN(
        n7044) );
  OAI22_X1 U24499 ( .A1(n27292), .A2(n27095), .B1(n9565), .B2(n27089), .ZN(
        n7045) );
  OAI22_X1 U24500 ( .A1(n27295), .A2(n27095), .B1(n9564), .B2(n27089), .ZN(
        n7046) );
  OAI22_X1 U24501 ( .A1(n27298), .A2(n27095), .B1(n9563), .B2(n27089), .ZN(
        n7047) );
  OAI22_X1 U24502 ( .A1(n27301), .A2(n27095), .B1(n9562), .B2(n27089), .ZN(
        n7048) );
  OAI22_X1 U24503 ( .A1(n27304), .A2(n27095), .B1(n9561), .B2(n27089), .ZN(
        n7049) );
  OAI22_X1 U24504 ( .A1(n27307), .A2(n27095), .B1(n9560), .B2(n27089), .ZN(
        n7050) );
  OAI22_X1 U24505 ( .A1(n27310), .A2(n27095), .B1(n9559), .B2(n27089), .ZN(
        n7051) );
  OAI22_X1 U24506 ( .A1(n27313), .A2(n27095), .B1(n9558), .B2(n27089), .ZN(
        n7052) );
  OAI22_X1 U24507 ( .A1(n27316), .A2(n27096), .B1(n9557), .B2(n27089), .ZN(
        n7053) );
  OAI22_X1 U24508 ( .A1(n27319), .A2(n27096), .B1(n9556), .B2(n27090), .ZN(
        n7054) );
  OAI22_X1 U24509 ( .A1(n27322), .A2(n27096), .B1(n9555), .B2(n27090), .ZN(
        n7055) );
  OAI22_X1 U24510 ( .A1(n27325), .A2(n27096), .B1(n9554), .B2(n27090), .ZN(
        n7056) );
  OAI22_X1 U24511 ( .A1(n27328), .A2(n27096), .B1(n9553), .B2(n27090), .ZN(
        n7057) );
  OAI22_X1 U24512 ( .A1(n27331), .A2(n27096), .B1(n9552), .B2(n27090), .ZN(
        n7058) );
  OAI22_X1 U24513 ( .A1(n27334), .A2(n27096), .B1(n9551), .B2(n27090), .ZN(
        n7059) );
  OAI22_X1 U24514 ( .A1(n27337), .A2(n27096), .B1(n9550), .B2(n27090), .ZN(
        n7060) );
  OAI22_X1 U24515 ( .A1(n27340), .A2(n27096), .B1(n9549), .B2(n27090), .ZN(
        n7061) );
  OAI22_X1 U24516 ( .A1(n27343), .A2(n27096), .B1(n9548), .B2(n27090), .ZN(
        n7062) );
  OAI22_X1 U24517 ( .A1(n27346), .A2(n27096), .B1(n9547), .B2(n27090), .ZN(
        n7063) );
  OAI22_X1 U24518 ( .A1(n27349), .A2(n27096), .B1(n9546), .B2(n27090), .ZN(
        n7064) );
  OAI22_X1 U24519 ( .A1(n27352), .A2(n27097), .B1(n9545), .B2(n27090), .ZN(
        n7065) );
  OAI22_X1 U24520 ( .A1(n27355), .A2(n27097), .B1(n9544), .B2(n27091), .ZN(
        n7066) );
  OAI22_X1 U24521 ( .A1(n27358), .A2(n27097), .B1(n9543), .B2(n27091), .ZN(
        n7067) );
  OAI22_X1 U24522 ( .A1(n27361), .A2(n27097), .B1(n9542), .B2(n27091), .ZN(
        n7068) );
  OAI22_X1 U24523 ( .A1(n27364), .A2(n27097), .B1(n9541), .B2(n27091), .ZN(
        n7069) );
  OAI22_X1 U24524 ( .A1(n27367), .A2(n27097), .B1(n9540), .B2(n27091), .ZN(
        n7070) );
  OAI22_X1 U24525 ( .A1(n27370), .A2(n27097), .B1(n9539), .B2(n27091), .ZN(
        n7071) );
  OAI22_X1 U24526 ( .A1(n27373), .A2(n27097), .B1(n9538), .B2(n27091), .ZN(
        n7072) );
  OAI22_X1 U24527 ( .A1(n27376), .A2(n27097), .B1(n9537), .B2(n27091), .ZN(
        n7073) );
  OAI22_X1 U24528 ( .A1(n27379), .A2(n27097), .B1(n9536), .B2(n27091), .ZN(
        n7074) );
  OAI22_X1 U24529 ( .A1(n27382), .A2(n27097), .B1(n9535), .B2(n27091), .ZN(
        n7075) );
  OAI22_X1 U24530 ( .A1(n27385), .A2(n27097), .B1(n9534), .B2(n27091), .ZN(
        n7076) );
  OAI22_X1 U24531 ( .A1(n27388), .A2(n27098), .B1(n9533), .B2(n27091), .ZN(
        n7077) );
  OAI22_X1 U24532 ( .A1(n27391), .A2(n27098), .B1(n9532), .B2(n27092), .ZN(
        n7078) );
  OAI22_X1 U24533 ( .A1(n27394), .A2(n27098), .B1(n9531), .B2(n27092), .ZN(
        n7079) );
  OAI22_X1 U24534 ( .A1(n27397), .A2(n27098), .B1(n9530), .B2(n27092), .ZN(
        n7080) );
  OAI22_X1 U24535 ( .A1(n27400), .A2(n27098), .B1(n9529), .B2(n27092), .ZN(
        n7081) );
  OAI22_X1 U24536 ( .A1(n27403), .A2(n27098), .B1(n9528), .B2(n27092), .ZN(
        n7082) );
  OAI22_X1 U24537 ( .A1(n27406), .A2(n27098), .B1(n9527), .B2(n27092), .ZN(
        n7083) );
  OAI22_X1 U24538 ( .A1(n27409), .A2(n27098), .B1(n9526), .B2(n27092), .ZN(
        n7084) );
  OAI22_X1 U24539 ( .A1(n27412), .A2(n27098), .B1(n9525), .B2(n27092), .ZN(
        n7085) );
  OAI22_X1 U24540 ( .A1(n27415), .A2(n27098), .B1(n9524), .B2(n27092), .ZN(
        n7086) );
  OAI22_X1 U24541 ( .A1(n27418), .A2(n27098), .B1(n9523), .B2(n27092), .ZN(
        n7087) );
  OAI22_X1 U24542 ( .A1(n27421), .A2(n27098), .B1(n9522), .B2(n27092), .ZN(
        n7088) );
  OAI22_X1 U24543 ( .A1(n27424), .A2(n27099), .B1(n9521), .B2(n27092), .ZN(
        n7089) );
  OAI22_X1 U24544 ( .A1(n27427), .A2(n27099), .B1(n9520), .B2(n27093), .ZN(
        n7090) );
  OAI22_X1 U24545 ( .A1(n27430), .A2(n27099), .B1(n9519), .B2(n27093), .ZN(
        n7091) );
  OAI22_X1 U24546 ( .A1(n27433), .A2(n27099), .B1(n9518), .B2(n27093), .ZN(
        n7092) );
  OAI22_X1 U24547 ( .A1(n27436), .A2(n27099), .B1(n9517), .B2(n27093), .ZN(
        n7093) );
  OAI22_X1 U24548 ( .A1(n27439), .A2(n27099), .B1(n9516), .B2(n27093), .ZN(
        n7094) );
  OAI22_X1 U24549 ( .A1(n27442), .A2(n27099), .B1(n9515), .B2(n27093), .ZN(
        n7095) );
  OAI22_X1 U24550 ( .A1(n27445), .A2(n27099), .B1(n9514), .B2(n27093), .ZN(
        n7096) );
  OAI22_X1 U24551 ( .A1(n27448), .A2(n27099), .B1(n9513), .B2(n27093), .ZN(
        n7097) );
  OAI22_X1 U24552 ( .A1(n27451), .A2(n27099), .B1(n9512), .B2(n27093), .ZN(
        n7098) );
  OAI22_X1 U24553 ( .A1(n27454), .A2(n27099), .B1(n9511), .B2(n27093), .ZN(
        n7099) );
  OAI22_X1 U24554 ( .A1(n27457), .A2(n27099), .B1(n9510), .B2(n27093), .ZN(
        n7100) );
  OAI22_X1 U24555 ( .A1(n27460), .A2(n27100), .B1(n9509), .B2(n27093), .ZN(
        n7101) );
  OAI22_X1 U24556 ( .A1(n27283), .A2(n27023), .B1(n9696), .B2(n27017), .ZN(
        n6658) );
  OAI22_X1 U24557 ( .A1(n27286), .A2(n27023), .B1(n9695), .B2(n27017), .ZN(
        n6659) );
  OAI22_X1 U24558 ( .A1(n27289), .A2(n27023), .B1(n9694), .B2(n27017), .ZN(
        n6660) );
  OAI22_X1 U24559 ( .A1(n27292), .A2(n27023), .B1(n9693), .B2(n27017), .ZN(
        n6661) );
  OAI22_X1 U24560 ( .A1(n27295), .A2(n27023), .B1(n9692), .B2(n27017), .ZN(
        n6662) );
  OAI22_X1 U24561 ( .A1(n27298), .A2(n27023), .B1(n9691), .B2(n27017), .ZN(
        n6663) );
  OAI22_X1 U24562 ( .A1(n27301), .A2(n27023), .B1(n9690), .B2(n27017), .ZN(
        n6664) );
  OAI22_X1 U24563 ( .A1(n27304), .A2(n27023), .B1(n9689), .B2(n27017), .ZN(
        n6665) );
  OAI22_X1 U24564 ( .A1(n27307), .A2(n27023), .B1(n9688), .B2(n27017), .ZN(
        n6666) );
  OAI22_X1 U24565 ( .A1(n27310), .A2(n27023), .B1(n9687), .B2(n27017), .ZN(
        n6667) );
  OAI22_X1 U24566 ( .A1(n27313), .A2(n27023), .B1(n9686), .B2(n27017), .ZN(
        n6668) );
  OAI22_X1 U24567 ( .A1(n27316), .A2(n27024), .B1(n9685), .B2(n27017), .ZN(
        n6669) );
  OAI22_X1 U24568 ( .A1(n27319), .A2(n27024), .B1(n9684), .B2(n27018), .ZN(
        n6670) );
  OAI22_X1 U24569 ( .A1(n27322), .A2(n27024), .B1(n9683), .B2(n27018), .ZN(
        n6671) );
  OAI22_X1 U24570 ( .A1(n27325), .A2(n27024), .B1(n9682), .B2(n27018), .ZN(
        n6672) );
  OAI22_X1 U24571 ( .A1(n27328), .A2(n27024), .B1(n9681), .B2(n27018), .ZN(
        n6673) );
  OAI22_X1 U24572 ( .A1(n27331), .A2(n27024), .B1(n9680), .B2(n27018), .ZN(
        n6674) );
  OAI22_X1 U24573 ( .A1(n27334), .A2(n27024), .B1(n9679), .B2(n27018), .ZN(
        n6675) );
  OAI22_X1 U24574 ( .A1(n27337), .A2(n27024), .B1(n9678), .B2(n27018), .ZN(
        n6676) );
  OAI22_X1 U24575 ( .A1(n27340), .A2(n27024), .B1(n9677), .B2(n27018), .ZN(
        n6677) );
  OAI22_X1 U24576 ( .A1(n27343), .A2(n27024), .B1(n9676), .B2(n27018), .ZN(
        n6678) );
  OAI22_X1 U24577 ( .A1(n27346), .A2(n27024), .B1(n9675), .B2(n27018), .ZN(
        n6679) );
  OAI22_X1 U24578 ( .A1(n27349), .A2(n27024), .B1(n9674), .B2(n27018), .ZN(
        n6680) );
  OAI22_X1 U24579 ( .A1(n27352), .A2(n27025), .B1(n9673), .B2(n27018), .ZN(
        n6681) );
  OAI22_X1 U24580 ( .A1(n27355), .A2(n27025), .B1(n9672), .B2(n27019), .ZN(
        n6682) );
  OAI22_X1 U24581 ( .A1(n27358), .A2(n27025), .B1(n9671), .B2(n27019), .ZN(
        n6683) );
  OAI22_X1 U24582 ( .A1(n27361), .A2(n27025), .B1(n9670), .B2(n27019), .ZN(
        n6684) );
  OAI22_X1 U24583 ( .A1(n27364), .A2(n27025), .B1(n9669), .B2(n27019), .ZN(
        n6685) );
  OAI22_X1 U24584 ( .A1(n27367), .A2(n27025), .B1(n9668), .B2(n27019), .ZN(
        n6686) );
  OAI22_X1 U24585 ( .A1(n27370), .A2(n27025), .B1(n9667), .B2(n27019), .ZN(
        n6687) );
  OAI22_X1 U24586 ( .A1(n27373), .A2(n27025), .B1(n9666), .B2(n27019), .ZN(
        n6688) );
  OAI22_X1 U24587 ( .A1(n27376), .A2(n27025), .B1(n9665), .B2(n27019), .ZN(
        n6689) );
  OAI22_X1 U24588 ( .A1(n27379), .A2(n27025), .B1(n9664), .B2(n27019), .ZN(
        n6690) );
  OAI22_X1 U24589 ( .A1(n27382), .A2(n27025), .B1(n9663), .B2(n27019), .ZN(
        n6691) );
  OAI22_X1 U24590 ( .A1(n27385), .A2(n27025), .B1(n9662), .B2(n27019), .ZN(
        n6692) );
  OAI22_X1 U24591 ( .A1(n27388), .A2(n27026), .B1(n9661), .B2(n27019), .ZN(
        n6693) );
  OAI22_X1 U24592 ( .A1(n27391), .A2(n27026), .B1(n9660), .B2(n27020), .ZN(
        n6694) );
  OAI22_X1 U24593 ( .A1(n27394), .A2(n27026), .B1(n9659), .B2(n27020), .ZN(
        n6695) );
  OAI22_X1 U24594 ( .A1(n27397), .A2(n27026), .B1(n9658), .B2(n27020), .ZN(
        n6696) );
  OAI22_X1 U24595 ( .A1(n27400), .A2(n27026), .B1(n9657), .B2(n27020), .ZN(
        n6697) );
  OAI22_X1 U24596 ( .A1(n27403), .A2(n27026), .B1(n9656), .B2(n27020), .ZN(
        n6698) );
  OAI22_X1 U24597 ( .A1(n27406), .A2(n27026), .B1(n9655), .B2(n27020), .ZN(
        n6699) );
  OAI22_X1 U24598 ( .A1(n27409), .A2(n27026), .B1(n9654), .B2(n27020), .ZN(
        n6700) );
  OAI22_X1 U24599 ( .A1(n27412), .A2(n27026), .B1(n9653), .B2(n27020), .ZN(
        n6701) );
  OAI22_X1 U24600 ( .A1(n27415), .A2(n27026), .B1(n9652), .B2(n27020), .ZN(
        n6702) );
  OAI22_X1 U24601 ( .A1(n27418), .A2(n27026), .B1(n9651), .B2(n27020), .ZN(
        n6703) );
  OAI22_X1 U24602 ( .A1(n27421), .A2(n27026), .B1(n9650), .B2(n27020), .ZN(
        n6704) );
  OAI22_X1 U24603 ( .A1(n27424), .A2(n27027), .B1(n9649), .B2(n27020), .ZN(
        n6705) );
  OAI22_X1 U24604 ( .A1(n27427), .A2(n27027), .B1(n9648), .B2(n27021), .ZN(
        n6706) );
  OAI22_X1 U24605 ( .A1(n27430), .A2(n27027), .B1(n9647), .B2(n27021), .ZN(
        n6707) );
  OAI22_X1 U24606 ( .A1(n27433), .A2(n27027), .B1(n9646), .B2(n27021), .ZN(
        n6708) );
  OAI22_X1 U24607 ( .A1(n27436), .A2(n27027), .B1(n9645), .B2(n27021), .ZN(
        n6709) );
  OAI22_X1 U24608 ( .A1(n27439), .A2(n27027), .B1(n9644), .B2(n27021), .ZN(
        n6710) );
  OAI22_X1 U24609 ( .A1(n27442), .A2(n27027), .B1(n9643), .B2(n27021), .ZN(
        n6711) );
  OAI22_X1 U24610 ( .A1(n27445), .A2(n27027), .B1(n9642), .B2(n27021), .ZN(
        n6712) );
  OAI22_X1 U24611 ( .A1(n27448), .A2(n27027), .B1(n9641), .B2(n27021), .ZN(
        n6713) );
  OAI22_X1 U24612 ( .A1(n27451), .A2(n27027), .B1(n9640), .B2(n27021), .ZN(
        n6714) );
  OAI22_X1 U24613 ( .A1(n27454), .A2(n27027), .B1(n9639), .B2(n27021), .ZN(
        n6715) );
  OAI22_X1 U24614 ( .A1(n27457), .A2(n27027), .B1(n9638), .B2(n27021), .ZN(
        n6716) );
  OAI22_X1 U24615 ( .A1(n27460), .A2(n27028), .B1(n9637), .B2(n27021), .ZN(
        n6717) );
  OAI22_X1 U24616 ( .A1(n27284), .A2(n26951), .B1(n26945), .B2(n22631), .ZN(
        n6274) );
  OAI22_X1 U24617 ( .A1(n27287), .A2(n26951), .B1(n26945), .B2(n22630), .ZN(
        n6275) );
  OAI22_X1 U24618 ( .A1(n27290), .A2(n26951), .B1(n26945), .B2(n22629), .ZN(
        n6276) );
  OAI22_X1 U24619 ( .A1(n27293), .A2(n26951), .B1(n26945), .B2(n22628), .ZN(
        n6277) );
  OAI22_X1 U24620 ( .A1(n27296), .A2(n26951), .B1(n26945), .B2(n22627), .ZN(
        n6278) );
  OAI22_X1 U24621 ( .A1(n27299), .A2(n26951), .B1(n26945), .B2(n22626), .ZN(
        n6279) );
  OAI22_X1 U24622 ( .A1(n27302), .A2(n26951), .B1(n26945), .B2(n22625), .ZN(
        n6280) );
  OAI22_X1 U24623 ( .A1(n27305), .A2(n26951), .B1(n26945), .B2(n22624), .ZN(
        n6281) );
  OAI22_X1 U24624 ( .A1(n27308), .A2(n26951), .B1(n26945), .B2(n22623), .ZN(
        n6282) );
  OAI22_X1 U24625 ( .A1(n27311), .A2(n26951), .B1(n26945), .B2(n22622), .ZN(
        n6283) );
  OAI22_X1 U24626 ( .A1(n27314), .A2(n26951), .B1(n26945), .B2(n22621), .ZN(
        n6284) );
  OAI22_X1 U24627 ( .A1(n27317), .A2(n26952), .B1(n26945), .B2(n22620), .ZN(
        n6285) );
  OAI22_X1 U24628 ( .A1(n27282), .A2(n27155), .B1(n27149), .B2(n22439), .ZN(
        n7362) );
  OAI22_X1 U24629 ( .A1(n27285), .A2(n27155), .B1(n27149), .B2(n22438), .ZN(
        n7363) );
  OAI22_X1 U24630 ( .A1(n27288), .A2(n27155), .B1(n27149), .B2(n22437), .ZN(
        n7364) );
  OAI22_X1 U24631 ( .A1(n27291), .A2(n27155), .B1(n27149), .B2(n22436), .ZN(
        n7365) );
  OAI22_X1 U24632 ( .A1(n27294), .A2(n27155), .B1(n27149), .B2(n22435), .ZN(
        n7366) );
  OAI22_X1 U24633 ( .A1(n27297), .A2(n27155), .B1(n27149), .B2(n22434), .ZN(
        n7367) );
  OAI22_X1 U24634 ( .A1(n27300), .A2(n27155), .B1(n27149), .B2(n22433), .ZN(
        n7368) );
  OAI22_X1 U24635 ( .A1(n27303), .A2(n27155), .B1(n27149), .B2(n22432), .ZN(
        n7369) );
  OAI22_X1 U24636 ( .A1(n27306), .A2(n27155), .B1(n27149), .B2(n22431), .ZN(
        n7370) );
  OAI22_X1 U24637 ( .A1(n27309), .A2(n27155), .B1(n27149), .B2(n22430), .ZN(
        n7371) );
  OAI22_X1 U24638 ( .A1(n27312), .A2(n27155), .B1(n27149), .B2(n22429), .ZN(
        n7372) );
  OAI22_X1 U24639 ( .A1(n27315), .A2(n27156), .B1(n27149), .B2(n22428), .ZN(
        n7373) );
  OAI22_X1 U24640 ( .A1(n27284), .A2(n26927), .B1(n26921), .B2(n22319), .ZN(
        n6146) );
  OAI22_X1 U24641 ( .A1(n27287), .A2(n26927), .B1(n26921), .B2(n22318), .ZN(
        n6147) );
  OAI22_X1 U24642 ( .A1(n27290), .A2(n26927), .B1(n26921), .B2(n22317), .ZN(
        n6148) );
  OAI22_X1 U24643 ( .A1(n27293), .A2(n26927), .B1(n26921), .B2(n22316), .ZN(
        n6149) );
  OAI22_X1 U24644 ( .A1(n27296), .A2(n26927), .B1(n26921), .B2(n22315), .ZN(
        n6150) );
  OAI22_X1 U24645 ( .A1(n27299), .A2(n26927), .B1(n26921), .B2(n22314), .ZN(
        n6151) );
  OAI22_X1 U24646 ( .A1(n27302), .A2(n26927), .B1(n26921), .B2(n22313), .ZN(
        n6152) );
  OAI22_X1 U24647 ( .A1(n27305), .A2(n26927), .B1(n26921), .B2(n22312), .ZN(
        n6153) );
  OAI22_X1 U24648 ( .A1(n27308), .A2(n26927), .B1(n26921), .B2(n22311), .ZN(
        n6154) );
  OAI22_X1 U24649 ( .A1(n27311), .A2(n26927), .B1(n26921), .B2(n22310), .ZN(
        n6155) );
  OAI22_X1 U24650 ( .A1(n27314), .A2(n26927), .B1(n26921), .B2(n22309), .ZN(
        n6156) );
  OAI22_X1 U24651 ( .A1(n27317), .A2(n26928), .B1(n26921), .B2(n22308), .ZN(
        n6157) );
  OAI22_X1 U24652 ( .A1(n27284), .A2(n26939), .B1(n26933), .B2(n22243), .ZN(
        n6210) );
  OAI22_X1 U24653 ( .A1(n27287), .A2(n26939), .B1(n26933), .B2(n22242), .ZN(
        n6211) );
  OAI22_X1 U24654 ( .A1(n27290), .A2(n26939), .B1(n26933), .B2(n22241), .ZN(
        n6212) );
  OAI22_X1 U24655 ( .A1(n27293), .A2(n26939), .B1(n26933), .B2(n22240), .ZN(
        n6213) );
  OAI22_X1 U24656 ( .A1(n27296), .A2(n26939), .B1(n26933), .B2(n22239), .ZN(
        n6214) );
  OAI22_X1 U24657 ( .A1(n27299), .A2(n26939), .B1(n26933), .B2(n22238), .ZN(
        n6215) );
  OAI22_X1 U24658 ( .A1(n27302), .A2(n26939), .B1(n26933), .B2(n22237), .ZN(
        n6216) );
  OAI22_X1 U24659 ( .A1(n27305), .A2(n26939), .B1(n26933), .B2(n22236), .ZN(
        n6217) );
  OAI22_X1 U24660 ( .A1(n27308), .A2(n26939), .B1(n26933), .B2(n22235), .ZN(
        n6218) );
  OAI22_X1 U24661 ( .A1(n27311), .A2(n26939), .B1(n26933), .B2(n22234), .ZN(
        n6219) );
  OAI22_X1 U24662 ( .A1(n27314), .A2(n26939), .B1(n26933), .B2(n22233), .ZN(
        n6220) );
  OAI22_X1 U24663 ( .A1(n27317), .A2(n26940), .B1(n26933), .B2(n22232), .ZN(
        n6221) );
  OAI22_X1 U24664 ( .A1(n27277), .A2(n27282), .B1(n27269), .B2(n22179), .ZN(
        n8002) );
  OAI22_X1 U24665 ( .A1(n27277), .A2(n27285), .B1(n27269), .B2(n22178), .ZN(
        n8003) );
  OAI22_X1 U24666 ( .A1(n27277), .A2(n27288), .B1(n27269), .B2(n22177), .ZN(
        n8004) );
  OAI22_X1 U24667 ( .A1(n27277), .A2(n27291), .B1(n27269), .B2(n22176), .ZN(
        n8005) );
  OAI22_X1 U24668 ( .A1(n27277), .A2(n27294), .B1(n27269), .B2(n22175), .ZN(
        n8006) );
  OAI22_X1 U24669 ( .A1(n27277), .A2(n27297), .B1(n27269), .B2(n22174), .ZN(
        n8007) );
  OAI22_X1 U24670 ( .A1(n27277), .A2(n27300), .B1(n27269), .B2(n22173), .ZN(
        n8008) );
  OAI22_X1 U24671 ( .A1(n27277), .A2(n27303), .B1(n27269), .B2(n22172), .ZN(
        n8009) );
  OAI22_X1 U24672 ( .A1(n27277), .A2(n27306), .B1(n27269), .B2(n22171), .ZN(
        n8010) );
  OAI22_X1 U24673 ( .A1(n27277), .A2(n27309), .B1(n27269), .B2(n22170), .ZN(
        n8011) );
  OAI22_X1 U24674 ( .A1(n27277), .A2(n27312), .B1(n27269), .B2(n22169), .ZN(
        n8012) );
  OAI22_X1 U24675 ( .A1(n27277), .A2(n27315), .B1(n27269), .B2(n22168), .ZN(
        n8013) );
  OAI22_X1 U24676 ( .A1(n27282), .A2(n27263), .B1(n27257), .B2(n22119), .ZN(
        n7938) );
  OAI22_X1 U24677 ( .A1(n27285), .A2(n27263), .B1(n27257), .B2(n22118), .ZN(
        n7939) );
  OAI22_X1 U24678 ( .A1(n27288), .A2(n27263), .B1(n27257), .B2(n22117), .ZN(
        n7940) );
  OAI22_X1 U24679 ( .A1(n27291), .A2(n27263), .B1(n27257), .B2(n22116), .ZN(
        n7941) );
  OAI22_X1 U24680 ( .A1(n27294), .A2(n27263), .B1(n27257), .B2(n22115), .ZN(
        n7942) );
  OAI22_X1 U24681 ( .A1(n27297), .A2(n27263), .B1(n27257), .B2(n22114), .ZN(
        n7943) );
  OAI22_X1 U24682 ( .A1(n27300), .A2(n27263), .B1(n27257), .B2(n22113), .ZN(
        n7944) );
  OAI22_X1 U24683 ( .A1(n27303), .A2(n27263), .B1(n27257), .B2(n22112), .ZN(
        n7945) );
  OAI22_X1 U24684 ( .A1(n27306), .A2(n27263), .B1(n27257), .B2(n22111), .ZN(
        n7946) );
  OAI22_X1 U24685 ( .A1(n27309), .A2(n27263), .B1(n27257), .B2(n22110), .ZN(
        n7947) );
  OAI22_X1 U24686 ( .A1(n27312), .A2(n27263), .B1(n27257), .B2(n22109), .ZN(
        n7948) );
  OAI22_X1 U24687 ( .A1(n27315), .A2(n27264), .B1(n27257), .B2(n22108), .ZN(
        n7949) );
  OAI22_X1 U24688 ( .A1(n27282), .A2(n27227), .B1(n27221), .B2(n21939), .ZN(
        n7746) );
  OAI22_X1 U24689 ( .A1(n27285), .A2(n27227), .B1(n27221), .B2(n21938), .ZN(
        n7747) );
  OAI22_X1 U24690 ( .A1(n27288), .A2(n27227), .B1(n27221), .B2(n21937), .ZN(
        n7748) );
  OAI22_X1 U24691 ( .A1(n27291), .A2(n27227), .B1(n27221), .B2(n21936), .ZN(
        n7749) );
  OAI22_X1 U24692 ( .A1(n27294), .A2(n27227), .B1(n27221), .B2(n21935), .ZN(
        n7750) );
  OAI22_X1 U24693 ( .A1(n27297), .A2(n27227), .B1(n27221), .B2(n21934), .ZN(
        n7751) );
  OAI22_X1 U24694 ( .A1(n27300), .A2(n27227), .B1(n27221), .B2(n21933), .ZN(
        n7752) );
  OAI22_X1 U24695 ( .A1(n27303), .A2(n27227), .B1(n27221), .B2(n21932), .ZN(
        n7753) );
  OAI22_X1 U24696 ( .A1(n27306), .A2(n27227), .B1(n27221), .B2(n21931), .ZN(
        n7754) );
  OAI22_X1 U24697 ( .A1(n27309), .A2(n27227), .B1(n27221), .B2(n21930), .ZN(
        n7755) );
  OAI22_X1 U24698 ( .A1(n27312), .A2(n27227), .B1(n27221), .B2(n21929), .ZN(
        n7756) );
  OAI22_X1 U24699 ( .A1(n27315), .A2(n27228), .B1(n27221), .B2(n21928), .ZN(
        n7757) );
  OAI22_X1 U24700 ( .A1(n27282), .A2(n27203), .B1(n27197), .B2(n21879), .ZN(
        n7618) );
  OAI22_X1 U24701 ( .A1(n27285), .A2(n27203), .B1(n27197), .B2(n21878), .ZN(
        n7619) );
  OAI22_X1 U24702 ( .A1(n27288), .A2(n27203), .B1(n27197), .B2(n21877), .ZN(
        n7620) );
  OAI22_X1 U24703 ( .A1(n27291), .A2(n27203), .B1(n27197), .B2(n21876), .ZN(
        n7621) );
  OAI22_X1 U24704 ( .A1(n27294), .A2(n27203), .B1(n27197), .B2(n21875), .ZN(
        n7622) );
  OAI22_X1 U24705 ( .A1(n27297), .A2(n27203), .B1(n27197), .B2(n21874), .ZN(
        n7623) );
  OAI22_X1 U24706 ( .A1(n27300), .A2(n27203), .B1(n27197), .B2(n21873), .ZN(
        n7624) );
  OAI22_X1 U24707 ( .A1(n27303), .A2(n27203), .B1(n27197), .B2(n21872), .ZN(
        n7625) );
  OAI22_X1 U24708 ( .A1(n27306), .A2(n27203), .B1(n27197), .B2(n21871), .ZN(
        n7626) );
  OAI22_X1 U24709 ( .A1(n27309), .A2(n27203), .B1(n27197), .B2(n21870), .ZN(
        n7627) );
  OAI22_X1 U24710 ( .A1(n27312), .A2(n27203), .B1(n27197), .B2(n21869), .ZN(
        n7628) );
  OAI22_X1 U24711 ( .A1(n27315), .A2(n27204), .B1(n27197), .B2(n21868), .ZN(
        n7629) );
  OAI22_X1 U24712 ( .A1(n27283), .A2(n27011), .B1(n27005), .B2(n21819), .ZN(
        n6594) );
  OAI22_X1 U24713 ( .A1(n27286), .A2(n27011), .B1(n27005), .B2(n21818), .ZN(
        n6595) );
  OAI22_X1 U24714 ( .A1(n27289), .A2(n27011), .B1(n27005), .B2(n21817), .ZN(
        n6596) );
  OAI22_X1 U24715 ( .A1(n27292), .A2(n27011), .B1(n27005), .B2(n21816), .ZN(
        n6597) );
  OAI22_X1 U24716 ( .A1(n27295), .A2(n27011), .B1(n27005), .B2(n21815), .ZN(
        n6598) );
  OAI22_X1 U24717 ( .A1(n27298), .A2(n27011), .B1(n27005), .B2(n21814), .ZN(
        n6599) );
  OAI22_X1 U24718 ( .A1(n27301), .A2(n27011), .B1(n27005), .B2(n21813), .ZN(
        n6600) );
  OAI22_X1 U24719 ( .A1(n27304), .A2(n27011), .B1(n27005), .B2(n21812), .ZN(
        n6601) );
  OAI22_X1 U24720 ( .A1(n27307), .A2(n27011), .B1(n27005), .B2(n21811), .ZN(
        n6602) );
  OAI22_X1 U24721 ( .A1(n27310), .A2(n27011), .B1(n27005), .B2(n21810), .ZN(
        n6603) );
  OAI22_X1 U24722 ( .A1(n27313), .A2(n27011), .B1(n27005), .B2(n21809), .ZN(
        n6604) );
  OAI22_X1 U24723 ( .A1(n27316), .A2(n27012), .B1(n27005), .B2(n21808), .ZN(
        n6605) );
  OAI22_X1 U24724 ( .A1(n27283), .A2(n27059), .B1(n27053), .B2(n21699), .ZN(
        n6850) );
  OAI22_X1 U24725 ( .A1(n27286), .A2(n27059), .B1(n27053), .B2(n21698), .ZN(
        n6851) );
  OAI22_X1 U24726 ( .A1(n27289), .A2(n27059), .B1(n27053), .B2(n21697), .ZN(
        n6852) );
  OAI22_X1 U24727 ( .A1(n27292), .A2(n27059), .B1(n27053), .B2(n21696), .ZN(
        n6853) );
  OAI22_X1 U24728 ( .A1(n27295), .A2(n27059), .B1(n27053), .B2(n21695), .ZN(
        n6854) );
  OAI22_X1 U24729 ( .A1(n27298), .A2(n27059), .B1(n27053), .B2(n21694), .ZN(
        n6855) );
  OAI22_X1 U24730 ( .A1(n27301), .A2(n27059), .B1(n27053), .B2(n21693), .ZN(
        n6856) );
  OAI22_X1 U24731 ( .A1(n27304), .A2(n27059), .B1(n27053), .B2(n21692), .ZN(
        n6857) );
  OAI22_X1 U24732 ( .A1(n27307), .A2(n27059), .B1(n27053), .B2(n21691), .ZN(
        n6858) );
  OAI22_X1 U24733 ( .A1(n27310), .A2(n27059), .B1(n27053), .B2(n21690), .ZN(
        n6859) );
  OAI22_X1 U24734 ( .A1(n27313), .A2(n27059), .B1(n27053), .B2(n21689), .ZN(
        n6860) );
  OAI22_X1 U24735 ( .A1(n27316), .A2(n27060), .B1(n27053), .B2(n21688), .ZN(
        n6861) );
  OAI22_X1 U24736 ( .A1(n27282), .A2(n27251), .B1(n27245), .B2(n21479), .ZN(
        n7874) );
  OAI22_X1 U24737 ( .A1(n27285), .A2(n27251), .B1(n27245), .B2(n21478), .ZN(
        n7875) );
  OAI22_X1 U24738 ( .A1(n27288), .A2(n27251), .B1(n27245), .B2(n21477), .ZN(
        n7876) );
  OAI22_X1 U24739 ( .A1(n27291), .A2(n27251), .B1(n27245), .B2(n21476), .ZN(
        n7877) );
  OAI22_X1 U24740 ( .A1(n27294), .A2(n27251), .B1(n27245), .B2(n21475), .ZN(
        n7878) );
  OAI22_X1 U24741 ( .A1(n27297), .A2(n27251), .B1(n27245), .B2(n21474), .ZN(
        n7879) );
  OAI22_X1 U24742 ( .A1(n27300), .A2(n27251), .B1(n27245), .B2(n21473), .ZN(
        n7880) );
  OAI22_X1 U24743 ( .A1(n27303), .A2(n27251), .B1(n27245), .B2(n21472), .ZN(
        n7881) );
  OAI22_X1 U24744 ( .A1(n27306), .A2(n27251), .B1(n27245), .B2(n21471), .ZN(
        n7882) );
  OAI22_X1 U24745 ( .A1(n27309), .A2(n27251), .B1(n27245), .B2(n21470), .ZN(
        n7883) );
  OAI22_X1 U24746 ( .A1(n27312), .A2(n27251), .B1(n27245), .B2(n21469), .ZN(
        n7884) );
  OAI22_X1 U24747 ( .A1(n27315), .A2(n27252), .B1(n27245), .B2(n21468), .ZN(
        n7885) );
  OAI22_X1 U24748 ( .A1(n27283), .A2(n27083), .B1(n27077), .B2(n21299), .ZN(
        n6978) );
  OAI22_X1 U24749 ( .A1(n27286), .A2(n27083), .B1(n27077), .B2(n21298), .ZN(
        n6979) );
  OAI22_X1 U24750 ( .A1(n27289), .A2(n27083), .B1(n27077), .B2(n21297), .ZN(
        n6980) );
  OAI22_X1 U24751 ( .A1(n27292), .A2(n27083), .B1(n27077), .B2(n21296), .ZN(
        n6981) );
  OAI22_X1 U24752 ( .A1(n27295), .A2(n27083), .B1(n27077), .B2(n21295), .ZN(
        n6982) );
  OAI22_X1 U24753 ( .A1(n27298), .A2(n27083), .B1(n27077), .B2(n21294), .ZN(
        n6983) );
  OAI22_X1 U24754 ( .A1(n27301), .A2(n27083), .B1(n27077), .B2(n21293), .ZN(
        n6984) );
  OAI22_X1 U24755 ( .A1(n27304), .A2(n27083), .B1(n27077), .B2(n21292), .ZN(
        n6985) );
  OAI22_X1 U24756 ( .A1(n27307), .A2(n27083), .B1(n27077), .B2(n21291), .ZN(
        n6986) );
  OAI22_X1 U24757 ( .A1(n27310), .A2(n27083), .B1(n27077), .B2(n21290), .ZN(
        n6987) );
  OAI22_X1 U24758 ( .A1(n27313), .A2(n27083), .B1(n27077), .B2(n21289), .ZN(
        n6988) );
  OAI22_X1 U24759 ( .A1(n27316), .A2(n27084), .B1(n27077), .B2(n21288), .ZN(
        n6989) );
  OAI22_X1 U24760 ( .A1(n27284), .A2(n26903), .B1(n26897), .B2(n20962), .ZN(
        n6018) );
  OAI22_X1 U24761 ( .A1(n27287), .A2(n26903), .B1(n26897), .B2(n20961), .ZN(
        n6019) );
  OAI22_X1 U24762 ( .A1(n27290), .A2(n26903), .B1(n26897), .B2(n20960), .ZN(
        n6020) );
  OAI22_X1 U24763 ( .A1(n27293), .A2(n26903), .B1(n26897), .B2(n20959), .ZN(
        n6021) );
  OAI22_X1 U24764 ( .A1(n27296), .A2(n26903), .B1(n26897), .B2(n20958), .ZN(
        n6022) );
  OAI22_X1 U24765 ( .A1(n27299), .A2(n26903), .B1(n26897), .B2(n20957), .ZN(
        n6023) );
  OAI22_X1 U24766 ( .A1(n27302), .A2(n26903), .B1(n26897), .B2(n20956), .ZN(
        n6024) );
  OAI22_X1 U24767 ( .A1(n27305), .A2(n26903), .B1(n26897), .B2(n20955), .ZN(
        n6025) );
  OAI22_X1 U24768 ( .A1(n27308), .A2(n26903), .B1(n26897), .B2(n20954), .ZN(
        n6026) );
  OAI22_X1 U24769 ( .A1(n27311), .A2(n26903), .B1(n26897), .B2(n20953), .ZN(
        n6027) );
  OAI22_X1 U24770 ( .A1(n27314), .A2(n26903), .B1(n26897), .B2(n20952), .ZN(
        n6028) );
  OAI22_X1 U24771 ( .A1(n27317), .A2(n26904), .B1(n26897), .B2(n20951), .ZN(
        n6029) );
  OAI22_X1 U24772 ( .A1(n27284), .A2(n26915), .B1(n26909), .B2(n20898), .ZN(
        n6082) );
  OAI22_X1 U24773 ( .A1(n27287), .A2(n26915), .B1(n26909), .B2(n20897), .ZN(
        n6083) );
  OAI22_X1 U24774 ( .A1(n27290), .A2(n26915), .B1(n26909), .B2(n20896), .ZN(
        n6084) );
  OAI22_X1 U24775 ( .A1(n27293), .A2(n26915), .B1(n26909), .B2(n20895), .ZN(
        n6085) );
  OAI22_X1 U24776 ( .A1(n27296), .A2(n26915), .B1(n26909), .B2(n20894), .ZN(
        n6086) );
  OAI22_X1 U24777 ( .A1(n27299), .A2(n26915), .B1(n26909), .B2(n20893), .ZN(
        n6087) );
  OAI22_X1 U24778 ( .A1(n27302), .A2(n26915), .B1(n26909), .B2(n20892), .ZN(
        n6088) );
  OAI22_X1 U24779 ( .A1(n27305), .A2(n26915), .B1(n26909), .B2(n20891), .ZN(
        n6089) );
  OAI22_X1 U24780 ( .A1(n27308), .A2(n26915), .B1(n26909), .B2(n20890), .ZN(
        n6090) );
  OAI22_X1 U24781 ( .A1(n27311), .A2(n26915), .B1(n26909), .B2(n20889), .ZN(
        n6091) );
  OAI22_X1 U24782 ( .A1(n27314), .A2(n26915), .B1(n26909), .B2(n20888), .ZN(
        n6092) );
  OAI22_X1 U24783 ( .A1(n27317), .A2(n26916), .B1(n26909), .B2(n20887), .ZN(
        n6093) );
  OAI21_X1 U24784 ( .B1(n26533), .B2(n19454), .A(ENABLE), .ZN(n19580) );
  OAI21_X1 U24785 ( .B1(n26533), .B2(n18553), .A(n27481), .ZN(n19507) );
  OAI21_X1 U24786 ( .B1(n26533), .B2(n18536), .A(n27481), .ZN(n19508) );
  OAI21_X1 U24787 ( .B1(n26533), .B2(n18519), .A(n27481), .ZN(n19509) );
  OAI21_X1 U24788 ( .B1(n26533), .B2(n18502), .A(n27481), .ZN(n19510) );
  OAI21_X1 U24789 ( .B1(n26533), .B2(n18485), .A(n27481), .ZN(n19511) );
  OAI21_X1 U24790 ( .B1(n26533), .B2(n18468), .A(n27481), .ZN(n19512) );
  OAI21_X1 U24791 ( .B1(n26533), .B2(n18451), .A(n27481), .ZN(n19513) );
  OAI21_X1 U24792 ( .B1(n26533), .B2(n18434), .A(n27481), .ZN(n19514) );
  OAI21_X1 U24793 ( .B1(n26533), .B2(n18417), .A(n27482), .ZN(n19515) );
  OAI21_X1 U24794 ( .B1(n26533), .B2(n18400), .A(n27482), .ZN(n19516) );
  OAI21_X1 U24795 ( .B1(n26533), .B2(n18383), .A(n27482), .ZN(n19517) );
  OAI21_X1 U24796 ( .B1(n26758), .B2(n18315), .A(n27486), .ZN(n19571) );
  OAI21_X1 U24797 ( .B1(n26758), .B2(n18314), .A(n27486), .ZN(n19570) );
  OAI21_X1 U24798 ( .B1(n26758), .B2(n18313), .A(n27486), .ZN(n19573) );
  OAI21_X1 U24799 ( .B1(n26758), .B2(n18312), .A(n27486), .ZN(n19572) );
  OAI21_X1 U24800 ( .B1(n26758), .B2(n18311), .A(ENABLE), .ZN(n19575) );
  OAI21_X1 U24801 ( .B1(n26758), .B2(n18310), .A(n27486), .ZN(n19574) );
  OAI21_X1 U24802 ( .B1(n26758), .B2(n18309), .A(ENABLE), .ZN(n19577) );
  OAI21_X1 U24803 ( .B1(n26758), .B2(n18307), .A(ENABLE), .ZN(n19579) );
  OAI21_X1 U24804 ( .B1(n26758), .B2(n18306), .A(ENABLE), .ZN(n19576) );
  OAI21_X1 U24805 ( .B1(n26758), .B2(n18305), .A(ENABLE), .ZN(n19581) );
  OAI21_X1 U24806 ( .B1(n26758), .B2(n18304), .A(ENABLE), .ZN(n19578) );
  OAI21_X1 U24807 ( .B1(n26758), .B2(n18303), .A(ENABLE), .ZN(n19582) );
  OAI21_X1 U24808 ( .B1(n26535), .B2(n19437), .A(n27477), .ZN(n19455) );
  OAI21_X1 U24809 ( .B1(n26535), .B2(n19420), .A(n27477), .ZN(n19456) );
  OAI21_X1 U24810 ( .B1(n26535), .B2(n19403), .A(n27477), .ZN(n19457) );
  OAI21_X1 U24811 ( .B1(n26535), .B2(n19386), .A(n27477), .ZN(n19458) );
  OAI21_X1 U24812 ( .B1(n26535), .B2(n19369), .A(n27477), .ZN(n19459) );
  OAI21_X1 U24813 ( .B1(n26535), .B2(n19352), .A(n27477), .ZN(n19460) );
  OAI21_X1 U24814 ( .B1(n26535), .B2(n19335), .A(n27477), .ZN(n19461) );
  OAI21_X1 U24815 ( .B1(n26535), .B2(n19318), .A(n27477), .ZN(n19462) );
  OAI21_X1 U24816 ( .B1(n26535), .B2(n19301), .A(n27477), .ZN(n19463) );
  OAI21_X1 U24817 ( .B1(n26535), .B2(n19284), .A(n27477), .ZN(n19464) );
  OAI21_X1 U24818 ( .B1(n26535), .B2(n19267), .A(n27477), .ZN(n19465) );
  OAI21_X1 U24819 ( .B1(n26535), .B2(n19250), .A(n27477), .ZN(n19466) );
  OAI21_X1 U24820 ( .B1(n26535), .B2(n19233), .A(n27478), .ZN(n19467) );
  OAI21_X1 U24821 ( .B1(n26534), .B2(n19216), .A(n27478), .ZN(n19468) );
  OAI21_X1 U24822 ( .B1(n26534), .B2(n19199), .A(n27478), .ZN(n19469) );
  OAI21_X1 U24823 ( .B1(n26534), .B2(n19182), .A(n27478), .ZN(n19470) );
  OAI21_X1 U24824 ( .B1(n26534), .B2(n19165), .A(n27478), .ZN(n19471) );
  OAI21_X1 U24825 ( .B1(n26534), .B2(n19148), .A(n27478), .ZN(n19472) );
  OAI21_X1 U24826 ( .B1(n26534), .B2(n19131), .A(n27478), .ZN(n19473) );
  OAI21_X1 U24827 ( .B1(n26534), .B2(n19114), .A(n27478), .ZN(n19474) );
  OAI21_X1 U24828 ( .B1(n26534), .B2(n19097), .A(n27478), .ZN(n19475) );
  OAI21_X1 U24829 ( .B1(n26534), .B2(n19080), .A(n27478), .ZN(n19476) );
  OAI21_X1 U24830 ( .B1(n26534), .B2(n19063), .A(n27478), .ZN(n19477) );
  OAI21_X1 U24831 ( .B1(n26534), .B2(n19046), .A(n27478), .ZN(n19478) );
  OAI21_X1 U24832 ( .B1(n26534), .B2(n19029), .A(n27479), .ZN(n19479) );
  OAI21_X1 U24833 ( .B1(n26534), .B2(n19012), .A(n27479), .ZN(n19480) );
  OAI21_X1 U24834 ( .B1(n26534), .B2(n18995), .A(n27479), .ZN(n19481) );
  OAI21_X1 U24835 ( .B1(n26533), .B2(n18978), .A(n27479), .ZN(n19482) );
  OAI21_X1 U24836 ( .B1(n26535), .B2(n18961), .A(n27479), .ZN(n19483) );
  OAI21_X1 U24837 ( .B1(n26534), .B2(n18944), .A(n27479), .ZN(n19484) );
  OAI21_X1 U24838 ( .B1(n26533), .B2(n18927), .A(n27479), .ZN(n19485) );
  OAI21_X1 U24839 ( .B1(n26535), .B2(n18910), .A(n27479), .ZN(n19486) );
  OAI21_X1 U24840 ( .B1(n26534), .B2(n18893), .A(n27479), .ZN(n19487) );
  OAI21_X1 U24841 ( .B1(n26533), .B2(n18876), .A(n27479), .ZN(n19488) );
  OAI21_X1 U24842 ( .B1(n26535), .B2(n18859), .A(n27479), .ZN(n19489) );
  OAI21_X1 U24843 ( .B1(n26534), .B2(n18842), .A(n27479), .ZN(n19490) );
  OAI21_X1 U24844 ( .B1(n26533), .B2(n18825), .A(n27480), .ZN(n19491) );
  OAI21_X1 U24845 ( .B1(n26535), .B2(n18808), .A(n27480), .ZN(n19492) );
  OAI21_X1 U24846 ( .B1(n26534), .B2(n18791), .A(n27480), .ZN(n19493) );
  OAI21_X1 U24847 ( .B1(n26535), .B2(n18774), .A(n27480), .ZN(n19494) );
  OAI21_X1 U24848 ( .B1(n26534), .B2(n18757), .A(n27480), .ZN(n19495) );
  OAI21_X1 U24849 ( .B1(n26534), .B2(n18740), .A(n27480), .ZN(n19496) );
  OAI21_X1 U24850 ( .B1(n26533), .B2(n18723), .A(n27480), .ZN(n19497) );
  OAI21_X1 U24851 ( .B1(n26535), .B2(n18706), .A(n27480), .ZN(n19498) );
  OAI21_X1 U24852 ( .B1(n26534), .B2(n18689), .A(n27480), .ZN(n19499) );
  OAI21_X1 U24853 ( .B1(n26533), .B2(n18672), .A(n27480), .ZN(n19500) );
  OAI21_X1 U24854 ( .B1(n26533), .B2(n18655), .A(n27480), .ZN(n19501) );
  OAI21_X1 U24855 ( .B1(n26535), .B2(n18638), .A(n27480), .ZN(n19502) );
  OAI21_X1 U24856 ( .B1(n26534), .B2(n18621), .A(n27481), .ZN(n19503) );
  OAI21_X1 U24857 ( .B1(n26535), .B2(n18604), .A(n27481), .ZN(n19504) );
  OAI21_X1 U24858 ( .B1(n26533), .B2(n18587), .A(n27481), .ZN(n19505) );
  OAI21_X1 U24859 ( .B1(n26535), .B2(n18570), .A(n27481), .ZN(n19506) );
  OAI21_X1 U24860 ( .B1(n26760), .B2(n18366), .A(n27482), .ZN(n19518) );
  OAI21_X1 U24861 ( .B1(n26758), .B2(n18365), .A(n27482), .ZN(n19521) );
  OAI21_X1 U24862 ( .B1(n26759), .B2(n18364), .A(n27482), .ZN(n19522) );
  OAI21_X1 U24863 ( .B1(n26760), .B2(n18363), .A(n27482), .ZN(n19523) );
  OAI21_X1 U24864 ( .B1(n26758), .B2(n18362), .A(n27482), .ZN(n19524) );
  OAI21_X1 U24865 ( .B1(n26759), .B2(n18361), .A(n27482), .ZN(n19525) );
  OAI21_X1 U24866 ( .B1(n26760), .B2(n18360), .A(n27482), .ZN(n19526) );
  OAI21_X1 U24867 ( .B1(n26758), .B2(n18359), .A(n27483), .ZN(n19527) );
  OAI21_X1 U24868 ( .B1(n26759), .B2(n18358), .A(n27483), .ZN(n19528) );
  OAI21_X1 U24869 ( .B1(n26760), .B2(n18357), .A(n27483), .ZN(n19529) );
  OAI21_X1 U24870 ( .B1(n26758), .B2(n18356), .A(n27483), .ZN(n19530) );
  OAI21_X1 U24871 ( .B1(n26760), .B2(n18355), .A(n27483), .ZN(n19531) );
  OAI21_X1 U24872 ( .B1(n26760), .B2(n18354), .A(n27483), .ZN(n19532) );
  OAI21_X1 U24873 ( .B1(n26760), .B2(n18353), .A(n27483), .ZN(n19533) );
  OAI21_X1 U24874 ( .B1(n26760), .B2(n18352), .A(n27483), .ZN(n19534) );
  OAI21_X1 U24875 ( .B1(n26760), .B2(n18351), .A(n27483), .ZN(n19535) );
  OAI21_X1 U24876 ( .B1(n26760), .B2(n18350), .A(n27483), .ZN(n19536) );
  OAI21_X1 U24877 ( .B1(n26760), .B2(n18349), .A(n27483), .ZN(n19537) );
  OAI21_X1 U24878 ( .B1(n26760), .B2(n18348), .A(n27483), .ZN(n19538) );
  OAI21_X1 U24879 ( .B1(n26760), .B2(n18347), .A(n27484), .ZN(n19539) );
  OAI21_X1 U24880 ( .B1(n26760), .B2(n18346), .A(n27484), .ZN(n19540) );
  OAI21_X1 U24881 ( .B1(n26760), .B2(n18345), .A(n27484), .ZN(n19541) );
  OAI21_X1 U24882 ( .B1(n26760), .B2(n18344), .A(n27484), .ZN(n19542) );
  OAI21_X1 U24883 ( .B1(n26760), .B2(n18343), .A(n27484), .ZN(n19543) );
  OAI21_X1 U24884 ( .B1(n26759), .B2(n18342), .A(n27484), .ZN(n19544) );
  OAI21_X1 U24885 ( .B1(n26760), .B2(n18341), .A(n27484), .ZN(n19545) );
  OAI21_X1 U24886 ( .B1(n26760), .B2(n18340), .A(n27484), .ZN(n19546) );
  OAI21_X1 U24887 ( .B1(n26758), .B2(n18339), .A(n27484), .ZN(n19547) );
  OAI21_X1 U24888 ( .B1(n26759), .B2(n18338), .A(n27484), .ZN(n19548) );
  OAI21_X1 U24889 ( .B1(n26759), .B2(n18337), .A(n27482), .ZN(n19520) );
  OAI21_X1 U24890 ( .B1(n26758), .B2(n18336), .A(n27484), .ZN(n19550) );
  OAI21_X1 U24891 ( .B1(n26760), .B2(n18335), .A(n27485), .ZN(n19551) );
  OAI21_X1 U24892 ( .B1(n26760), .B2(n18334), .A(n27482), .ZN(n19519) );
  OAI21_X1 U24893 ( .B1(n26758), .B2(n18333), .A(n27485), .ZN(n19553) );
  OAI21_X1 U24894 ( .B1(n26759), .B2(n18332), .A(n27485), .ZN(n19552) );
  OAI21_X1 U24895 ( .B1(n26759), .B2(n18331), .A(n27485), .ZN(n19555) );
  OAI21_X1 U24896 ( .B1(n26760), .B2(n18330), .A(n27485), .ZN(n19554) );
  OAI21_X1 U24897 ( .B1(n26759), .B2(n18329), .A(n27485), .ZN(n19557) );
  OAI21_X1 U24898 ( .B1(n26758), .B2(n18328), .A(n27485), .ZN(n19556) );
  OAI21_X1 U24899 ( .B1(n26759), .B2(n18327), .A(n27485), .ZN(n19559) );
  OAI21_X1 U24900 ( .B1(n26759), .B2(n18326), .A(n27485), .ZN(n19558) );
  OAI21_X1 U24901 ( .B1(n26759), .B2(n18325), .A(n27485), .ZN(n19561) );
  OAI21_X1 U24902 ( .B1(n26759), .B2(n18324), .A(n27485), .ZN(n19560) );
  OAI21_X1 U24903 ( .B1(n26759), .B2(n18323), .A(n27486), .ZN(n19563) );
  OAI21_X1 U24904 ( .B1(n26759), .B2(n18322), .A(n27485), .ZN(n19562) );
  OAI21_X1 U24905 ( .B1(n26759), .B2(n18321), .A(n27486), .ZN(n19565) );
  OAI21_X1 U24906 ( .B1(n26759), .B2(n18320), .A(n27486), .ZN(n19564) );
  OAI21_X1 U24907 ( .B1(n26759), .B2(n18319), .A(n27486), .ZN(n19567) );
  OAI21_X1 U24908 ( .B1(n26759), .B2(n18318), .A(n27486), .ZN(n19566) );
  OAI21_X1 U24909 ( .B1(n26759), .B2(n18317), .A(n27486), .ZN(n19569) );
  OAI21_X1 U24910 ( .B1(n26759), .B2(n18316), .A(n27486), .ZN(n19568) );
  OAI21_X1 U24911 ( .B1(n26759), .B2(n18308), .A(n27484), .ZN(n19549) );
  NOR3_X1 U24912 ( .A1(ADD_WR[1]), .A2(ADD_WR[2]), .A3(ADD_WR[0]), .ZN(n22694)
         );
  NOR3_X1 U24913 ( .A1(n20633), .A2(ADD_WR[2]), .A3(n20632), .ZN(n22704) );
  NOR3_X1 U24914 ( .A1(ADD_WR[0]), .A2(ADD_WR[2]), .A3(n20632), .ZN(n22701) );
  NOR3_X1 U24915 ( .A1(ADD_WR[1]), .A2(ADD_WR[2]), .A3(n20633), .ZN(n22698) );
  NOR3_X1 U24916 ( .A1(n20643), .A2(ADD_RD2[3]), .A3(n20639), .ZN(n25147) );
  NOR3_X1 U24917 ( .A1(n20638), .A2(ADD_RD1[3]), .A3(n20634), .ZN(n23948) );
  NOR3_X1 U24918 ( .A1(ADD_RD2[0]), .A2(ADD_RD2[4]), .A3(n20640), .ZN(n25153)
         );
  NOR3_X1 U24919 ( .A1(ADD_RD1[0]), .A2(ADD_RD1[4]), .A3(n20635), .ZN(n23954)
         );
  NOR3_X1 U24920 ( .A1(n20643), .A2(ADD_RD2[4]), .A3(n20640), .ZN(n25155) );
  NOR3_X1 U24921 ( .A1(n20638), .A2(ADD_RD1[4]), .A3(n20635), .ZN(n23956) );
  NOR3_X1 U24922 ( .A1(n20640), .A2(ADD_RD2[0]), .A3(n20639), .ZN(n25146) );
  NOR3_X1 U24923 ( .A1(n20635), .A2(ADD_RD1[0]), .A3(n20634), .ZN(n23947) );
  NOR3_X1 U24924 ( .A1(ADD_RD2[0]), .A2(ADD_RD2[3]), .A3(n20639), .ZN(n25150)
         );
  NOR3_X1 U24925 ( .A1(ADD_RD1[0]), .A2(ADD_RD1[3]), .A3(n20634), .ZN(n23951)
         );
  NOR3_X1 U24926 ( .A1(ADD_RD2[3]), .A2(ADD_RD2[4]), .A3(ADD_RD2[0]), .ZN(
        n25163) );
  NOR3_X1 U24927 ( .A1(ADD_RD1[3]), .A2(ADD_RD1[4]), .A3(ADD_RD1[0]), .ZN(
        n23964) );
  AND3_X1 U24928 ( .A1(n22717), .A2(n20631), .A3(ADD_WR[4]), .ZN(n22737) );
  AND3_X1 U24929 ( .A1(ADD_WR[3]), .A2(n22717), .A3(ADD_WR[4]), .ZN(n22754) );
  AND3_X1 U24930 ( .A1(n22717), .A2(n20630), .A3(ADD_WR[3]), .ZN(n22720) );
  NOR2_X1 U24931 ( .A1(n26536), .A2(WR), .ZN(n25164) );
  NOR2_X1 U24932 ( .A1(n26761), .A2(WR), .ZN(n23965) );
  NAND2_X1 U24933 ( .A1(WR), .A2(n26533), .ZN(n24015) );
  NAND2_X1 U24934 ( .A1(WR), .A2(n26758), .ZN(n22816) );
  AND3_X1 U24935 ( .A1(n25164), .A2(n20641), .A3(ADD_RD2[1]), .ZN(n25144) );
  AND3_X1 U24936 ( .A1(n23965), .A2(n20636), .A3(ADD_RD1[1]), .ZN(n23945) );
  AND3_X1 U24937 ( .A1(ADD_RD2[1]), .A2(n25164), .A3(ADD_RD2[2]), .ZN(n25148)
         );
  AND3_X1 U24938 ( .A1(ADD_RD1[1]), .A2(n23965), .A3(ADD_RD1[2]), .ZN(n23949)
         );
  AND3_X1 U24939 ( .A1(n25164), .A2(n20642), .A3(ADD_RD2[2]), .ZN(n25145) );
  AND3_X1 U24940 ( .A1(n23965), .A2(n20637), .A3(ADD_RD1[2]), .ZN(n23946) );
  INV_X1 U24941 ( .A(ADD_RD2[4]), .ZN(n20639) );
  INV_X1 U24942 ( .A(ADD_RD1[4]), .ZN(n20634) );
  INV_X1 U24943 ( .A(ADD_RD2[3]), .ZN(n20640) );
  INV_X1 U24944 ( .A(ADD_RD1[3]), .ZN(n20635) );
  AND3_X1 U24945 ( .A1(n20633), .A2(n20632), .A3(ADD_WR[2]), .ZN(n22707) );
  AND3_X1 U24946 ( .A1(ADD_WR[0]), .A2(n20632), .A3(ADD_WR[2]), .ZN(n22710) );
  AND3_X1 U24947 ( .A1(ADD_WR[1]), .A2(n20633), .A3(ADD_WR[2]), .ZN(n22713) );
  AND3_X1 U24948 ( .A1(ADD_WR[1]), .A2(ADD_WR[0]), .A3(ADD_WR[2]), .ZN(n22716)
         );
  INV_X1 U24949 ( .A(ADD_WR[1]), .ZN(n20632) );
  INV_X1 U24950 ( .A(ADD_WR[0]), .ZN(n20633) );
  NOR2_X1 U24951 ( .A1(RD2), .A2(n27487), .ZN(n24003) );
  NOR2_X1 U24952 ( .A1(RD1), .A2(n27487), .ZN(n22804) );
  INV_X1 U24953 ( .A(ADD_RD2[0]), .ZN(n20643) );
  INV_X1 U24954 ( .A(ADD_RD1[0]), .ZN(n20638) );
  AND2_X1 U24955 ( .A1(WR), .A2(ENABLE), .ZN(n22717) );
  INV_X1 U24956 ( .A(RESET), .ZN(n20626) );
  INV_X1 U24957 ( .A(DATAIN[0]), .ZN(n20707) );
  INV_X1 U24958 ( .A(DATAIN[1]), .ZN(n20706) );
  INV_X1 U24959 ( .A(DATAIN[2]), .ZN(n20705) );
  INV_X1 U24960 ( .A(DATAIN[3]), .ZN(n20704) );
  INV_X1 U24961 ( .A(DATAIN[4]), .ZN(n20703) );
  INV_X1 U24962 ( .A(DATAIN[5]), .ZN(n20702) );
  INV_X1 U24963 ( .A(DATAIN[6]), .ZN(n20701) );
  INV_X1 U24964 ( .A(DATAIN[7]), .ZN(n20700) );
  INV_X1 U24965 ( .A(DATAIN[8]), .ZN(n20699) );
  INV_X1 U24966 ( .A(DATAIN[9]), .ZN(n20698) );
  INV_X1 U24967 ( .A(DATAIN[10]), .ZN(n20697) );
  INV_X1 U24968 ( .A(DATAIN[11]), .ZN(n20696) );
  INV_X1 U24969 ( .A(DATAIN[12]), .ZN(n20695) );
  INV_X1 U24970 ( .A(DATAIN[13]), .ZN(n20694) );
  INV_X1 U24971 ( .A(DATAIN[14]), .ZN(n20693) );
  INV_X1 U24972 ( .A(DATAIN[15]), .ZN(n20692) );
  INV_X1 U24973 ( .A(DATAIN[16]), .ZN(n20691) );
  INV_X1 U24974 ( .A(DATAIN[17]), .ZN(n20690) );
  INV_X1 U24975 ( .A(DATAIN[18]), .ZN(n20689) );
  INV_X1 U24976 ( .A(DATAIN[19]), .ZN(n20688) );
  INV_X1 U24977 ( .A(DATAIN[20]), .ZN(n20687) );
  INV_X1 U24978 ( .A(DATAIN[21]), .ZN(n20686) );
  INV_X1 U24979 ( .A(DATAIN[22]), .ZN(n20685) );
  INV_X1 U24980 ( .A(DATAIN[23]), .ZN(n20684) );
  INV_X1 U24981 ( .A(DATAIN[24]), .ZN(n20683) );
  INV_X1 U24982 ( .A(DATAIN[25]), .ZN(n20682) );
  INV_X1 U24983 ( .A(DATAIN[26]), .ZN(n20681) );
  INV_X1 U24984 ( .A(DATAIN[27]), .ZN(n20680) );
  INV_X1 U24985 ( .A(DATAIN[28]), .ZN(n20679) );
  INV_X1 U24986 ( .A(DATAIN[29]), .ZN(n20678) );
  INV_X1 U24987 ( .A(DATAIN[30]), .ZN(n20677) );
  INV_X1 U24988 ( .A(DATAIN[31]), .ZN(n20676) );
  INV_X1 U24989 ( .A(DATAIN[32]), .ZN(n20675) );
  INV_X1 U24990 ( .A(DATAIN[33]), .ZN(n20674) );
  INV_X1 U24991 ( .A(DATAIN[34]), .ZN(n20673) );
  INV_X1 U24992 ( .A(DATAIN[35]), .ZN(n20672) );
  INV_X1 U24993 ( .A(DATAIN[36]), .ZN(n20671) );
  INV_X1 U24994 ( .A(DATAIN[37]), .ZN(n20670) );
  INV_X1 U24995 ( .A(DATAIN[38]), .ZN(n20669) );
  INV_X1 U24996 ( .A(DATAIN[39]), .ZN(n20668) );
  INV_X1 U24997 ( .A(DATAIN[40]), .ZN(n20667) );
  INV_X1 U24998 ( .A(DATAIN[41]), .ZN(n20666) );
  INV_X1 U24999 ( .A(DATAIN[42]), .ZN(n20665) );
  INV_X1 U25000 ( .A(DATAIN[43]), .ZN(n20664) );
  INV_X1 U25001 ( .A(DATAIN[44]), .ZN(n20663) );
  INV_X1 U25002 ( .A(DATAIN[45]), .ZN(n20662) );
  INV_X1 U25003 ( .A(DATAIN[46]), .ZN(n20661) );
  INV_X1 U25004 ( .A(DATAIN[47]), .ZN(n20660) );
  INV_X1 U25005 ( .A(DATAIN[48]), .ZN(n20659) );
  INV_X1 U25006 ( .A(DATAIN[49]), .ZN(n20658) );
  INV_X1 U25007 ( .A(DATAIN[50]), .ZN(n20657) );
  INV_X1 U25008 ( .A(DATAIN[51]), .ZN(n20656) );
  INV_X1 U25009 ( .A(DATAIN[52]), .ZN(n20655) );
  INV_X1 U25010 ( .A(DATAIN[53]), .ZN(n20654) );
  INV_X1 U25011 ( .A(DATAIN[54]), .ZN(n20653) );
  INV_X1 U25012 ( .A(DATAIN[55]), .ZN(n20652) );
  INV_X1 U25013 ( .A(DATAIN[56]), .ZN(n20651) );
  INV_X1 U25014 ( .A(DATAIN[57]), .ZN(n20650) );
  INV_X1 U25015 ( .A(DATAIN[58]), .ZN(n20649) );
  INV_X1 U25016 ( .A(DATAIN[59]), .ZN(n20648) );
  INV_X1 U25017 ( .A(DATAIN[60]), .ZN(n20647) );
  INV_X1 U25018 ( .A(DATAIN[61]), .ZN(n20646) );
  INV_X1 U25019 ( .A(DATAIN[62]), .ZN(n20645) );
  INV_X1 U25020 ( .A(DATAIN[63]), .ZN(n20644) );
  AND4_X1 U25021 ( .A1(n25164), .A2(ADD_RD2[0]), .A3(n20640), .A4(n20639), 
        .ZN(n25165) );
  AND4_X1 U25022 ( .A1(n23965), .A2(ADD_RD1[0]), .A3(n20635), .A4(n20634), 
        .ZN(n23966) );
  INV_X1 U25023 ( .A(ADD_RD2[2]), .ZN(n20641) );
  INV_X1 U25024 ( .A(ADD_RD1[2]), .ZN(n20636) );
  INV_X1 U25025 ( .A(ADD_RD2[1]), .ZN(n20642) );
  INV_X1 U25026 ( .A(ADD_RD1[1]), .ZN(n20637) );
  INV_X1 U25027 ( .A(ADD_WR[4]), .ZN(n20630) );
  INV_X1 U25028 ( .A(ADD_WR[3]), .ZN(n20631) );
  CLKBUF_X1 U25029 ( .A(n24019), .Z(n26452) );
  CLKBUF_X1 U25030 ( .A(n24018), .Z(n26458) );
  CLKBUF_X1 U25031 ( .A(n24017), .Z(n26464) );
  CLKBUF_X1 U25032 ( .A(n24015), .Z(n26470) );
  CLKBUF_X1 U25033 ( .A(n24014), .Z(n26476) );
  CLKBUF_X1 U25034 ( .A(n24013), .Z(n26482) );
  CLKBUF_X1 U25035 ( .A(n24012), .Z(n26488) );
  CLKBUF_X1 U25036 ( .A(n24010), .Z(n26494) );
  CLKBUF_X1 U25037 ( .A(n24009), .Z(n26500) );
  CLKBUF_X1 U25038 ( .A(n24008), .Z(n26506) );
  CLKBUF_X1 U25039 ( .A(n24007), .Z(n26512) );
  CLKBUF_X1 U25040 ( .A(n24005), .Z(n26518) );
  CLKBUF_X1 U25041 ( .A(n24004), .Z(n26524) );
  CLKBUF_X1 U25042 ( .A(n24002), .Z(n26557) );
  CLKBUF_X1 U25043 ( .A(n24000), .Z(n26563) );
  CLKBUF_X1 U25044 ( .A(n23999), .Z(n26569) );
  CLKBUF_X1 U25045 ( .A(n23994), .Z(n26575) );
  CLKBUF_X1 U25046 ( .A(n23993), .Z(n26581) );
  CLKBUF_X1 U25047 ( .A(n23992), .Z(n26587) );
  CLKBUF_X1 U25048 ( .A(n23990), .Z(n26593) );
  CLKBUF_X1 U25049 ( .A(n23989), .Z(n26599) );
  CLKBUF_X1 U25050 ( .A(n23988), .Z(n26605) );
  CLKBUF_X1 U25051 ( .A(n23987), .Z(n26611) );
  CLKBUF_X1 U25052 ( .A(n23985), .Z(n26617) );
  CLKBUF_X1 U25053 ( .A(n23984), .Z(n26623) );
  CLKBUF_X1 U25054 ( .A(n23983), .Z(n26629) );
  CLKBUF_X1 U25055 ( .A(n23982), .Z(n26635) );
  CLKBUF_X1 U25056 ( .A(n23980), .Z(n26641) );
  CLKBUF_X1 U25057 ( .A(n23979), .Z(n26647) );
  CLKBUF_X1 U25058 ( .A(n23978), .Z(n26653) );
  CLKBUF_X1 U25059 ( .A(n23977), .Z(n26659) );
  CLKBUF_X1 U25060 ( .A(n23975), .Z(n26665) );
  CLKBUF_X1 U25061 ( .A(n23974), .Z(n26671) );
  CLKBUF_X1 U25062 ( .A(n22820), .Z(n26677) );
  CLKBUF_X1 U25063 ( .A(n22819), .Z(n26683) );
  CLKBUF_X1 U25064 ( .A(n22818), .Z(n26689) );
  CLKBUF_X1 U25065 ( .A(n22816), .Z(n26695) );
  CLKBUF_X1 U25066 ( .A(n22815), .Z(n26701) );
  CLKBUF_X1 U25067 ( .A(n22814), .Z(n26707) );
  CLKBUF_X1 U25068 ( .A(n22813), .Z(n26713) );
  CLKBUF_X1 U25069 ( .A(n22811), .Z(n26719) );
  CLKBUF_X1 U25070 ( .A(n22810), .Z(n26725) );
  CLKBUF_X1 U25071 ( .A(n22809), .Z(n26731) );
  CLKBUF_X1 U25072 ( .A(n22808), .Z(n26737) );
  CLKBUF_X1 U25073 ( .A(n22806), .Z(n26743) );
  CLKBUF_X1 U25074 ( .A(n22805), .Z(n26749) );
  CLKBUF_X1 U25075 ( .A(n22803), .Z(n26782) );
  CLKBUF_X1 U25076 ( .A(n22801), .Z(n26788) );
  CLKBUF_X1 U25077 ( .A(n22800), .Z(n26794) );
  CLKBUF_X1 U25078 ( .A(n22795), .Z(n26800) );
  CLKBUF_X1 U25079 ( .A(n22794), .Z(n26806) );
  CLKBUF_X1 U25080 ( .A(n22793), .Z(n26812) );
  CLKBUF_X1 U25081 ( .A(n22791), .Z(n26818) );
  CLKBUF_X1 U25082 ( .A(n22790), .Z(n26824) );
  CLKBUF_X1 U25083 ( .A(n22789), .Z(n26830) );
  CLKBUF_X1 U25084 ( .A(n22788), .Z(n26836) );
  CLKBUF_X1 U25085 ( .A(n22786), .Z(n26842) );
  CLKBUF_X1 U25086 ( .A(n22785), .Z(n26848) );
  CLKBUF_X1 U25087 ( .A(n22784), .Z(n26854) );
  CLKBUF_X1 U25088 ( .A(n22783), .Z(n26860) );
  CLKBUF_X1 U25089 ( .A(n22781), .Z(n26866) );
  CLKBUF_X1 U25090 ( .A(n22780), .Z(n26872) );
  CLKBUF_X1 U25091 ( .A(n22779), .Z(n26878) );
  CLKBUF_X1 U25092 ( .A(n22778), .Z(n26884) );
  CLKBUF_X1 U25093 ( .A(n22776), .Z(n26890) );
  CLKBUF_X1 U25094 ( .A(n22775), .Z(n26896) );
  CLKBUF_X1 U25095 ( .A(n22768), .Z(n26902) );
  CLKBUF_X1 U25096 ( .A(n22767), .Z(n26908) );
  CLKBUF_X1 U25097 ( .A(n22766), .Z(n26914) );
  CLKBUF_X1 U25098 ( .A(n22765), .Z(n26920) );
  CLKBUF_X1 U25099 ( .A(n22764), .Z(n26926) );
  CLKBUF_X1 U25100 ( .A(n22763), .Z(n26932) );
  CLKBUF_X1 U25101 ( .A(n22762), .Z(n26938) );
  CLKBUF_X1 U25102 ( .A(n22761), .Z(n26944) );
  CLKBUF_X1 U25103 ( .A(n22760), .Z(n26950) );
  CLKBUF_X1 U25104 ( .A(n22759), .Z(n26956) );
  CLKBUF_X1 U25105 ( .A(n22758), .Z(n26962) );
  CLKBUF_X1 U25106 ( .A(n22757), .Z(n26968) );
  CLKBUF_X1 U25107 ( .A(n22756), .Z(n26974) );
  CLKBUF_X1 U25108 ( .A(n22755), .Z(n26980) );
  CLKBUF_X1 U25109 ( .A(n22753), .Z(n26986) );
  CLKBUF_X1 U25110 ( .A(n22752), .Z(n26992) );
  CLKBUF_X1 U25111 ( .A(n22751), .Z(n26998) );
  CLKBUF_X1 U25112 ( .A(n22750), .Z(n27004) );
  CLKBUF_X1 U25113 ( .A(n22749), .Z(n27010) );
  CLKBUF_X1 U25114 ( .A(n22748), .Z(n27016) );
  CLKBUF_X1 U25115 ( .A(n22747), .Z(n27022) );
  CLKBUF_X1 U25116 ( .A(n22746), .Z(n27028) );
  CLKBUF_X1 U25117 ( .A(n22745), .Z(n27034) );
  CLKBUF_X1 U25118 ( .A(n22744), .Z(n27040) );
  CLKBUF_X1 U25119 ( .A(n22743), .Z(n27046) );
  CLKBUF_X1 U25120 ( .A(n22742), .Z(n27052) );
  CLKBUF_X1 U25121 ( .A(n22741), .Z(n27058) );
  CLKBUF_X1 U25122 ( .A(n22740), .Z(n27064) );
  CLKBUF_X1 U25123 ( .A(n22739), .Z(n27070) );
  CLKBUF_X1 U25124 ( .A(n22738), .Z(n27076) );
  CLKBUF_X1 U25125 ( .A(n22736), .Z(n27082) );
  CLKBUF_X1 U25126 ( .A(n22735), .Z(n27088) );
  CLKBUF_X1 U25127 ( .A(n22734), .Z(n27094) );
  CLKBUF_X1 U25128 ( .A(n22733), .Z(n27100) );
  CLKBUF_X1 U25129 ( .A(n22732), .Z(n27106) );
  CLKBUF_X1 U25130 ( .A(n22731), .Z(n27112) );
  CLKBUF_X1 U25131 ( .A(n22730), .Z(n27118) );
  CLKBUF_X1 U25132 ( .A(n22729), .Z(n27124) );
  CLKBUF_X1 U25133 ( .A(n22728), .Z(n27130) );
  CLKBUF_X1 U25134 ( .A(n22727), .Z(n27136) );
  CLKBUF_X1 U25135 ( .A(n22726), .Z(n27142) );
  CLKBUF_X1 U25136 ( .A(n22725), .Z(n27148) );
  CLKBUF_X1 U25137 ( .A(n22724), .Z(n27154) );
  CLKBUF_X1 U25138 ( .A(n22723), .Z(n27160) );
  CLKBUF_X1 U25139 ( .A(n22722), .Z(n27166) );
  CLKBUF_X1 U25140 ( .A(n22721), .Z(n27172) );
  CLKBUF_X1 U25141 ( .A(n22719), .Z(n27178) );
  CLKBUF_X1 U25142 ( .A(n22718), .Z(n27184) );
  CLKBUF_X1 U25143 ( .A(n22715), .Z(n27190) );
  CLKBUF_X1 U25144 ( .A(n22714), .Z(n27196) );
  CLKBUF_X1 U25145 ( .A(n22712), .Z(n27202) );
  CLKBUF_X1 U25146 ( .A(n22711), .Z(n27208) );
  CLKBUF_X1 U25147 ( .A(n22709), .Z(n27214) );
  CLKBUF_X1 U25148 ( .A(n22708), .Z(n27220) );
  CLKBUF_X1 U25149 ( .A(n22706), .Z(n27226) );
  CLKBUF_X1 U25150 ( .A(n22705), .Z(n27232) );
  CLKBUF_X1 U25151 ( .A(n22703), .Z(n27238) );
  CLKBUF_X1 U25152 ( .A(n22702), .Z(n27244) );
  CLKBUF_X1 U25153 ( .A(n22700), .Z(n27250) );
  CLKBUF_X1 U25154 ( .A(n22699), .Z(n27256) );
  CLKBUF_X1 U25155 ( .A(n22697), .Z(n27262) );
  CLKBUF_X1 U25156 ( .A(n22696), .Z(n27268) );
  CLKBUF_X1 U25157 ( .A(n22693), .Z(n27274) );
  INV_X1 U25158 ( .A(ENABLE), .ZN(n27487) );
endmodule

