package constants is

  constant numBit : integer := 4;

end package constants;
