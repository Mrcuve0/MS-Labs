package constants is

  constant numBit : integer := 32;
  constant radixN : integer := 3;

end package constants;
