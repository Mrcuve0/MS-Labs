

package constants is

--library ieee;
--use ieee.math_real."log2";
  
  
  constant radixN : integer := 4;
  constant numBit : integer := 64;
  --constant rows : integer := integer(log2(real(numBit)));
  --constant rows : integer := 5;

end package constants;
