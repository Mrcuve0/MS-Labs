package constants is

  constant numBit : integer := 8;

end package constants;
