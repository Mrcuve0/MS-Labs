
module registers_N32_0 ( Clk, Rst, A, B, A_out, B_out );
  input [31:0] A;
  input [31:0] B;
  output [31:0] A_out;
  output [31:0] B_out;
  input Clk, Rst;
  wire   n128, n129, n130, n131, n132, n133, n134, n135, n136, n137;

  SDFF_X1 \B_out_reg[31]  ( .D(1'b0), .SI(n131), .SE(B[31]), .CK(Clk), .Q(
        B_out[31]) );
  SDFF_X1 \B_out_reg[30]  ( .D(1'b0), .SI(n131), .SE(B[30]), .CK(Clk), .Q(
        B_out[30]) );
  SDFF_X1 \B_out_reg[29]  ( .D(1'b0), .SI(n131), .SE(B[29]), .CK(Clk), .Q(
        B_out[29]) );
  SDFF_X1 \B_out_reg[28]  ( .D(1'b0), .SI(n130), .SE(B[28]), .CK(Clk), .Q(
        B_out[28]) );
  SDFF_X1 \B_out_reg[27]  ( .D(1'b0), .SI(n130), .SE(B[27]), .CK(Clk), .Q(
        B_out[27]) );
  SDFF_X1 \B_out_reg[26]  ( .D(1'b0), .SI(n130), .SE(B[26]), .CK(Clk), .Q(
        B_out[26]) );
  SDFF_X1 \B_out_reg[25]  ( .D(1'b0), .SI(n130), .SE(B[25]), .CK(Clk), .Q(
        B_out[25]) );
  SDFF_X1 \B_out_reg[24]  ( .D(1'b0), .SI(n130), .SE(B[24]), .CK(Clk), .Q(
        B_out[24]) );
  SDFF_X1 \B_out_reg[23]  ( .D(1'b0), .SI(n130), .SE(B[23]), .CK(Clk), .Q(
        B_out[23]) );
  SDFF_X1 \B_out_reg[22]  ( .D(1'b0), .SI(n130), .SE(B[22]), .CK(Clk), .Q(
        B_out[22]) );
  SDFF_X1 \B_out_reg[21]  ( .D(1'b0), .SI(n130), .SE(B[21]), .CK(Clk), .Q(
        B_out[21]) );
  SDFF_X1 \B_out_reg[20]  ( .D(1'b0), .SI(n130), .SE(B[20]), .CK(Clk), .Q(
        B_out[20]) );
  SDFF_X1 \B_out_reg[19]  ( .D(1'b0), .SI(n130), .SE(B[19]), .CK(Clk), .Q(
        B_out[19]) );
  SDFF_X1 \B_out_reg[18]  ( .D(1'b0), .SI(n129), .SE(B[18]), .CK(Clk), .Q(
        B_out[18]) );
  SDFF_X1 \B_out_reg[17]  ( .D(1'b0), .SI(n129), .SE(B[17]), .CK(Clk), .Q(
        B_out[17]) );
  SDFF_X1 \B_out_reg[16]  ( .D(1'b0), .SI(n129), .SE(B[16]), .CK(Clk), .Q(
        B_out[16]) );
  SDFF_X1 \B_out_reg[15]  ( .D(1'b0), .SI(n129), .SE(B[15]), .CK(Clk), .Q(
        B_out[15]) );
  SDFF_X1 \B_out_reg[14]  ( .D(1'b0), .SI(n129), .SE(B[14]), .CK(Clk), .Q(
        B_out[14]) );
  SDFF_X1 \B_out_reg[13]  ( .D(1'b0), .SI(n129), .SE(B[13]), .CK(Clk), .Q(
        B_out[13]) );
  SDFF_X1 \B_out_reg[12]  ( .D(1'b0), .SI(n129), .SE(B[12]), .CK(Clk), .Q(
        B_out[12]) );
  SDFF_X1 \B_out_reg[11]  ( .D(1'b0), .SI(n129), .SE(B[11]), .CK(Clk), .Q(
        B_out[11]) );
  SDFF_X1 \B_out_reg[10]  ( .D(1'b0), .SI(n129), .SE(B[10]), .CK(Clk), .Q(
        B_out[10]) );
  SDFF_X1 \B_out_reg[9]  ( .D(1'b0), .SI(n129), .SE(B[9]), .CK(Clk), .Q(
        B_out[9]) );
  SDFF_X1 \B_out_reg[8]  ( .D(1'b0), .SI(n128), .SE(B[8]), .CK(Clk), .Q(
        B_out[8]) );
  SDFF_X1 \B_out_reg[7]  ( .D(1'b0), .SI(n128), .SE(B[7]), .CK(Clk), .Q(
        B_out[7]) );
  SDFF_X1 \B_out_reg[6]  ( .D(1'b0), .SI(n128), .SE(B[6]), .CK(Clk), .Q(
        B_out[6]) );
  SDFF_X1 \B_out_reg[5]  ( .D(1'b0), .SI(n128), .SE(B[5]), .CK(Clk), .Q(
        B_out[5]) );
  SDFF_X1 \B_out_reg[4]  ( .D(1'b0), .SI(n128), .SE(B[4]), .CK(Clk), .Q(
        B_out[4]) );
  SDFF_X1 \B_out_reg[3]  ( .D(1'b0), .SI(n128), .SE(B[3]), .CK(Clk), .Q(
        B_out[3]) );
  SDFF_X1 \B_out_reg[2]  ( .D(1'b0), .SI(n128), .SE(B[2]), .CK(Clk), .Q(
        B_out[2]) );
  SDFF_X1 \B_out_reg[1]  ( .D(1'b0), .SI(n128), .SE(B[1]), .CK(Clk), .Q(
        B_out[1]) );
  SDFF_X1 \B_out_reg[0]  ( .D(1'b0), .SI(n128), .SE(B[0]), .CK(Clk), .Q(
        B_out[0]) );
  SDFF_X1 \A_out_reg[31]  ( .D(1'b0), .SI(n128), .SE(A[31]), .CK(Clk), .Q(
        A_out[31]) );
  SDFF_X1 \A_out_reg[0]  ( .D(1'b0), .SI(n131), .SE(A[0]), .CK(Clk), .Q(
        A_out[0]) );
  SDFF_X1 \A_out_reg[6]  ( .D(1'b0), .SI(n131), .SE(A[6]), .CK(Clk), .Q(
        A_out[6]) );
  SDFF_X1 \A_out_reg[4]  ( .D(1'b0), .SI(n131), .SE(A[4]), .CK(Clk), .Q(
        A_out[4]) );
  SDFF_X1 \A_out_reg[2]  ( .D(1'b0), .SI(n131), .SE(A[2]), .CK(Clk), .Q(
        A_out[2]) );
  SDFF_X1 \A_out_reg[7]  ( .D(1'b0), .SI(n131), .SE(A[7]), .CK(Clk), .Q(
        A_out[7]) );
  SDFF_X1 \A_out_reg[10]  ( .D(1'b0), .SI(n131), .SE(A[10]), .CK(Clk), .Q(
        A_out[10]) );
  SDFF_X1 \A_out_reg[5]  ( .D(1'b0), .SI(n131), .SE(A[5]), .CK(Clk), .Q(
        A_out[5]) );
  SDFF_X1 \A_out_reg[3]  ( .D(1'b0), .SI(n132), .SE(A[3]), .CK(Clk), .Q(
        A_out[3]) );
  SDFF_X1 \A_out_reg[1]  ( .D(1'b0), .SI(n132), .SE(A[1]), .CK(Clk), .Q(
        A_out[1]) );
  SDFF_X1 \A_out_reg[9]  ( .D(1'b0), .SI(n132), .SE(A[9]), .CK(Clk), .Q(
        A_out[9]) );
  SDFF_X1 \A_out_reg[8]  ( .D(1'b0), .SI(n132), .SE(A[8]), .CK(Clk), .Q(
        A_out[8]) );
  SDFF_X1 \A_out_reg[30]  ( .D(1'b0), .SI(n132), .SE(A[30]), .CK(Clk), .Q(
        A_out[30]) );
  SDFF_X1 \A_out_reg[29]  ( .D(1'b0), .SI(n132), .SE(A[29]), .CK(Clk), .Q(
        A_out[29]) );
  SDFF_X1 \A_out_reg[28]  ( .D(1'b0), .SI(n132), .SE(A[28]), .CK(Clk), .Q(
        A_out[28]) );
  SDFF_X1 \A_out_reg[27]  ( .D(1'b0), .SI(n132), .SE(A[27]), .CK(Clk), .Q(
        A_out[27]) );
  SDFF_X1 \A_out_reg[26]  ( .D(1'b0), .SI(n132), .SE(A[26]), .CK(Clk), .Q(
        A_out[26]) );
  SDFF_X1 \A_out_reg[25]  ( .D(1'b0), .SI(n132), .SE(A[25]), .CK(Clk), .Q(
        A_out[25]) );
  SDFF_X1 \A_out_reg[24]  ( .D(1'b0), .SI(n133), .SE(A[24]), .CK(Clk), .Q(
        A_out[24]) );
  SDFF_X1 \A_out_reg[23]  ( .D(1'b0), .SI(n133), .SE(A[23]), .CK(Clk), .Q(
        A_out[23]) );
  SDFF_X1 \A_out_reg[22]  ( .D(1'b0), .SI(n133), .SE(A[22]), .CK(Clk), .Q(
        A_out[22]) );
  SDFF_X1 \A_out_reg[21]  ( .D(1'b0), .SI(n133), .SE(A[21]), .CK(Clk), .Q(
        A_out[21]) );
  SDFF_X1 \A_out_reg[20]  ( .D(1'b0), .SI(n133), .SE(A[20]), .CK(Clk), .Q(
        A_out[20]) );
  SDFF_X1 \A_out_reg[19]  ( .D(1'b0), .SI(n133), .SE(A[19]), .CK(Clk), .Q(
        A_out[19]) );
  SDFF_X1 \A_out_reg[11]  ( .D(1'b0), .SI(n133), .SE(A[11]), .CK(Clk), .Q(
        A_out[11]) );
  SDFF_X1 \A_out_reg[12]  ( .D(1'b0), .SI(n133), .SE(A[12]), .CK(Clk), .Q(
        A_out[12]) );
  SDFF_X1 \A_out_reg[13]  ( .D(1'b0), .SI(n133), .SE(A[13]), .CK(Clk), .Q(
        A_out[13]) );
  SDFF_X1 \A_out_reg[14]  ( .D(1'b0), .SI(n133), .SE(A[14]), .CK(Clk), .Q(
        A_out[14]) );
  SDFF_X1 \A_out_reg[15]  ( .D(1'b0), .SI(n134), .SE(A[15]), .CK(Clk), .Q(
        A_out[15]) );
  SDFF_X1 \A_out_reg[16]  ( .D(1'b0), .SI(n134), .SE(A[16]), .CK(Clk), .Q(
        A_out[16]) );
  SDFF_X1 \A_out_reg[17]  ( .D(1'b0), .SI(n134), .SE(A[17]), .CK(Clk), .Q(
        A_out[17]) );
  SDFF_X1 \A_out_reg[18]  ( .D(1'b0), .SI(n134), .SE(A[18]), .CK(Clk), .Q(
        A_out[18]) );
  BUF_X1 U67 ( .A(n135), .Z(n133) );
  BUF_X1 U68 ( .A(n135), .Z(n132) );
  BUF_X1 U69 ( .A(n135), .Z(n131) );
  BUF_X1 U70 ( .A(n136), .Z(n128) );
  BUF_X1 U71 ( .A(n136), .Z(n129) );
  BUF_X1 U72 ( .A(n136), .Z(n130) );
  BUF_X1 U73 ( .A(n137), .Z(n135) );
  BUF_X1 U74 ( .A(n137), .Z(n136) );
  INV_X1 U75 ( .A(Rst), .ZN(n137) );
  CLKBUF_X1 U76 ( .A(n135), .Z(n134) );
endmodule


module encoder_N64_RADIX3_0 ( X, Z );
  input [2:0] X;
  output [2:0] Z;
  wire   n2, n3, n5;

  OAI21_X1 U1 ( .B1(X[1]), .B2(X[0]), .A(n3), .ZN(n2) );
  NAND2_X1 U2 ( .A1(X[1]), .A2(X[0]), .ZN(n3) );
  OAI22_X1 U3 ( .A1(n2), .A2(n5), .B1(X[2]), .B2(n3), .ZN(Z[1]) );
  AOI21_X1 U4 ( .B1(n2), .B2(n3), .A(X[2]), .ZN(Z[0]) );
  AND3_X1 U5 ( .A1(X[2]), .A2(n3), .A3(n2), .ZN(Z[2]) );
  INV_X1 U6 ( .A(X[2]), .ZN(n5) );
endmodule


module shifter_N64_0 ( \input , shiftLeftOnePos );
  input [63:0] \input ;
  output [63:0] shiftLeftOnePos;
  wire   \input[62] , \input[61] , \input[60] , \input[59] , \input[58] ,
         \input[57] , \input[56] , \input[55] , \input[54] , \input[53] ,
         \input[52] , \input[51] , \input[50] , \input[49] , \input[48] ,
         \input[47] , \input[46] , \input[45] , \input[44] , \input[43] ,
         \input[42] , \input[41] , \input[40] , \input[39] , \input[38] ,
         \input[37] , \input[36] , \input[35] , \input[34] , \input[33] ,
         \input[32] , \input[31] , \input[30] , \input[29] , \input[28] ,
         \input[27] , \input[26] , \input[25] , \input[24] , \input[23] ,
         \input[22] , \input[21] , \input[20] , \input[19] , \input[18] ,
         \input[17] , \input[16] , \input[15] , \input[14] , \input[13] ,
         \input[12] , \input[11] , \input[10] , \input[9] , \input[8] ,
         \input[7] , \input[6] , \input[5] , \input[4] , \input[3] ,
         \input[2] , \input[1] , \input[0] ;
  assign shiftLeftOnePos[0] = 1'b0;
  assign shiftLeftOnePos[63] = \input[62] ;
  assign \input[62]  = \input  [62];
  assign shiftLeftOnePos[62] = \input[61] ;
  assign \input[61]  = \input  [61];
  assign shiftLeftOnePos[61] = \input[60] ;
  assign \input[60]  = \input  [60];
  assign shiftLeftOnePos[60] = \input[59] ;
  assign \input[59]  = \input  [59];
  assign shiftLeftOnePos[59] = \input[58] ;
  assign \input[58]  = \input  [58];
  assign shiftLeftOnePos[58] = \input[57] ;
  assign \input[57]  = \input  [57];
  assign shiftLeftOnePos[57] = \input[56] ;
  assign \input[56]  = \input  [56];
  assign shiftLeftOnePos[56] = \input[55] ;
  assign \input[55]  = \input  [55];
  assign shiftLeftOnePos[55] = \input[54] ;
  assign \input[54]  = \input  [54];
  assign shiftLeftOnePos[54] = \input[53] ;
  assign \input[53]  = \input  [53];
  assign shiftLeftOnePos[53] = \input[52] ;
  assign \input[52]  = \input  [52];
  assign shiftLeftOnePos[52] = \input[51] ;
  assign \input[51]  = \input  [51];
  assign shiftLeftOnePos[51] = \input[50] ;
  assign \input[50]  = \input  [50];
  assign shiftLeftOnePos[50] = \input[49] ;
  assign \input[49]  = \input  [49];
  assign shiftLeftOnePos[49] = \input[48] ;
  assign \input[48]  = \input  [48];
  assign shiftLeftOnePos[48] = \input[47] ;
  assign \input[47]  = \input  [47];
  assign shiftLeftOnePos[47] = \input[46] ;
  assign \input[46]  = \input  [46];
  assign shiftLeftOnePos[46] = \input[45] ;
  assign \input[45]  = \input  [45];
  assign shiftLeftOnePos[45] = \input[44] ;
  assign \input[44]  = \input  [44];
  assign shiftLeftOnePos[44] = \input[43] ;
  assign \input[43]  = \input  [43];
  assign shiftLeftOnePos[43] = \input[42] ;
  assign \input[42]  = \input  [42];
  assign shiftLeftOnePos[42] = \input[41] ;
  assign \input[41]  = \input  [41];
  assign shiftLeftOnePos[41] = \input[40] ;
  assign \input[40]  = \input  [40];
  assign shiftLeftOnePos[40] = \input[39] ;
  assign \input[39]  = \input  [39];
  assign shiftLeftOnePos[39] = \input[38] ;
  assign \input[38]  = \input  [38];
  assign shiftLeftOnePos[38] = \input[37] ;
  assign \input[37]  = \input  [37];
  assign shiftLeftOnePos[37] = \input[36] ;
  assign \input[36]  = \input  [36];
  assign shiftLeftOnePos[36] = \input[35] ;
  assign \input[35]  = \input  [35];
  assign shiftLeftOnePos[35] = \input[34] ;
  assign \input[34]  = \input  [34];
  assign shiftLeftOnePos[34] = \input[33] ;
  assign \input[33]  = \input  [33];
  assign shiftLeftOnePos[33] = \input[32] ;
  assign \input[32]  = \input  [32];
  assign shiftLeftOnePos[32] = \input[31] ;
  assign \input[31]  = \input  [31];
  assign shiftLeftOnePos[31] = \input[30] ;
  assign \input[30]  = \input  [30];
  assign shiftLeftOnePos[30] = \input[29] ;
  assign \input[29]  = \input  [29];
  assign shiftLeftOnePos[29] = \input[28] ;
  assign \input[28]  = \input  [28];
  assign shiftLeftOnePos[28] = \input[27] ;
  assign \input[27]  = \input  [27];
  assign shiftLeftOnePos[27] = \input[26] ;
  assign \input[26]  = \input  [26];
  assign shiftLeftOnePos[26] = \input[25] ;
  assign \input[25]  = \input  [25];
  assign shiftLeftOnePos[25] = \input[24] ;
  assign \input[24]  = \input  [24];
  assign shiftLeftOnePos[24] = \input[23] ;
  assign \input[23]  = \input  [23];
  assign shiftLeftOnePos[23] = \input[22] ;
  assign \input[22]  = \input  [22];
  assign shiftLeftOnePos[22] = \input[21] ;
  assign \input[21]  = \input  [21];
  assign shiftLeftOnePos[21] = \input[20] ;
  assign \input[20]  = \input  [20];
  assign shiftLeftOnePos[20] = \input[19] ;
  assign \input[19]  = \input  [19];
  assign shiftLeftOnePos[19] = \input[18] ;
  assign \input[18]  = \input  [18];
  assign shiftLeftOnePos[18] = \input[17] ;
  assign \input[17]  = \input  [17];
  assign shiftLeftOnePos[17] = \input[16] ;
  assign \input[16]  = \input  [16];
  assign shiftLeftOnePos[16] = \input[15] ;
  assign \input[15]  = \input  [15];
  assign shiftLeftOnePos[15] = \input[14] ;
  assign \input[14]  = \input  [14];
  assign shiftLeftOnePos[14] = \input[13] ;
  assign \input[13]  = \input  [13];
  assign shiftLeftOnePos[13] = \input[12] ;
  assign \input[12]  = \input  [12];
  assign shiftLeftOnePos[12] = \input[11] ;
  assign \input[11]  = \input  [11];
  assign shiftLeftOnePos[11] = \input[10] ;
  assign \input[10]  = \input  [10];
  assign shiftLeftOnePos[10] = \input[9] ;
  assign \input[9]  = \input  [9];
  assign shiftLeftOnePos[9] = \input[8] ;
  assign \input[8]  = \input  [8];
  assign shiftLeftOnePos[8] = \input[7] ;
  assign \input[7]  = \input  [7];
  assign shiftLeftOnePos[7] = \input[6] ;
  assign \input[6]  = \input  [6];
  assign shiftLeftOnePos[6] = \input[5] ;
  assign \input[5]  = \input  [5];
  assign shiftLeftOnePos[5] = \input[4] ;
  assign \input[4]  = \input  [4];
  assign shiftLeftOnePos[4] = \input[3] ;
  assign \input[3]  = \input  [3];
  assign shiftLeftOnePos[3] = \input[2] ;
  assign \input[2]  = \input  [2];
  assign shiftLeftOnePos[2] = \input[1] ;
  assign \input[1]  = \input  [1];
  assign shiftLeftOnePos[1] = \input[0] ;
  assign \input[0]  = \input  [0];

endmodule


module complementer_N64_0_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n190, n191, n192, n194, n196, n197, n198, n199, n200, n202,
         n203, n204, n206, n207, n208, n210, n211, n212, n213, n214, n216,
         n217, n218, n220, n221, n222, n224, n225, n226, n228, n229, n230,
         n232, n233, n234, n235, n237, n238, n239, n241, n242, n243, n245,
         n246, n247, n249, n250, n189, n193, n195, n201, n205, n209, n215,
         n219, n223, n227, n231, n236, n240, n244, n248, n251;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U81 ( .A(n190), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U82 ( .A(n192), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U85 ( .A(n196), .B(B[62]), .Z(DIFF[62]) );
  XOR2_X1 U86 ( .A(n194), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U87 ( .A(n198), .B(B[59]), .Z(DIFF[59]) );
  XOR2_X1 U89 ( .A(n200), .B(B[57]), .Z(DIFF[57]) );
  XOR2_X1 U90 ( .A(n202), .B(B[55]), .Z(DIFF[55]) );
  XOR2_X1 U92 ( .A(n204), .B(B[53]), .Z(DIFF[53]) );
  XOR2_X1 U93 ( .A(n206), .B(B[51]), .Z(DIFF[51]) );
  XOR2_X1 U95 ( .A(n208), .B(B[49]), .Z(DIFF[49]) );
  XOR2_X1 U96 ( .A(n212), .B(B[47]), .Z(DIFF[47]) );
  XOR2_X1 U98 ( .A(n214), .B(B[45]), .Z(DIFF[45]) );
  XOR2_X1 U99 ( .A(n216), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U101 ( .A(n218), .B(B[41]), .Z(DIFF[41]) );
  XOR2_X1 U102 ( .A(n211), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U103 ( .A(n220), .B(B[39]), .Z(DIFF[39]) );
  XOR2_X1 U105 ( .A(n222), .B(B[37]), .Z(DIFF[37]) );
  XOR2_X1 U106 ( .A(n224), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U108 ( .A(n226), .B(B[33]), .Z(DIFF[33]) );
  XOR2_X1 U109 ( .A(n228), .B(B[31]), .Z(DIFF[31]) );
  XOR2_X1 U111 ( .A(n230), .B(B[29]), .Z(DIFF[29]) );
  XOR2_X1 U112 ( .A(n233), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U114 ( .A(n235), .B(B[25]), .Z(DIFF[25]) );
  XOR2_X1 U115 ( .A(n237), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U117 ( .A(n239), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U118 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U119 ( .A(n241), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U121 ( .A(n243), .B(B[17]), .Z(DIFF[17]) );
  XOR2_X1 U122 ( .A(n245), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U124 ( .A(n247), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U125 ( .A(n249), .B(B[11]), .Z(DIFF[11]) );
  XOR2_X1 U1 ( .A(n197), .B(n251), .Z(DIFF[61]) );
  NAND2_X1 U2 ( .A1(n197), .A2(n251), .ZN(n196) );
  XNOR2_X1 U3 ( .A(n189), .B(B[34]), .ZN(DIFF[34]) );
  NOR2_X1 U4 ( .A1(n226), .A2(B[33]), .ZN(n189) );
  XNOR2_X1 U5 ( .A(B[36]), .B(n225), .ZN(DIFF[36]) );
  NOR2_X1 U6 ( .A1(B[35]), .A2(n224), .ZN(n225) );
  XNOR2_X1 U7 ( .A(B[40]), .B(n221), .ZN(DIFF[40]) );
  NOR2_X1 U8 ( .A1(B[39]), .A2(n220), .ZN(n221) );
  XNOR2_X1 U9 ( .A(B[44]), .B(n217), .ZN(DIFF[44]) );
  NOR2_X1 U10 ( .A1(B[43]), .A2(n216), .ZN(n217) );
  XNOR2_X1 U11 ( .A(n193), .B(B[38]), .ZN(DIFF[38]) );
  NOR2_X1 U12 ( .A1(n222), .A2(B[37]), .ZN(n193) );
  OR3_X1 U13 ( .A1(B[37]), .A2(B[38]), .A3(n222), .ZN(n220) );
  OR3_X1 U14 ( .A1(B[41]), .A2(B[42]), .A3(n218), .ZN(n216) );
  OR3_X1 U15 ( .A1(B[35]), .A2(B[36]), .A3(n224), .ZN(n222) );
  OR3_X1 U16 ( .A1(B[39]), .A2(B[40]), .A3(n220), .ZN(n218) );
  OR3_X1 U17 ( .A1(B[33]), .A2(B[34]), .A3(n226), .ZN(n224) );
  OR3_X1 U18 ( .A1(B[43]), .A2(B[44]), .A3(n216), .ZN(n214) );
  XNOR2_X1 U19 ( .A(n195), .B(B[42]), .ZN(DIFF[42]) );
  NOR2_X1 U20 ( .A1(n218), .A2(B[41]), .ZN(n195) );
  NOR3_X1 U21 ( .A1(B[59]), .A2(B[60]), .A3(n198), .ZN(n197) );
  XNOR2_X1 U22 ( .A(B[56]), .B(n203), .ZN(DIFF[56]) );
  NOR2_X1 U23 ( .A1(B[55]), .A2(n202), .ZN(n203) );
  XNOR2_X1 U24 ( .A(B[60]), .B(n199), .ZN(DIFF[60]) );
  NOR2_X1 U25 ( .A1(B[59]), .A2(n198), .ZN(n199) );
  XNOR2_X1 U26 ( .A(n201), .B(B[58]), .ZN(DIFF[58]) );
  NOR2_X1 U27 ( .A1(n200), .A2(B[57]), .ZN(n201) );
  XNOR2_X1 U28 ( .A(B[48]), .B(n213), .ZN(DIFF[48]) );
  NOR2_X1 U29 ( .A1(B[47]), .A2(n212), .ZN(n213) );
  XNOR2_X1 U30 ( .A(B[52]), .B(n207), .ZN(DIFF[52]) );
  NOR2_X1 U31 ( .A1(B[51]), .A2(n206), .ZN(n207) );
  OR3_X1 U32 ( .A1(B[45]), .A2(B[46]), .A3(n214), .ZN(n212) );
  OR3_X1 U33 ( .A1(B[49]), .A2(B[50]), .A3(n208), .ZN(n206) );
  OR3_X1 U34 ( .A1(B[47]), .A2(B[48]), .A3(n212), .ZN(n208) );
  OR3_X1 U35 ( .A1(B[51]), .A2(B[52]), .A3(n206), .ZN(n204) );
  OR3_X1 U36 ( .A1(B[55]), .A2(B[56]), .A3(n202), .ZN(n200) );
  OR3_X1 U37 ( .A1(B[53]), .A2(B[54]), .A3(n204), .ZN(n202) );
  OR3_X1 U38 ( .A1(B[57]), .A2(B[58]), .A3(n200), .ZN(n198) );
  XNOR2_X1 U39 ( .A(n205), .B(B[63]), .ZN(DIFF[63]) );
  NOR2_X1 U40 ( .A1(n196), .A2(B[62]), .ZN(n205) );
  XNOR2_X1 U41 ( .A(n209), .B(B[50]), .ZN(DIFF[50]) );
  NOR2_X1 U42 ( .A1(n208), .A2(B[49]), .ZN(n209) );
  XNOR2_X1 U43 ( .A(n215), .B(B[46]), .ZN(DIFF[46]) );
  NOR2_X1 U44 ( .A1(n214), .A2(B[45]), .ZN(n215) );
  XNOR2_X1 U45 ( .A(n219), .B(B[54]), .ZN(DIFF[54]) );
  NOR2_X1 U46 ( .A1(n204), .A2(B[53]), .ZN(n219) );
  XNOR2_X1 U47 ( .A(B[32]), .B(n229), .ZN(DIFF[32]) );
  NOR2_X1 U48 ( .A1(B[31]), .A2(n228), .ZN(n229) );
  OR3_X1 U49 ( .A1(B[31]), .A2(B[32]), .A3(n228), .ZN(n226) );
  XNOR2_X1 U50 ( .A(n223), .B(B[18]), .ZN(DIFF[18]) );
  NOR2_X1 U51 ( .A1(n243), .A2(B[17]), .ZN(n223) );
  XNOR2_X1 U52 ( .A(n227), .B(B[14]), .ZN(DIFF[14]) );
  NOR2_X1 U53 ( .A1(n247), .A2(B[13]), .ZN(n227) );
  XNOR2_X1 U54 ( .A(n231), .B(B[10]), .ZN(DIFF[10]) );
  NOR2_X1 U55 ( .A1(n190), .A2(B[9]), .ZN(n231) );
  XNOR2_X1 U56 ( .A(n236), .B(B[6]), .ZN(DIFF[6]) );
  NOR2_X1 U57 ( .A1(n194), .A2(B[5]), .ZN(n236) );
  XNOR2_X1 U58 ( .A(B[2]), .B(n232), .ZN(DIFF[2]) );
  NOR2_X1 U59 ( .A1(\B[0] ), .A2(B[1]), .ZN(n232) );
  XNOR2_X1 U60 ( .A(B[16]), .B(n246), .ZN(DIFF[16]) );
  NOR2_X1 U61 ( .A1(B[15]), .A2(n245), .ZN(n246) );
  XNOR2_X1 U62 ( .A(B[12]), .B(n250), .ZN(DIFF[12]) );
  NOR2_X1 U63 ( .A1(B[11]), .A2(n249), .ZN(n250) );
  XNOR2_X1 U64 ( .A(B[8]), .B(n191), .ZN(DIFF[8]) );
  NOR2_X1 U65 ( .A1(B[7]), .A2(n192), .ZN(n191) );
  XNOR2_X1 U66 ( .A(B[4]), .B(n210), .ZN(DIFF[4]) );
  NOR2_X1 U67 ( .A1(B[3]), .A2(n211), .ZN(n210) );
  OR3_X1 U68 ( .A1(B[1]), .A2(B[2]), .A3(\B[0] ), .ZN(n211) );
  OR3_X1 U69 ( .A1(B[5]), .A2(B[6]), .A3(n194), .ZN(n192) );
  OR3_X1 U70 ( .A1(B[13]), .A2(B[14]), .A3(n247), .ZN(n245) );
  OR3_X1 U71 ( .A1(B[17]), .A2(B[18]), .A3(n243), .ZN(n241) );
  OR3_X1 U72 ( .A1(B[10]), .A2(B[9]), .A3(n190), .ZN(n249) );
  OR3_X1 U73 ( .A1(B[3]), .A2(B[4]), .A3(n211), .ZN(n194) );
  OR3_X1 U74 ( .A1(B[7]), .A2(B[8]), .A3(n192), .ZN(n190) );
  OR3_X1 U75 ( .A1(B[11]), .A2(B[12]), .A3(n249), .ZN(n247) );
  OR3_X1 U76 ( .A1(B[15]), .A2(B[16]), .A3(n245), .ZN(n243) );
  XNOR2_X1 U77 ( .A(n240), .B(B[26]), .ZN(DIFF[26]) );
  NOR2_X1 U78 ( .A1(n235), .A2(B[25]), .ZN(n240) );
  XNOR2_X1 U79 ( .A(n244), .B(B[22]), .ZN(DIFF[22]) );
  NOR2_X1 U80 ( .A1(n239), .A2(B[21]), .ZN(n244) );
  XNOR2_X1 U83 ( .A(n248), .B(B[30]), .ZN(DIFF[30]) );
  NOR2_X1 U84 ( .A1(n230), .A2(B[29]), .ZN(n248) );
  XNOR2_X1 U88 ( .A(B[28]), .B(n234), .ZN(DIFF[28]) );
  NOR2_X1 U91 ( .A1(B[27]), .A2(n233), .ZN(n234) );
  XNOR2_X1 U94 ( .A(B[24]), .B(n238), .ZN(DIFF[24]) );
  NOR2_X1 U97 ( .A1(B[23]), .A2(n237), .ZN(n238) );
  XNOR2_X1 U100 ( .A(B[20]), .B(n242), .ZN(DIFF[20]) );
  NOR2_X1 U104 ( .A1(B[19]), .A2(n241), .ZN(n242) );
  OR3_X1 U107 ( .A1(B[21]), .A2(B[22]), .A3(n239), .ZN(n237) );
  OR3_X1 U110 ( .A1(B[25]), .A2(B[26]), .A3(n235), .ZN(n233) );
  OR3_X1 U113 ( .A1(B[29]), .A2(B[30]), .A3(n230), .ZN(n228) );
  OR3_X1 U116 ( .A1(B[19]), .A2(B[20]), .A3(n241), .ZN(n239) );
  OR3_X1 U120 ( .A1(B[23]), .A2(B[24]), .A3(n237), .ZN(n235) );
  OR3_X1 U123 ( .A1(B[27]), .A2(B[28]), .A3(n233), .ZN(n230) );
  INV_X1 U126 ( .A(B[61]), .ZN(n251) );
endmodule


module complementer_N64_0 ( \input , complement2 );
  input [63:0] \input ;
  output [63:0] complement2;


  complementer_N64_0_DW01_sub_0 sub_add_31_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(\input ), .CI(1'b0), .DIFF(complement2) );
endmodule


module complementer_N64_31_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n189;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U81 ( .A(n190), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U82 ( .A(n192), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U83 ( .A(n193), .B(B[6]), .Z(DIFF[6]) );
  XOR2_X1 U84 ( .A(n195), .B(B[63]), .Z(DIFF[63]) );
  XOR2_X1 U85 ( .A(n196), .B(B[62]), .Z(DIFF[62]) );
  XOR2_X1 U86 ( .A(n194), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U87 ( .A(n198), .B(B[59]), .Z(DIFF[59]) );
  XOR2_X1 U88 ( .A(n201), .B(B[58]), .Z(DIFF[58]) );
  XOR2_X1 U89 ( .A(n200), .B(B[57]), .Z(DIFF[57]) );
  XOR2_X1 U90 ( .A(n202), .B(B[55]), .Z(DIFF[55]) );
  XOR2_X1 U91 ( .A(n205), .B(B[54]), .Z(DIFF[54]) );
  XOR2_X1 U92 ( .A(n204), .B(B[53]), .Z(DIFF[53]) );
  XOR2_X1 U93 ( .A(n206), .B(B[51]), .Z(DIFF[51]) );
  XOR2_X1 U94 ( .A(n209), .B(B[50]), .Z(DIFF[50]) );
  XOR2_X1 U95 ( .A(n208), .B(B[49]), .Z(DIFF[49]) );
  XOR2_X1 U96 ( .A(n212), .B(B[47]), .Z(DIFF[47]) );
  XOR2_X1 U97 ( .A(n215), .B(B[46]), .Z(DIFF[46]) );
  XOR2_X1 U98 ( .A(n214), .B(B[45]), .Z(DIFF[45]) );
  XOR2_X1 U99 ( .A(n216), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U100 ( .A(n219), .B(B[42]), .Z(DIFF[42]) );
  XOR2_X1 U101 ( .A(n218), .B(B[41]), .Z(DIFF[41]) );
  XOR2_X1 U102 ( .A(n211), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U103 ( .A(n220), .B(B[39]), .Z(DIFF[39]) );
  XOR2_X1 U104 ( .A(n223), .B(B[38]), .Z(DIFF[38]) );
  XOR2_X1 U105 ( .A(n222), .B(B[37]), .Z(DIFF[37]) );
  XOR2_X1 U106 ( .A(n224), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U107 ( .A(n227), .B(B[34]), .Z(DIFF[34]) );
  XOR2_X1 U108 ( .A(n226), .B(B[33]), .Z(DIFF[33]) );
  XOR2_X1 U109 ( .A(n228), .B(B[31]), .Z(DIFF[31]) );
  XOR2_X1 U110 ( .A(n231), .B(B[30]), .Z(DIFF[30]) );
  XOR2_X1 U111 ( .A(n230), .B(B[29]), .Z(DIFF[29]) );
  XOR2_X1 U112 ( .A(n233), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U113 ( .A(n236), .B(B[26]), .Z(DIFF[26]) );
  XOR2_X1 U114 ( .A(n235), .B(B[25]), .Z(DIFF[25]) );
  XOR2_X1 U115 ( .A(n237), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U116 ( .A(n240), .B(B[22]), .Z(DIFF[22]) );
  XOR2_X1 U117 ( .A(n239), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U118 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U119 ( .A(n241), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U120 ( .A(n244), .B(B[18]), .Z(DIFF[18]) );
  XOR2_X1 U121 ( .A(n243), .B(B[17]), .Z(DIFF[17]) );
  XOR2_X1 U122 ( .A(n245), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U123 ( .A(n248), .B(B[14]), .Z(DIFF[14]) );
  XOR2_X1 U124 ( .A(n247), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U125 ( .A(n249), .B(B[11]), .Z(DIFF[11]) );
  XOR2_X1 U126 ( .A(n251), .B(B[10]), .Z(DIFF[10]) );
  NOR2_X1 U1 ( .A1(B[43]), .A2(n216), .ZN(n217) );
  NOR2_X1 U2 ( .A1(B[39]), .A2(n220), .ZN(n221) );
  NOR2_X1 U3 ( .A1(B[59]), .A2(n198), .ZN(n199) );
  NAND2_X1 U4 ( .A1(n197), .A2(n189), .ZN(n196) );
  OR3_X1 U5 ( .A1(B[53]), .A2(B[54]), .A3(n204), .ZN(n202) );
  OR3_X1 U6 ( .A1(B[43]), .A2(B[44]), .A3(n216), .ZN(n214) );
  XNOR2_X1 U7 ( .A(B[48]), .B(n213), .ZN(DIFF[48]) );
  OR2_X1 U8 ( .A1(n204), .A2(B[53]), .ZN(n205) );
  OR2_X1 U9 ( .A1(n208), .A2(B[49]), .ZN(n209) );
  NOR2_X1 U10 ( .A1(B[35]), .A2(n224), .ZN(n225) );
  XNOR2_X1 U11 ( .A(B[32]), .B(n229), .ZN(DIFF[32]) );
  OR3_X1 U12 ( .A1(B[37]), .A2(B[38]), .A3(n222), .ZN(n220) );
  OR3_X1 U13 ( .A1(B[41]), .A2(B[42]), .A3(n218), .ZN(n216) );
  OR3_X1 U14 ( .A1(B[35]), .A2(B[36]), .A3(n224), .ZN(n222) );
  OR3_X1 U15 ( .A1(B[39]), .A2(B[40]), .A3(n220), .ZN(n218) );
  XNOR2_X1 U16 ( .A(B[36]), .B(n225), .ZN(DIFF[36]) );
  XNOR2_X1 U17 ( .A(B[40]), .B(n221), .ZN(DIFF[40]) );
  XNOR2_X1 U18 ( .A(B[44]), .B(n217), .ZN(DIFF[44]) );
  OR3_X1 U19 ( .A1(B[33]), .A2(B[34]), .A3(n226), .ZN(n224) );
  OR2_X1 U20 ( .A1(n222), .A2(B[37]), .ZN(n223) );
  OR2_X1 U21 ( .A1(n218), .A2(B[41]), .ZN(n219) );
  OR2_X1 U22 ( .A1(n226), .A2(B[33]), .ZN(n227) );
  NOR3_X1 U23 ( .A1(B[59]), .A2(B[60]), .A3(n198), .ZN(n197) );
  NOR2_X1 U24 ( .A1(B[47]), .A2(n212), .ZN(n213) );
  NOR2_X1 U25 ( .A1(B[51]), .A2(n206), .ZN(n207) );
  NOR2_X1 U26 ( .A1(B[55]), .A2(n202), .ZN(n203) );
  OR3_X1 U27 ( .A1(B[57]), .A2(B[58]), .A3(n200), .ZN(n198) );
  OR3_X1 U28 ( .A1(B[45]), .A2(B[46]), .A3(n214), .ZN(n212) );
  OR3_X1 U29 ( .A1(B[47]), .A2(B[48]), .A3(n212), .ZN(n208) );
  OR3_X1 U30 ( .A1(B[51]), .A2(B[52]), .A3(n206), .ZN(n204) );
  OR3_X1 U31 ( .A1(B[55]), .A2(B[56]), .A3(n202), .ZN(n200) );
  OR3_X1 U32 ( .A1(B[49]), .A2(B[50]), .A3(n208), .ZN(n206) );
  XNOR2_X1 U33 ( .A(n197), .B(B[61]), .ZN(DIFF[61]) );
  XNOR2_X1 U34 ( .A(B[52]), .B(n207), .ZN(DIFF[52]) );
  XNOR2_X1 U35 ( .A(B[56]), .B(n203), .ZN(DIFF[56]) );
  XNOR2_X1 U36 ( .A(B[60]), .B(n199), .ZN(DIFF[60]) );
  OR2_X1 U37 ( .A1(n200), .A2(B[57]), .ZN(n201) );
  OR2_X1 U38 ( .A1(n196), .A2(B[62]), .ZN(n195) );
  OR2_X1 U39 ( .A1(n214), .A2(B[45]), .ZN(n215) );
  NOR2_X1 U40 ( .A1(B[31]), .A2(n228), .ZN(n229) );
  OR3_X1 U41 ( .A1(B[31]), .A2(B[32]), .A3(n228), .ZN(n226) );
  XNOR2_X1 U42 ( .A(B[16]), .B(n246), .ZN(DIFF[16]) );
  NOR2_X1 U43 ( .A1(B[3]), .A2(n211), .ZN(n210) );
  NOR2_X1 U44 ( .A1(B[15]), .A2(n245), .ZN(n246) );
  NOR2_X1 U45 ( .A1(B[11]), .A2(n249), .ZN(n250) );
  NOR2_X1 U46 ( .A1(B[7]), .A2(n192), .ZN(n191) );
  NOR2_X1 U47 ( .A1(\B[0] ), .A2(B[1]), .ZN(n232) );
  OR3_X1 U48 ( .A1(B[1]), .A2(B[2]), .A3(\B[0] ), .ZN(n211) );
  OR3_X1 U49 ( .A1(B[10]), .A2(B[9]), .A3(n190), .ZN(n249) );
  OR3_X1 U50 ( .A1(B[17]), .A2(B[18]), .A3(n243), .ZN(n241) );
  OR3_X1 U51 ( .A1(B[13]), .A2(B[14]), .A3(n247), .ZN(n245) );
  OR3_X1 U52 ( .A1(B[5]), .A2(B[6]), .A3(n194), .ZN(n192) );
  OR3_X1 U53 ( .A1(B[15]), .A2(B[16]), .A3(n245), .ZN(n243) );
  OR3_X1 U54 ( .A1(B[11]), .A2(B[12]), .A3(n249), .ZN(n247) );
  OR3_X1 U55 ( .A1(B[7]), .A2(B[8]), .A3(n192), .ZN(n190) );
  OR3_X1 U56 ( .A1(B[3]), .A2(B[4]), .A3(n211), .ZN(n194) );
  XNOR2_X1 U57 ( .A(B[12]), .B(n250), .ZN(DIFF[12]) );
  XNOR2_X1 U58 ( .A(B[8]), .B(n191), .ZN(DIFF[8]) );
  XNOR2_X1 U59 ( .A(B[4]), .B(n210), .ZN(DIFF[4]) );
  XNOR2_X1 U60 ( .A(B[2]), .B(n232), .ZN(DIFF[2]) );
  OR2_X1 U61 ( .A1(n243), .A2(B[17]), .ZN(n244) );
  OR2_X1 U62 ( .A1(n247), .A2(B[13]), .ZN(n248) );
  OR2_X1 U63 ( .A1(n190), .A2(B[9]), .ZN(n251) );
  OR2_X1 U64 ( .A1(n194), .A2(B[5]), .ZN(n193) );
  XNOR2_X1 U65 ( .A(B[28]), .B(n234), .ZN(DIFF[28]) );
  XNOR2_X1 U66 ( .A(B[24]), .B(n238), .ZN(DIFF[24]) );
  XNOR2_X1 U67 ( .A(B[20]), .B(n242), .ZN(DIFF[20]) );
  NOR2_X1 U68 ( .A1(B[27]), .A2(n233), .ZN(n234) );
  NOR2_X1 U69 ( .A1(B[23]), .A2(n237), .ZN(n238) );
  NOR2_X1 U70 ( .A1(B[19]), .A2(n241), .ZN(n242) );
  OR3_X1 U71 ( .A1(B[29]), .A2(B[30]), .A3(n230), .ZN(n228) );
  OR3_X1 U72 ( .A1(B[25]), .A2(B[26]), .A3(n235), .ZN(n233) );
  OR3_X1 U73 ( .A1(B[21]), .A2(B[22]), .A3(n239), .ZN(n237) );
  OR3_X1 U74 ( .A1(B[27]), .A2(B[28]), .A3(n233), .ZN(n230) );
  OR3_X1 U75 ( .A1(B[23]), .A2(B[24]), .A3(n237), .ZN(n235) );
  OR3_X1 U76 ( .A1(B[19]), .A2(B[20]), .A3(n241), .ZN(n239) );
  OR2_X1 U77 ( .A1(n230), .A2(B[29]), .ZN(n231) );
  OR2_X1 U78 ( .A1(n235), .A2(B[25]), .ZN(n236) );
  OR2_X1 U79 ( .A1(n239), .A2(B[21]), .ZN(n240) );
  INV_X1 U80 ( .A(B[61]), .ZN(n189) );
endmodule


module complementer_N64_31 ( \input , complement2 );
  input [63:0] \input ;
  output [63:0] complement2;


  complementer_N64_31_DW01_sub_0 sub_add_31_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(\input ), .CI(1'b0), .DIFF(complement2) );
endmodule


module ShiftnCompl_special_N64 ( plusA, plusA_out, minusA_out, plus2A_out, 
        minus2A_out );
  input [63:0] plusA;
  output [63:0] plusA_out;
  output [63:0] minusA_out;
  output [63:0] plus2A_out;
  output [63:0] minus2A_out;
  wire   n17, n18, n19, n20, n21, n22, n23, n24;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign plusA_out[63] = plusA[63];
  assign plusA_out[62] = plusA[62];
  assign plusA_out[61] = plusA[61];
  assign plusA_out[60] = plusA[60];
  assign plusA_out[59] = plusA[59];
  assign plusA_out[57] = plusA[57];
  assign plusA_out[56] = plusA[56];
  assign plusA_out[55] = plusA[55];
  assign plusA_out[54] = plusA[54];
  assign plusA_out[52] = plusA[52];
  assign plusA_out[51] = plusA[51];
  assign plusA_out[50] = plusA[50];
  assign plusA_out[49] = plusA[49];
  assign plusA_out[47] = plusA[47];
  assign plusA_out[46] = plusA[46];
  assign plusA_out[45] = plusA[45];
  assign plusA_out[44] = plusA[44];
  assign plusA_out[42] = plusA[42];
  assign plusA_out[41] = plusA[41];
  assign plusA_out[40] = plusA[40];
  assign plusA_out[39] = plusA[39];
  assign plusA_out[37] = plusA[37];
  assign plusA_out[36] = plusA[36];
  assign plusA_out[35] = plusA[35];
  assign plusA_out[34] = plusA[34];
  assign plusA_out[32] = plusA[32];
  assign plusA_out[31] = plusA[31];
  assign plusA_out[30] = plusA[30];
  assign plusA_out[29] = plusA[29];
  assign plusA_out[28] = plusA[28];
  assign plusA_out[27] = plusA[27];
  assign plusA_out[26] = plusA[26];
  assign plusA_out[25] = plusA[25];
  assign plusA_out[24] = plusA[24];
  assign plusA_out[23] = plusA[23];
  assign plusA_out[22] = plusA[22];
  assign plusA_out[21] = plusA[21];
  assign plusA_out[20] = plusA[20];
  assign plusA_out[19] = plusA[19];
  assign plusA_out[18] = plusA[18];
  assign plusA_out[17] = plusA[17];
  assign plusA_out[16] = plusA[16];
  assign plusA_out[15] = plusA[15];
  assign plusA_out[14] = plusA[14];
  assign plusA_out[13] = plusA[13];
  assign plusA_out[12] = plusA[12];
  assign plusA_out[11] = plusA[11];
  assign plusA_out[10] = plusA[10];
  assign plusA_out[9] = plusA[9];
  assign plusA_out[8] = plusA[8];
  assign plusA_out[7] = plusA[7];
  assign plusA_out[6] = plusA[6];
  assign plusA_out[5] = plusA[5];
  assign plusA_out[4] = plusA[4];
  assign plusA_out[3] = plusA[3];
  assign plusA_out[2] = plusA[2];
  assign plusA_out[1] = plusA[1];
  assign plusA_out[0] = plusA[0];
  assign plus2A_out[0] = 1'b0;

  shifter_N64_0 shifter_1 ( .\input ({plusA[63:59], plusA_out[58], 
        plusA[57:54], plusA_out[53], plusA[52:49], plusA_out[48], plusA[47:44], 
        plusA_out[43], plusA[42:39], plusA_out[38], plusA[37:34], 
        plusA_out[33], plusA[32:0]}), .shiftLeftOnePos({plus2A_out[63:59], n17, 
        plus2A_out[57:54], n18, plus2A_out[52:49], n19, plus2A_out[47:44], n20, 
        plus2A_out[42:39], n21, plus2A_out[37:34], n22, n23, n24, 
        plus2A_out[30:1], SYNOPSYS_UNCONNECTED__0}) );
  complementer_N64_0 complementer_1 ( .\input ({plusA[63:59], plusA_out[58], 
        plusA[57:54], plusA_out[53], plusA[52:49], plusA_out[48], plusA[47:44], 
        plusA_out[43], plusA[42:39], plusA_out[38], plusA[37:34], 
        plusA_out[33], plusA[32:0]}), .complement2(minusA_out) );
  complementer_N64_31 complementer_2 ( .\input ({plus2A_out[63:1], 1'b0}), 
        .complement2(minus2A_out) );
  BUF_X1 U1 ( .A(plusA[43]), .Z(plusA_out[43]) );
  BUF_X1 U2 ( .A(plusA[33]), .Z(plusA_out[33]) );
  BUF_X1 U4 ( .A(n22), .Z(plus2A_out[33]) );
  BUF_X1 U5 ( .A(n21), .Z(plus2A_out[38]) );
  BUF_X1 U6 ( .A(plusA[38]), .Z(plusA_out[38]) );
  BUF_X1 U7 ( .A(plusA[53]), .Z(plusA_out[53]) );
  BUF_X1 U8 ( .A(n20), .Z(plus2A_out[43]) );
  BUF_X1 U9 ( .A(n19), .Z(plus2A_out[48]) );
  BUF_X1 U10 ( .A(plusA[48]), .Z(plusA_out[48]) );
  BUF_X1 U11 ( .A(n18), .Z(plus2A_out[53]) );
  BUF_X1 U12 ( .A(plusA[58]), .Z(plusA_out[58]) );
  BUF_X1 U13 ( .A(n17), .Z(plus2A_out[58]) );
  BUF_X1 U14 ( .A(n24), .Z(plus2A_out[31]) );
  BUF_X1 U15 ( .A(n23), .Z(plus2A_out[32]) );
endmodule


module MUX_GENERIC_N64_RADIX3_0 ( plusA, minusA, plus2A, minus2A, SEL, Y );
  input [63:0] plusA;
  input [63:0] minusA;
  input [63:0] plus2A;
  input [63:0] minus2A;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304;
  tri   [63:0] Y;

  TBUF_X1 \Y_tri[1]  ( .A(n208), .EN(n296), .Z(Y[1]) );
  TBUF_X1 \Y_tri[55]  ( .A(n263), .EN(n301), .Z(Y[55]) );
  TBUF_X1 \Y_tri[56]  ( .A(n264), .EN(n301), .Z(Y[56]) );
  TBUF_X1 \Y_tri[57]  ( .A(n265), .EN(n301), .Z(Y[57]) );
  TBUF_X1 \Y_tri[58]  ( .A(n266), .EN(n301), .Z(Y[58]) );
  TBUF_X1 \Y_tri[59]  ( .A(n267), .EN(n301), .Z(Y[59]) );
  TBUF_X1 \Y_tri[60]  ( .A(n268), .EN(n301), .Z(Y[60]) );
  TBUF_X1 \Y_tri[61]  ( .A(n269), .EN(n301), .Z(Y[61]) );
  TBUF_X1 \Y_tri[62]  ( .A(n270), .EN(n301), .Z(Y[62]) );
  TBUF_X1 \Y_tri[63]  ( .A(n271), .EN(n301), .Z(Y[63]) );
  TBUF_X1 \Y_tri[46]  ( .A(n254), .EN(n300), .Z(Y[46]) );
  TBUF_X1 \Y_tri[47]  ( .A(n255), .EN(n300), .Z(Y[47]) );
  TBUF_X1 \Y_tri[48]  ( .A(n256), .EN(n300), .Z(Y[48]) );
  TBUF_X1 \Y_tri[49]  ( .A(n257), .EN(n300), .Z(Y[49]) );
  TBUF_X1 \Y_tri[50]  ( .A(n258), .EN(n300), .Z(Y[50]) );
  TBUF_X1 \Y_tri[51]  ( .A(n259), .EN(n300), .Z(Y[51]) );
  TBUF_X1 \Y_tri[52]  ( .A(n260), .EN(n300), .Z(Y[52]) );
  TBUF_X1 \Y_tri[53]  ( .A(n261), .EN(n300), .Z(Y[53]) );
  TBUF_X1 \Y_tri[54]  ( .A(n262), .EN(n300), .Z(Y[54]) );
  TBUF_X1 \Y_tri[20]  ( .A(n228), .EN(n297), .Z(Y[20]) );
  TBUF_X1 \Y_tri[21]  ( .A(n229), .EN(n297), .Z(Y[21]) );
  TBUF_X1 \Y_tri[22]  ( .A(n230), .EN(n298), .Z(Y[22]) );
  TBUF_X1 \Y_tri[23]  ( .A(n231), .EN(n298), .Z(Y[23]) );
  TBUF_X1 \Y_tri[24]  ( .A(n232), .EN(n298), .Z(Y[24]) );
  TBUF_X1 \Y_tri[25]  ( .A(n233), .EN(n298), .Z(Y[25]) );
  TBUF_X1 \Y_tri[26]  ( .A(n234), .EN(n298), .Z(Y[26]) );
  TBUF_X1 \Y_tri[27]  ( .A(n235), .EN(n298), .Z(Y[27]) );
  TBUF_X1 \Y_tri[28]  ( .A(n236), .EN(n298), .Z(Y[28]) );
  TBUF_X1 \Y_tri[29]  ( .A(n237), .EN(n298), .Z(Y[29]) );
  TBUF_X1 \Y_tri[30]  ( .A(n238), .EN(n298), .Z(Y[30]) );
  TBUF_X1 \Y_tri[31]  ( .A(n239), .EN(n298), .Z(Y[31]) );
  TBUF_X1 \Y_tri[32]  ( .A(n240), .EN(n298), .Z(Y[32]) );
  TBUF_X1 \Y_tri[33]  ( .A(n241), .EN(n299), .Z(Y[33]) );
  TBUF_X1 \Y_tri[34]  ( .A(n242), .EN(n299), .Z(Y[34]) );
  TBUF_X1 \Y_tri[35]  ( .A(n243), .EN(n299), .Z(Y[35]) );
  TBUF_X1 \Y_tri[36]  ( .A(n244), .EN(n299), .Z(Y[36]) );
  TBUF_X1 \Y_tri[37]  ( .A(n245), .EN(n299), .Z(Y[37]) );
  TBUF_X1 \Y_tri[38]  ( .A(n246), .EN(n299), .Z(Y[38]) );
  TBUF_X1 \Y_tri[39]  ( .A(n247), .EN(n299), .Z(Y[39]) );
  TBUF_X1 \Y_tri[40]  ( .A(n248), .EN(n299), .Z(Y[40]) );
  TBUF_X1 \Y_tri[41]  ( .A(n249), .EN(n299), .Z(Y[41]) );
  TBUF_X1 \Y_tri[42]  ( .A(n250), .EN(n299), .Z(Y[42]) );
  TBUF_X1 \Y_tri[43]  ( .A(n251), .EN(n299), .Z(Y[43]) );
  TBUF_X1 \Y_tri[44]  ( .A(n252), .EN(n300), .Z(Y[44]) );
  TBUF_X1 \Y_tri[45]  ( .A(n253), .EN(n300), .Z(Y[45]) );
  TBUF_X1 \Y_tri[4]  ( .A(n211), .EN(n296), .Z(Y[4]) );
  TBUF_X1 \Y_tri[5]  ( .A(n212), .EN(n296), .Z(Y[5]) );
  TBUF_X1 \Y_tri[6]  ( .A(n213), .EN(n296), .Z(Y[6]) );
  TBUF_X1 \Y_tri[7]  ( .A(n214), .EN(n296), .Z(Y[7]) );
  TBUF_X1 \Y_tri[8]  ( .A(n215), .EN(n296), .Z(Y[8]) );
  TBUF_X1 \Y_tri[9]  ( .A(n217), .EN(n296), .Z(Y[9]) );
  TBUF_X1 \Y_tri[10]  ( .A(n218), .EN(n296), .Z(Y[10]) );
  TBUF_X1 \Y_tri[2]  ( .A(n209), .EN(n296), .Z(Y[2]) );
  TBUF_X1 \Y_tri[0]  ( .A(n207), .EN(n296), .Z(Y[0]) );
  TBUF_X1 \Y_tri[3]  ( .A(n210), .EN(n296), .Z(Y[3]) );
  TBUF_X1 \Y_tri[11]  ( .A(n219), .EN(n297), .Z(Y[11]) );
  TBUF_X1 \Y_tri[12]  ( .A(n220), .EN(n297), .Z(Y[12]) );
  TBUF_X1 \Y_tri[13]  ( .A(n221), .EN(n297), .Z(Y[13]) );
  TBUF_X1 \Y_tri[14]  ( .A(n222), .EN(n297), .Z(Y[14]) );
  TBUF_X1 \Y_tri[15]  ( .A(n223), .EN(n297), .Z(Y[15]) );
  TBUF_X1 \Y_tri[16]  ( .A(n224), .EN(n297), .Z(Y[16]) );
  TBUF_X1 \Y_tri[17]  ( .A(n225), .EN(n297), .Z(Y[17]) );
  TBUF_X1 \Y_tri[18]  ( .A(n226), .EN(n297), .Z(Y[18]) );
  TBUF_X1 \Y_tri[19]  ( .A(n227), .EN(n297), .Z(Y[19]) );
  NAND2_X1 U2 ( .A1(n48), .A2(n49), .ZN(n251) );
  AOI22_X1 U3 ( .A1(plusA[43]), .A2(n281), .B1(plus2A[43]), .B2(n275), .ZN(n48) );
  AOI22_X1 U4 ( .A1(minus2A[43]), .A2(n293), .B1(minusA[43]), .B2(n287), .ZN(
        n49) );
  NAND2_X1 U5 ( .A1(n58), .A2(n59), .ZN(n246) );
  AOI22_X1 U6 ( .A1(plusA[38]), .A2(n281), .B1(plus2A[38]), .B2(n275), .ZN(n58) );
  AOI22_X1 U7 ( .A1(minus2A[38]), .A2(n293), .B1(minusA[38]), .B2(n287), .ZN(
        n59) );
  NAND2_X1 U8 ( .A1(n28), .A2(n29), .ZN(n261) );
  AOI22_X1 U9 ( .A1(plusA[53]), .A2(n282), .B1(plus2A[53]), .B2(n276), .ZN(n28) );
  AOI22_X1 U10 ( .A1(minus2A[53]), .A2(n294), .B1(minusA[53]), .B2(n288), .ZN(
        n29) );
  NAND2_X1 U11 ( .A1(n38), .A2(n39), .ZN(n256) );
  AOI22_X1 U12 ( .A1(plusA[48]), .A2(n282), .B1(plus2A[48]), .B2(n276), .ZN(
        n38) );
  AOI22_X1 U13 ( .A1(minus2A[48]), .A2(n294), .B1(minusA[48]), .B2(n288), .ZN(
        n39) );
  NAND2_X1 U14 ( .A1(n18), .A2(n19), .ZN(n266) );
  AOI22_X1 U15 ( .A1(plusA[58]), .A2(n282), .B1(plus2A[58]), .B2(n276), .ZN(
        n18) );
  AOI22_X1 U16 ( .A1(minus2A[58]), .A2(n294), .B1(minusA[58]), .B2(n288), .ZN(
        n19) );
  BUF_X1 U17 ( .A(n8), .Z(n278) );
  BUF_X1 U18 ( .A(n8), .Z(n279) );
  BUF_X1 U19 ( .A(n6), .Z(n291) );
  BUF_X1 U20 ( .A(n7), .Z(n285) );
  BUF_X1 U21 ( .A(n9), .Z(n272) );
  BUF_X1 U22 ( .A(n9), .Z(n273) );
  BUF_X1 U23 ( .A(n7), .Z(n284) );
  BUF_X1 U24 ( .A(n216), .Z(n297) );
  BUF_X1 U25 ( .A(n216), .Z(n296) );
  BUF_X1 U26 ( .A(n6), .Z(n290) );
  NAND2_X1 U27 ( .A1(n70), .A2(n71), .ZN(n240) );
  AOI22_X1 U28 ( .A1(plusA[32]), .A2(n280), .B1(plus2A[32]), .B2(n274), .ZN(
        n70) );
  AOI22_X1 U29 ( .A1(minus2A[32]), .A2(n292), .B1(minusA[32]), .B2(n286), .ZN(
        n71) );
  NAND2_X1 U30 ( .A1(n50), .A2(n51), .ZN(n250) );
  AOI22_X1 U31 ( .A1(plusA[42]), .A2(n281), .B1(plus2A[42]), .B2(n275), .ZN(
        n50) );
  AOI22_X1 U32 ( .A1(minus2A[42]), .A2(n293), .B1(minusA[42]), .B2(n287), .ZN(
        n51) );
  NAND2_X1 U33 ( .A1(n60), .A2(n61), .ZN(n245) );
  AOI22_X1 U34 ( .A1(plusA[37]), .A2(n281), .B1(plus2A[37]), .B2(n275), .ZN(
        n60) );
  AOI22_X1 U35 ( .A1(minus2A[37]), .A2(n293), .B1(minusA[37]), .B2(n287), .ZN(
        n61) );
  NAND2_X1 U36 ( .A1(n52), .A2(n53), .ZN(n249) );
  AOI22_X1 U37 ( .A1(plusA[41]), .A2(n281), .B1(plus2A[41]), .B2(n275), .ZN(
        n52) );
  AOI22_X1 U38 ( .A1(minus2A[41]), .A2(n293), .B1(minusA[41]), .B2(n287), .ZN(
        n53) );
  NAND2_X1 U39 ( .A1(n62), .A2(n63), .ZN(n244) );
  AOI22_X1 U40 ( .A1(plusA[36]), .A2(n281), .B1(plus2A[36]), .B2(n275), .ZN(
        n62) );
  AOI22_X1 U41 ( .A1(minus2A[36]), .A2(n293), .B1(minusA[36]), .B2(n287), .ZN(
        n63) );
  NAND2_X1 U42 ( .A1(n44), .A2(n45), .ZN(n253) );
  AOI22_X1 U43 ( .A1(plusA[45]), .A2(n281), .B1(plus2A[45]), .B2(n275), .ZN(
        n44) );
  AOI22_X1 U44 ( .A1(minus2A[45]), .A2(n293), .B1(minusA[45]), .B2(n287), .ZN(
        n45) );
  NAND2_X1 U45 ( .A1(n54), .A2(n55), .ZN(n248) );
  AOI22_X1 U46 ( .A1(plusA[40]), .A2(n281), .B1(plus2A[40]), .B2(n275), .ZN(
        n54) );
  AOI22_X1 U47 ( .A1(minus2A[40]), .A2(n293), .B1(minusA[40]), .B2(n287), .ZN(
        n55) );
  NAND2_X1 U48 ( .A1(n64), .A2(n65), .ZN(n243) );
  AOI22_X1 U49 ( .A1(plusA[35]), .A2(n280), .B1(plus2A[35]), .B2(n274), .ZN(
        n64) );
  AOI22_X1 U50 ( .A1(minus2A[35]), .A2(n292), .B1(minusA[35]), .B2(n286), .ZN(
        n65) );
  NAND2_X1 U51 ( .A1(n46), .A2(n47), .ZN(n252) );
  AOI22_X1 U52 ( .A1(plusA[44]), .A2(n281), .B1(plus2A[44]), .B2(n275), .ZN(
        n46) );
  AOI22_X1 U53 ( .A1(minus2A[44]), .A2(n293), .B1(minusA[44]), .B2(n287), .ZN(
        n47) );
  NAND2_X1 U54 ( .A1(n56), .A2(n57), .ZN(n247) );
  AOI22_X1 U55 ( .A1(plusA[39]), .A2(n281), .B1(plus2A[39]), .B2(n275), .ZN(
        n56) );
  AOI22_X1 U56 ( .A1(minus2A[39]), .A2(n293), .B1(minusA[39]), .B2(n287), .ZN(
        n57) );
  NAND2_X1 U57 ( .A1(n66), .A2(n67), .ZN(n242) );
  AOI22_X1 U58 ( .A1(plusA[34]), .A2(n280), .B1(plus2A[34]), .B2(n274), .ZN(
        n66) );
  AOI22_X1 U59 ( .A1(minus2A[34]), .A2(n292), .B1(minusA[34]), .B2(n286), .ZN(
        n67) );
  NAND2_X1 U60 ( .A1(n68), .A2(n69), .ZN(n241) );
  AOI22_X1 U61 ( .A1(plusA[33]), .A2(n280), .B1(plus2A[33]), .B2(n274), .ZN(
        n68) );
  AOI22_X1 U62 ( .A1(minus2A[33]), .A2(n292), .B1(minusA[33]), .B2(n286), .ZN(
        n69) );
  BUF_X1 U63 ( .A(n8), .Z(n280) );
  BUF_X1 U64 ( .A(n6), .Z(n292) );
  BUF_X1 U65 ( .A(n7), .Z(n286) );
  BUF_X1 U66 ( .A(n9), .Z(n274) );
  BUF_X1 U67 ( .A(n216), .Z(n298) );
  NAND2_X1 U68 ( .A1(n4), .A2(n5), .ZN(n271) );
  AOI22_X1 U69 ( .A1(plusA[63]), .A2(n283), .B1(plus2A[63]), .B2(n277), .ZN(n4) );
  AOI22_X1 U70 ( .A1(minus2A[63]), .A2(n295), .B1(minusA[63]), .B2(n289), .ZN(
        n5) );
  NAND2_X1 U71 ( .A1(n20), .A2(n21), .ZN(n265) );
  AOI22_X1 U72 ( .A1(plusA[57]), .A2(n282), .B1(plus2A[57]), .B2(n276), .ZN(
        n20) );
  AOI22_X1 U73 ( .A1(minus2A[57]), .A2(n294), .B1(minusA[57]), .B2(n288), .ZN(
        n21) );
  NAND2_X1 U74 ( .A1(n40), .A2(n41), .ZN(n255) );
  AOI22_X1 U75 ( .A1(plusA[47]), .A2(n281), .B1(plus2A[47]), .B2(n275), .ZN(
        n40) );
  AOI22_X1 U76 ( .A1(minus2A[47]), .A2(n293), .B1(minusA[47]), .B2(n287), .ZN(
        n41) );
  NAND2_X1 U77 ( .A1(n12), .A2(n13), .ZN(n269) );
  AOI22_X1 U78 ( .A1(plusA[61]), .A2(n283), .B1(plus2A[61]), .B2(n277), .ZN(
        n12) );
  AOI22_X1 U79 ( .A1(minus2A[61]), .A2(n295), .B1(minusA[61]), .B2(n289), .ZN(
        n13) );
  NAND2_X1 U80 ( .A1(n30), .A2(n31), .ZN(n260) );
  AOI22_X1 U81 ( .A1(plusA[52]), .A2(n282), .B1(plus2A[52]), .B2(n276), .ZN(
        n30) );
  AOI22_X1 U82 ( .A1(minus2A[52]), .A2(n294), .B1(minusA[52]), .B2(n288), .ZN(
        n31) );
  NAND2_X1 U83 ( .A1(n32), .A2(n33), .ZN(n259) );
  AOI22_X1 U84 ( .A1(plusA[51]), .A2(n282), .B1(plus2A[51]), .B2(n276), .ZN(
        n32) );
  AOI22_X1 U85 ( .A1(minus2A[51]), .A2(n294), .B1(minusA[51]), .B2(n288), .ZN(
        n33) );
  NAND2_X1 U86 ( .A1(n10), .A2(n11), .ZN(n270) );
  AOI22_X1 U87 ( .A1(plusA[62]), .A2(n283), .B1(plus2A[62]), .B2(n277), .ZN(
        n10) );
  AOI22_X1 U88 ( .A1(minus2A[62]), .A2(n295), .B1(minusA[62]), .B2(n289), .ZN(
        n11) );
  NAND2_X1 U89 ( .A1(n34), .A2(n35), .ZN(n258) );
  AOI22_X1 U90 ( .A1(plusA[50]), .A2(n282), .B1(plus2A[50]), .B2(n276), .ZN(
        n34) );
  AOI22_X1 U91 ( .A1(minus2A[50]), .A2(n294), .B1(minusA[50]), .B2(n288), .ZN(
        n35) );
  NAND2_X1 U92 ( .A1(n42), .A2(n43), .ZN(n254) );
  AOI22_X1 U93 ( .A1(plusA[46]), .A2(n281), .B1(plus2A[46]), .B2(n275), .ZN(
        n42) );
  AOI22_X1 U94 ( .A1(minus2A[46]), .A2(n293), .B1(minusA[46]), .B2(n287), .ZN(
        n43) );
  NAND2_X1 U95 ( .A1(n22), .A2(n23), .ZN(n264) );
  AOI22_X1 U96 ( .A1(plusA[56]), .A2(n282), .B1(plus2A[56]), .B2(n276), .ZN(
        n22) );
  AOI22_X1 U97 ( .A1(minus2A[56]), .A2(n294), .B1(minusA[56]), .B2(n288), .ZN(
        n23) );
  NAND2_X1 U98 ( .A1(n14), .A2(n15), .ZN(n268) );
  AOI22_X1 U99 ( .A1(plusA[60]), .A2(n283), .B1(plus2A[60]), .B2(n277), .ZN(
        n14) );
  AOI22_X1 U100 ( .A1(minus2A[60]), .A2(n295), .B1(minusA[60]), .B2(n289), 
        .ZN(n15) );
  NAND2_X1 U101 ( .A1(n24), .A2(n25), .ZN(n263) );
  AOI22_X1 U102 ( .A1(plusA[55]), .A2(n282), .B1(plus2A[55]), .B2(n276), .ZN(
        n24) );
  AOI22_X1 U103 ( .A1(minus2A[55]), .A2(n294), .B1(minusA[55]), .B2(n288), 
        .ZN(n25) );
  NAND2_X1 U104 ( .A1(n36), .A2(n37), .ZN(n257) );
  AOI22_X1 U105 ( .A1(plusA[49]), .A2(n282), .B1(plus2A[49]), .B2(n276), .ZN(
        n36) );
  AOI22_X1 U106 ( .A1(minus2A[49]), .A2(n294), .B1(minusA[49]), .B2(n288), 
        .ZN(n37) );
  NAND2_X1 U107 ( .A1(n16), .A2(n17), .ZN(n267) );
  AOI22_X1 U108 ( .A1(plusA[59]), .A2(n282), .B1(plus2A[59]), .B2(n276), .ZN(
        n16) );
  AOI22_X1 U109 ( .A1(minus2A[59]), .A2(n294), .B1(minusA[59]), .B2(n288), 
        .ZN(n17) );
  NAND2_X1 U110 ( .A1(n26), .A2(n27), .ZN(n262) );
  AOI22_X1 U111 ( .A1(plusA[54]), .A2(n282), .B1(plus2A[54]), .B2(n276), .ZN(
        n26) );
  AOI22_X1 U112 ( .A1(minus2A[54]), .A2(n294), .B1(minusA[54]), .B2(n288), 
        .ZN(n27) );
  BUF_X1 U113 ( .A(n8), .Z(n281) );
  BUF_X1 U114 ( .A(n6), .Z(n293) );
  BUF_X1 U115 ( .A(n7), .Z(n287) );
  BUF_X1 U116 ( .A(n9), .Z(n275) );
  BUF_X1 U117 ( .A(n216), .Z(n299) );
  BUF_X1 U118 ( .A(n8), .Z(n282) );
  BUF_X1 U119 ( .A(n6), .Z(n294) );
  BUF_X1 U120 ( .A(n7), .Z(n288) );
  BUF_X1 U121 ( .A(n9), .Z(n276) );
  BUF_X1 U122 ( .A(n216), .Z(n300) );
  BUF_X1 U123 ( .A(n216), .Z(n301) );
  NOR3_X1 U124 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n302), .ZN(n7) );
  NOR3_X1 U125 ( .A1(n302), .A2(SEL[2]), .A3(n303), .ZN(n9) );
  NOR3_X1 U126 ( .A1(SEL[1]), .A2(SEL[2]), .A3(n303), .ZN(n8) );
  NOR2_X1 U127 ( .A1(n118), .A2(n304), .ZN(n216) );
  INV_X1 U128 ( .A(SEL[2]), .ZN(n304) );
  AND2_X1 U129 ( .A1(SEL[2]), .A2(n118), .ZN(n6) );
  INV_X1 U130 ( .A(SEL[1]), .ZN(n302) );
  NAND2_X1 U131 ( .A1(n72), .A2(n73), .ZN(n239) );
  AOI22_X1 U132 ( .A1(plusA[31]), .A2(n280), .B1(plus2A[31]), .B2(n274), .ZN(
        n72) );
  AOI22_X1 U133 ( .A1(minus2A[31]), .A2(n292), .B1(minusA[31]), .B2(n286), 
        .ZN(n73) );
  NAND2_X1 U134 ( .A1(n96), .A2(n97), .ZN(n227) );
  AOI22_X1 U135 ( .A1(plusA[19]), .A2(n279), .B1(plus2A[19]), .B2(n273), .ZN(
        n96) );
  AOI22_X1 U136 ( .A1(minus2A[19]), .A2(n291), .B1(minusA[19]), .B2(n285), 
        .ZN(n97) );
  NAND2_X1 U137 ( .A1(n98), .A2(n99), .ZN(n226) );
  AOI22_X1 U138 ( .A1(plusA[18]), .A2(n279), .B1(plus2A[18]), .B2(n273), .ZN(
        n98) );
  AOI22_X1 U139 ( .A1(minus2A[18]), .A2(n291), .B1(minusA[18]), .B2(n285), 
        .ZN(n99) );
  NAND2_X1 U140 ( .A1(n100), .A2(n101), .ZN(n225) );
  AOI22_X1 U141 ( .A1(plusA[17]), .A2(n279), .B1(plus2A[17]), .B2(n273), .ZN(
        n100) );
  AOI22_X1 U142 ( .A1(minus2A[17]), .A2(n291), .B1(minusA[17]), .B2(n285), 
        .ZN(n101) );
  NAND2_X1 U143 ( .A1(n102), .A2(n103), .ZN(n224) );
  AOI22_X1 U144 ( .A1(plusA[16]), .A2(n279), .B1(plus2A[16]), .B2(n273), .ZN(
        n102) );
  AOI22_X1 U145 ( .A1(minus2A[16]), .A2(n291), .B1(minusA[16]), .B2(n285), 
        .ZN(n103) );
  NAND2_X1 U146 ( .A1(n135), .A2(n136), .ZN(n207) );
  AOI22_X1 U147 ( .A1(plusA[0]), .A2(n278), .B1(plus2A[0]), .B2(n272), .ZN(
        n135) );
  AOI22_X1 U148 ( .A1(plusA[1]), .A2(n278), .B1(plus2A[1]), .B2(n272), .ZN(
        n133) );
  NAND2_X1 U149 ( .A1(n129), .A2(n130), .ZN(n210) );
  AOI22_X1 U150 ( .A1(plusA[3]), .A2(n278), .B1(plus2A[3]), .B2(n272), .ZN(
        n129) );
  NAND2_X1 U151 ( .A1(n110), .A2(n111), .ZN(n220) );
  AOI22_X1 U152 ( .A1(plusA[12]), .A2(n279), .B1(plus2A[12]), .B2(n273), .ZN(
        n110) );
  AOI22_X1 U153 ( .A1(minus2A[12]), .A2(n291), .B1(minusA[12]), .B2(n285), 
        .ZN(n111) );
  NAND2_X1 U154 ( .A1(n119), .A2(n120), .ZN(n215) );
  AOI22_X1 U155 ( .A1(plusA[8]), .A2(n278), .B1(plus2A[8]), .B2(n272), .ZN(
        n119) );
  NAND2_X1 U156 ( .A1(n127), .A2(n128), .ZN(n211) );
  AOI22_X1 U157 ( .A1(plusA[4]), .A2(n278), .B1(plus2A[4]), .B2(n272), .ZN(
        n127) );
  NAND2_X1 U158 ( .A1(n131), .A2(n132), .ZN(n209) );
  AOI22_X1 U159 ( .A1(plusA[2]), .A2(n278), .B1(plus2A[2]), .B2(n272), .ZN(
        n131) );
  NAND2_X1 U160 ( .A1(n104), .A2(n105), .ZN(n223) );
  AOI22_X1 U161 ( .A1(plusA[15]), .A2(n279), .B1(plus2A[15]), .B2(n273), .ZN(
        n104) );
  AOI22_X1 U162 ( .A1(minus2A[15]), .A2(n291), .B1(minusA[15]), .B2(n285), 
        .ZN(n105) );
  NAND2_X1 U163 ( .A1(n121), .A2(n122), .ZN(n214) );
  AOI22_X1 U164 ( .A1(plusA[7]), .A2(n278), .B1(plus2A[7]), .B2(n272), .ZN(
        n121) );
  NAND2_X1 U165 ( .A1(n112), .A2(n113), .ZN(n219) );
  AOI22_X1 U166 ( .A1(plusA[11]), .A2(n278), .B1(plus2A[11]), .B2(n272), .ZN(
        n112) );
  NAND2_X1 U167 ( .A1(n116), .A2(n117), .ZN(n217) );
  AOI22_X1 U168 ( .A1(plusA[9]), .A2(n278), .B1(plus2A[9]), .B2(n272), .ZN(
        n116) );
  NAND2_X1 U169 ( .A1(n108), .A2(n109), .ZN(n221) );
  AOI22_X1 U170 ( .A1(plusA[13]), .A2(n279), .B1(plus2A[13]), .B2(n273), .ZN(
        n108) );
  AOI22_X1 U171 ( .A1(minus2A[13]), .A2(n291), .B1(minusA[13]), .B2(n285), 
        .ZN(n109) );
  NAND2_X1 U172 ( .A1(n125), .A2(n126), .ZN(n212) );
  AOI22_X1 U173 ( .A1(plusA[5]), .A2(n278), .B1(plus2A[5]), .B2(n272), .ZN(
        n125) );
  NAND2_X1 U174 ( .A1(n106), .A2(n107), .ZN(n222) );
  AOI22_X1 U175 ( .A1(plusA[14]), .A2(n279), .B1(plus2A[14]), .B2(n273), .ZN(
        n106) );
  AOI22_X1 U176 ( .A1(minus2A[14]), .A2(n291), .B1(minusA[14]), .B2(n285), 
        .ZN(n107) );
  NAND2_X1 U177 ( .A1(n114), .A2(n115), .ZN(n218) );
  AOI22_X1 U178 ( .A1(plusA[10]), .A2(n278), .B1(plus2A[10]), .B2(n272), .ZN(
        n114) );
  NAND2_X1 U179 ( .A1(n123), .A2(n124), .ZN(n213) );
  AOI22_X1 U180 ( .A1(plusA[6]), .A2(n278), .B1(plus2A[6]), .B2(n272), .ZN(
        n123) );
  NAND2_X1 U181 ( .A1(n74), .A2(n75), .ZN(n238) );
  AOI22_X1 U182 ( .A1(plusA[30]), .A2(n280), .B1(plus2A[30]), .B2(n274), .ZN(
        n74) );
  AOI22_X1 U183 ( .A1(minus2A[30]), .A2(n292), .B1(minusA[30]), .B2(n286), 
        .ZN(n75) );
  NAND2_X1 U184 ( .A1(n76), .A2(n77), .ZN(n237) );
  AOI22_X1 U185 ( .A1(plusA[29]), .A2(n280), .B1(plus2A[29]), .B2(n274), .ZN(
        n76) );
  AOI22_X1 U186 ( .A1(minus2A[29]), .A2(n292), .B1(minusA[29]), .B2(n286), 
        .ZN(n77) );
  NAND2_X1 U187 ( .A1(n78), .A2(n79), .ZN(n236) );
  AOI22_X1 U188 ( .A1(plusA[28]), .A2(n280), .B1(plus2A[28]), .B2(n274), .ZN(
        n78) );
  AOI22_X1 U189 ( .A1(minus2A[28]), .A2(n292), .B1(minusA[28]), .B2(n286), 
        .ZN(n79) );
  NAND2_X1 U190 ( .A1(n80), .A2(n81), .ZN(n235) );
  AOI22_X1 U191 ( .A1(plusA[27]), .A2(n280), .B1(plus2A[27]), .B2(n274), .ZN(
        n80) );
  AOI22_X1 U192 ( .A1(minus2A[27]), .A2(n292), .B1(minusA[27]), .B2(n286), 
        .ZN(n81) );
  NAND2_X1 U193 ( .A1(n82), .A2(n83), .ZN(n234) );
  AOI22_X1 U194 ( .A1(plusA[26]), .A2(n280), .B1(plus2A[26]), .B2(n274), .ZN(
        n82) );
  AOI22_X1 U195 ( .A1(minus2A[26]), .A2(n292), .B1(minusA[26]), .B2(n286), 
        .ZN(n83) );
  NAND2_X1 U196 ( .A1(n84), .A2(n85), .ZN(n233) );
  AOI22_X1 U197 ( .A1(plusA[25]), .A2(n280), .B1(plus2A[25]), .B2(n274), .ZN(
        n84) );
  AOI22_X1 U198 ( .A1(minus2A[25]), .A2(n292), .B1(minusA[25]), .B2(n286), 
        .ZN(n85) );
  NAND2_X1 U199 ( .A1(n86), .A2(n87), .ZN(n232) );
  AOI22_X1 U200 ( .A1(plusA[24]), .A2(n280), .B1(plus2A[24]), .B2(n274), .ZN(
        n86) );
  AOI22_X1 U201 ( .A1(minus2A[24]), .A2(n292), .B1(minusA[24]), .B2(n286), 
        .ZN(n87) );
  NAND2_X1 U202 ( .A1(n88), .A2(n89), .ZN(n231) );
  AOI22_X1 U203 ( .A1(plusA[23]), .A2(n279), .B1(plus2A[23]), .B2(n273), .ZN(
        n88) );
  AOI22_X1 U204 ( .A1(minus2A[23]), .A2(n291), .B1(minusA[23]), .B2(n285), 
        .ZN(n89) );
  NAND2_X1 U205 ( .A1(n90), .A2(n91), .ZN(n230) );
  AOI22_X1 U206 ( .A1(plusA[22]), .A2(n279), .B1(plus2A[22]), .B2(n273), .ZN(
        n90) );
  AOI22_X1 U207 ( .A1(minus2A[22]), .A2(n291), .B1(minusA[22]), .B2(n285), 
        .ZN(n91) );
  NAND2_X1 U208 ( .A1(n92), .A2(n93), .ZN(n229) );
  AOI22_X1 U209 ( .A1(plusA[21]), .A2(n279), .B1(plus2A[21]), .B2(n273), .ZN(
        n92) );
  AOI22_X1 U210 ( .A1(minus2A[21]), .A2(n291), .B1(minusA[21]), .B2(n285), 
        .ZN(n93) );
  NAND2_X1 U211 ( .A1(n94), .A2(n95), .ZN(n228) );
  AOI22_X1 U212 ( .A1(plusA[20]), .A2(n279), .B1(plus2A[20]), .B2(n273), .ZN(
        n94) );
  AOI22_X1 U213 ( .A1(minus2A[20]), .A2(n291), .B1(minusA[20]), .B2(n285), 
        .ZN(n95) );
  NAND2_X1 U214 ( .A1(n133), .A2(n134), .ZN(n208) );
  NOR2_X1 U215 ( .A1(SEL[1]), .A2(SEL[0]), .ZN(n118) );
  INV_X1 U216 ( .A(SEL[0]), .ZN(n303) );
  AOI22_X1 U217 ( .A1(minus2A[11]), .A2(n290), .B1(minusA[11]), .B2(n284), 
        .ZN(n113) );
  AOI22_X1 U218 ( .A1(minus2A[10]), .A2(n290), .B1(minusA[10]), .B2(n284), 
        .ZN(n115) );
  AOI22_X1 U219 ( .A1(minus2A[9]), .A2(n290), .B1(minusA[9]), .B2(n284), .ZN(
        n117) );
  AOI22_X1 U220 ( .A1(minus2A[8]), .A2(n290), .B1(minusA[8]), .B2(n284), .ZN(
        n120) );
  AOI22_X1 U221 ( .A1(minus2A[7]), .A2(n290), .B1(minusA[7]), .B2(n284), .ZN(
        n122) );
  AOI22_X1 U222 ( .A1(minus2A[6]), .A2(n290), .B1(minusA[6]), .B2(n284), .ZN(
        n124) );
  AOI22_X1 U223 ( .A1(minus2A[5]), .A2(n290), .B1(minusA[5]), .B2(n284), .ZN(
        n126) );
  AOI22_X1 U224 ( .A1(minus2A[4]), .A2(n290), .B1(minusA[4]), .B2(n284), .ZN(
        n128) );
  AOI22_X1 U225 ( .A1(minus2A[3]), .A2(n290), .B1(minusA[3]), .B2(n284), .ZN(
        n130) );
  AOI22_X1 U226 ( .A1(minus2A[2]), .A2(n290), .B1(minusA[2]), .B2(n284), .ZN(
        n132) );
  AOI22_X1 U227 ( .A1(minus2A[1]), .A2(n290), .B1(minusA[1]), .B2(n284), .ZN(
        n134) );
  AOI22_X1 U228 ( .A1(minus2A[0]), .A2(n290), .B1(minusA[0]), .B2(n284), .ZN(
        n136) );
  CLKBUF_X1 U229 ( .A(n9), .Z(n277) );
  CLKBUF_X1 U230 ( .A(n8), .Z(n283) );
  CLKBUF_X1 U231 ( .A(n7), .Z(n289) );
  CLKBUF_X1 U232 ( .A(n6), .Z(n295) );
endmodule


module booth_mul_row_special_N64_RADIX3 ( A, encoderIn, nextA, nextSum );
  input [63:0] A;
  input [2:0] encoderIn;
  output [63:0] nextA;
  output [63:0] nextSum;
  wire   n4, n5;
  wire   [2:0] encoder_to_mux;
  wire   [63:0] plusA_s;
  wire   [63:0] minusA_s;
  wire   [63:0] minus2A_s;
  tri   [63:0] nextSum;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign nextA[51] = n4;
  assign nextA[39] = n5;
  assign nextA[0] = 1'b0;

  encoder_N64_RADIX3_0 encoder_1 ( .X(encoderIn), .Z(encoder_to_mux) );
  ShiftnCompl_special_N64 ShiftnCompl_special_1 ( .plusA(A), .plusA_out(
        plusA_s), .minusA_out(minusA_s), .plus2A_out({nextA[63:52], n4, 
        nextA[50:40], n5, nextA[38:1], SYNOPSYS_UNCONNECTED__0}), 
        .minus2A_out(minus2A_s) );
  MUX_GENERIC_N64_RADIX3_0 mux_1 ( .plusA(plusA_s), .minusA(minusA_s), 
        .plus2A({nextA[63:52], n4, nextA[50:40], n5, nextA[38:1], 1'b0}), 
        .minus2A(minus2A_s), .SEL(encoder_to_mux), .Y(nextSum) );
endmodule


module encoder_N64_RADIX3_15 ( X, Z );
  input [2:0] X;
  output [2:0] Z;
  wire   n5, n7, n8;

  INV_X1 U1 ( .A(X[2]), .ZN(n5) );
  OAI22_X1 U2 ( .A1(n8), .A2(n5), .B1(X[2]), .B2(n7), .ZN(Z[1]) );
  AOI21_X1 U3 ( .B1(n8), .B2(n7), .A(X[2]), .ZN(Z[0]) );
  AND3_X1 U4 ( .A1(X[2]), .A2(n7), .A3(n8), .ZN(Z[2]) );
  OAI21_X1 U5 ( .B1(X[1]), .B2(X[0]), .A(n7), .ZN(n8) );
  NAND2_X1 U6 ( .A1(X[1]), .A2(X[0]), .ZN(n7) );
endmodule


module shifter_N64_30 ( \input , shiftLeftOnePos );
  input [63:0] \input ;
  output [63:0] shiftLeftOnePos;
  wire   \input[62] , \input[61] , \input[60] , \input[59] , \input[58] ,
         \input[57] , \input[56] , \input[55] , \input[54] , \input[53] ,
         \input[52] , \input[51] , \input[50] , \input[49] , \input[48] ,
         \input[47] , \input[46] , \input[45] , \input[44] , \input[43] ,
         \input[42] , \input[41] , \input[40] , \input[39] , \input[38] ,
         \input[37] , \input[36] , \input[35] , \input[34] , \input[33] ,
         \input[32] , \input[31] , \input[30] , \input[29] , \input[28] ,
         \input[27] , \input[26] , \input[25] , \input[24] , \input[23] ,
         \input[22] , \input[21] , \input[20] , \input[19] , \input[18] ,
         \input[17] , \input[16] , \input[15] , \input[14] , \input[13] ,
         \input[12] , \input[11] , \input[10] , \input[9] , \input[8] ,
         \input[7] , \input[6] , \input[5] , \input[4] , \input[3] ,
         \input[2] , \input[1] , \input[0] ;
  assign shiftLeftOnePos[0] = 1'b0;
  assign shiftLeftOnePos[63] = \input[62] ;
  assign \input[62]  = \input  [62];
  assign shiftLeftOnePos[62] = \input[61] ;
  assign \input[61]  = \input  [61];
  assign shiftLeftOnePos[61] = \input[60] ;
  assign \input[60]  = \input  [60];
  assign shiftLeftOnePos[60] = \input[59] ;
  assign \input[59]  = \input  [59];
  assign shiftLeftOnePos[59] = \input[58] ;
  assign \input[58]  = \input  [58];
  assign shiftLeftOnePos[58] = \input[57] ;
  assign \input[57]  = \input  [57];
  assign shiftLeftOnePos[57] = \input[56] ;
  assign \input[56]  = \input  [56];
  assign shiftLeftOnePos[56] = \input[55] ;
  assign \input[55]  = \input  [55];
  assign shiftLeftOnePos[55] = \input[54] ;
  assign \input[54]  = \input  [54];
  assign shiftLeftOnePos[54] = \input[53] ;
  assign \input[53]  = \input  [53];
  assign shiftLeftOnePos[53] = \input[52] ;
  assign \input[52]  = \input  [52];
  assign shiftLeftOnePos[52] = \input[51] ;
  assign \input[51]  = \input  [51];
  assign shiftLeftOnePos[51] = \input[50] ;
  assign \input[50]  = \input  [50];
  assign shiftLeftOnePos[50] = \input[49] ;
  assign \input[49]  = \input  [49];
  assign shiftLeftOnePos[49] = \input[48] ;
  assign \input[48]  = \input  [48];
  assign shiftLeftOnePos[48] = \input[47] ;
  assign \input[47]  = \input  [47];
  assign shiftLeftOnePos[47] = \input[46] ;
  assign \input[46]  = \input  [46];
  assign shiftLeftOnePos[46] = \input[45] ;
  assign \input[45]  = \input  [45];
  assign shiftLeftOnePos[45] = \input[44] ;
  assign \input[44]  = \input  [44];
  assign shiftLeftOnePos[44] = \input[43] ;
  assign \input[43]  = \input  [43];
  assign shiftLeftOnePos[43] = \input[42] ;
  assign \input[42]  = \input  [42];
  assign shiftLeftOnePos[42] = \input[41] ;
  assign \input[41]  = \input  [41];
  assign shiftLeftOnePos[41] = \input[40] ;
  assign \input[40]  = \input  [40];
  assign shiftLeftOnePos[40] = \input[39] ;
  assign \input[39]  = \input  [39];
  assign shiftLeftOnePos[39] = \input[38] ;
  assign \input[38]  = \input  [38];
  assign shiftLeftOnePos[38] = \input[37] ;
  assign \input[37]  = \input  [37];
  assign shiftLeftOnePos[37] = \input[36] ;
  assign \input[36]  = \input  [36];
  assign shiftLeftOnePos[36] = \input[35] ;
  assign \input[35]  = \input  [35];
  assign shiftLeftOnePos[35] = \input[34] ;
  assign \input[34]  = \input  [34];
  assign shiftLeftOnePos[34] = \input[33] ;
  assign \input[33]  = \input  [33];
  assign shiftLeftOnePos[33] = \input[32] ;
  assign \input[32]  = \input  [32];
  assign shiftLeftOnePos[32] = \input[31] ;
  assign \input[31]  = \input  [31];
  assign shiftLeftOnePos[31] = \input[30] ;
  assign \input[30]  = \input  [30];
  assign shiftLeftOnePos[30] = \input[29] ;
  assign \input[29]  = \input  [29];
  assign shiftLeftOnePos[29] = \input[28] ;
  assign \input[28]  = \input  [28];
  assign shiftLeftOnePos[28] = \input[27] ;
  assign \input[27]  = \input  [27];
  assign shiftLeftOnePos[27] = \input[26] ;
  assign \input[26]  = \input  [26];
  assign shiftLeftOnePos[26] = \input[25] ;
  assign \input[25]  = \input  [25];
  assign shiftLeftOnePos[25] = \input[24] ;
  assign \input[24]  = \input  [24];
  assign shiftLeftOnePos[24] = \input[23] ;
  assign \input[23]  = \input  [23];
  assign shiftLeftOnePos[23] = \input[22] ;
  assign \input[22]  = \input  [22];
  assign shiftLeftOnePos[22] = \input[21] ;
  assign \input[21]  = \input  [21];
  assign shiftLeftOnePos[21] = \input[20] ;
  assign \input[20]  = \input  [20];
  assign shiftLeftOnePos[20] = \input[19] ;
  assign \input[19]  = \input  [19];
  assign shiftLeftOnePos[19] = \input[18] ;
  assign \input[18]  = \input  [18];
  assign shiftLeftOnePos[18] = \input[17] ;
  assign \input[17]  = \input  [17];
  assign shiftLeftOnePos[17] = \input[16] ;
  assign \input[16]  = \input  [16];
  assign shiftLeftOnePos[16] = \input[15] ;
  assign \input[15]  = \input  [15];
  assign shiftLeftOnePos[15] = \input[14] ;
  assign \input[14]  = \input  [14];
  assign shiftLeftOnePos[14] = \input[13] ;
  assign \input[13]  = \input  [13];
  assign shiftLeftOnePos[13] = \input[12] ;
  assign \input[12]  = \input  [12];
  assign shiftLeftOnePos[12] = \input[11] ;
  assign \input[11]  = \input  [11];
  assign shiftLeftOnePos[11] = \input[10] ;
  assign \input[10]  = \input  [10];
  assign shiftLeftOnePos[10] = \input[9] ;
  assign \input[9]  = \input  [9];
  assign shiftLeftOnePos[9] = \input[8] ;
  assign \input[8]  = \input  [8];
  assign shiftLeftOnePos[8] = \input[7] ;
  assign \input[7]  = \input  [7];
  assign shiftLeftOnePos[7] = \input[6] ;
  assign \input[6]  = \input  [6];
  assign shiftLeftOnePos[6] = \input[5] ;
  assign \input[5]  = \input  [5];
  assign shiftLeftOnePos[5] = \input[4] ;
  assign \input[4]  = \input  [4];
  assign shiftLeftOnePos[4] = \input[3] ;
  assign \input[3]  = \input  [3];
  assign shiftLeftOnePos[3] = \input[2] ;
  assign \input[2]  = \input  [2];
  assign shiftLeftOnePos[2] = \input[1] ;
  assign \input[1]  = \input  [1];
  assign shiftLeftOnePos[1] = \input[0] ;
  assign \input[0]  = \input  [0];

endmodule


module shifter_N64_29 ( \input , shiftLeftOnePos );
  input [63:0] \input ;
  output [63:0] shiftLeftOnePos;
  wire   \input[62] , \input[61] , \input[60] , \input[59] , \input[58] ,
         \input[57] , \input[56] , \input[55] , \input[54] , \input[53] ,
         \input[52] , \input[51] , \input[50] , \input[49] , \input[48] ,
         \input[47] , \input[46] , \input[45] , \input[44] , \input[43] ,
         \input[42] , \input[41] , \input[40] , \input[39] , \input[38] ,
         \input[37] , \input[36] , \input[35] , \input[34] , \input[33] ,
         \input[32] , \input[31] , \input[30] , \input[29] , \input[28] ,
         \input[27] , \input[26] , \input[25] , \input[24] , \input[23] ,
         \input[22] , \input[21] , \input[20] , \input[19] , \input[18] ,
         \input[17] , \input[16] , \input[15] , \input[14] , \input[13] ,
         \input[12] , \input[11] , \input[10] , \input[9] , \input[8] ,
         \input[7] , \input[6] , \input[5] , \input[4] , \input[3] ,
         \input[2] , \input[1] , \input[0] ;
  assign shiftLeftOnePos[0] = 1'b0;
  assign shiftLeftOnePos[63] = \input[62] ;
  assign \input[62]  = \input  [62];
  assign shiftLeftOnePos[62] = \input[61] ;
  assign \input[61]  = \input  [61];
  assign shiftLeftOnePos[61] = \input[60] ;
  assign \input[60]  = \input  [60];
  assign shiftLeftOnePos[60] = \input[59] ;
  assign \input[59]  = \input  [59];
  assign shiftLeftOnePos[59] = \input[58] ;
  assign \input[58]  = \input  [58];
  assign shiftLeftOnePos[58] = \input[57] ;
  assign \input[57]  = \input  [57];
  assign shiftLeftOnePos[57] = \input[56] ;
  assign \input[56]  = \input  [56];
  assign shiftLeftOnePos[56] = \input[55] ;
  assign \input[55]  = \input  [55];
  assign shiftLeftOnePos[55] = \input[54] ;
  assign \input[54]  = \input  [54];
  assign shiftLeftOnePos[54] = \input[53] ;
  assign \input[53]  = \input  [53];
  assign shiftLeftOnePos[53] = \input[52] ;
  assign \input[52]  = \input  [52];
  assign shiftLeftOnePos[52] = \input[51] ;
  assign \input[51]  = \input  [51];
  assign shiftLeftOnePos[51] = \input[50] ;
  assign \input[50]  = \input  [50];
  assign shiftLeftOnePos[50] = \input[49] ;
  assign \input[49]  = \input  [49];
  assign shiftLeftOnePos[49] = \input[48] ;
  assign \input[48]  = \input  [48];
  assign shiftLeftOnePos[48] = \input[47] ;
  assign \input[47]  = \input  [47];
  assign shiftLeftOnePos[47] = \input[46] ;
  assign \input[46]  = \input  [46];
  assign shiftLeftOnePos[46] = \input[45] ;
  assign \input[45]  = \input  [45];
  assign shiftLeftOnePos[45] = \input[44] ;
  assign \input[44]  = \input  [44];
  assign shiftLeftOnePos[44] = \input[43] ;
  assign \input[43]  = \input  [43];
  assign shiftLeftOnePos[43] = \input[42] ;
  assign \input[42]  = \input  [42];
  assign shiftLeftOnePos[42] = \input[41] ;
  assign \input[41]  = \input  [41];
  assign shiftLeftOnePos[41] = \input[40] ;
  assign \input[40]  = \input  [40];
  assign shiftLeftOnePos[40] = \input[39] ;
  assign \input[39]  = \input  [39];
  assign shiftLeftOnePos[39] = \input[38] ;
  assign \input[38]  = \input  [38];
  assign shiftLeftOnePos[38] = \input[37] ;
  assign \input[37]  = \input  [37];
  assign shiftLeftOnePos[37] = \input[36] ;
  assign \input[36]  = \input  [36];
  assign shiftLeftOnePos[36] = \input[35] ;
  assign \input[35]  = \input  [35];
  assign shiftLeftOnePos[35] = \input[34] ;
  assign \input[34]  = \input  [34];
  assign shiftLeftOnePos[34] = \input[33] ;
  assign \input[33]  = \input  [33];
  assign shiftLeftOnePos[33] = \input[32] ;
  assign \input[32]  = \input  [32];
  assign shiftLeftOnePos[32] = \input[31] ;
  assign \input[31]  = \input  [31];
  assign shiftLeftOnePos[31] = \input[30] ;
  assign \input[30]  = \input  [30];
  assign shiftLeftOnePos[30] = \input[29] ;
  assign \input[29]  = \input  [29];
  assign shiftLeftOnePos[29] = \input[28] ;
  assign \input[28]  = \input  [28];
  assign shiftLeftOnePos[28] = \input[27] ;
  assign \input[27]  = \input  [27];
  assign shiftLeftOnePos[27] = \input[26] ;
  assign \input[26]  = \input  [26];
  assign shiftLeftOnePos[26] = \input[25] ;
  assign \input[25]  = \input  [25];
  assign shiftLeftOnePos[25] = \input[24] ;
  assign \input[24]  = \input  [24];
  assign shiftLeftOnePos[24] = \input[23] ;
  assign \input[23]  = \input  [23];
  assign shiftLeftOnePos[23] = \input[22] ;
  assign \input[22]  = \input  [22];
  assign shiftLeftOnePos[22] = \input[21] ;
  assign \input[21]  = \input  [21];
  assign shiftLeftOnePos[21] = \input[20] ;
  assign \input[20]  = \input  [20];
  assign shiftLeftOnePos[20] = \input[19] ;
  assign \input[19]  = \input  [19];
  assign shiftLeftOnePos[19] = \input[18] ;
  assign \input[18]  = \input  [18];
  assign shiftLeftOnePos[18] = \input[17] ;
  assign \input[17]  = \input  [17];
  assign shiftLeftOnePos[17] = \input[16] ;
  assign \input[16]  = \input  [16];
  assign shiftLeftOnePos[16] = \input[15] ;
  assign \input[15]  = \input  [15];
  assign shiftLeftOnePos[15] = \input[14] ;
  assign \input[14]  = \input  [14];
  assign shiftLeftOnePos[14] = \input[13] ;
  assign \input[13]  = \input  [13];
  assign shiftLeftOnePos[13] = \input[12] ;
  assign \input[12]  = \input  [12];
  assign shiftLeftOnePos[12] = \input[11] ;
  assign \input[11]  = \input  [11];
  assign shiftLeftOnePos[11] = \input[10] ;
  assign \input[10]  = \input  [10];
  assign shiftLeftOnePos[10] = \input[9] ;
  assign \input[9]  = \input  [9];
  assign shiftLeftOnePos[9] = \input[8] ;
  assign \input[8]  = \input  [8];
  assign shiftLeftOnePos[8] = \input[7] ;
  assign \input[7]  = \input  [7];
  assign shiftLeftOnePos[7] = \input[6] ;
  assign \input[6]  = \input  [6];
  assign shiftLeftOnePos[6] = \input[5] ;
  assign \input[5]  = \input  [5];
  assign shiftLeftOnePos[5] = \input[4] ;
  assign \input[4]  = \input  [4];
  assign shiftLeftOnePos[4] = \input[3] ;
  assign \input[3]  = \input  [3];
  assign shiftLeftOnePos[3] = \input[2] ;
  assign \input[2]  = \input  [2];
  assign shiftLeftOnePos[2] = \input[1] ;
  assign \input[1]  = \input  [1];
  assign shiftLeftOnePos[1] = \input[0] ;
  assign \input[0]  = \input  [0];

endmodule


module complementer_N64_30_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n190, n191, n192, n194, n196, n197, n198, n199, n200, n202,
         n203, n204, n206, n207, n208, n210, n211, n212, n213, n214, n216,
         n217, n218, n220, n221, n222, n224, n225, n226, n228, n229, n230,
         n232, n233, n234, n235, n237, n238, n239, n241, n242, n243, n245,
         n246, n247, n249, n250, n189, n193, n195, n201, n205, n209, n215,
         n219, n223, n227, n231, n236, n240, n244, n248, n251;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U81 ( .A(n190), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U82 ( .A(n192), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U85 ( .A(n196), .B(B[62]), .Z(DIFF[62]) );
  XOR2_X1 U86 ( .A(n194), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U87 ( .A(n198), .B(B[59]), .Z(DIFF[59]) );
  XOR2_X1 U89 ( .A(n200), .B(B[57]), .Z(DIFF[57]) );
  XOR2_X1 U90 ( .A(n202), .B(B[55]), .Z(DIFF[55]) );
  XOR2_X1 U92 ( .A(n204), .B(B[53]), .Z(DIFF[53]) );
  XOR2_X1 U93 ( .A(n206), .B(B[51]), .Z(DIFF[51]) );
  XOR2_X1 U95 ( .A(n208), .B(B[49]), .Z(DIFF[49]) );
  XOR2_X1 U96 ( .A(n212), .B(B[47]), .Z(DIFF[47]) );
  XOR2_X1 U98 ( .A(n214), .B(B[45]), .Z(DIFF[45]) );
  XOR2_X1 U99 ( .A(n216), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U101 ( .A(n218), .B(B[41]), .Z(DIFF[41]) );
  XOR2_X1 U102 ( .A(n211), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U103 ( .A(n220), .B(B[39]), .Z(DIFF[39]) );
  XOR2_X1 U105 ( .A(n222), .B(B[37]), .Z(DIFF[37]) );
  XOR2_X1 U106 ( .A(n224), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U108 ( .A(n226), .B(B[33]), .Z(DIFF[33]) );
  XOR2_X1 U109 ( .A(n228), .B(B[31]), .Z(DIFF[31]) );
  XOR2_X1 U111 ( .A(n230), .B(B[29]), .Z(DIFF[29]) );
  XOR2_X1 U112 ( .A(n233), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U114 ( .A(n235), .B(B[25]), .Z(DIFF[25]) );
  XOR2_X1 U115 ( .A(n237), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U117 ( .A(n239), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U118 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U119 ( .A(n241), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U121 ( .A(n243), .B(B[17]), .Z(DIFF[17]) );
  XOR2_X1 U122 ( .A(n245), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U124 ( .A(n247), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U125 ( .A(n249), .B(B[11]), .Z(DIFF[11]) );
  XNOR2_X1 U1 ( .A(B[44]), .B(n217), .ZN(DIFF[44]) );
  NOR2_X1 U2 ( .A1(B[43]), .A2(n216), .ZN(n217) );
  XNOR2_X1 U3 ( .A(B[40]), .B(n221), .ZN(DIFF[40]) );
  NOR2_X1 U4 ( .A1(B[39]), .A2(n220), .ZN(n221) );
  OR3_X1 U5 ( .A1(B[43]), .A2(B[44]), .A3(n216), .ZN(n214) );
  OR3_X1 U6 ( .A1(B[39]), .A2(B[40]), .A3(n220), .ZN(n218) );
  NOR3_X1 U7 ( .A1(B[59]), .A2(B[60]), .A3(n198), .ZN(n197) );
  XNOR2_X1 U8 ( .A(n189), .B(B[54]), .ZN(DIFF[54]) );
  NOR2_X1 U9 ( .A1(n204), .A2(B[53]), .ZN(n189) );
  XNOR2_X1 U10 ( .A(B[60]), .B(n199), .ZN(DIFF[60]) );
  NOR2_X1 U11 ( .A1(B[59]), .A2(n198), .ZN(n199) );
  XOR2_X1 U12 ( .A(n197), .B(n251), .Z(DIFF[61]) );
  NAND2_X1 U13 ( .A1(n197), .A2(n251), .ZN(n196) );
  OR3_X1 U14 ( .A1(B[53]), .A2(B[54]), .A3(n204), .ZN(n202) );
  OR3_X1 U15 ( .A1(B[49]), .A2(B[50]), .A3(n208), .ZN(n206) );
  XNOR2_X1 U16 ( .A(n193), .B(B[50]), .ZN(DIFF[50]) );
  NOR2_X1 U17 ( .A1(n208), .A2(B[49]), .ZN(n193) );
  XNOR2_X1 U18 ( .A(B[36]), .B(n225), .ZN(DIFF[36]) );
  NOR2_X1 U19 ( .A1(B[35]), .A2(n224), .ZN(n225) );
  XNOR2_X1 U20 ( .A(n195), .B(B[34]), .ZN(DIFF[34]) );
  NOR2_X1 U21 ( .A1(n226), .A2(B[33]), .ZN(n195) );
  XNOR2_X1 U22 ( .A(n201), .B(B[38]), .ZN(DIFF[38]) );
  NOR2_X1 U23 ( .A1(n222), .A2(B[37]), .ZN(n201) );
  XNOR2_X1 U24 ( .A(B[48]), .B(n213), .ZN(DIFF[48]) );
  NOR2_X1 U25 ( .A1(B[47]), .A2(n212), .ZN(n213) );
  OR3_X1 U26 ( .A1(B[37]), .A2(B[38]), .A3(n222), .ZN(n220) );
  OR3_X1 U27 ( .A1(B[41]), .A2(B[42]), .A3(n218), .ZN(n216) );
  OR3_X1 U28 ( .A1(B[45]), .A2(B[46]), .A3(n214), .ZN(n212) );
  OR3_X1 U29 ( .A1(B[35]), .A2(B[36]), .A3(n224), .ZN(n222) );
  OR3_X1 U30 ( .A1(B[33]), .A2(B[34]), .A3(n226), .ZN(n224) );
  XNOR2_X1 U31 ( .A(n205), .B(B[42]), .ZN(DIFF[42]) );
  NOR2_X1 U32 ( .A1(n218), .A2(B[41]), .ZN(n205) );
  XNOR2_X1 U33 ( .A(n209), .B(B[46]), .ZN(DIFF[46]) );
  NOR2_X1 U34 ( .A1(n214), .A2(B[45]), .ZN(n209) );
  XNOR2_X1 U35 ( .A(B[52]), .B(n207), .ZN(DIFF[52]) );
  NOR2_X1 U36 ( .A1(B[51]), .A2(n206), .ZN(n207) );
  XNOR2_X1 U37 ( .A(B[56]), .B(n203), .ZN(DIFF[56]) );
  NOR2_X1 U38 ( .A1(B[55]), .A2(n202), .ZN(n203) );
  OR3_X1 U39 ( .A1(B[57]), .A2(B[58]), .A3(n200), .ZN(n198) );
  OR3_X1 U40 ( .A1(B[47]), .A2(B[48]), .A3(n212), .ZN(n208) );
  OR3_X1 U41 ( .A1(B[51]), .A2(B[52]), .A3(n206), .ZN(n204) );
  OR3_X1 U42 ( .A1(B[55]), .A2(B[56]), .A3(n202), .ZN(n200) );
  XNOR2_X1 U43 ( .A(n215), .B(B[63]), .ZN(DIFF[63]) );
  NOR2_X1 U44 ( .A1(n196), .A2(B[62]), .ZN(n215) );
  XNOR2_X1 U45 ( .A(n219), .B(B[58]), .ZN(DIFF[58]) );
  NOR2_X1 U46 ( .A1(n200), .A2(B[57]), .ZN(n219) );
  XNOR2_X1 U47 ( .A(n223), .B(B[22]), .ZN(DIFF[22]) );
  NOR2_X1 U48 ( .A1(n239), .A2(B[21]), .ZN(n223) );
  XNOR2_X1 U49 ( .A(n227), .B(B[18]), .ZN(DIFF[18]) );
  NOR2_X1 U50 ( .A1(n243), .A2(B[17]), .ZN(n227) );
  XNOR2_X1 U51 ( .A(n231), .B(B[14]), .ZN(DIFF[14]) );
  NOR2_X1 U52 ( .A1(n247), .A2(B[13]), .ZN(n231) );
  XNOR2_X1 U53 ( .A(n236), .B(B[10]), .ZN(DIFF[10]) );
  NOR2_X1 U54 ( .A1(n190), .A2(B[9]), .ZN(n236) );
  XNOR2_X1 U55 ( .A(n240), .B(B[6]), .ZN(DIFF[6]) );
  NOR2_X1 U56 ( .A1(n194), .A2(B[5]), .ZN(n240) );
  XNOR2_X1 U57 ( .A(B[20]), .B(n242), .ZN(DIFF[20]) );
  NOR2_X1 U58 ( .A1(B[19]), .A2(n241), .ZN(n242) );
  XNOR2_X1 U59 ( .A(B[16]), .B(n246), .ZN(DIFF[16]) );
  NOR2_X1 U60 ( .A1(B[15]), .A2(n245), .ZN(n246) );
  XNOR2_X1 U61 ( .A(B[12]), .B(n250), .ZN(DIFF[12]) );
  NOR2_X1 U62 ( .A1(B[11]), .A2(n249), .ZN(n250) );
  XNOR2_X1 U63 ( .A(B[8]), .B(n191), .ZN(DIFF[8]) );
  NOR2_X1 U64 ( .A1(B[7]), .A2(n192), .ZN(n191) );
  XNOR2_X1 U65 ( .A(B[4]), .B(n210), .ZN(DIFF[4]) );
  NOR2_X1 U66 ( .A1(B[3]), .A2(n211), .ZN(n210) );
  OR3_X1 U67 ( .A1(B[5]), .A2(B[6]), .A3(n194), .ZN(n192) );
  OR3_X1 U68 ( .A1(B[13]), .A2(B[14]), .A3(n247), .ZN(n245) );
  OR3_X1 U69 ( .A1(B[17]), .A2(B[18]), .A3(n243), .ZN(n241) );
  OR3_X1 U70 ( .A1(B[21]), .A2(B[22]), .A3(n239), .ZN(n237) );
  OR3_X1 U71 ( .A1(B[10]), .A2(B[9]), .A3(n190), .ZN(n249) );
  OR3_X1 U72 ( .A1(B[3]), .A2(B[4]), .A3(n211), .ZN(n194) );
  OR3_X1 U73 ( .A1(B[7]), .A2(B[8]), .A3(n192), .ZN(n190) );
  OR3_X1 U74 ( .A1(B[11]), .A2(B[12]), .A3(n249), .ZN(n247) );
  OR3_X1 U75 ( .A1(B[15]), .A2(B[16]), .A3(n245), .ZN(n243) );
  OR3_X1 U76 ( .A1(B[19]), .A2(B[20]), .A3(n241), .ZN(n239) );
  XNOR2_X1 U77 ( .A(n244), .B(B[30]), .ZN(DIFF[30]) );
  NOR2_X1 U78 ( .A1(n230), .A2(B[29]), .ZN(n244) );
  XNOR2_X1 U79 ( .A(n248), .B(B[26]), .ZN(DIFF[26]) );
  NOR2_X1 U80 ( .A1(n235), .A2(B[25]), .ZN(n248) );
  XNOR2_X1 U83 ( .A(B[32]), .B(n229), .ZN(DIFF[32]) );
  NOR2_X1 U84 ( .A1(B[31]), .A2(n228), .ZN(n229) );
  XNOR2_X1 U88 ( .A(B[28]), .B(n234), .ZN(DIFF[28]) );
  NOR2_X1 U91 ( .A1(B[27]), .A2(n233), .ZN(n234) );
  XNOR2_X1 U94 ( .A(B[24]), .B(n238), .ZN(DIFF[24]) );
  NOR2_X1 U97 ( .A1(B[23]), .A2(n237), .ZN(n238) );
  OR3_X1 U100 ( .A1(B[25]), .A2(B[26]), .A3(n235), .ZN(n233) );
  OR3_X1 U104 ( .A1(B[29]), .A2(B[30]), .A3(n230), .ZN(n228) );
  OR3_X1 U107 ( .A1(B[23]), .A2(B[24]), .A3(n237), .ZN(n235) );
  OR3_X1 U110 ( .A1(B[27]), .A2(B[28]), .A3(n233), .ZN(n230) );
  OR3_X1 U113 ( .A1(B[31]), .A2(B[32]), .A3(n228), .ZN(n226) );
  OR3_X1 U116 ( .A1(B[1]), .A2(B[2]), .A3(\B[0] ), .ZN(n211) );
  XNOR2_X1 U120 ( .A(B[2]), .B(n232), .ZN(DIFF[2]) );
  NOR2_X1 U123 ( .A1(\B[0] ), .A2(B[1]), .ZN(n232) );
  INV_X1 U126 ( .A(B[61]), .ZN(n251) );
endmodule


module complementer_N64_30 ( \input , complement2 );
  input [63:0] \input ;
  output [63:0] complement2;


  complementer_N64_30_DW01_sub_0 sub_add_31_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(\input ), .CI(1'b0), .DIFF(complement2) );
endmodule


module complementer_N64_29_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n189;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U81 ( .A(n190), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U82 ( .A(n192), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U83 ( .A(n193), .B(B[6]), .Z(DIFF[6]) );
  XOR2_X1 U84 ( .A(n195), .B(B[63]), .Z(DIFF[63]) );
  XOR2_X1 U85 ( .A(n196), .B(B[62]), .Z(DIFF[62]) );
  XOR2_X1 U86 ( .A(n194), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U87 ( .A(n198), .B(B[59]), .Z(DIFF[59]) );
  XOR2_X1 U88 ( .A(n201), .B(B[58]), .Z(DIFF[58]) );
  XOR2_X1 U89 ( .A(n200), .B(B[57]), .Z(DIFF[57]) );
  XOR2_X1 U90 ( .A(n202), .B(B[55]), .Z(DIFF[55]) );
  XOR2_X1 U91 ( .A(n205), .B(B[54]), .Z(DIFF[54]) );
  XOR2_X1 U92 ( .A(n204), .B(B[53]), .Z(DIFF[53]) );
  XOR2_X1 U93 ( .A(n206), .B(B[51]), .Z(DIFF[51]) );
  XOR2_X1 U94 ( .A(n209), .B(B[50]), .Z(DIFF[50]) );
  XOR2_X1 U95 ( .A(n208), .B(B[49]), .Z(DIFF[49]) );
  XOR2_X1 U96 ( .A(n212), .B(B[47]), .Z(DIFF[47]) );
  XOR2_X1 U97 ( .A(n215), .B(B[46]), .Z(DIFF[46]) );
  XOR2_X1 U98 ( .A(n214), .B(B[45]), .Z(DIFF[45]) );
  XOR2_X1 U99 ( .A(n216), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U100 ( .A(n219), .B(B[42]), .Z(DIFF[42]) );
  XOR2_X1 U101 ( .A(n218), .B(B[41]), .Z(DIFF[41]) );
  XOR2_X1 U102 ( .A(n211), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U103 ( .A(n220), .B(B[39]), .Z(DIFF[39]) );
  XOR2_X1 U104 ( .A(n223), .B(B[38]), .Z(DIFF[38]) );
  XOR2_X1 U105 ( .A(n222), .B(B[37]), .Z(DIFF[37]) );
  XOR2_X1 U106 ( .A(n224), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U107 ( .A(n227), .B(B[34]), .Z(DIFF[34]) );
  XOR2_X1 U108 ( .A(n226), .B(B[33]), .Z(DIFF[33]) );
  XOR2_X1 U109 ( .A(n228), .B(B[31]), .Z(DIFF[31]) );
  XOR2_X1 U110 ( .A(n231), .B(B[30]), .Z(DIFF[30]) );
  XOR2_X1 U111 ( .A(n230), .B(B[29]), .Z(DIFF[29]) );
  XOR2_X1 U112 ( .A(n233), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U113 ( .A(n236), .B(B[26]), .Z(DIFF[26]) );
  XOR2_X1 U114 ( .A(n235), .B(B[25]), .Z(DIFF[25]) );
  XOR2_X1 U115 ( .A(n237), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U116 ( .A(n240), .B(B[22]), .Z(DIFF[22]) );
  XOR2_X1 U117 ( .A(n239), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U118 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U119 ( .A(n241), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U120 ( .A(n244), .B(B[18]), .Z(DIFF[18]) );
  XOR2_X1 U121 ( .A(n243), .B(B[17]), .Z(DIFF[17]) );
  XOR2_X1 U122 ( .A(n245), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U123 ( .A(n248), .B(B[14]), .Z(DIFF[14]) );
  XOR2_X1 U124 ( .A(n247), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U125 ( .A(n249), .B(B[11]), .Z(DIFF[11]) );
  XOR2_X1 U126 ( .A(n251), .B(B[10]), .Z(DIFF[10]) );
  NAND2_X1 U1 ( .A1(n197), .A2(n189), .ZN(n196) );
  NOR2_X1 U2 ( .A1(B[43]), .A2(n216), .ZN(n217) );
  NOR2_X1 U3 ( .A1(B[39]), .A2(n220), .ZN(n221) );
  OR3_X1 U4 ( .A1(B[43]), .A2(B[44]), .A3(n216), .ZN(n214) );
  OR3_X1 U5 ( .A1(B[39]), .A2(B[40]), .A3(n220), .ZN(n218) );
  XNOR2_X1 U6 ( .A(B[44]), .B(n217), .ZN(DIFF[44]) );
  XNOR2_X1 U7 ( .A(B[48]), .B(n213), .ZN(DIFF[48]) );
  XNOR2_X1 U8 ( .A(B[40]), .B(n221), .ZN(DIFF[40]) );
  OR2_X1 U9 ( .A1(n218), .A2(B[41]), .ZN(n219) );
  NOR3_X1 U10 ( .A1(B[59]), .A2(B[60]), .A3(n198), .ZN(n197) );
  NOR2_X1 U11 ( .A1(B[55]), .A2(n202), .ZN(n203) );
  NOR2_X1 U12 ( .A1(B[51]), .A2(n206), .ZN(n207) );
  NOR2_X1 U13 ( .A1(B[59]), .A2(n198), .ZN(n199) );
  OR3_X1 U14 ( .A1(B[45]), .A2(B[46]), .A3(n214), .ZN(n212) );
  OR3_X1 U15 ( .A1(B[53]), .A2(B[54]), .A3(n204), .ZN(n202) );
  OR3_X1 U16 ( .A1(B[49]), .A2(B[50]), .A3(n208), .ZN(n206) );
  OR3_X1 U17 ( .A1(B[55]), .A2(B[56]), .A3(n202), .ZN(n200) );
  XNOR2_X1 U18 ( .A(B[60]), .B(n199), .ZN(DIFF[60]) );
  OR2_X1 U19 ( .A1(n214), .A2(B[45]), .ZN(n215) );
  OR2_X1 U20 ( .A1(n204), .A2(B[53]), .ZN(n205) );
  OR2_X1 U21 ( .A1(n208), .A2(B[49]), .ZN(n209) );
  NOR2_X1 U22 ( .A1(B[35]), .A2(n224), .ZN(n225) );
  OR3_X1 U23 ( .A1(B[37]), .A2(B[38]), .A3(n222), .ZN(n220) );
  OR3_X1 U24 ( .A1(B[41]), .A2(B[42]), .A3(n218), .ZN(n216) );
  XNOR2_X1 U25 ( .A(B[36]), .B(n225), .ZN(DIFF[36]) );
  OR3_X1 U26 ( .A1(B[35]), .A2(B[36]), .A3(n224), .ZN(n222) );
  OR2_X1 U27 ( .A1(n222), .A2(B[37]), .ZN(n223) );
  NOR2_X1 U28 ( .A1(B[47]), .A2(n212), .ZN(n213) );
  OR3_X1 U29 ( .A1(B[57]), .A2(B[58]), .A3(n200), .ZN(n198) );
  OR3_X1 U30 ( .A1(B[47]), .A2(B[48]), .A3(n212), .ZN(n208) );
  OR3_X1 U31 ( .A1(B[51]), .A2(B[52]), .A3(n206), .ZN(n204) );
  XNOR2_X1 U32 ( .A(B[52]), .B(n207), .ZN(DIFF[52]) );
  XNOR2_X1 U33 ( .A(n197), .B(B[61]), .ZN(DIFF[61]) );
  XNOR2_X1 U34 ( .A(B[56]), .B(n203), .ZN(DIFF[56]) );
  OR2_X1 U35 ( .A1(n196), .A2(B[62]), .ZN(n195) );
  OR2_X1 U36 ( .A1(n200), .A2(B[57]), .ZN(n201) );
  NOR2_X1 U37 ( .A1(B[3]), .A2(n211), .ZN(n210) );
  NOR2_X1 U38 ( .A1(B[19]), .A2(n241), .ZN(n242) );
  NOR2_X1 U39 ( .A1(B[15]), .A2(n245), .ZN(n246) );
  NOR2_X1 U40 ( .A1(B[11]), .A2(n249), .ZN(n250) );
  NOR2_X1 U41 ( .A1(B[7]), .A2(n192), .ZN(n191) );
  OR3_X1 U42 ( .A1(B[10]), .A2(B[9]), .A3(n190), .ZN(n249) );
  OR3_X1 U43 ( .A1(B[5]), .A2(B[6]), .A3(n194), .ZN(n192) );
  OR3_X1 U44 ( .A1(B[13]), .A2(B[14]), .A3(n247), .ZN(n245) );
  OR3_X1 U45 ( .A1(B[17]), .A2(B[18]), .A3(n243), .ZN(n241) );
  OR3_X1 U46 ( .A1(B[7]), .A2(B[8]), .A3(n192), .ZN(n190) );
  OR3_X1 U47 ( .A1(B[3]), .A2(B[4]), .A3(n211), .ZN(n194) );
  OR3_X1 U48 ( .A1(B[11]), .A2(B[12]), .A3(n249), .ZN(n247) );
  OR3_X1 U49 ( .A1(B[15]), .A2(B[16]), .A3(n245), .ZN(n243) );
  XNOR2_X1 U50 ( .A(B[4]), .B(n210), .ZN(DIFF[4]) );
  XNOR2_X1 U51 ( .A(B[20]), .B(n242), .ZN(DIFF[20]) );
  XNOR2_X1 U52 ( .A(B[16]), .B(n246), .ZN(DIFF[16]) );
  XNOR2_X1 U53 ( .A(B[12]), .B(n250), .ZN(DIFF[12]) );
  XNOR2_X1 U54 ( .A(B[8]), .B(n191), .ZN(DIFF[8]) );
  OR2_X1 U55 ( .A1(n243), .A2(B[17]), .ZN(n244) );
  OR2_X1 U56 ( .A1(n247), .A2(B[13]), .ZN(n248) );
  OR2_X1 U57 ( .A1(n190), .A2(B[9]), .ZN(n251) );
  OR2_X1 U58 ( .A1(n194), .A2(B[5]), .ZN(n193) );
  NOR2_X1 U59 ( .A1(B[31]), .A2(n228), .ZN(n229) );
  NOR2_X1 U60 ( .A1(B[27]), .A2(n233), .ZN(n234) );
  NOR2_X1 U61 ( .A1(B[23]), .A2(n237), .ZN(n238) );
  OR3_X1 U62 ( .A1(B[33]), .A2(B[34]), .A3(n226), .ZN(n224) );
  OR3_X1 U63 ( .A1(B[29]), .A2(B[30]), .A3(n230), .ZN(n228) );
  OR3_X1 U64 ( .A1(B[25]), .A2(B[26]), .A3(n235), .ZN(n233) );
  OR3_X1 U65 ( .A1(B[21]), .A2(B[22]), .A3(n239), .ZN(n237) );
  OR3_X1 U66 ( .A1(B[31]), .A2(B[32]), .A3(n228), .ZN(n226) );
  OR3_X1 U67 ( .A1(B[27]), .A2(B[28]), .A3(n233), .ZN(n230) );
  OR3_X1 U68 ( .A1(B[23]), .A2(B[24]), .A3(n237), .ZN(n235) );
  OR3_X1 U69 ( .A1(B[19]), .A2(B[20]), .A3(n241), .ZN(n239) );
  XNOR2_X1 U70 ( .A(B[32]), .B(n229), .ZN(DIFF[32]) );
  XNOR2_X1 U71 ( .A(B[28]), .B(n234), .ZN(DIFF[28]) );
  XNOR2_X1 U72 ( .A(B[24]), .B(n238), .ZN(DIFF[24]) );
  OR2_X1 U73 ( .A1(n226), .A2(B[33]), .ZN(n227) );
  OR2_X1 U74 ( .A1(n230), .A2(B[29]), .ZN(n231) );
  OR2_X1 U75 ( .A1(n235), .A2(B[25]), .ZN(n236) );
  OR2_X1 U76 ( .A1(n239), .A2(B[21]), .ZN(n240) );
  XNOR2_X1 U77 ( .A(B[2]), .B(n232), .ZN(DIFF[2]) );
  OR3_X1 U78 ( .A1(B[1]), .A2(B[2]), .A3(\B[0] ), .ZN(n211) );
  NOR2_X1 U79 ( .A1(\B[0] ), .A2(B[1]), .ZN(n232) );
  INV_X1 U80 ( .A(B[61]), .ZN(n189) );
endmodule


module complementer_N64_29 ( \input , complement2 );
  input [63:0] \input ;
  output [63:0] complement2;


  complementer_N64_29_DW01_sub_0 sub_add_31_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(\input ), .CI(1'b0), .DIFF(complement2) );
endmodule


module ShiftnCompl_N64_0 ( plusA, plus2A_out, minus2A_out, plus4A_out, 
        minus4A_out );
  input [63:0] plusA;
  output [63:0] plus2A_out;
  output [63:0] minus2A_out;
  output [63:0] plus4A_out;
  output [63:0] minus4A_out;
  wire   n45, n46, n3, n47, n48, n4, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign plus2A_out[0] = 1'b0;
  assign plus2A_out[51] = n3;
  assign plus2A_out[39] = n4;
  assign plus4A_out[0] = 1'b0;

  shifter_N64_30 shifter_1 ( .\input (plusA), .shiftLeftOnePos({
        plus2A_out[63:59], n45, plus2A_out[57:54], n46, plus2A_out[52], n3, 
        plus2A_out[50:49], n47, plus2A_out[47:44], n48, plus2A_out[42:40], n4, 
        n49, plus2A_out[37:32], n50, n51, n52, n53, n54, n55, n56, n57, n58, 
        n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, 
        n73, n74, n75, n76, n77, n78, n79, plus2A_out[1], 
        SYNOPSYS_UNCONNECTED__0}) );
  shifter_N64_29 shifter_2 ( .\input ({plus2A_out[63:52], n3, 
        plus2A_out[50:40], n4, plus2A_out[38:1], 1'b0}), .shiftLeftOnePos({
        plus4A_out[63:59], n80, plus4A_out[57:54], n81, plus4A_out[52:49], n82, 
        plus4A_out[47:44], n83, plus4A_out[42:39], n84, plus4A_out[37:1], 
        SYNOPSYS_UNCONNECTED__1}) );
  complementer_N64_30 complementer_1 ( .\input ({plus2A_out[63:52], n3, 
        plus2A_out[50:40], n4, plus2A_out[38:1], 1'b0}), .complement2(
        minus2A_out) );
  complementer_N64_29 complementer_2 ( .\input ({plus4A_out[63:1], 1'b0}), 
        .complement2(minus4A_out) );
  BUF_X1 U1 ( .A(n48), .Z(plus2A_out[43]) );
  BUF_X1 U2 ( .A(n83), .Z(plus4A_out[43]) );
  BUF_X1 U5 ( .A(n49), .Z(plus2A_out[38]) );
  BUF_X1 U6 ( .A(n84), .Z(plus4A_out[38]) );
  BUF_X1 U7 ( .A(n81), .Z(plus4A_out[53]) );
  BUF_X1 U8 ( .A(n46), .Z(plus2A_out[53]) );
  BUF_X1 U9 ( .A(n82), .Z(plus4A_out[48]) );
  BUF_X1 U10 ( .A(n47), .Z(plus2A_out[48]) );
  BUF_X1 U11 ( .A(n80), .Z(plus4A_out[58]) );
  BUF_X1 U12 ( .A(n45), .Z(plus2A_out[58]) );
  BUF_X1 U13 ( .A(n74), .Z(plus2A_out[7]) );
  BUF_X1 U14 ( .A(n72), .Z(plus2A_out[9]) );
  BUF_X1 U15 ( .A(n76), .Z(plus2A_out[5]) );
  BUF_X1 U16 ( .A(n75), .Z(plus2A_out[6]) );
  BUF_X1 U17 ( .A(n73), .Z(plus2A_out[8]) );
  BUF_X1 U18 ( .A(n77), .Z(plus2A_out[4]) );
  BUF_X1 U19 ( .A(n62), .Z(plus2A_out[19]) );
  BUF_X1 U20 ( .A(n66), .Z(plus2A_out[15]) );
  BUF_X1 U21 ( .A(n70), .Z(plus2A_out[11]) );
  BUF_X1 U22 ( .A(n64), .Z(plus2A_out[17]) );
  BUF_X1 U23 ( .A(n68), .Z(plus2A_out[13]) );
  BUF_X1 U24 ( .A(n71), .Z(plus2A_out[10]) );
  BUF_X1 U25 ( .A(n63), .Z(plus2A_out[18]) );
  BUF_X1 U26 ( .A(n67), .Z(plus2A_out[14]) );
  BUF_X1 U27 ( .A(n65), .Z(plus2A_out[16]) );
  BUF_X1 U28 ( .A(n69), .Z(plus2A_out[12]) );
  BUF_X1 U29 ( .A(n54), .Z(plus2A_out[27]) );
  BUF_X1 U30 ( .A(n58), .Z(plus2A_out[23]) );
  BUF_X1 U31 ( .A(n52), .Z(plus2A_out[29]) );
  BUF_X1 U32 ( .A(n56), .Z(plus2A_out[25]) );
  BUF_X1 U33 ( .A(n60), .Z(plus2A_out[21]) );
  BUF_X1 U34 ( .A(n51), .Z(plus2A_out[30]) );
  BUF_X1 U35 ( .A(n55), .Z(plus2A_out[26]) );
  BUF_X1 U36 ( .A(n59), .Z(plus2A_out[22]) );
  BUF_X1 U37 ( .A(n53), .Z(plus2A_out[28]) );
  BUF_X1 U38 ( .A(n57), .Z(plus2A_out[24]) );
  BUF_X1 U39 ( .A(n61), .Z(plus2A_out[20]) );
  BUF_X1 U40 ( .A(n50), .Z(plus2A_out[31]) );
  BUF_X2 U41 ( .A(n78), .Z(plus2A_out[3]) );
  BUF_X1 U42 ( .A(n79), .Z(plus2A_out[2]) );
endmodule


module MUX_GENERIC_N64_RADIX3_15 ( plusA, minusA, plus2A, minus2A, SEL, Y );
  input [63:0] plusA;
  input [63:0] minusA;
  input [63:0] plus2A;
  input [63:0] minus2A;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498;
  tri   [63:0] Y;

  TBUF_X1 \Y_tri[0]  ( .A(n498), .EN(n293), .Z(Y[0]) );
  TBUF_X1 \Y_tri[1]  ( .A(n497), .EN(n293), .Z(Y[1]) );
  TBUF_X1 \Y_tri[55]  ( .A(n442), .EN(n297), .Z(Y[55]) );
  TBUF_X1 \Y_tri[56]  ( .A(n441), .EN(n296), .Z(Y[56]) );
  TBUF_X1 \Y_tri[57]  ( .A(n440), .EN(n295), .Z(Y[57]) );
  TBUF_X1 \Y_tri[58]  ( .A(n439), .EN(n294), .Z(Y[58]) );
  TBUF_X1 \Y_tri[59]  ( .A(n438), .EN(n298), .Z(Y[59]) );
  TBUF_X1 \Y_tri[60]  ( .A(n437), .EN(n297), .Z(Y[60]) );
  TBUF_X1 \Y_tri[61]  ( .A(n436), .EN(n296), .Z(Y[61]) );
  TBUF_X1 \Y_tri[62]  ( .A(n435), .EN(n295), .Z(Y[62]) );
  TBUF_X1 \Y_tri[63]  ( .A(n434), .EN(n294), .Z(Y[63]) );
  TBUF_X1 \Y_tri[49]  ( .A(n448), .EN(n298), .Z(Y[49]) );
  TBUF_X1 \Y_tri[50]  ( .A(n447), .EN(n297), .Z(Y[50]) );
  TBUF_X1 \Y_tri[51]  ( .A(n446), .EN(n296), .Z(Y[51]) );
  TBUF_X1 \Y_tri[52]  ( .A(n445), .EN(n295), .Z(Y[52]) );
  TBUF_X1 \Y_tri[53]  ( .A(n444), .EN(n294), .Z(Y[53]) );
  TBUF_X1 \Y_tri[54]  ( .A(n443), .EN(n298), .Z(Y[54]) );
  TBUF_X1 \Y_tri[24]  ( .A(n473), .EN(n298), .Z(Y[24]) );
  TBUF_X1 \Y_tri[25]  ( .A(n472), .EN(n297), .Z(Y[25]) );
  TBUF_X1 \Y_tri[26]  ( .A(n471), .EN(n296), .Z(Y[26]) );
  TBUF_X1 \Y_tri[27]  ( .A(n470), .EN(n295), .Z(Y[27]) );
  TBUF_X1 \Y_tri[28]  ( .A(n469), .EN(n294), .Z(Y[28]) );
  TBUF_X1 \Y_tri[29]  ( .A(n468), .EN(n298), .Z(Y[29]) );
  TBUF_X1 \Y_tri[30]  ( .A(n467), .EN(n297), .Z(Y[30]) );
  TBUF_X1 \Y_tri[31]  ( .A(n466), .EN(n296), .Z(Y[31]) );
  TBUF_X1 \Y_tri[32]  ( .A(n465), .EN(n295), .Z(Y[32]) );
  TBUF_X1 \Y_tri[33]  ( .A(n464), .EN(n294), .Z(Y[33]) );
  TBUF_X1 \Y_tri[34]  ( .A(n463), .EN(n298), .Z(Y[34]) );
  TBUF_X1 \Y_tri[35]  ( .A(n462), .EN(n297), .Z(Y[35]) );
  TBUF_X1 \Y_tri[36]  ( .A(n461), .EN(n296), .Z(Y[36]) );
  TBUF_X1 \Y_tri[37]  ( .A(n460), .EN(n295), .Z(Y[37]) );
  TBUF_X1 \Y_tri[38]  ( .A(n459), .EN(n294), .Z(Y[38]) );
  TBUF_X1 \Y_tri[39]  ( .A(n458), .EN(n298), .Z(Y[39]) );
  TBUF_X1 \Y_tri[40]  ( .A(n457), .EN(n297), .Z(Y[40]) );
  TBUF_X1 \Y_tri[41]  ( .A(n456), .EN(n296), .Z(Y[41]) );
  TBUF_X1 \Y_tri[42]  ( .A(n455), .EN(n295), .Z(Y[42]) );
  TBUF_X1 \Y_tri[43]  ( .A(n454), .EN(n294), .Z(Y[43]) );
  TBUF_X1 \Y_tri[44]  ( .A(n453), .EN(n298), .Z(Y[44]) );
  TBUF_X1 \Y_tri[45]  ( .A(n452), .EN(n297), .Z(Y[45]) );
  TBUF_X1 \Y_tri[46]  ( .A(n451), .EN(n296), .Z(Y[46]) );
  TBUF_X1 \Y_tri[47]  ( .A(n450), .EN(n295), .Z(Y[47]) );
  TBUF_X1 \Y_tri[48]  ( .A(n449), .EN(n294), .Z(Y[48]) );
  TBUF_X1 \Y_tri[5]  ( .A(n493), .EN(n297), .Z(Y[5]) );
  TBUF_X1 \Y_tri[6]  ( .A(n492), .EN(n296), .Z(Y[6]) );
  TBUF_X1 \Y_tri[7]  ( .A(n491), .EN(n295), .Z(Y[7]) );
  TBUF_X1 \Y_tri[8]  ( .A(n490), .EN(n294), .Z(Y[8]) );
  TBUF_X1 \Y_tri[9]  ( .A(n488), .EN(n298), .Z(Y[9]) );
  TBUF_X1 \Y_tri[10]  ( .A(n487), .EN(n297), .Z(Y[10]) );
  TBUF_X1 \Y_tri[2]  ( .A(n496), .EN(n295), .Z(Y[2]) );
  TBUF_X1 \Y_tri[3]  ( .A(n495), .EN(n294), .Z(Y[3]) );
  TBUF_X1 \Y_tri[4]  ( .A(n494), .EN(n298), .Z(Y[4]) );
  TBUF_X1 \Y_tri[11]  ( .A(n486), .EN(n296), .Z(Y[11]) );
  TBUF_X1 \Y_tri[12]  ( .A(n485), .EN(n295), .Z(Y[12]) );
  TBUF_X1 \Y_tri[13]  ( .A(n484), .EN(n294), .Z(Y[13]) );
  TBUF_X1 \Y_tri[14]  ( .A(n483), .EN(n298), .Z(Y[14]) );
  TBUF_X1 \Y_tri[16]  ( .A(n481), .EN(n296), .Z(Y[16]) );
  TBUF_X1 \Y_tri[17]  ( .A(n480), .EN(n295), .Z(Y[17]) );
  TBUF_X1 \Y_tri[18]  ( .A(n479), .EN(n294), .Z(Y[18]) );
  TBUF_X1 \Y_tri[19]  ( .A(n478), .EN(n298), .Z(Y[19]) );
  TBUF_X1 \Y_tri[20]  ( .A(n477), .EN(n297), .Z(Y[20]) );
  TBUF_X1 \Y_tri[21]  ( .A(n476), .EN(n296), .Z(Y[21]) );
  TBUF_X1 \Y_tri[22]  ( .A(n475), .EN(n295), .Z(Y[22]) );
  TBUF_X1 \Y_tri[23]  ( .A(n474), .EN(n294), .Z(Y[23]) );
  TBUF_X1 \Y_tri[15]  ( .A(n482), .EN(n297), .Z(Y[15]) );
  BUF_X2 U2 ( .A(n272), .Z(n280) );
  NAND2_X1 U3 ( .A1(n392), .A2(n391), .ZN(n453) );
  AOI22_X1 U4 ( .A1(plusA[44]), .A2(n280), .B1(plus2A[44]), .B2(n276), .ZN(
        n392) );
  AOI22_X1 U5 ( .A1(minus2A[44]), .A2(n290), .B1(minusA[44]), .B2(n284), .ZN(
        n391) );
  NAND2_X1 U6 ( .A1(n390), .A2(n389), .ZN(n454) );
  AOI22_X1 U7 ( .A1(plusA[43]), .A2(n280), .B1(plus2A[43]), .B2(n276), .ZN(
        n390) );
  AOI22_X1 U8 ( .A1(minus2A[43]), .A2(n290), .B1(minusA[43]), .B2(n284), .ZN(
        n389) );
  NAND2_X1 U9 ( .A1(n394), .A2(n393), .ZN(n452) );
  AOI22_X1 U10 ( .A1(plusA[45]), .A2(n280), .B1(plus2A[45]), .B2(n276), .ZN(
        n394) );
  AOI22_X1 U11 ( .A1(minus2A[45]), .A2(n290), .B1(minusA[45]), .B2(n284), .ZN(
        n393) );
  NAND2_X1 U12 ( .A1(n400), .A2(n399), .ZN(n449) );
  AOI22_X1 U13 ( .A1(plusA[48]), .A2(n280), .B1(plus2A[48]), .B2(n277), .ZN(
        n400) );
  AOI22_X1 U14 ( .A1(minus2A[48]), .A2(n291), .B1(minusA[48]), .B2(n285), .ZN(
        n399) );
  NAND2_X1 U15 ( .A1(n382), .A2(n381), .ZN(n458) );
  AOI22_X1 U16 ( .A1(plusA[39]), .A2(n280), .B1(plus2A[39]), .B2(n276), .ZN(
        n382) );
  AOI22_X1 U17 ( .A1(minus2A[39]), .A2(n290), .B1(minusA[39]), .B2(n284), .ZN(
        n381) );
  NAND2_X1 U18 ( .A1(n384), .A2(n383), .ZN(n457) );
  AOI22_X1 U19 ( .A1(plusA[40]), .A2(n280), .B1(plus2A[40]), .B2(n276), .ZN(
        n384) );
  AOI22_X1 U20 ( .A1(minus2A[40]), .A2(n290), .B1(minusA[40]), .B2(n284), .ZN(
        n383) );
  NAND2_X1 U21 ( .A1(n380), .A2(n379), .ZN(n459) );
  AOI22_X1 U22 ( .A1(plusA[38]), .A2(n280), .B1(plus2A[38]), .B2(n276), .ZN(
        n380) );
  AOI22_X1 U23 ( .A1(minus2A[38]), .A2(n290), .B1(minusA[38]), .B2(n284), .ZN(
        n379) );
  NAND2_X1 U24 ( .A1(n422), .A2(n421), .ZN(n438) );
  AOI22_X1 U25 ( .A1(plusA[59]), .A2(n279), .B1(plus2A[59]), .B2(n277), .ZN(
        n422) );
  AOI22_X1 U26 ( .A1(minus2A[59]), .A2(n291), .B1(minusA[59]), .B2(n285), .ZN(
        n421) );
  NAND2_X1 U27 ( .A1(n414), .A2(n413), .ZN(n442) );
  AOI22_X1 U28 ( .A1(plusA[55]), .A2(n279), .B1(plus2A[55]), .B2(n277), .ZN(
        n414) );
  AOI22_X1 U29 ( .A1(minus2A[55]), .A2(n291), .B1(minusA[55]), .B2(n285), .ZN(
        n413) );
  NAND2_X1 U30 ( .A1(n412), .A2(n411), .ZN(n443) );
  AOI22_X1 U31 ( .A1(plusA[54]), .A2(n280), .B1(plus2A[54]), .B2(n277), .ZN(
        n412) );
  AOI22_X1 U32 ( .A1(minus2A[54]), .A2(n291), .B1(minusA[54]), .B2(n285), .ZN(
        n411) );
  NAND2_X1 U33 ( .A1(n410), .A2(n409), .ZN(n444) );
  AOI22_X1 U34 ( .A1(plusA[53]), .A2(n280), .B1(plus2A[53]), .B2(n277), .ZN(
        n410) );
  AOI22_X1 U35 ( .A1(minus2A[53]), .A2(n291), .B1(minusA[53]), .B2(n285), .ZN(
        n409) );
  NAND2_X1 U36 ( .A1(n402), .A2(n401), .ZN(n448) );
  AOI22_X1 U37 ( .A1(plusA[49]), .A2(n280), .B1(plus2A[49]), .B2(n277), .ZN(
        n402) );
  AOI22_X1 U38 ( .A1(minus2A[49]), .A2(n291), .B1(minusA[49]), .B2(n285), .ZN(
        n401) );
  NAND2_X1 U39 ( .A1(n404), .A2(n403), .ZN(n447) );
  AOI22_X1 U40 ( .A1(plusA[50]), .A2(n280), .B1(plus2A[50]), .B2(n277), .ZN(
        n404) );
  AOI22_X1 U41 ( .A1(minus2A[50]), .A2(n291), .B1(minusA[50]), .B2(n285), .ZN(
        n403) );
  NAND2_X1 U42 ( .A1(n420), .A2(n419), .ZN(n439) );
  AOI22_X1 U43 ( .A1(plusA[58]), .A2(n280), .B1(plus2A[58]), .B2(n277), .ZN(
        n420) );
  AOI22_X1 U44 ( .A1(minus2A[58]), .A2(n291), .B1(minusA[58]), .B2(n285), .ZN(
        n419) );
  NAND2_X1 U45 ( .A1(n424), .A2(n423), .ZN(n437) );
  AOI22_X1 U46 ( .A1(plusA[60]), .A2(n280), .B1(plus2A[60]), .B2(n278), .ZN(
        n424) );
  AOI22_X1 U47 ( .A1(minus2A[60]), .A2(n292), .B1(minusA[60]), .B2(n286), .ZN(
        n423) );
  BUF_X1 U48 ( .A(n272), .Z(n279) );
  BUF_X1 U49 ( .A(n429), .Z(n273) );
  BUF_X1 U50 ( .A(n429), .Z(n274) );
  BUF_X1 U51 ( .A(n431), .Z(n287) );
  BUF_X1 U52 ( .A(n431), .Z(n288) );
  BUF_X1 U53 ( .A(n430), .Z(n281) );
  BUF_X1 U54 ( .A(n430), .Z(n282) );
  BUF_X1 U55 ( .A(n489), .Z(n294) );
  BUF_X1 U56 ( .A(n489), .Z(n293) );
  BUF_X1 U57 ( .A(n489), .Z(n295) );
  NAND2_X1 U58 ( .A1(n398), .A2(n397), .ZN(n450) );
  AOI22_X1 U59 ( .A1(plusA[47]), .A2(n280), .B1(plus2A[47]), .B2(n276), .ZN(
        n398) );
  AOI22_X1 U60 ( .A1(minus2A[47]), .A2(n290), .B1(minusA[47]), .B2(n284), .ZN(
        n397) );
  NAND2_X1 U61 ( .A1(n388), .A2(n387), .ZN(n455) );
  AOI22_X1 U62 ( .A1(plusA[42]), .A2(n280), .B1(plus2A[42]), .B2(n276), .ZN(
        n388) );
  AOI22_X1 U63 ( .A1(minus2A[42]), .A2(n290), .B1(minusA[42]), .B2(n284), .ZN(
        n387) );
  NAND2_X1 U64 ( .A1(n378), .A2(n377), .ZN(n460) );
  AOI22_X1 U65 ( .A1(plusA[37]), .A2(n280), .B1(plus2A[37]), .B2(n276), .ZN(
        n378) );
  AOI22_X1 U66 ( .A1(minus2A[37]), .A2(n290), .B1(minusA[37]), .B2(n284), .ZN(
        n377) );
  NAND2_X1 U67 ( .A1(n396), .A2(n395), .ZN(n451) );
  AOI22_X1 U68 ( .A1(plusA[46]), .A2(n280), .B1(plus2A[46]), .B2(n276), .ZN(
        n396) );
  AOI22_X1 U69 ( .A1(minus2A[46]), .A2(n290), .B1(minusA[46]), .B2(n284), .ZN(
        n395) );
  NAND2_X1 U70 ( .A1(n386), .A2(n385), .ZN(n456) );
  AOI22_X1 U71 ( .A1(plusA[41]), .A2(n280), .B1(plus2A[41]), .B2(n276), .ZN(
        n386) );
  AOI22_X1 U72 ( .A1(minus2A[41]), .A2(n290), .B1(minusA[41]), .B2(n284), .ZN(
        n385) );
  NAND2_X1 U73 ( .A1(n376), .A2(n375), .ZN(n461) );
  AOI22_X1 U74 ( .A1(plusA[36]), .A2(n280), .B1(plus2A[36]), .B2(n276), .ZN(
        n376) );
  AOI22_X1 U75 ( .A1(minus2A[36]), .A2(n290), .B1(minusA[36]), .B2(n284), .ZN(
        n375) );
  NAND2_X1 U76 ( .A1(n374), .A2(n373), .ZN(n462) );
  AOI22_X1 U77 ( .A1(plusA[35]), .A2(n280), .B1(plus2A[35]), .B2(n275), .ZN(
        n374) );
  AOI22_X1 U78 ( .A1(minus2A[35]), .A2(n289), .B1(minusA[35]), .B2(n283), .ZN(
        n373) );
  NAND2_X1 U79 ( .A1(n372), .A2(n371), .ZN(n463) );
  AOI22_X1 U80 ( .A1(plusA[34]), .A2(n280), .B1(plus2A[34]), .B2(n275), .ZN(
        n372) );
  AOI22_X1 U81 ( .A1(minus2A[34]), .A2(n289), .B1(minusA[34]), .B2(n283), .ZN(
        n371) );
  BUF_X1 U82 ( .A(n429), .Z(n275) );
  BUF_X1 U83 ( .A(n431), .Z(n289) );
  BUF_X1 U84 ( .A(n430), .Z(n283) );
  NAND2_X1 U85 ( .A1(n433), .A2(n432), .ZN(n434) );
  AOI22_X1 U86 ( .A1(plusA[63]), .A2(n280), .B1(plus2A[63]), .B2(n278), .ZN(
        n433) );
  AOI22_X1 U87 ( .A1(minus2A[63]), .A2(n292), .B1(minusA[63]), .B2(n286), .ZN(
        n432) );
  NAND2_X1 U88 ( .A1(n408), .A2(n407), .ZN(n445) );
  AOI22_X1 U89 ( .A1(plusA[52]), .A2(n280), .B1(plus2A[52]), .B2(n277), .ZN(
        n408) );
  AOI22_X1 U90 ( .A1(minus2A[52]), .A2(n291), .B1(minusA[52]), .B2(n285), .ZN(
        n407) );
  NAND2_X1 U91 ( .A1(n428), .A2(n427), .ZN(n435) );
  AOI22_X1 U92 ( .A1(plusA[62]), .A2(n279), .B1(plus2A[62]), .B2(n278), .ZN(
        n428) );
  AOI22_X1 U93 ( .A1(minus2A[62]), .A2(n292), .B1(minusA[62]), .B2(n286), .ZN(
        n427) );
  NAND2_X1 U94 ( .A1(n418), .A2(n417), .ZN(n440) );
  AOI22_X1 U95 ( .A1(plusA[57]), .A2(n279), .B1(plus2A[57]), .B2(n277), .ZN(
        n418) );
  AOI22_X1 U96 ( .A1(minus2A[57]), .A2(n291), .B1(minusA[57]), .B2(n285), .ZN(
        n417) );
  NAND2_X1 U97 ( .A1(n406), .A2(n405), .ZN(n446) );
  AOI22_X1 U98 ( .A1(plusA[51]), .A2(n280), .B1(plus2A[51]), .B2(n277), .ZN(
        n406) );
  AOI22_X1 U99 ( .A1(minus2A[51]), .A2(n291), .B1(minusA[51]), .B2(n285), .ZN(
        n405) );
  NAND2_X1 U100 ( .A1(n426), .A2(n425), .ZN(n436) );
  AOI22_X1 U101 ( .A1(plusA[61]), .A2(n280), .B1(plus2A[61]), .B2(n278), .ZN(
        n426) );
  AOI22_X1 U102 ( .A1(minus2A[61]), .A2(n292), .B1(minusA[61]), .B2(n286), 
        .ZN(n425) );
  NAND2_X1 U103 ( .A1(n416), .A2(n415), .ZN(n441) );
  AOI22_X1 U104 ( .A1(plusA[56]), .A2(n280), .B1(plus2A[56]), .B2(n277), .ZN(
        n416) );
  AOI22_X1 U105 ( .A1(minus2A[56]), .A2(n291), .B1(minusA[56]), .B2(n285), 
        .ZN(n415) );
  BUF_X1 U106 ( .A(n429), .Z(n276) );
  BUF_X1 U107 ( .A(n431), .Z(n290) );
  BUF_X1 U108 ( .A(n430), .Z(n284) );
  BUF_X1 U109 ( .A(n489), .Z(n296) );
  BUF_X1 U110 ( .A(n429), .Z(n277) );
  BUF_X1 U111 ( .A(n431), .Z(n291) );
  BUF_X1 U112 ( .A(n430), .Z(n285) );
  BUF_X1 U113 ( .A(n489), .Z(n297) );
  BUF_X1 U114 ( .A(n489), .Z(n298) );
  NOR3_X1 U115 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n299), .ZN(n430) );
  NOR2_X1 U116 ( .A1(n320), .A2(n301), .ZN(n489) );
  NAND2_X1 U117 ( .A1(n350), .A2(n349), .ZN(n474) );
  AOI22_X1 U118 ( .A1(plusA[23]), .A2(n279), .B1(plus2A[23]), .B2(n274), .ZN(
        n350) );
  AOI22_X1 U119 ( .A1(minus2A[23]), .A2(n288), .B1(minusA[23]), .B2(n282), 
        .ZN(n349) );
  NAND2_X1 U120 ( .A1(n348), .A2(n347), .ZN(n475) );
  AOI22_X1 U121 ( .A1(plusA[22]), .A2(n279), .B1(plus2A[22]), .B2(n274), .ZN(
        n348) );
  AOI22_X1 U122 ( .A1(minus2A[22]), .A2(n288), .B1(minusA[22]), .B2(n282), 
        .ZN(n347) );
  NAND2_X1 U123 ( .A1(n346), .A2(n345), .ZN(n476) );
  AOI22_X1 U124 ( .A1(plusA[21]), .A2(n279), .B1(plus2A[21]), .B2(n274), .ZN(
        n346) );
  AOI22_X1 U125 ( .A1(minus2A[21]), .A2(n288), .B1(minusA[21]), .B2(n282), 
        .ZN(n345) );
  NAND2_X1 U126 ( .A1(n342), .A2(n341), .ZN(n478) );
  AOI22_X1 U127 ( .A1(plusA[19]), .A2(n279), .B1(plus2A[19]), .B2(n274), .ZN(
        n342) );
  AOI22_X1 U128 ( .A1(minus2A[19]), .A2(n288), .B1(minusA[19]), .B2(n282), 
        .ZN(n341) );
  NAND2_X1 U129 ( .A1(n340), .A2(n339), .ZN(n479) );
  AOI22_X1 U130 ( .A1(plusA[18]), .A2(n279), .B1(plus2A[18]), .B2(n274), .ZN(
        n340) );
  AOI22_X1 U131 ( .A1(minus2A[18]), .A2(n288), .B1(minusA[18]), .B2(n282), 
        .ZN(n339) );
  NAND2_X1 U132 ( .A1(n338), .A2(n337), .ZN(n480) );
  AOI22_X1 U133 ( .A1(plusA[17]), .A2(n279), .B1(plus2A[17]), .B2(n274), .ZN(
        n338) );
  AOI22_X1 U134 ( .A1(minus2A[17]), .A2(n288), .B1(minusA[17]), .B2(n282), 
        .ZN(n337) );
  NOR3_X1 U135 ( .A1(SEL[1]), .A2(SEL[2]), .A3(n300), .ZN(n272) );
  INV_X1 U136 ( .A(SEL[1]), .ZN(n299) );
  NAND2_X1 U137 ( .A1(n334), .A2(n333), .ZN(n482) );
  AOI22_X1 U138 ( .A1(plusA[15]), .A2(n279), .B1(plus2A[15]), .B2(n274), .ZN(
        n334) );
  AOI22_X1 U139 ( .A1(minus2A[15]), .A2(n288), .B1(minusA[15]), .B2(n282), 
        .ZN(n333) );
  NAND2_X1 U140 ( .A1(n311), .A2(n310), .ZN(n494) );
  AOI22_X1 U141 ( .A1(minus2A[4]), .A2(n287), .B1(minusA[4]), .B2(n281), .ZN(
        n310) );
  AOI22_X1 U142 ( .A1(plusA[4]), .A2(n279), .B1(plus2A[4]), .B2(n273), .ZN(
        n311) );
  NAND2_X1 U143 ( .A1(n344), .A2(n343), .ZN(n477) );
  AOI22_X1 U144 ( .A1(plusA[20]), .A2(n279), .B1(plus2A[20]), .B2(n274), .ZN(
        n344) );
  AOI22_X1 U145 ( .A1(minus2A[20]), .A2(n288), .B1(minusA[20]), .B2(n282), 
        .ZN(n343) );
  NAND2_X1 U146 ( .A1(n336), .A2(n335), .ZN(n481) );
  AOI22_X1 U147 ( .A1(plusA[16]), .A2(n279), .B1(plus2A[16]), .B2(n274), .ZN(
        n336) );
  AOI22_X1 U148 ( .A1(minus2A[16]), .A2(n288), .B1(minusA[16]), .B2(n282), 
        .ZN(n335) );
  NAND2_X1 U149 ( .A1(n332), .A2(n331), .ZN(n483) );
  AOI22_X1 U150 ( .A1(plusA[14]), .A2(n279), .B1(plus2A[14]), .B2(n274), .ZN(
        n332) );
  AOI22_X1 U151 ( .A1(minus2A[14]), .A2(n288), .B1(minusA[14]), .B2(n282), 
        .ZN(n331) );
  NAND2_X1 U152 ( .A1(n330), .A2(n329), .ZN(n484) );
  AOI22_X1 U153 ( .A1(plusA[13]), .A2(n279), .B1(plus2A[13]), .B2(n274), .ZN(
        n330) );
  AOI22_X1 U154 ( .A1(minus2A[13]), .A2(n288), .B1(minusA[13]), .B2(n282), 
        .ZN(n329) );
  NAND2_X1 U155 ( .A1(n328), .A2(n327), .ZN(n485) );
  AOI22_X1 U156 ( .A1(plusA[12]), .A2(n279), .B1(plus2A[12]), .B2(n274), .ZN(
        n328) );
  AOI22_X1 U157 ( .A1(minus2A[12]), .A2(n288), .B1(minusA[12]), .B2(n282), 
        .ZN(n327) );
  NAND2_X1 U158 ( .A1(n319), .A2(n318), .ZN(n490) );
  AOI22_X1 U159 ( .A1(plusA[8]), .A2(n280), .B1(plus2A[8]), .B2(n273), .ZN(
        n319) );
  AOI22_X1 U160 ( .A1(minus2A[8]), .A2(n287), .B1(minusA[8]), .B2(n281), .ZN(
        n318) );
  NAND2_X1 U161 ( .A1(n324), .A2(n323), .ZN(n487) );
  AOI22_X1 U162 ( .A1(plusA[10]), .A2(n280), .B1(plus2A[10]), .B2(n273), .ZN(
        n324) );
  AOI22_X1 U163 ( .A1(minus2A[10]), .A2(n287), .B1(minusA[10]), .B2(n281), 
        .ZN(n323) );
  NAND2_X1 U164 ( .A1(n315), .A2(n314), .ZN(n492) );
  AOI22_X1 U165 ( .A1(minus2A[6]), .A2(n287), .B1(minusA[6]), .B2(n281), .ZN(
        n314) );
  AOI22_X1 U166 ( .A1(plusA[6]), .A2(n280), .B1(plus2A[6]), .B2(n273), .ZN(
        n315) );
  NAND2_X1 U167 ( .A1(n309), .A2(n308), .ZN(n495) );
  AOI22_X1 U168 ( .A1(minus2A[3]), .A2(n287), .B1(minusA[3]), .B2(n281), .ZN(
        n308) );
  AOI22_X1 U169 ( .A1(plusA[3]), .A2(n272), .B1(plus2A[3]), .B2(n273), .ZN(
        n309) );
  NAND2_X1 U170 ( .A1(n313), .A2(n312), .ZN(n493) );
  AOI22_X1 U171 ( .A1(minus2A[5]), .A2(n287), .B1(minusA[5]), .B2(n281), .ZN(
        n312) );
  AOI22_X1 U172 ( .A1(plusA[5]), .A2(n280), .B1(plus2A[5]), .B2(n273), .ZN(
        n313) );
  NAND2_X1 U173 ( .A1(n322), .A2(n321), .ZN(n488) );
  AOI22_X1 U174 ( .A1(plusA[9]), .A2(n280), .B1(plus2A[9]), .B2(n273), .ZN(
        n322) );
  AOI22_X1 U175 ( .A1(minus2A[9]), .A2(n287), .B1(minusA[9]), .B2(n281), .ZN(
        n321) );
  NAND2_X1 U176 ( .A1(n326), .A2(n325), .ZN(n486) );
  AOI22_X1 U177 ( .A1(plusA[11]), .A2(n280), .B1(plus2A[11]), .B2(n273), .ZN(
        n326) );
  AOI22_X1 U178 ( .A1(minus2A[11]), .A2(n287), .B1(minusA[11]), .B2(n281), 
        .ZN(n325) );
  NAND2_X1 U179 ( .A1(n317), .A2(n316), .ZN(n491) );
  AOI22_X1 U180 ( .A1(plusA[7]), .A2(n280), .B1(plus2A[7]), .B2(n273), .ZN(
        n317) );
  AOI22_X1 U181 ( .A1(minus2A[7]), .A2(n287), .B1(minusA[7]), .B2(n281), .ZN(
        n316) );
  NAND2_X1 U182 ( .A1(n362), .A2(n361), .ZN(n468) );
  AOI22_X1 U183 ( .A1(plusA[29]), .A2(n280), .B1(plus2A[29]), .B2(n275), .ZN(
        n362) );
  AOI22_X1 U184 ( .A1(minus2A[29]), .A2(n289), .B1(minusA[29]), .B2(n283), 
        .ZN(n361) );
  NAND2_X1 U185 ( .A1(n358), .A2(n357), .ZN(n470) );
  AOI22_X1 U186 ( .A1(plusA[27]), .A2(n280), .B1(plus2A[27]), .B2(n275), .ZN(
        n358) );
  AOI22_X1 U187 ( .A1(minus2A[27]), .A2(n289), .B1(minusA[27]), .B2(n283), 
        .ZN(n357) );
  NAND2_X1 U188 ( .A1(n356), .A2(n355), .ZN(n471) );
  AOI22_X1 U189 ( .A1(plusA[26]), .A2(n280), .B1(plus2A[26]), .B2(n275), .ZN(
        n356) );
  AOI22_X1 U190 ( .A1(minus2A[26]), .A2(n289), .B1(minusA[26]), .B2(n283), 
        .ZN(n355) );
  NAND2_X1 U191 ( .A1(n354), .A2(n353), .ZN(n472) );
  AOI22_X1 U192 ( .A1(plusA[25]), .A2(n280), .B1(plus2A[25]), .B2(n275), .ZN(
        n354) );
  AOI22_X1 U193 ( .A1(minus2A[25]), .A2(n289), .B1(minusA[25]), .B2(n283), 
        .ZN(n353) );
  NAND2_X1 U194 ( .A1(n368), .A2(n367), .ZN(n465) );
  AOI22_X1 U195 ( .A1(plusA[32]), .A2(n280), .B1(plus2A[32]), .B2(n275), .ZN(
        n368) );
  AOI22_X1 U196 ( .A1(minus2A[32]), .A2(n289), .B1(minusA[32]), .B2(n283), 
        .ZN(n367) );
  NAND2_X1 U197 ( .A1(n360), .A2(n359), .ZN(n469) );
  AOI22_X1 U198 ( .A1(plusA[28]), .A2(n280), .B1(plus2A[28]), .B2(n275), .ZN(
        n360) );
  AOI22_X1 U199 ( .A1(minus2A[28]), .A2(n289), .B1(minusA[28]), .B2(n283), 
        .ZN(n359) );
  NAND2_X1 U200 ( .A1(n352), .A2(n351), .ZN(n473) );
  AOI22_X1 U201 ( .A1(plusA[24]), .A2(n280), .B1(plus2A[24]), .B2(n275), .ZN(
        n352) );
  AOI22_X1 U202 ( .A1(minus2A[24]), .A2(n289), .B1(minusA[24]), .B2(n283), 
        .ZN(n351) );
  NAND2_X1 U203 ( .A1(n370), .A2(n369), .ZN(n464) );
  AOI22_X1 U204 ( .A1(plusA[33]), .A2(n280), .B1(plus2A[33]), .B2(n275), .ZN(
        n370) );
  AOI22_X1 U205 ( .A1(minus2A[33]), .A2(n289), .B1(minusA[33]), .B2(n283), 
        .ZN(n369) );
  NAND2_X1 U206 ( .A1(n364), .A2(n363), .ZN(n467) );
  AOI22_X1 U207 ( .A1(plusA[30]), .A2(n280), .B1(plus2A[30]), .B2(n275), .ZN(
        n364) );
  AOI22_X1 U208 ( .A1(minus2A[30]), .A2(n289), .B1(minusA[30]), .B2(n283), 
        .ZN(n363) );
  NAND2_X1 U209 ( .A1(n366), .A2(n365), .ZN(n466) );
  AOI22_X1 U210 ( .A1(plusA[31]), .A2(n280), .B1(plus2A[31]), .B2(n275), .ZN(
        n366) );
  AOI22_X1 U211 ( .A1(minus2A[31]), .A2(n289), .B1(minusA[31]), .B2(n283), 
        .ZN(n365) );
  NAND2_X1 U212 ( .A1(n307), .A2(n306), .ZN(n496) );
  AOI22_X1 U213 ( .A1(plusA[2]), .A2(n272), .B1(plus2A[2]), .B2(n273), .ZN(
        n307) );
  AOI22_X1 U214 ( .A1(minus2A[2]), .A2(n287), .B1(minusA[2]), .B2(n281), .ZN(
        n306) );
  AOI22_X1 U215 ( .A1(plusA[1]), .A2(n279), .B1(plus2A[1]), .B2(n273), .ZN(
        n305) );
  AOI22_X1 U216 ( .A1(minus2A[1]), .A2(n287), .B1(minusA[1]), .B2(n281), .ZN(
        n304) );
  AOI22_X1 U217 ( .A1(plusA[0]), .A2(n280), .B1(plus2A[0]), .B2(n273), .ZN(
        n303) );
  AOI22_X1 U218 ( .A1(minus2A[0]), .A2(n287), .B1(minusA[0]), .B2(n281), .ZN(
        n302) );
  NAND2_X1 U219 ( .A1(n305), .A2(n304), .ZN(n497) );
  INV_X1 U220 ( .A(SEL[0]), .ZN(n300) );
  NOR2_X1 U221 ( .A1(SEL[1]), .A2(SEL[0]), .ZN(n320) );
  AND2_X1 U222 ( .A1(SEL[2]), .A2(n320), .ZN(n431) );
  NOR3_X1 U223 ( .A1(n299), .A2(SEL[2]), .A3(n300), .ZN(n429) );
  INV_X1 U224 ( .A(SEL[2]), .ZN(n301) );
  NAND2_X1 U225 ( .A1(n303), .A2(n302), .ZN(n498) );
  CLKBUF_X1 U226 ( .A(n429), .Z(n278) );
  CLKBUF_X1 U227 ( .A(n430), .Z(n286) );
  CLKBUF_X1 U228 ( .A(n431), .Z(n292) );
endmodule


module FA_0 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;
  tri   A;
  tri   B;

  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  XOR2_X1 U1 ( .A(Ci), .B(n3), .Z(S) );
  INV_X1 U2 ( .A(n2), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n2) );
endmodule


module FA_959 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_958 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_957 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_956 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_955 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_954 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_953 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_952 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_951 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_950 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_949 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_948 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_947 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_946 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_945 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  XOR2_X1 U1 ( .A(Ci), .B(n5), .Z(S) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U3 ( .A(n6), .ZN(Co) );
endmodule


module FA_944 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_943 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_942 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_941 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_940 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_939 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_938 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_937 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_936 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_935 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_934 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_933 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_932 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_931 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_930 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_929 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_928 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_927 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_926 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_925 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_924 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_923 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_922 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_921 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_920 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_919 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_918 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_917 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_916 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_915 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_914 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_913 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_912 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_911 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_910 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_909 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_908 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_907 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_906 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_905 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_904 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_903 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_902 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_901 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_900 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_899 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_898 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_897 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;
  tri   B;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N64_0 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Ci;
  output Co;

  wire   [63:1] CTMP;
  tri   [63:0] A;
  tri   [63:0] B;

  FA_0 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_959 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_958 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_957 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(CTMP[4]) );
  FA_956 FAI_5 ( .A(A[4]), .B(B[4]), .Ci(CTMP[4]), .S(S[4]), .Co(CTMP[5]) );
  FA_955 FAI_6 ( .A(A[5]), .B(B[5]), .Ci(CTMP[5]), .S(S[5]), .Co(CTMP[6]) );
  FA_954 FAI_7 ( .A(A[6]), .B(B[6]), .Ci(CTMP[6]), .S(S[6]), .Co(CTMP[7]) );
  FA_953 FAI_8 ( .A(A[7]), .B(B[7]), .Ci(CTMP[7]), .S(S[7]), .Co(CTMP[8]) );
  FA_952 FAI_9 ( .A(A[8]), .B(B[8]), .Ci(CTMP[8]), .S(S[8]), .Co(CTMP[9]) );
  FA_951 FAI_10 ( .A(A[9]), .B(B[9]), .Ci(CTMP[9]), .S(S[9]), .Co(CTMP[10]) );
  FA_950 FAI_11 ( .A(A[10]), .B(B[10]), .Ci(CTMP[10]), .S(S[10]), .Co(CTMP[11]) );
  FA_949 FAI_12 ( .A(A[11]), .B(B[11]), .Ci(CTMP[11]), .S(S[11]), .Co(CTMP[12]) );
  FA_948 FAI_13 ( .A(A[12]), .B(B[12]), .Ci(CTMP[12]), .S(S[12]), .Co(CTMP[13]) );
  FA_947 FAI_14 ( .A(A[13]), .B(B[13]), .Ci(CTMP[13]), .S(S[13]), .Co(CTMP[14]) );
  FA_946 FAI_15 ( .A(A[14]), .B(B[14]), .Ci(CTMP[14]), .S(S[14]), .Co(CTMP[15]) );
  FA_945 FAI_16 ( .A(A[15]), .B(B[15]), .Ci(CTMP[15]), .S(S[15]), .Co(CTMP[16]) );
  FA_944 FAI_17 ( .A(A[16]), .B(B[16]), .Ci(CTMP[16]), .S(S[16]), .Co(CTMP[17]) );
  FA_943 FAI_18 ( .A(A[17]), .B(B[17]), .Ci(CTMP[17]), .S(S[17]), .Co(CTMP[18]) );
  FA_942 FAI_19 ( .A(A[18]), .B(B[18]), .Ci(CTMP[18]), .S(S[18]), .Co(CTMP[19]) );
  FA_941 FAI_20 ( .A(A[19]), .B(B[19]), .Ci(CTMP[19]), .S(S[19]), .Co(CTMP[20]) );
  FA_940 FAI_21 ( .A(A[20]), .B(B[20]), .Ci(CTMP[20]), .S(S[20]), .Co(CTMP[21]) );
  FA_939 FAI_22 ( .A(A[21]), .B(B[21]), .Ci(CTMP[21]), .S(S[21]), .Co(CTMP[22]) );
  FA_938 FAI_23 ( .A(A[22]), .B(B[22]), .Ci(CTMP[22]), .S(S[22]), .Co(CTMP[23]) );
  FA_937 FAI_24 ( .A(A[23]), .B(B[23]), .Ci(CTMP[23]), .S(S[23]), .Co(CTMP[24]) );
  FA_936 FAI_25 ( .A(A[24]), .B(B[24]), .Ci(CTMP[24]), .S(S[24]), .Co(CTMP[25]) );
  FA_935 FAI_26 ( .A(A[25]), .B(B[25]), .Ci(CTMP[25]), .S(S[25]), .Co(CTMP[26]) );
  FA_934 FAI_27 ( .A(A[26]), .B(B[26]), .Ci(CTMP[26]), .S(S[26]), .Co(CTMP[27]) );
  FA_933 FAI_28 ( .A(A[27]), .B(B[27]), .Ci(CTMP[27]), .S(S[27]), .Co(CTMP[28]) );
  FA_932 FAI_29 ( .A(A[28]), .B(B[28]), .Ci(CTMP[28]), .S(S[28]), .Co(CTMP[29]) );
  FA_931 FAI_30 ( .A(A[29]), .B(B[29]), .Ci(CTMP[29]), .S(S[29]), .Co(CTMP[30]) );
  FA_930 FAI_31 ( .A(A[30]), .B(B[30]), .Ci(CTMP[30]), .S(S[30]), .Co(CTMP[31]) );
  FA_929 FAI_32 ( .A(A[31]), .B(B[31]), .Ci(CTMP[31]), .S(S[31]), .Co(CTMP[32]) );
  FA_928 FAI_33 ( .A(A[32]), .B(B[32]), .Ci(CTMP[32]), .S(S[32]), .Co(CTMP[33]) );
  FA_927 FAI_34 ( .A(A[33]), .B(B[33]), .Ci(CTMP[33]), .S(S[33]), .Co(CTMP[34]) );
  FA_926 FAI_35 ( .A(A[34]), .B(B[34]), .Ci(CTMP[34]), .S(S[34]), .Co(CTMP[35]) );
  FA_925 FAI_36 ( .A(A[35]), .B(B[35]), .Ci(CTMP[35]), .S(S[35]), .Co(CTMP[36]) );
  FA_924 FAI_37 ( .A(A[36]), .B(B[36]), .Ci(CTMP[36]), .S(S[36]), .Co(CTMP[37]) );
  FA_923 FAI_38 ( .A(A[37]), .B(B[37]), .Ci(CTMP[37]), .S(S[37]), .Co(CTMP[38]) );
  FA_922 FAI_39 ( .A(A[38]), .B(B[38]), .Ci(CTMP[38]), .S(S[38]), .Co(CTMP[39]) );
  FA_921 FAI_40 ( .A(A[39]), .B(B[39]), .Ci(CTMP[39]), .S(S[39]), .Co(CTMP[40]) );
  FA_920 FAI_41 ( .A(A[40]), .B(B[40]), .Ci(CTMP[40]), .S(S[40]), .Co(CTMP[41]) );
  FA_919 FAI_42 ( .A(A[41]), .B(B[41]), .Ci(CTMP[41]), .S(S[41]), .Co(CTMP[42]) );
  FA_918 FAI_43 ( .A(A[42]), .B(B[42]), .Ci(CTMP[42]), .S(S[42]), .Co(CTMP[43]) );
  FA_917 FAI_44 ( .A(A[43]), .B(B[43]), .Ci(CTMP[43]), .S(S[43]), .Co(CTMP[44]) );
  FA_916 FAI_45 ( .A(A[44]), .B(B[44]), .Ci(CTMP[44]), .S(S[44]), .Co(CTMP[45]) );
  FA_915 FAI_46 ( .A(A[45]), .B(B[45]), .Ci(CTMP[45]), .S(S[45]), .Co(CTMP[46]) );
  FA_914 FAI_47 ( .A(A[46]), .B(B[46]), .Ci(CTMP[46]), .S(S[46]), .Co(CTMP[47]) );
  FA_913 FAI_48 ( .A(A[47]), .B(B[47]), .Ci(CTMP[47]), .S(S[47]), .Co(CTMP[48]) );
  FA_912 FAI_49 ( .A(A[48]), .B(B[48]), .Ci(CTMP[48]), .S(S[48]), .Co(CTMP[49]) );
  FA_911 FAI_50 ( .A(A[49]), .B(B[49]), .Ci(CTMP[49]), .S(S[49]), .Co(CTMP[50]) );
  FA_910 FAI_51 ( .A(A[50]), .B(B[50]), .Ci(CTMP[50]), .S(S[50]), .Co(CTMP[51]) );
  FA_909 FAI_52 ( .A(A[51]), .B(B[51]), .Ci(CTMP[51]), .S(S[51]), .Co(CTMP[52]) );
  FA_908 FAI_53 ( .A(A[52]), .B(B[52]), .Ci(CTMP[52]), .S(S[52]), .Co(CTMP[53]) );
  FA_907 FAI_54 ( .A(A[53]), .B(B[53]), .Ci(CTMP[53]), .S(S[53]), .Co(CTMP[54]) );
  FA_906 FAI_55 ( .A(A[54]), .B(B[54]), .Ci(CTMP[54]), .S(S[54]), .Co(CTMP[55]) );
  FA_905 FAI_56 ( .A(A[55]), .B(B[55]), .Ci(CTMP[55]), .S(S[55]), .Co(CTMP[56]) );
  FA_904 FAI_57 ( .A(A[56]), .B(B[56]), .Ci(CTMP[56]), .S(S[56]), .Co(CTMP[57]) );
  FA_903 FAI_58 ( .A(A[57]), .B(B[57]), .Ci(CTMP[57]), .S(S[57]), .Co(CTMP[58]) );
  FA_902 FAI_59 ( .A(A[58]), .B(B[58]), .Ci(CTMP[58]), .S(S[58]), .Co(CTMP[59]) );
  FA_901 FAI_60 ( .A(A[59]), .B(B[59]), .Ci(CTMP[59]), .S(S[59]), .Co(CTMP[60]) );
  FA_900 FAI_61 ( .A(A[60]), .B(B[60]), .Ci(CTMP[60]), .S(S[60]), .Co(CTMP[61]) );
  FA_899 FAI_62 ( .A(A[61]), .B(B[61]), .Ci(CTMP[61]), .S(S[61]), .Co(CTMP[62]) );
  FA_898 FAI_63 ( .A(A[62]), .B(B[62]), .Ci(CTMP[62]), .S(S[62]), .Co(CTMP[63]) );
  FA_897 FAI_64 ( .A(A[63]), .B(B[63]), .Ci(CTMP[63]), .S(S[63]), .Co(Co) );
endmodule


module booth_mul_row_N64_RADIX3_0 ( prevA, prevSum, encoderIn, nextA, nextSum
 );
  input [63:0] prevA;
  input [63:0] prevSum;
  input [2:0] encoderIn;
  output [63:0] nextA;
  output [63:0] nextSum;
  wire   n4, n5;
  wire   [2:0] encoder_to_mux;
  wire   [63:0] plus2A_s;
  wire   [63:0] minus2A_s;
  wire   [63:0] minus4A_s;
  tri   [63:0] prevSum;
  tri   [63:0] mux_to_adder;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign nextA[51] = n4;
  assign nextA[39] = n5;
  assign nextA[0] = 1'b0;

  encoder_N64_RADIX3_15 encoder_1 ( .X(encoderIn), .Z(encoder_to_mux) );
  ShiftnCompl_N64_0 ShiftnCompl_1 ( .plusA(prevA), .plus2A_out({plus2A_s[63:1], 
        SYNOPSYS_UNCONNECTED__0}), .minus2A_out(minus2A_s), .plus4A_out({
        nextA[63:52], n4, nextA[50:40], n5, nextA[38:1], 
        SYNOPSYS_UNCONNECTED__1}), .minus4A_out(minus4A_s) );
  MUX_GENERIC_N64_RADIX3_15 mux_1 ( .plusA({plus2A_s[63:1], 1'b0}), .minusA(
        minus2A_s), .plus2A({nextA[63:52], n4, nextA[50:40], n5, nextA[38:1], 
        1'b0}), .minus2A(minus4A_s), .SEL(encoder_to_mux), .Y(mux_to_adder) );
  RCA_N64_0 rca_1 ( .A(mux_to_adder), .B(prevSum), .Ci(1'b0), .S(nextSum) );
endmodule


module encoder_N64_RADIX3_14 ( X, Z );
  input [2:0] X;
  output [2:0] Z;
  wire   n5, n7, n8;

  OAI22_X1 U1 ( .A1(n8), .A2(n5), .B1(X[2]), .B2(n7), .ZN(Z[1]) );
  INV_X1 U2 ( .A(X[2]), .ZN(n5) );
  AOI21_X1 U3 ( .B1(n8), .B2(n7), .A(X[2]), .ZN(Z[0]) );
  OAI21_X1 U4 ( .B1(X[1]), .B2(X[0]), .A(n7), .ZN(n8) );
  AND3_X1 U5 ( .A1(X[2]), .A2(n7), .A3(n8), .ZN(Z[2]) );
  NAND2_X1 U6 ( .A1(X[1]), .A2(X[0]), .ZN(n7) );
endmodule


module shifter_N64_28 ( \input , shiftLeftOnePos );
  input [63:0] \input ;
  output [63:0] shiftLeftOnePos;
  wire   \input[62] , \input[61] , \input[60] , \input[59] , \input[58] ,
         \input[57] , \input[56] , \input[55] , \input[54] , \input[53] ,
         \input[52] , \input[51] , \input[50] , \input[49] , \input[48] ,
         \input[47] , \input[46] , \input[45] , \input[44] , \input[43] ,
         \input[42] , \input[41] , \input[40] , \input[39] , \input[38] ,
         \input[37] , \input[36] , \input[35] , \input[34] , \input[33] ,
         \input[32] , \input[31] , \input[30] , \input[29] , \input[28] ,
         \input[27] , \input[26] , \input[25] , \input[24] , \input[23] ,
         \input[22] , \input[21] , \input[20] , \input[19] , \input[18] ,
         \input[17] , \input[16] , \input[15] , \input[14] , \input[13] ,
         \input[12] , \input[11] , \input[10] , \input[9] , \input[8] ,
         \input[7] , \input[6] , \input[5] , \input[4] , \input[3] ,
         \input[2] , \input[1] , \input[0] ;
  assign shiftLeftOnePos[0] = 1'b0;
  assign shiftLeftOnePos[63] = \input[62] ;
  assign \input[62]  = \input  [62];
  assign shiftLeftOnePos[62] = \input[61] ;
  assign \input[61]  = \input  [61];
  assign shiftLeftOnePos[61] = \input[60] ;
  assign \input[60]  = \input  [60];
  assign shiftLeftOnePos[60] = \input[59] ;
  assign \input[59]  = \input  [59];
  assign shiftLeftOnePos[59] = \input[58] ;
  assign \input[58]  = \input  [58];
  assign shiftLeftOnePos[58] = \input[57] ;
  assign \input[57]  = \input  [57];
  assign shiftLeftOnePos[57] = \input[56] ;
  assign \input[56]  = \input  [56];
  assign shiftLeftOnePos[56] = \input[55] ;
  assign \input[55]  = \input  [55];
  assign shiftLeftOnePos[55] = \input[54] ;
  assign \input[54]  = \input  [54];
  assign shiftLeftOnePos[54] = \input[53] ;
  assign \input[53]  = \input  [53];
  assign shiftLeftOnePos[53] = \input[52] ;
  assign \input[52]  = \input  [52];
  assign shiftLeftOnePos[52] = \input[51] ;
  assign \input[51]  = \input  [51];
  assign shiftLeftOnePos[51] = \input[50] ;
  assign \input[50]  = \input  [50];
  assign shiftLeftOnePos[50] = \input[49] ;
  assign \input[49]  = \input  [49];
  assign shiftLeftOnePos[49] = \input[48] ;
  assign \input[48]  = \input  [48];
  assign shiftLeftOnePos[48] = \input[47] ;
  assign \input[47]  = \input  [47];
  assign shiftLeftOnePos[47] = \input[46] ;
  assign \input[46]  = \input  [46];
  assign shiftLeftOnePos[46] = \input[45] ;
  assign \input[45]  = \input  [45];
  assign shiftLeftOnePos[45] = \input[44] ;
  assign \input[44]  = \input  [44];
  assign shiftLeftOnePos[44] = \input[43] ;
  assign \input[43]  = \input  [43];
  assign shiftLeftOnePos[43] = \input[42] ;
  assign \input[42]  = \input  [42];
  assign shiftLeftOnePos[42] = \input[41] ;
  assign \input[41]  = \input  [41];
  assign shiftLeftOnePos[41] = \input[40] ;
  assign \input[40]  = \input  [40];
  assign shiftLeftOnePos[40] = \input[39] ;
  assign \input[39]  = \input  [39];
  assign shiftLeftOnePos[39] = \input[38] ;
  assign \input[38]  = \input  [38];
  assign shiftLeftOnePos[38] = \input[37] ;
  assign \input[37]  = \input  [37];
  assign shiftLeftOnePos[37] = \input[36] ;
  assign \input[36]  = \input  [36];
  assign shiftLeftOnePos[36] = \input[35] ;
  assign \input[35]  = \input  [35];
  assign shiftLeftOnePos[35] = \input[34] ;
  assign \input[34]  = \input  [34];
  assign shiftLeftOnePos[34] = \input[33] ;
  assign \input[33]  = \input  [33];
  assign shiftLeftOnePos[33] = \input[32] ;
  assign \input[32]  = \input  [32];
  assign shiftLeftOnePos[32] = \input[31] ;
  assign \input[31]  = \input  [31];
  assign shiftLeftOnePos[31] = \input[30] ;
  assign \input[30]  = \input  [30];
  assign shiftLeftOnePos[30] = \input[29] ;
  assign \input[29]  = \input  [29];
  assign shiftLeftOnePos[29] = \input[28] ;
  assign \input[28]  = \input  [28];
  assign shiftLeftOnePos[28] = \input[27] ;
  assign \input[27]  = \input  [27];
  assign shiftLeftOnePos[27] = \input[26] ;
  assign \input[26]  = \input  [26];
  assign shiftLeftOnePos[26] = \input[25] ;
  assign \input[25]  = \input  [25];
  assign shiftLeftOnePos[25] = \input[24] ;
  assign \input[24]  = \input  [24];
  assign shiftLeftOnePos[24] = \input[23] ;
  assign \input[23]  = \input  [23];
  assign shiftLeftOnePos[23] = \input[22] ;
  assign \input[22]  = \input  [22];
  assign shiftLeftOnePos[22] = \input[21] ;
  assign \input[21]  = \input  [21];
  assign shiftLeftOnePos[21] = \input[20] ;
  assign \input[20]  = \input  [20];
  assign shiftLeftOnePos[20] = \input[19] ;
  assign \input[19]  = \input  [19];
  assign shiftLeftOnePos[19] = \input[18] ;
  assign \input[18]  = \input  [18];
  assign shiftLeftOnePos[18] = \input[17] ;
  assign \input[17]  = \input  [17];
  assign shiftLeftOnePos[17] = \input[16] ;
  assign \input[16]  = \input  [16];
  assign shiftLeftOnePos[16] = \input[15] ;
  assign \input[15]  = \input  [15];
  assign shiftLeftOnePos[15] = \input[14] ;
  assign \input[14]  = \input  [14];
  assign shiftLeftOnePos[14] = \input[13] ;
  assign \input[13]  = \input  [13];
  assign shiftLeftOnePos[13] = \input[12] ;
  assign \input[12]  = \input  [12];
  assign shiftLeftOnePos[12] = \input[11] ;
  assign \input[11]  = \input  [11];
  assign shiftLeftOnePos[11] = \input[10] ;
  assign \input[10]  = \input  [10];
  assign shiftLeftOnePos[10] = \input[9] ;
  assign \input[9]  = \input  [9];
  assign shiftLeftOnePos[9] = \input[8] ;
  assign \input[8]  = \input  [8];
  assign shiftLeftOnePos[8] = \input[7] ;
  assign \input[7]  = \input  [7];
  assign shiftLeftOnePos[7] = \input[6] ;
  assign \input[6]  = \input  [6];
  assign shiftLeftOnePos[6] = \input[5] ;
  assign \input[5]  = \input  [5];
  assign shiftLeftOnePos[5] = \input[4] ;
  assign \input[4]  = \input  [4];
  assign shiftLeftOnePos[4] = \input[3] ;
  assign \input[3]  = \input  [3];
  assign shiftLeftOnePos[3] = \input[2] ;
  assign \input[2]  = \input  [2];
  assign shiftLeftOnePos[2] = \input[1] ;
  assign \input[1]  = \input  [1];
  assign shiftLeftOnePos[1] = \input[0] ;
  assign \input[0]  = \input  [0];

endmodule


module shifter_N64_27 ( \input , shiftLeftOnePos );
  input [63:0] \input ;
  output [63:0] shiftLeftOnePos;
  wire   \input[62] , \input[61] , \input[60] , \input[59] , \input[58] ,
         \input[57] , \input[56] , \input[55] , \input[54] , \input[53] ,
         \input[52] , \input[51] , \input[50] , \input[49] , \input[48] ,
         \input[47] , \input[46] , \input[45] , \input[44] , \input[43] ,
         \input[42] , \input[41] , \input[40] , \input[39] , \input[38] ,
         \input[37] , \input[36] , \input[35] , \input[34] , \input[33] ,
         \input[32] , \input[31] , \input[30] , \input[29] , \input[28] ,
         \input[27] , \input[26] , \input[25] , \input[24] , \input[23] ,
         \input[22] , \input[21] , \input[20] , \input[19] , \input[18] ,
         \input[17] , \input[16] , \input[15] , \input[14] , \input[13] ,
         \input[12] , \input[11] , \input[10] , \input[9] , \input[8] ,
         \input[7] , \input[6] , \input[5] , \input[4] , \input[3] ,
         \input[2] , \input[1] , \input[0] ;
  assign shiftLeftOnePos[0] = 1'b0;
  assign shiftLeftOnePos[63] = \input[62] ;
  assign \input[62]  = \input  [62];
  assign shiftLeftOnePos[62] = \input[61] ;
  assign \input[61]  = \input  [61];
  assign shiftLeftOnePos[61] = \input[60] ;
  assign \input[60]  = \input  [60];
  assign shiftLeftOnePos[60] = \input[59] ;
  assign \input[59]  = \input  [59];
  assign shiftLeftOnePos[59] = \input[58] ;
  assign \input[58]  = \input  [58];
  assign shiftLeftOnePos[58] = \input[57] ;
  assign \input[57]  = \input  [57];
  assign shiftLeftOnePos[57] = \input[56] ;
  assign \input[56]  = \input  [56];
  assign shiftLeftOnePos[56] = \input[55] ;
  assign \input[55]  = \input  [55];
  assign shiftLeftOnePos[55] = \input[54] ;
  assign \input[54]  = \input  [54];
  assign shiftLeftOnePos[54] = \input[53] ;
  assign \input[53]  = \input  [53];
  assign shiftLeftOnePos[53] = \input[52] ;
  assign \input[52]  = \input  [52];
  assign shiftLeftOnePos[52] = \input[51] ;
  assign \input[51]  = \input  [51];
  assign shiftLeftOnePos[51] = \input[50] ;
  assign \input[50]  = \input  [50];
  assign shiftLeftOnePos[50] = \input[49] ;
  assign \input[49]  = \input  [49];
  assign shiftLeftOnePos[49] = \input[48] ;
  assign \input[48]  = \input  [48];
  assign shiftLeftOnePos[48] = \input[47] ;
  assign \input[47]  = \input  [47];
  assign shiftLeftOnePos[47] = \input[46] ;
  assign \input[46]  = \input  [46];
  assign shiftLeftOnePos[46] = \input[45] ;
  assign \input[45]  = \input  [45];
  assign shiftLeftOnePos[45] = \input[44] ;
  assign \input[44]  = \input  [44];
  assign shiftLeftOnePos[44] = \input[43] ;
  assign \input[43]  = \input  [43];
  assign shiftLeftOnePos[43] = \input[42] ;
  assign \input[42]  = \input  [42];
  assign shiftLeftOnePos[42] = \input[41] ;
  assign \input[41]  = \input  [41];
  assign shiftLeftOnePos[41] = \input[40] ;
  assign \input[40]  = \input  [40];
  assign shiftLeftOnePos[40] = \input[39] ;
  assign \input[39]  = \input  [39];
  assign shiftLeftOnePos[39] = \input[38] ;
  assign \input[38]  = \input  [38];
  assign shiftLeftOnePos[38] = \input[37] ;
  assign \input[37]  = \input  [37];
  assign shiftLeftOnePos[37] = \input[36] ;
  assign \input[36]  = \input  [36];
  assign shiftLeftOnePos[36] = \input[35] ;
  assign \input[35]  = \input  [35];
  assign shiftLeftOnePos[35] = \input[34] ;
  assign \input[34]  = \input  [34];
  assign shiftLeftOnePos[34] = \input[33] ;
  assign \input[33]  = \input  [33];
  assign shiftLeftOnePos[33] = \input[32] ;
  assign \input[32]  = \input  [32];
  assign shiftLeftOnePos[32] = \input[31] ;
  assign \input[31]  = \input  [31];
  assign shiftLeftOnePos[31] = \input[30] ;
  assign \input[30]  = \input  [30];
  assign shiftLeftOnePos[30] = \input[29] ;
  assign \input[29]  = \input  [29];
  assign shiftLeftOnePos[29] = \input[28] ;
  assign \input[28]  = \input  [28];
  assign shiftLeftOnePos[28] = \input[27] ;
  assign \input[27]  = \input  [27];
  assign shiftLeftOnePos[27] = \input[26] ;
  assign \input[26]  = \input  [26];
  assign shiftLeftOnePos[26] = \input[25] ;
  assign \input[25]  = \input  [25];
  assign shiftLeftOnePos[25] = \input[24] ;
  assign \input[24]  = \input  [24];
  assign shiftLeftOnePos[24] = \input[23] ;
  assign \input[23]  = \input  [23];
  assign shiftLeftOnePos[23] = \input[22] ;
  assign \input[22]  = \input  [22];
  assign shiftLeftOnePos[22] = \input[21] ;
  assign \input[21]  = \input  [21];
  assign shiftLeftOnePos[21] = \input[20] ;
  assign \input[20]  = \input  [20];
  assign shiftLeftOnePos[20] = \input[19] ;
  assign \input[19]  = \input  [19];
  assign shiftLeftOnePos[19] = \input[18] ;
  assign \input[18]  = \input  [18];
  assign shiftLeftOnePos[18] = \input[17] ;
  assign \input[17]  = \input  [17];
  assign shiftLeftOnePos[17] = \input[16] ;
  assign \input[16]  = \input  [16];
  assign shiftLeftOnePos[16] = \input[15] ;
  assign \input[15]  = \input  [15];
  assign shiftLeftOnePos[15] = \input[14] ;
  assign \input[14]  = \input  [14];
  assign shiftLeftOnePos[14] = \input[13] ;
  assign \input[13]  = \input  [13];
  assign shiftLeftOnePos[13] = \input[12] ;
  assign \input[12]  = \input  [12];
  assign shiftLeftOnePos[12] = \input[11] ;
  assign \input[11]  = \input  [11];
  assign shiftLeftOnePos[11] = \input[10] ;
  assign \input[10]  = \input  [10];
  assign shiftLeftOnePos[10] = \input[9] ;
  assign \input[9]  = \input  [9];
  assign shiftLeftOnePos[9] = \input[8] ;
  assign \input[8]  = \input  [8];
  assign shiftLeftOnePos[8] = \input[7] ;
  assign \input[7]  = \input  [7];
  assign shiftLeftOnePos[7] = \input[6] ;
  assign \input[6]  = \input  [6];
  assign shiftLeftOnePos[6] = \input[5] ;
  assign \input[5]  = \input  [5];
  assign shiftLeftOnePos[5] = \input[4] ;
  assign \input[4]  = \input  [4];
  assign shiftLeftOnePos[4] = \input[3] ;
  assign \input[3]  = \input  [3];
  assign shiftLeftOnePos[3] = \input[2] ;
  assign \input[2]  = \input  [2];
  assign shiftLeftOnePos[2] = \input[1] ;
  assign \input[1]  = \input  [1];
  assign shiftLeftOnePos[1] = \input[0] ;
  assign \input[0]  = \input  [0];

endmodule


module complementer_N64_28_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n190, n191, n192, n194, n196, n197, n198, n199, n200, n202,
         n203, n204, n206, n207, n208, n210, n211, n212, n213, n214, n216,
         n217, n218, n220, n221, n222, n224, n225, n226, n228, n229, n230,
         n232, n233, n234, n235, n237, n238, n239, n241, n242, n243, n245,
         n246, n247, n249, n250, n189, n193, n195, n201, n205, n209, n215,
         n219, n223, n227, n231, n236, n240, n244, n248, n251;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U81 ( .A(n190), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U82 ( .A(n192), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U85 ( .A(n196), .B(B[62]), .Z(DIFF[62]) );
  XOR2_X1 U86 ( .A(n194), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U87 ( .A(n198), .B(B[59]), .Z(DIFF[59]) );
  XOR2_X1 U89 ( .A(n200), .B(B[57]), .Z(DIFF[57]) );
  XOR2_X1 U90 ( .A(n202), .B(B[55]), .Z(DIFF[55]) );
  XOR2_X1 U92 ( .A(n204), .B(B[53]), .Z(DIFF[53]) );
  XOR2_X1 U93 ( .A(n206), .B(B[51]), .Z(DIFF[51]) );
  XOR2_X1 U95 ( .A(n208), .B(B[49]), .Z(DIFF[49]) );
  XOR2_X1 U96 ( .A(n212), .B(B[47]), .Z(DIFF[47]) );
  XOR2_X1 U98 ( .A(n214), .B(B[45]), .Z(DIFF[45]) );
  XOR2_X1 U99 ( .A(n216), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U101 ( .A(n218), .B(B[41]), .Z(DIFF[41]) );
  XOR2_X1 U102 ( .A(n211), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U103 ( .A(n220), .B(B[39]), .Z(DIFF[39]) );
  XOR2_X1 U105 ( .A(n222), .B(B[37]), .Z(DIFF[37]) );
  XOR2_X1 U106 ( .A(n224), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U108 ( .A(n226), .B(B[33]), .Z(DIFF[33]) );
  XOR2_X1 U109 ( .A(n228), .B(B[31]), .Z(DIFF[31]) );
  XOR2_X1 U111 ( .A(n230), .B(B[29]), .Z(DIFF[29]) );
  XOR2_X1 U112 ( .A(n233), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U114 ( .A(n235), .B(B[25]), .Z(DIFF[25]) );
  XOR2_X1 U115 ( .A(n237), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U117 ( .A(n239), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U118 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U119 ( .A(n241), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U121 ( .A(n243), .B(B[17]), .Z(DIFF[17]) );
  XOR2_X1 U122 ( .A(n245), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U124 ( .A(n247), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U125 ( .A(n249), .B(B[11]), .Z(DIFF[11]) );
  XOR2_X1 U1 ( .A(n197), .B(n251), .Z(DIFF[61]) );
  NAND2_X1 U2 ( .A1(n197), .A2(n251), .ZN(n196) );
  XNOR2_X1 U3 ( .A(B[40]), .B(n221), .ZN(DIFF[40]) );
  NOR2_X1 U4 ( .A1(B[39]), .A2(n220), .ZN(n221) );
  OR3_X1 U5 ( .A1(B[37]), .A2(B[38]), .A3(n222), .ZN(n220) );
  OR3_X1 U6 ( .A1(B[39]), .A2(B[40]), .A3(n220), .ZN(n218) );
  XNOR2_X1 U7 ( .A(n189), .B(B[38]), .ZN(DIFF[38]) );
  NOR2_X1 U8 ( .A1(n222), .A2(B[37]), .ZN(n189) );
  NOR3_X1 U9 ( .A1(B[59]), .A2(B[60]), .A3(n198), .ZN(n197) );
  XNOR2_X1 U10 ( .A(n193), .B(B[46]), .ZN(DIFF[46]) );
  NOR2_X1 U11 ( .A1(n214), .A2(B[45]), .ZN(n193) );
  XNOR2_X1 U12 ( .A(n195), .B(B[54]), .ZN(DIFF[54]) );
  NOR2_X1 U13 ( .A1(n204), .A2(B[53]), .ZN(n195) );
  XNOR2_X1 U14 ( .A(B[44]), .B(n217), .ZN(DIFF[44]) );
  NOR2_X1 U15 ( .A1(B[43]), .A2(n216), .ZN(n217) );
  XNOR2_X1 U16 ( .A(B[48]), .B(n213), .ZN(DIFF[48]) );
  NOR2_X1 U17 ( .A1(B[47]), .A2(n212), .ZN(n213) );
  XNOR2_X1 U18 ( .A(B[56]), .B(n203), .ZN(DIFF[56]) );
  NOR2_X1 U19 ( .A1(B[55]), .A2(n202), .ZN(n203) );
  XNOR2_X1 U20 ( .A(B[52]), .B(n207), .ZN(DIFF[52]) );
  NOR2_X1 U21 ( .A1(B[51]), .A2(n206), .ZN(n207) );
  XNOR2_X1 U22 ( .A(B[60]), .B(n199), .ZN(DIFF[60]) );
  NOR2_X1 U23 ( .A1(B[59]), .A2(n198), .ZN(n199) );
  OR3_X1 U24 ( .A1(B[45]), .A2(B[46]), .A3(n214), .ZN(n212) );
  OR3_X1 U25 ( .A1(B[57]), .A2(B[58]), .A3(n200), .ZN(n198) );
  OR3_X1 U26 ( .A1(B[53]), .A2(B[54]), .A3(n204), .ZN(n202) );
  OR3_X1 U27 ( .A1(B[49]), .A2(B[50]), .A3(n208), .ZN(n206) );
  OR3_X1 U28 ( .A1(B[41]), .A2(B[42]), .A3(n218), .ZN(n216) );
  OR3_X1 U29 ( .A1(B[43]), .A2(B[44]), .A3(n216), .ZN(n214) );
  OR3_X1 U30 ( .A1(B[47]), .A2(B[48]), .A3(n212), .ZN(n208) );
  OR3_X1 U31 ( .A1(B[55]), .A2(B[56]), .A3(n202), .ZN(n200) );
  OR3_X1 U32 ( .A1(B[51]), .A2(B[52]), .A3(n206), .ZN(n204) );
  XNOR2_X1 U33 ( .A(n201), .B(B[58]), .ZN(DIFF[58]) );
  NOR2_X1 U34 ( .A1(n200), .A2(B[57]), .ZN(n201) );
  XNOR2_X1 U35 ( .A(n205), .B(B[50]), .ZN(DIFF[50]) );
  NOR2_X1 U36 ( .A1(n208), .A2(B[49]), .ZN(n205) );
  XNOR2_X1 U37 ( .A(n209), .B(B[42]), .ZN(DIFF[42]) );
  NOR2_X1 U38 ( .A1(n218), .A2(B[41]), .ZN(n209) );
  XNOR2_X1 U39 ( .A(B[36]), .B(n225), .ZN(DIFF[36]) );
  NOR2_X1 U40 ( .A1(B[35]), .A2(n224), .ZN(n225) );
  OR3_X1 U41 ( .A1(B[35]), .A2(B[36]), .A3(n224), .ZN(n222) );
  XNOR2_X1 U42 ( .A(n215), .B(B[63]), .ZN(DIFF[63]) );
  NOR2_X1 U43 ( .A1(n196), .A2(B[62]), .ZN(n215) );
  XNOR2_X1 U44 ( .A(n219), .B(B[14]), .ZN(DIFF[14]) );
  NOR2_X1 U45 ( .A1(n247), .A2(B[13]), .ZN(n219) );
  XNOR2_X1 U46 ( .A(n223), .B(B[10]), .ZN(DIFF[10]) );
  NOR2_X1 U47 ( .A1(n190), .A2(B[9]), .ZN(n223) );
  XNOR2_X1 U48 ( .A(n227), .B(B[6]), .ZN(DIFF[6]) );
  NOR2_X1 U49 ( .A1(n194), .A2(B[5]), .ZN(n227) );
  XNOR2_X1 U50 ( .A(B[12]), .B(n250), .ZN(DIFF[12]) );
  NOR2_X1 U51 ( .A1(B[11]), .A2(n249), .ZN(n250) );
  XNOR2_X1 U52 ( .A(B[8]), .B(n191), .ZN(DIFF[8]) );
  NOR2_X1 U53 ( .A1(B[7]), .A2(n192), .ZN(n191) );
  XNOR2_X1 U54 ( .A(B[16]), .B(n246), .ZN(DIFF[16]) );
  NOR2_X1 U55 ( .A1(B[15]), .A2(n245), .ZN(n246) );
  OR3_X1 U56 ( .A1(B[5]), .A2(B[6]), .A3(n194), .ZN(n192) );
  OR3_X1 U57 ( .A1(B[13]), .A2(B[14]), .A3(n247), .ZN(n245) );
  OR3_X1 U58 ( .A1(B[17]), .A2(B[18]), .A3(n243), .ZN(n241) );
  OR3_X1 U59 ( .A1(B[21]), .A2(B[22]), .A3(n239), .ZN(n237) );
  OR3_X1 U60 ( .A1(B[10]), .A2(B[9]), .A3(n190), .ZN(n249) );
  OR3_X1 U61 ( .A1(B[7]), .A2(B[8]), .A3(n192), .ZN(n190) );
  OR3_X1 U62 ( .A1(B[11]), .A2(B[12]), .A3(n249), .ZN(n247) );
  OR3_X1 U63 ( .A1(B[15]), .A2(B[16]), .A3(n245), .ZN(n243) );
  OR3_X1 U64 ( .A1(B[19]), .A2(B[20]), .A3(n241), .ZN(n239) );
  XNOR2_X1 U65 ( .A(n231), .B(B[34]), .ZN(DIFF[34]) );
  NOR2_X1 U66 ( .A1(n226), .A2(B[33]), .ZN(n231) );
  XNOR2_X1 U67 ( .A(n236), .B(B[30]), .ZN(DIFF[30]) );
  NOR2_X1 U68 ( .A1(n230), .A2(B[29]), .ZN(n236) );
  XNOR2_X1 U69 ( .A(n240), .B(B[26]), .ZN(DIFF[26]) );
  NOR2_X1 U70 ( .A1(n235), .A2(B[25]), .ZN(n240) );
  XNOR2_X1 U71 ( .A(n244), .B(B[22]), .ZN(DIFF[22]) );
  NOR2_X1 U72 ( .A1(n239), .A2(B[21]), .ZN(n244) );
  XNOR2_X1 U73 ( .A(n248), .B(B[18]), .ZN(DIFF[18]) );
  NOR2_X1 U74 ( .A1(n243), .A2(B[17]), .ZN(n248) );
  XNOR2_X1 U75 ( .A(B[28]), .B(n234), .ZN(DIFF[28]) );
  NOR2_X1 U76 ( .A1(B[27]), .A2(n233), .ZN(n234) );
  XNOR2_X1 U77 ( .A(B[20]), .B(n242), .ZN(DIFF[20]) );
  NOR2_X1 U78 ( .A1(B[19]), .A2(n241), .ZN(n242) );
  XNOR2_X1 U79 ( .A(B[32]), .B(n229), .ZN(DIFF[32]) );
  NOR2_X1 U80 ( .A1(B[31]), .A2(n228), .ZN(n229) );
  XNOR2_X1 U83 ( .A(B[24]), .B(n238), .ZN(DIFF[24]) );
  NOR2_X1 U84 ( .A1(B[23]), .A2(n237), .ZN(n238) );
  OR3_X1 U88 ( .A1(B[25]), .A2(B[26]), .A3(n235), .ZN(n233) );
  OR3_X1 U91 ( .A1(B[29]), .A2(B[30]), .A3(n230), .ZN(n228) );
  OR3_X1 U94 ( .A1(B[33]), .A2(B[34]), .A3(n226), .ZN(n224) );
  OR3_X1 U97 ( .A1(B[23]), .A2(B[24]), .A3(n237), .ZN(n235) );
  OR3_X1 U100 ( .A1(B[27]), .A2(B[28]), .A3(n233), .ZN(n230) );
  OR3_X1 U104 ( .A1(B[31]), .A2(B[32]), .A3(n228), .ZN(n226) );
  OR3_X1 U107 ( .A1(B[3]), .A2(B[4]), .A3(n211), .ZN(n194) );
  XNOR2_X1 U110 ( .A(B[4]), .B(n210), .ZN(DIFF[4]) );
  NOR2_X1 U113 ( .A1(B[3]), .A2(n211), .ZN(n210) );
  XNOR2_X1 U116 ( .A(B[2]), .B(n232), .ZN(DIFF[2]) );
  OR3_X1 U120 ( .A1(B[1]), .A2(B[2]), .A3(\B[0] ), .ZN(n211) );
  NOR2_X1 U123 ( .A1(\B[0] ), .A2(B[1]), .ZN(n232) );
  INV_X1 U126 ( .A(B[61]), .ZN(n251) );
endmodule


module complementer_N64_28 ( \input , complement2 );
  input [63:0] \input ;
  output [63:0] complement2;


  complementer_N64_28_DW01_sub_0 sub_add_31_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(\input ), .CI(1'b0), .DIFF(complement2) );
endmodule


module complementer_N64_27_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n189;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U81 ( .A(n190), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U82 ( .A(n192), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U83 ( .A(n193), .B(B[6]), .Z(DIFF[6]) );
  XOR2_X1 U84 ( .A(n195), .B(B[63]), .Z(DIFF[63]) );
  XOR2_X1 U85 ( .A(n196), .B(B[62]), .Z(DIFF[62]) );
  XOR2_X1 U86 ( .A(n194), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U87 ( .A(n198), .B(B[59]), .Z(DIFF[59]) );
  XOR2_X1 U88 ( .A(n201), .B(B[58]), .Z(DIFF[58]) );
  XOR2_X1 U89 ( .A(n200), .B(B[57]), .Z(DIFF[57]) );
  XOR2_X1 U90 ( .A(n202), .B(B[55]), .Z(DIFF[55]) );
  XOR2_X1 U91 ( .A(n205), .B(B[54]), .Z(DIFF[54]) );
  XOR2_X1 U92 ( .A(n204), .B(B[53]), .Z(DIFF[53]) );
  XOR2_X1 U93 ( .A(n206), .B(B[51]), .Z(DIFF[51]) );
  XOR2_X1 U94 ( .A(n209), .B(B[50]), .Z(DIFF[50]) );
  XOR2_X1 U95 ( .A(n208), .B(B[49]), .Z(DIFF[49]) );
  XOR2_X1 U96 ( .A(n212), .B(B[47]), .Z(DIFF[47]) );
  XOR2_X1 U97 ( .A(n215), .B(B[46]), .Z(DIFF[46]) );
  XOR2_X1 U98 ( .A(n214), .B(B[45]), .Z(DIFF[45]) );
  XOR2_X1 U99 ( .A(n216), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U100 ( .A(n219), .B(B[42]), .Z(DIFF[42]) );
  XOR2_X1 U101 ( .A(n218), .B(B[41]), .Z(DIFF[41]) );
  XOR2_X1 U102 ( .A(n211), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U103 ( .A(n220), .B(B[39]), .Z(DIFF[39]) );
  XOR2_X1 U104 ( .A(n223), .B(B[38]), .Z(DIFF[38]) );
  XOR2_X1 U105 ( .A(n222), .B(B[37]), .Z(DIFF[37]) );
  XOR2_X1 U106 ( .A(n224), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U107 ( .A(n227), .B(B[34]), .Z(DIFF[34]) );
  XOR2_X1 U108 ( .A(n226), .B(B[33]), .Z(DIFF[33]) );
  XOR2_X1 U109 ( .A(n228), .B(B[31]), .Z(DIFF[31]) );
  XOR2_X1 U110 ( .A(n231), .B(B[30]), .Z(DIFF[30]) );
  XOR2_X1 U111 ( .A(n230), .B(B[29]), .Z(DIFF[29]) );
  XOR2_X1 U112 ( .A(n233), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U113 ( .A(n236), .B(B[26]), .Z(DIFF[26]) );
  XOR2_X1 U114 ( .A(n235), .B(B[25]), .Z(DIFF[25]) );
  XOR2_X1 U115 ( .A(n237), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U116 ( .A(n240), .B(B[22]), .Z(DIFF[22]) );
  XOR2_X1 U117 ( .A(n239), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U118 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U119 ( .A(n241), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U120 ( .A(n244), .B(B[18]), .Z(DIFF[18]) );
  XOR2_X1 U121 ( .A(n243), .B(B[17]), .Z(DIFF[17]) );
  XOR2_X1 U122 ( .A(n245), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U123 ( .A(n248), .B(B[14]), .Z(DIFF[14]) );
  XOR2_X1 U124 ( .A(n247), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U125 ( .A(n249), .B(B[11]), .Z(DIFF[11]) );
  XOR2_X1 U126 ( .A(n251), .B(B[10]), .Z(DIFF[10]) );
  NOR2_X1 U1 ( .A1(B[43]), .A2(n216), .ZN(n217) );
  NAND2_X1 U2 ( .A1(n197), .A2(n189), .ZN(n196) );
  OR2_X1 U3 ( .A1(n204), .A2(B[53]), .ZN(n205) );
  XNOR2_X1 U4 ( .A(B[40]), .B(n221), .ZN(DIFF[40]) );
  NOR3_X1 U5 ( .A1(B[59]), .A2(B[60]), .A3(n198), .ZN(n197) );
  NOR2_X1 U6 ( .A1(B[47]), .A2(n212), .ZN(n213) );
  NOR2_X1 U7 ( .A1(B[55]), .A2(n202), .ZN(n203) );
  NOR2_X1 U8 ( .A1(B[51]), .A2(n206), .ZN(n207) );
  NOR2_X1 U9 ( .A1(B[39]), .A2(n220), .ZN(n221) );
  NOR2_X1 U10 ( .A1(B[59]), .A2(n198), .ZN(n199) );
  OR3_X1 U11 ( .A1(B[45]), .A2(B[46]), .A3(n214), .ZN(n212) );
  OR3_X1 U12 ( .A1(B[57]), .A2(B[58]), .A3(n200), .ZN(n198) );
  OR3_X1 U13 ( .A1(B[53]), .A2(B[54]), .A3(n204), .ZN(n202) );
  OR3_X1 U14 ( .A1(B[49]), .A2(B[50]), .A3(n208), .ZN(n206) );
  OR3_X1 U15 ( .A1(B[41]), .A2(B[42]), .A3(n218), .ZN(n216) );
  OR3_X1 U16 ( .A1(B[43]), .A2(B[44]), .A3(n216), .ZN(n214) );
  OR3_X1 U17 ( .A1(B[47]), .A2(B[48]), .A3(n212), .ZN(n208) );
  OR3_X1 U18 ( .A1(B[55]), .A2(B[56]), .A3(n202), .ZN(n200) );
  OR3_X1 U19 ( .A1(B[51]), .A2(B[52]), .A3(n206), .ZN(n204) );
  OR3_X1 U20 ( .A1(B[39]), .A2(B[40]), .A3(n220), .ZN(n218) );
  XNOR2_X1 U21 ( .A(B[44]), .B(n217), .ZN(DIFF[44]) );
  XNOR2_X1 U22 ( .A(B[56]), .B(n203), .ZN(DIFF[56]) );
  XNOR2_X1 U23 ( .A(B[52]), .B(n207), .ZN(DIFF[52]) );
  XNOR2_X1 U24 ( .A(B[48]), .B(n213), .ZN(DIFF[48]) );
  XNOR2_X1 U25 ( .A(n197), .B(B[61]), .ZN(DIFF[61]) );
  XNOR2_X1 U26 ( .A(B[60]), .B(n199), .ZN(DIFF[60]) );
  OR2_X1 U27 ( .A1(n214), .A2(B[45]), .ZN(n215) );
  OR2_X1 U28 ( .A1(n208), .A2(B[49]), .ZN(n209) );
  OR2_X1 U29 ( .A1(n200), .A2(B[57]), .ZN(n201) );
  OR2_X1 U30 ( .A1(n218), .A2(B[41]), .ZN(n219) );
  OR2_X1 U31 ( .A1(n196), .A2(B[62]), .ZN(n195) );
  XNOR2_X1 U32 ( .A(B[36]), .B(n225), .ZN(DIFF[36]) );
  OR2_X1 U33 ( .A1(n222), .A2(B[37]), .ZN(n223) );
  OR3_X1 U34 ( .A1(B[37]), .A2(B[38]), .A3(n222), .ZN(n220) );
  NOR2_X1 U35 ( .A1(B[15]), .A2(n245), .ZN(n246) );
  NOR2_X1 U36 ( .A1(B[11]), .A2(n249), .ZN(n250) );
  NOR2_X1 U37 ( .A1(B[7]), .A2(n192), .ZN(n191) );
  OR3_X1 U38 ( .A1(B[10]), .A2(B[9]), .A3(n190), .ZN(n249) );
  OR3_X1 U39 ( .A1(B[21]), .A2(B[22]), .A3(n239), .ZN(n237) );
  OR3_X1 U40 ( .A1(B[17]), .A2(B[18]), .A3(n243), .ZN(n241) );
  OR3_X1 U41 ( .A1(B[13]), .A2(B[14]), .A3(n247), .ZN(n245) );
  OR3_X1 U42 ( .A1(B[5]), .A2(B[6]), .A3(n194), .ZN(n192) );
  OR3_X1 U43 ( .A1(B[19]), .A2(B[20]), .A3(n241), .ZN(n239) );
  OR3_X1 U44 ( .A1(B[15]), .A2(B[16]), .A3(n245), .ZN(n243) );
  OR3_X1 U45 ( .A1(B[11]), .A2(B[12]), .A3(n249), .ZN(n247) );
  OR3_X1 U46 ( .A1(B[7]), .A2(B[8]), .A3(n192), .ZN(n190) );
  XNOR2_X1 U47 ( .A(B[16]), .B(n246), .ZN(DIFF[16]) );
  XNOR2_X1 U48 ( .A(B[12]), .B(n250), .ZN(DIFF[12]) );
  XNOR2_X1 U49 ( .A(B[8]), .B(n191), .ZN(DIFF[8]) );
  OR2_X1 U50 ( .A1(n194), .A2(B[5]), .ZN(n193) );
  OR2_X1 U51 ( .A1(n190), .A2(B[9]), .ZN(n251) );
  NOR2_X1 U52 ( .A1(B[35]), .A2(n224), .ZN(n225) );
  NOR2_X1 U53 ( .A1(B[31]), .A2(n228), .ZN(n229) );
  NOR2_X1 U54 ( .A1(B[27]), .A2(n233), .ZN(n234) );
  NOR2_X1 U55 ( .A1(B[23]), .A2(n237), .ZN(n238) );
  NOR2_X1 U56 ( .A1(B[19]), .A2(n241), .ZN(n242) );
  OR3_X1 U57 ( .A1(B[33]), .A2(B[34]), .A3(n226), .ZN(n224) );
  OR3_X1 U58 ( .A1(B[29]), .A2(B[30]), .A3(n230), .ZN(n228) );
  OR3_X1 U59 ( .A1(B[25]), .A2(B[26]), .A3(n235), .ZN(n233) );
  OR3_X1 U60 ( .A1(B[35]), .A2(B[36]), .A3(n224), .ZN(n222) );
  OR3_X1 U61 ( .A1(B[31]), .A2(B[32]), .A3(n228), .ZN(n226) );
  OR3_X1 U62 ( .A1(B[27]), .A2(B[28]), .A3(n233), .ZN(n230) );
  OR3_X1 U63 ( .A1(B[23]), .A2(B[24]), .A3(n237), .ZN(n235) );
  XNOR2_X1 U64 ( .A(B[32]), .B(n229), .ZN(DIFF[32]) );
  XNOR2_X1 U65 ( .A(B[28]), .B(n234), .ZN(DIFF[28]) );
  XNOR2_X1 U66 ( .A(B[24]), .B(n238), .ZN(DIFF[24]) );
  XNOR2_X1 U67 ( .A(B[20]), .B(n242), .ZN(DIFF[20]) );
  OR2_X1 U68 ( .A1(n226), .A2(B[33]), .ZN(n227) );
  OR2_X1 U69 ( .A1(n230), .A2(B[29]), .ZN(n231) );
  OR2_X1 U70 ( .A1(n235), .A2(B[25]), .ZN(n236) );
  OR2_X1 U71 ( .A1(n239), .A2(B[21]), .ZN(n240) );
  OR2_X1 U72 ( .A1(n243), .A2(B[17]), .ZN(n244) );
  OR2_X1 U73 ( .A1(n247), .A2(B[13]), .ZN(n248) );
  XNOR2_X1 U74 ( .A(B[4]), .B(n210), .ZN(DIFF[4]) );
  NOR2_X1 U75 ( .A1(B[3]), .A2(n211), .ZN(n210) );
  XNOR2_X1 U76 ( .A(B[2]), .B(n232), .ZN(DIFF[2]) );
  NOR2_X1 U77 ( .A1(\B[0] ), .A2(B[1]), .ZN(n232) );
  OR3_X1 U78 ( .A1(B[3]), .A2(B[4]), .A3(n211), .ZN(n194) );
  OR3_X1 U79 ( .A1(B[1]), .A2(B[2]), .A3(\B[0] ), .ZN(n211) );
  INV_X1 U80 ( .A(B[61]), .ZN(n189) );
endmodule


module complementer_N64_27 ( \input , complement2 );
  input [63:0] \input ;
  output [63:0] complement2;


  complementer_N64_27_DW01_sub_0 sub_add_31_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(\input ), .CI(1'b0), .DIFF(complement2) );
endmodule


module ShiftnCompl_N64_14 ( plusA, plus2A_out, minus2A_out, plus4A_out, 
        minus4A_out );
  input [63:0] plusA;
  output [63:0] plus2A_out;
  output [63:0] minus2A_out;
  output [63:0] plus4A_out;
  output [63:0] minus4A_out;
  wire   n15, n16, n3, n17, n18, n4, n19, n20, n21, n22, n23, n24;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign plus2A_out[0] = 1'b0;
  assign plus2A_out[51] = n3;
  assign plus2A_out[39] = n4;
  assign plus4A_out[0] = 1'b0;

  shifter_N64_28 shifter_1 ( .\input (plusA), .shiftLeftOnePos({
        plus2A_out[63:59], n15, plus2A_out[57:54], n16, plus2A_out[52], n3, 
        plus2A_out[50:49], n17, plus2A_out[47:44], n18, plus2A_out[42:40], n4, 
        n19, plus2A_out[37:1], SYNOPSYS_UNCONNECTED__0}) );
  shifter_N64_27 shifter_2 ( .\input ({plus2A_out[63:52], n3, 
        plus2A_out[50:40], n4, plus2A_out[38:1], 1'b0}), .shiftLeftOnePos({
        plus4A_out[63:59], n20, plus4A_out[57:54], n21, plus4A_out[52:49], n22, 
        plus4A_out[47:44], n23, plus4A_out[42:39], n24, plus4A_out[37:1], 
        SYNOPSYS_UNCONNECTED__1}) );
  complementer_N64_28 complementer_1 ( .\input ({plus2A_out[63:52], n3, 
        plus2A_out[50:40], n4, plus2A_out[38:1], 1'b0}), .complement2(
        minus2A_out) );
  complementer_N64_27 complementer_2 ( .\input ({plus4A_out[63:1], 1'b0}), 
        .complement2(minus4A_out) );
  BUF_X1 U1 ( .A(n24), .Z(plus4A_out[38]) );
  BUF_X1 U2 ( .A(n23), .Z(plus4A_out[43]) );
  BUF_X1 U5 ( .A(n22), .Z(plus4A_out[48]) );
  BUF_X1 U6 ( .A(n21), .Z(plus4A_out[53]) );
  BUF_X1 U7 ( .A(n20), .Z(plus4A_out[58]) );
  BUF_X1 U8 ( .A(n19), .Z(plus2A_out[38]) );
  BUF_X1 U9 ( .A(n18), .Z(plus2A_out[43]) );
  BUF_X1 U10 ( .A(n17), .Z(plus2A_out[48]) );
  BUF_X1 U11 ( .A(n16), .Z(plus2A_out[53]) );
  BUF_X1 U12 ( .A(n15), .Z(plus2A_out[58]) );
endmodule


module MUX_GENERIC_N64_RADIX3_14 ( plusA, minusA, plus2A, minus2A, SEL, Y );
  input [63:0] plusA;
  input [63:0] minusA;
  input [63:0] plus2A;
  input [63:0] minus2A;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304;
  tri   [63:0] Y;

  TBUF_X1 \Y_tri[55]  ( .A(n263), .EN(n301), .Z(Y[55]) );
  TBUF_X1 \Y_tri[56]  ( .A(n264), .EN(n301), .Z(Y[56]) );
  TBUF_X1 \Y_tri[57]  ( .A(n265), .EN(n301), .Z(Y[57]) );
  TBUF_X1 \Y_tri[58]  ( .A(n266), .EN(n301), .Z(Y[58]) );
  TBUF_X1 \Y_tri[59]  ( .A(n267), .EN(n301), .Z(Y[59]) );
  TBUF_X1 \Y_tri[60]  ( .A(n268), .EN(n301), .Z(Y[60]) );
  TBUF_X1 \Y_tri[61]  ( .A(n269), .EN(n301), .Z(Y[61]) );
  TBUF_X1 \Y_tri[63]  ( .A(n271), .EN(n301), .Z(Y[63]) );
  TBUF_X1 \Y_tri[42]  ( .A(n250), .EN(n299), .Z(Y[42]) );
  TBUF_X1 \Y_tri[43]  ( .A(n251), .EN(n299), .Z(Y[43]) );
  TBUF_X1 \Y_tri[44]  ( .A(n252), .EN(n300), .Z(Y[44]) );
  TBUF_X1 \Y_tri[45]  ( .A(n253), .EN(n300), .Z(Y[45]) );
  TBUF_X1 \Y_tri[46]  ( .A(n254), .EN(n300), .Z(Y[46]) );
  TBUF_X1 \Y_tri[47]  ( .A(n255), .EN(n300), .Z(Y[47]) );
  TBUF_X1 \Y_tri[48]  ( .A(n256), .EN(n300), .Z(Y[48]) );
  TBUF_X1 \Y_tri[49]  ( .A(n257), .EN(n300), .Z(Y[49]) );
  TBUF_X1 \Y_tri[50]  ( .A(n258), .EN(n300), .Z(Y[50]) );
  TBUF_X1 \Y_tri[51]  ( .A(n259), .EN(n300), .Z(Y[51]) );
  TBUF_X1 \Y_tri[52]  ( .A(n260), .EN(n300), .Z(Y[52]) );
  TBUF_X1 \Y_tri[53]  ( .A(n261), .EN(n300), .Z(Y[53]) );
  TBUF_X1 \Y_tri[54]  ( .A(n262), .EN(n300), .Z(Y[54]) );
  TBUF_X1 \Y_tri[17]  ( .A(n225), .EN(n297), .Z(Y[17]) );
  TBUF_X1 \Y_tri[18]  ( .A(n226), .EN(n297), .Z(Y[18]) );
  TBUF_X1 \Y_tri[19]  ( .A(n227), .EN(n297), .Z(Y[19]) );
  TBUF_X1 \Y_tri[20]  ( .A(n228), .EN(n297), .Z(Y[20]) );
  TBUF_X1 \Y_tri[21]  ( .A(n229), .EN(n297), .Z(Y[21]) );
  TBUF_X1 \Y_tri[22]  ( .A(n230), .EN(n298), .Z(Y[22]) );
  TBUF_X1 \Y_tri[24]  ( .A(n232), .EN(n298), .Z(Y[24]) );
  TBUF_X1 \Y_tri[25]  ( .A(n233), .EN(n298), .Z(Y[25]) );
  TBUF_X1 \Y_tri[26]  ( .A(n234), .EN(n298), .Z(Y[26]) );
  TBUF_X1 \Y_tri[27]  ( .A(n235), .EN(n298), .Z(Y[27]) );
  TBUF_X1 \Y_tri[28]  ( .A(n236), .EN(n298), .Z(Y[28]) );
  TBUF_X1 \Y_tri[29]  ( .A(n237), .EN(n298), .Z(Y[29]) );
  TBUF_X1 \Y_tri[30]  ( .A(n238), .EN(n298), .Z(Y[30]) );
  TBUF_X1 \Y_tri[31]  ( .A(n239), .EN(n298), .Z(Y[31]) );
  TBUF_X1 \Y_tri[32]  ( .A(n240), .EN(n298), .Z(Y[32]) );
  TBUF_X1 \Y_tri[33]  ( .A(n241), .EN(n299), .Z(Y[33]) );
  TBUF_X1 \Y_tri[34]  ( .A(n242), .EN(n299), .Z(Y[34]) );
  TBUF_X1 \Y_tri[35]  ( .A(n243), .EN(n299), .Z(Y[35]) );
  TBUF_X1 \Y_tri[36]  ( .A(n244), .EN(n299), .Z(Y[36]) );
  TBUF_X1 \Y_tri[37]  ( .A(n245), .EN(n299), .Z(Y[37]) );
  TBUF_X1 \Y_tri[38]  ( .A(n246), .EN(n299), .Z(Y[38]) );
  TBUF_X1 \Y_tri[39]  ( .A(n247), .EN(n299), .Z(Y[39]) );
  TBUF_X1 \Y_tri[40]  ( .A(n248), .EN(n299), .Z(Y[40]) );
  TBUF_X1 \Y_tri[41]  ( .A(n249), .EN(n299), .Z(Y[41]) );
  TBUF_X1 \Y_tri[2]  ( .A(n209), .EN(n296), .Z(Y[2]) );
  TBUF_X1 \Y_tri[3]  ( .A(n210), .EN(n296), .Z(Y[3]) );
  TBUF_X1 \Y_tri[4]  ( .A(n211), .EN(n296), .Z(Y[4]) );
  TBUF_X1 \Y_tri[5]  ( .A(n212), .EN(n296), .Z(Y[5]) );
  TBUF_X1 \Y_tri[6]  ( .A(n213), .EN(n296), .Z(Y[6]) );
  TBUF_X1 \Y_tri[8]  ( .A(n215), .EN(n296), .Z(Y[8]) );
  TBUF_X1 \Y_tri[9]  ( .A(n217), .EN(n296), .Z(Y[9]) );
  TBUF_X1 \Y_tri[10]  ( .A(n218), .EN(n296), .Z(Y[10]) );
  TBUF_X1 \Y_tri[11]  ( .A(n219), .EN(n297), .Z(Y[11]) );
  TBUF_X1 \Y_tri[12]  ( .A(n220), .EN(n297), .Z(Y[12]) );
  TBUF_X1 \Y_tri[13]  ( .A(n221), .EN(n297), .Z(Y[13]) );
  TBUF_X1 \Y_tri[14]  ( .A(n222), .EN(n297), .Z(Y[14]) );
  TBUF_X1 \Y_tri[15]  ( .A(n223), .EN(n297), .Z(Y[15]) );
  TBUF_X1 \Y_tri[1]  ( .A(n208), .EN(n296), .Z(Y[1]) );
  TBUF_X1 \Y_tri[0]  ( .A(n207), .EN(n296), .Z(Y[0]) );
  TBUF_X1 \Y_tri[7]  ( .A(n214), .EN(n296), .Z(Y[7]) );
  TBUF_X1 \Y_tri[16]  ( .A(n224), .EN(n297), .Z(Y[16]) );
  TBUF_X1 \Y_tri[23]  ( .A(n231), .EN(n298), .Z(Y[23]) );
  TBUF_X1 \Y_tri[62]  ( .A(n270), .EN(n301), .Z(Y[62]) );
  NAND2_X1 U2 ( .A1(n52), .A2(n53), .ZN(n249) );
  AOI22_X1 U3 ( .A1(plusA[41]), .A2(n281), .B1(plus2A[41]), .B2(n275), .ZN(n52) );
  AOI22_X1 U4 ( .A1(minus2A[41]), .A2(n293), .B1(minusA[41]), .B2(n287), .ZN(
        n53) );
  NAND2_X1 U5 ( .A1(n56), .A2(n57), .ZN(n247) );
  AOI22_X1 U6 ( .A1(plusA[39]), .A2(n281), .B1(plus2A[39]), .B2(n275), .ZN(n56) );
  AOI22_X1 U7 ( .A1(minus2A[39]), .A2(n293), .B1(minusA[39]), .B2(n287), .ZN(
        n57) );
  NAND2_X1 U8 ( .A1(n54), .A2(n55), .ZN(n248) );
  AOI22_X1 U9 ( .A1(plusA[40]), .A2(n281), .B1(plus2A[40]), .B2(n275), .ZN(n54) );
  AOI22_X1 U10 ( .A1(minus2A[40]), .A2(n293), .B1(minusA[40]), .B2(n287), .ZN(
        n55) );
  NAND2_X1 U11 ( .A1(n58), .A2(n59), .ZN(n246) );
  AOI22_X1 U12 ( .A1(plusA[38]), .A2(n281), .B1(plus2A[38]), .B2(n275), .ZN(
        n58) );
  AOI22_X1 U13 ( .A1(minus2A[38]), .A2(n293), .B1(minusA[38]), .B2(n287), .ZN(
        n59) );
  NAND2_X1 U14 ( .A1(n42), .A2(n43), .ZN(n254) );
  AOI22_X1 U15 ( .A1(plusA[46]), .A2(n281), .B1(plus2A[46]), .B2(n275), .ZN(
        n42) );
  AOI22_X1 U16 ( .A1(minus2A[46]), .A2(n293), .B1(minusA[46]), .B2(n287), .ZN(
        n43) );
  NAND2_X1 U17 ( .A1(n46), .A2(n47), .ZN(n252) );
  AOI22_X1 U18 ( .A1(plusA[44]), .A2(n281), .B1(plus2A[44]), .B2(n275), .ZN(
        n46) );
  AOI22_X1 U19 ( .A1(minus2A[44]), .A2(n293), .B1(minusA[44]), .B2(n287), .ZN(
        n47) );
  NAND2_X1 U20 ( .A1(n44), .A2(n45), .ZN(n253) );
  AOI22_X1 U21 ( .A1(plusA[45]), .A2(n281), .B1(plus2A[45]), .B2(n275), .ZN(
        n44) );
  AOI22_X1 U22 ( .A1(minus2A[45]), .A2(n293), .B1(minusA[45]), .B2(n287), .ZN(
        n45) );
  NAND2_X1 U23 ( .A1(n40), .A2(n41), .ZN(n255) );
  AOI22_X1 U24 ( .A1(plusA[47]), .A2(n281), .B1(plus2A[47]), .B2(n275), .ZN(
        n40) );
  AOI22_X1 U25 ( .A1(minus2A[47]), .A2(n293), .B1(minusA[47]), .B2(n287), .ZN(
        n41) );
  NAND2_X1 U26 ( .A1(n48), .A2(n49), .ZN(n251) );
  AOI22_X1 U27 ( .A1(plusA[43]), .A2(n281), .B1(plus2A[43]), .B2(n275), .ZN(
        n48) );
  AOI22_X1 U28 ( .A1(minus2A[43]), .A2(n293), .B1(minusA[43]), .B2(n287), .ZN(
        n49) );
  NAND2_X1 U29 ( .A1(n22), .A2(n23), .ZN(n264) );
  AOI22_X1 U30 ( .A1(plusA[56]), .A2(n282), .B1(plus2A[56]), .B2(n276), .ZN(
        n22) );
  AOI22_X1 U31 ( .A1(minus2A[56]), .A2(n294), .B1(minusA[56]), .B2(n288), .ZN(
        n23) );
  NAND2_X1 U32 ( .A1(n26), .A2(n27), .ZN(n262) );
  AOI22_X1 U33 ( .A1(plusA[54]), .A2(n282), .B1(plus2A[54]), .B2(n276), .ZN(
        n26) );
  AOI22_X1 U34 ( .A1(minus2A[54]), .A2(n294), .B1(minusA[54]), .B2(n288), .ZN(
        n27) );
  NAND2_X1 U35 ( .A1(n24), .A2(n25), .ZN(n263) );
  AOI22_X1 U36 ( .A1(plusA[55]), .A2(n282), .B1(plus2A[55]), .B2(n276), .ZN(
        n24) );
  AOI22_X1 U37 ( .A1(minus2A[55]), .A2(n294), .B1(minusA[55]), .B2(n288), .ZN(
        n25) );
  NAND2_X1 U38 ( .A1(n28), .A2(n29), .ZN(n261) );
  AOI22_X1 U39 ( .A1(plusA[53]), .A2(n282), .B1(plus2A[53]), .B2(n276), .ZN(
        n28) );
  AOI22_X1 U40 ( .A1(minus2A[53]), .A2(n294), .B1(minusA[53]), .B2(n288), .ZN(
        n29) );
  NAND2_X1 U41 ( .A1(n20), .A2(n21), .ZN(n265) );
  AOI22_X1 U42 ( .A1(plusA[57]), .A2(n282), .B1(plus2A[57]), .B2(n276), .ZN(
        n20) );
  AOI22_X1 U43 ( .A1(minus2A[57]), .A2(n294), .B1(minusA[57]), .B2(n288), .ZN(
        n21) );
  NAND2_X1 U44 ( .A1(n32), .A2(n33), .ZN(n259) );
  AOI22_X1 U45 ( .A1(plusA[51]), .A2(n282), .B1(plus2A[51]), .B2(n276), .ZN(
        n32) );
  AOI22_X1 U46 ( .A1(minus2A[51]), .A2(n294), .B1(minusA[51]), .B2(n288), .ZN(
        n33) );
  NAND2_X1 U47 ( .A1(n36), .A2(n37), .ZN(n257) );
  AOI22_X1 U48 ( .A1(plusA[49]), .A2(n282), .B1(plus2A[49]), .B2(n276), .ZN(
        n36) );
  AOI22_X1 U49 ( .A1(minus2A[49]), .A2(n294), .B1(minusA[49]), .B2(n288), .ZN(
        n37) );
  NAND2_X1 U50 ( .A1(n30), .A2(n31), .ZN(n260) );
  AOI22_X1 U51 ( .A1(plusA[52]), .A2(n282), .B1(plus2A[52]), .B2(n276), .ZN(
        n30) );
  AOI22_X1 U52 ( .A1(minus2A[52]), .A2(n294), .B1(minusA[52]), .B2(n288), .ZN(
        n31) );
  NAND2_X1 U53 ( .A1(n34), .A2(n35), .ZN(n258) );
  AOI22_X1 U54 ( .A1(plusA[50]), .A2(n282), .B1(plus2A[50]), .B2(n276), .ZN(
        n34) );
  AOI22_X1 U55 ( .A1(minus2A[50]), .A2(n294), .B1(minusA[50]), .B2(n288), .ZN(
        n35) );
  NAND2_X1 U56 ( .A1(n38), .A2(n39), .ZN(n256) );
  AOI22_X1 U57 ( .A1(plusA[48]), .A2(n282), .B1(plus2A[48]), .B2(n276), .ZN(
        n38) );
  AOI22_X1 U58 ( .A1(minus2A[48]), .A2(n294), .B1(minusA[48]), .B2(n288), .ZN(
        n39) );
  NAND2_X1 U59 ( .A1(n50), .A2(n51), .ZN(n250) );
  AOI22_X1 U60 ( .A1(plusA[42]), .A2(n281), .B1(plus2A[42]), .B2(n275), .ZN(
        n50) );
  AOI22_X1 U61 ( .A1(minus2A[42]), .A2(n293), .B1(minusA[42]), .B2(n287), .ZN(
        n51) );
  NAND2_X1 U62 ( .A1(n12), .A2(n13), .ZN(n269) );
  AOI22_X1 U63 ( .A1(plusA[61]), .A2(n283), .B1(plus2A[61]), .B2(n277), .ZN(
        n12) );
  AOI22_X1 U64 ( .A1(minus2A[61]), .A2(n295), .B1(minusA[61]), .B2(n289), .ZN(
        n13) );
  NAND2_X1 U65 ( .A1(n14), .A2(n15), .ZN(n268) );
  AOI22_X1 U66 ( .A1(plusA[60]), .A2(n283), .B1(plus2A[60]), .B2(n277), .ZN(
        n14) );
  AOI22_X1 U67 ( .A1(minus2A[60]), .A2(n295), .B1(minusA[60]), .B2(n289), .ZN(
        n15) );
  NAND2_X1 U68 ( .A1(n16), .A2(n17), .ZN(n267) );
  AOI22_X1 U69 ( .A1(plusA[59]), .A2(n282), .B1(plus2A[59]), .B2(n276), .ZN(
        n16) );
  AOI22_X1 U70 ( .A1(minus2A[59]), .A2(n294), .B1(minusA[59]), .B2(n288), .ZN(
        n17) );
  NAND2_X1 U71 ( .A1(n18), .A2(n19), .ZN(n266) );
  AOI22_X1 U72 ( .A1(plusA[58]), .A2(n282), .B1(plus2A[58]), .B2(n276), .ZN(
        n18) );
  AOI22_X1 U73 ( .A1(minus2A[58]), .A2(n294), .B1(minusA[58]), .B2(n288), .ZN(
        n19) );
  NAND2_X1 U74 ( .A1(n10), .A2(n11), .ZN(n270) );
  AOI22_X1 U75 ( .A1(plusA[62]), .A2(n283), .B1(plus2A[62]), .B2(n277), .ZN(
        n10) );
  AOI22_X1 U76 ( .A1(minus2A[62]), .A2(n295), .B1(minusA[62]), .B2(n289), .ZN(
        n11) );
  BUF_X1 U77 ( .A(n8), .Z(n278) );
  BUF_X1 U78 ( .A(n6), .Z(n290) );
  BUF_X1 U79 ( .A(n7), .Z(n284) );
  BUF_X1 U80 ( .A(n9), .Z(n272) );
  BUF_X1 U81 ( .A(n216), .Z(n296) );
  BUF_X1 U82 ( .A(n8), .Z(n279) );
  BUF_X1 U83 ( .A(n6), .Z(n291) );
  BUF_X1 U84 ( .A(n7), .Z(n285) );
  BUF_X1 U85 ( .A(n9), .Z(n273) );
  BUF_X1 U86 ( .A(n216), .Z(n298) );
  BUF_X1 U87 ( .A(n216), .Z(n297) );
  NAND2_X1 U88 ( .A1(n60), .A2(n61), .ZN(n245) );
  AOI22_X1 U89 ( .A1(plusA[37]), .A2(n281), .B1(plus2A[37]), .B2(n275), .ZN(
        n60) );
  AOI22_X1 U90 ( .A1(minus2A[37]), .A2(n293), .B1(minusA[37]), .B2(n287), .ZN(
        n61) );
  NAND2_X1 U91 ( .A1(n62), .A2(n63), .ZN(n244) );
  AOI22_X1 U92 ( .A1(plusA[36]), .A2(n281), .B1(plus2A[36]), .B2(n275), .ZN(
        n62) );
  AOI22_X1 U93 ( .A1(minus2A[36]), .A2(n293), .B1(minusA[36]), .B2(n287), .ZN(
        n63) );
  BUF_X1 U94 ( .A(n8), .Z(n280) );
  BUF_X1 U95 ( .A(n6), .Z(n292) );
  BUF_X1 U96 ( .A(n7), .Z(n286) );
  BUF_X1 U97 ( .A(n9), .Z(n274) );
  NAND2_X1 U98 ( .A1(n4), .A2(n5), .ZN(n271) );
  AOI22_X1 U99 ( .A1(plusA[63]), .A2(n283), .B1(plus2A[63]), .B2(n277), .ZN(n4) );
  AOI22_X1 U100 ( .A1(minus2A[63]), .A2(n295), .B1(minusA[63]), .B2(n289), 
        .ZN(n5) );
  BUF_X1 U101 ( .A(n8), .Z(n281) );
  BUF_X1 U102 ( .A(n6), .Z(n293) );
  BUF_X1 U103 ( .A(n7), .Z(n287) );
  BUF_X1 U104 ( .A(n9), .Z(n275) );
  BUF_X1 U105 ( .A(n216), .Z(n299) );
  BUF_X1 U106 ( .A(n8), .Z(n282) );
  BUF_X1 U107 ( .A(n6), .Z(n294) );
  BUF_X1 U108 ( .A(n7), .Z(n288) );
  BUF_X1 U109 ( .A(n9), .Z(n276) );
  BUF_X1 U110 ( .A(n216), .Z(n300) );
  BUF_X1 U111 ( .A(n216), .Z(n301) );
  NOR3_X1 U112 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n302), .ZN(n7) );
  NOR3_X1 U113 ( .A1(n302), .A2(SEL[2]), .A3(n303), .ZN(n9) );
  NOR3_X1 U114 ( .A1(SEL[1]), .A2(SEL[2]), .A3(n303), .ZN(n8) );
  NOR2_X1 U115 ( .A1(n118), .A2(n304), .ZN(n216) );
  INV_X1 U116 ( .A(SEL[2]), .ZN(n304) );
  NAND2_X1 U117 ( .A1(n88), .A2(n89), .ZN(n231) );
  AOI22_X1 U118 ( .A1(plusA[23]), .A2(n279), .B1(plus2A[23]), .B2(n273), .ZN(
        n88) );
  AOI22_X1 U119 ( .A1(minus2A[23]), .A2(n291), .B1(minusA[23]), .B2(n285), 
        .ZN(n89) );
  NAND2_X1 U120 ( .A1(n104), .A2(n105), .ZN(n223) );
  AOI22_X1 U121 ( .A1(plusA[15]), .A2(n279), .B1(plus2A[15]), .B2(n273), .ZN(
        n104) );
  AOI22_X1 U122 ( .A1(minus2A[15]), .A2(n291), .B1(minusA[15]), .B2(n285), 
        .ZN(n105) );
  NOR2_X1 U123 ( .A1(SEL[1]), .A2(SEL[0]), .ZN(n118) );
  AND2_X1 U124 ( .A1(SEL[2]), .A2(n118), .ZN(n6) );
  INV_X1 U125 ( .A(SEL[1]), .ZN(n302) );
  INV_X1 U126 ( .A(SEL[0]), .ZN(n303) );
  NAND2_X1 U127 ( .A1(n123), .A2(n124), .ZN(n213) );
  AOI22_X1 U128 ( .A1(plusA[6]), .A2(n278), .B1(plus2A[6]), .B2(n272), .ZN(
        n123) );
  AOI22_X1 U129 ( .A1(minus2A[6]), .A2(n290), .B1(minusA[6]), .B2(n284), .ZN(
        n124) );
  NAND2_X1 U130 ( .A1(n106), .A2(n107), .ZN(n222) );
  AOI22_X1 U131 ( .A1(plusA[14]), .A2(n279), .B1(plus2A[14]), .B2(n273), .ZN(
        n106) );
  AOI22_X1 U132 ( .A1(minus2A[14]), .A2(n291), .B1(minusA[14]), .B2(n285), 
        .ZN(n107) );
  NAND2_X1 U133 ( .A1(n114), .A2(n115), .ZN(n218) );
  AOI22_X1 U134 ( .A1(plusA[10]), .A2(n278), .B1(plus2A[10]), .B2(n272), .ZN(
        n114) );
  AOI22_X1 U135 ( .A1(minus2A[10]), .A2(n290), .B1(minusA[10]), .B2(n284), 
        .ZN(n115) );
  NAND2_X1 U136 ( .A1(n102), .A2(n103), .ZN(n224) );
  AOI22_X1 U137 ( .A1(plusA[16]), .A2(n279), .B1(plus2A[16]), .B2(n273), .ZN(
        n102) );
  AOI22_X1 U138 ( .A1(minus2A[16]), .A2(n291), .B1(minusA[16]), .B2(n285), 
        .ZN(n103) );
  NAND2_X1 U139 ( .A1(n110), .A2(n111), .ZN(n220) );
  AOI22_X1 U140 ( .A1(plusA[12]), .A2(n279), .B1(plus2A[12]), .B2(n273), .ZN(
        n110) );
  AOI22_X1 U141 ( .A1(minus2A[12]), .A2(n291), .B1(minusA[12]), .B2(n285), 
        .ZN(n111) );
  NAND2_X1 U142 ( .A1(n119), .A2(n120), .ZN(n215) );
  AOI22_X1 U143 ( .A1(plusA[8]), .A2(n278), .B1(plus2A[8]), .B2(n272), .ZN(
        n119) );
  AOI22_X1 U144 ( .A1(minus2A[8]), .A2(n290), .B1(minusA[8]), .B2(n284), .ZN(
        n120) );
  NAND2_X1 U145 ( .A1(n125), .A2(n126), .ZN(n212) );
  AOI22_X1 U146 ( .A1(plusA[5]), .A2(n278), .B1(plus2A[5]), .B2(n272), .ZN(
        n125) );
  AOI22_X1 U147 ( .A1(minus2A[5]), .A2(n290), .B1(minusA[5]), .B2(n284), .ZN(
        n126) );
  NAND2_X1 U148 ( .A1(n121), .A2(n122), .ZN(n214) );
  AOI22_X1 U149 ( .A1(plusA[7]), .A2(n278), .B1(plus2A[7]), .B2(n272), .ZN(
        n121) );
  AOI22_X1 U150 ( .A1(minus2A[7]), .A2(n290), .B1(minusA[7]), .B2(n284), .ZN(
        n122) );
  NAND2_X1 U151 ( .A1(n112), .A2(n113), .ZN(n219) );
  AOI22_X1 U152 ( .A1(plusA[11]), .A2(n278), .B1(plus2A[11]), .B2(n272), .ZN(
        n112) );
  AOI22_X1 U153 ( .A1(minus2A[11]), .A2(n290), .B1(minusA[11]), .B2(n284), 
        .ZN(n113) );
  NAND2_X1 U154 ( .A1(n108), .A2(n109), .ZN(n221) );
  AOI22_X1 U155 ( .A1(plusA[13]), .A2(n279), .B1(plus2A[13]), .B2(n273), .ZN(
        n108) );
  AOI22_X1 U156 ( .A1(minus2A[13]), .A2(n291), .B1(minusA[13]), .B2(n285), 
        .ZN(n109) );
  NAND2_X1 U157 ( .A1(n116), .A2(n117), .ZN(n217) );
  AOI22_X1 U158 ( .A1(plusA[9]), .A2(n278), .B1(plus2A[9]), .B2(n272), .ZN(
        n116) );
  AOI22_X1 U159 ( .A1(minus2A[9]), .A2(n290), .B1(minusA[9]), .B2(n284), .ZN(
        n117) );
  NAND2_X1 U160 ( .A1(n72), .A2(n73), .ZN(n239) );
  AOI22_X1 U161 ( .A1(plusA[31]), .A2(n280), .B1(plus2A[31]), .B2(n274), .ZN(
        n72) );
  AOI22_X1 U162 ( .A1(minus2A[31]), .A2(n292), .B1(minusA[31]), .B2(n286), 
        .ZN(n73) );
  NAND2_X1 U163 ( .A1(n74), .A2(n75), .ZN(n238) );
  AOI22_X1 U164 ( .A1(plusA[30]), .A2(n280), .B1(plus2A[30]), .B2(n274), .ZN(
        n74) );
  AOI22_X1 U165 ( .A1(minus2A[30]), .A2(n292), .B1(minusA[30]), .B2(n286), 
        .ZN(n75) );
  NAND2_X1 U166 ( .A1(n76), .A2(n77), .ZN(n237) );
  AOI22_X1 U167 ( .A1(plusA[29]), .A2(n280), .B1(plus2A[29]), .B2(n274), .ZN(
        n76) );
  AOI22_X1 U168 ( .A1(minus2A[29]), .A2(n292), .B1(minusA[29]), .B2(n286), 
        .ZN(n77) );
  NAND2_X1 U169 ( .A1(n80), .A2(n81), .ZN(n235) );
  AOI22_X1 U170 ( .A1(plusA[27]), .A2(n280), .B1(plus2A[27]), .B2(n274), .ZN(
        n80) );
  AOI22_X1 U171 ( .A1(minus2A[27]), .A2(n292), .B1(minusA[27]), .B2(n286), 
        .ZN(n81) );
  NAND2_X1 U172 ( .A1(n82), .A2(n83), .ZN(n234) );
  AOI22_X1 U173 ( .A1(plusA[26]), .A2(n280), .B1(plus2A[26]), .B2(n274), .ZN(
        n82) );
  AOI22_X1 U174 ( .A1(minus2A[26]), .A2(n292), .B1(minusA[26]), .B2(n286), 
        .ZN(n83) );
  NAND2_X1 U175 ( .A1(n84), .A2(n85), .ZN(n233) );
  AOI22_X1 U176 ( .A1(plusA[25]), .A2(n280), .B1(plus2A[25]), .B2(n274), .ZN(
        n84) );
  AOI22_X1 U177 ( .A1(minus2A[25]), .A2(n292), .B1(minusA[25]), .B2(n286), 
        .ZN(n85) );
  NAND2_X1 U178 ( .A1(n90), .A2(n91), .ZN(n230) );
  AOI22_X1 U179 ( .A1(plusA[22]), .A2(n279), .B1(plus2A[22]), .B2(n273), .ZN(
        n90) );
  AOI22_X1 U180 ( .A1(minus2A[22]), .A2(n291), .B1(minusA[22]), .B2(n285), 
        .ZN(n91) );
  NAND2_X1 U181 ( .A1(n92), .A2(n93), .ZN(n229) );
  AOI22_X1 U182 ( .A1(plusA[21]), .A2(n279), .B1(plus2A[21]), .B2(n273), .ZN(
        n92) );
  AOI22_X1 U183 ( .A1(minus2A[21]), .A2(n291), .B1(minusA[21]), .B2(n285), 
        .ZN(n93) );
  NAND2_X1 U184 ( .A1(n96), .A2(n97), .ZN(n227) );
  AOI22_X1 U185 ( .A1(plusA[19]), .A2(n279), .B1(plus2A[19]), .B2(n273), .ZN(
        n96) );
  AOI22_X1 U186 ( .A1(minus2A[19]), .A2(n291), .B1(minusA[19]), .B2(n285), 
        .ZN(n97) );
  NAND2_X1 U187 ( .A1(n98), .A2(n99), .ZN(n226) );
  AOI22_X1 U188 ( .A1(plusA[18]), .A2(n279), .B1(plus2A[18]), .B2(n273), .ZN(
        n98) );
  AOI22_X1 U189 ( .A1(minus2A[18]), .A2(n291), .B1(minusA[18]), .B2(n285), 
        .ZN(n99) );
  NAND2_X1 U190 ( .A1(n100), .A2(n101), .ZN(n225) );
  AOI22_X1 U191 ( .A1(plusA[17]), .A2(n279), .B1(plus2A[17]), .B2(n273), .ZN(
        n100) );
  AOI22_X1 U192 ( .A1(minus2A[17]), .A2(n291), .B1(minusA[17]), .B2(n285), 
        .ZN(n101) );
  NAND2_X1 U193 ( .A1(n66), .A2(n67), .ZN(n242) );
  AOI22_X1 U194 ( .A1(plusA[34]), .A2(n280), .B1(plus2A[34]), .B2(n274), .ZN(
        n66) );
  AOI22_X1 U195 ( .A1(minus2A[34]), .A2(n292), .B1(minusA[34]), .B2(n286), 
        .ZN(n67) );
  NAND2_X1 U196 ( .A1(n64), .A2(n65), .ZN(n243) );
  AOI22_X1 U197 ( .A1(plusA[35]), .A2(n280), .B1(plus2A[35]), .B2(n274), .ZN(
        n64) );
  AOI22_X1 U198 ( .A1(minus2A[35]), .A2(n292), .B1(minusA[35]), .B2(n286), 
        .ZN(n65) );
  NAND2_X1 U199 ( .A1(n70), .A2(n71), .ZN(n240) );
  AOI22_X1 U200 ( .A1(plusA[32]), .A2(n280), .B1(plus2A[32]), .B2(n274), .ZN(
        n70) );
  AOI22_X1 U201 ( .A1(minus2A[32]), .A2(n292), .B1(minusA[32]), .B2(n286), 
        .ZN(n71) );
  NAND2_X1 U202 ( .A1(n78), .A2(n79), .ZN(n236) );
  AOI22_X1 U203 ( .A1(plusA[28]), .A2(n280), .B1(plus2A[28]), .B2(n274), .ZN(
        n78) );
  AOI22_X1 U204 ( .A1(minus2A[28]), .A2(n292), .B1(minusA[28]), .B2(n286), 
        .ZN(n79) );
  NAND2_X1 U205 ( .A1(n86), .A2(n87), .ZN(n232) );
  AOI22_X1 U206 ( .A1(plusA[24]), .A2(n280), .B1(plus2A[24]), .B2(n274), .ZN(
        n86) );
  AOI22_X1 U207 ( .A1(minus2A[24]), .A2(n292), .B1(minusA[24]), .B2(n286), 
        .ZN(n87) );
  NAND2_X1 U208 ( .A1(n94), .A2(n95), .ZN(n228) );
  AOI22_X1 U209 ( .A1(plusA[20]), .A2(n279), .B1(plus2A[20]), .B2(n273), .ZN(
        n94) );
  AOI22_X1 U210 ( .A1(minus2A[20]), .A2(n291), .B1(minusA[20]), .B2(n285), 
        .ZN(n95) );
  NAND2_X1 U211 ( .A1(n68), .A2(n69), .ZN(n241) );
  AOI22_X1 U212 ( .A1(plusA[33]), .A2(n280), .B1(plus2A[33]), .B2(n274), .ZN(
        n68) );
  AOI22_X1 U213 ( .A1(minus2A[33]), .A2(n292), .B1(minusA[33]), .B2(n286), 
        .ZN(n69) );
  NAND2_X1 U214 ( .A1(n127), .A2(n128), .ZN(n211) );
  AOI22_X1 U215 ( .A1(plusA[4]), .A2(n278), .B1(plus2A[4]), .B2(n272), .ZN(
        n127) );
  AOI22_X1 U216 ( .A1(minus2A[4]), .A2(n290), .B1(minusA[4]), .B2(n284), .ZN(
        n128) );
  NAND2_X1 U217 ( .A1(n129), .A2(n130), .ZN(n210) );
  AOI22_X1 U218 ( .A1(plusA[3]), .A2(n278), .B1(plus2A[3]), .B2(n272), .ZN(
        n129) );
  AOI22_X1 U219 ( .A1(minus2A[3]), .A2(n290), .B1(minusA[3]), .B2(n284), .ZN(
        n130) );
  NAND2_X1 U220 ( .A1(n131), .A2(n132), .ZN(n209) );
  AOI22_X1 U221 ( .A1(plusA[2]), .A2(n278), .B1(plus2A[2]), .B2(n272), .ZN(
        n131) );
  AOI22_X1 U222 ( .A1(minus2A[2]), .A2(n290), .B1(minusA[2]), .B2(n284), .ZN(
        n132) );
  NAND2_X1 U223 ( .A1(n133), .A2(n134), .ZN(n208) );
  AOI22_X1 U224 ( .A1(plusA[1]), .A2(n278), .B1(plus2A[1]), .B2(n272), .ZN(
        n133) );
  AOI22_X1 U225 ( .A1(minus2A[1]), .A2(n290), .B1(minusA[1]), .B2(n284), .ZN(
        n134) );
  NAND2_X1 U226 ( .A1(n135), .A2(n136), .ZN(n207) );
  AOI22_X1 U227 ( .A1(plusA[0]), .A2(n278), .B1(plus2A[0]), .B2(n272), .ZN(
        n135) );
  AOI22_X1 U228 ( .A1(minus2A[0]), .A2(n290), .B1(minusA[0]), .B2(n284), .ZN(
        n136) );
  CLKBUF_X1 U229 ( .A(n9), .Z(n277) );
  CLKBUF_X1 U230 ( .A(n8), .Z(n283) );
  CLKBUF_X1 U231 ( .A(n7), .Z(n289) );
  CLKBUF_X1 U232 ( .A(n6), .Z(n295) );
endmodule


module FA_896 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_895 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_894 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_893 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_892 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_891 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_890 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_889 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  AOI22_X1 U4 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
  INV_X1 U5 ( .A(n7), .ZN(Co) );
endmodule


module FA_888 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_887 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_886 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_885 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_884 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_883 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_882 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_881 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_880 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  AOI22_X1 U4 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
  INV_X1 U5 ( .A(n7), .ZN(Co) );
endmodule


module FA_879 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_878 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_877 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_876 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_875 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_874 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_873 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  XNOR2_X1 U4 ( .A(n4), .B(B), .ZN(n6) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_872 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_871 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_870 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_869 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_868 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_867 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_866 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_865 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_864 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_863 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_862 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_861 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_860 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_859 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_858 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_857 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_856 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_855 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_854 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_853 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_852 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_851 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_850 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_849 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_848 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_847 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_846 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_845 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_844 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_843 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_842 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_841 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_840 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_839 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_838 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_837 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_836 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_835 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_834 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  XNOR2_X1 U4 ( .A(n4), .B(B), .ZN(n6) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_833 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N64_14 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Ci;
  output Co;

  wire   [63:1] CTMP;
  tri   [63:0] A;

  FA_896 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_895 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_894 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_893 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(CTMP[4]) );
  FA_892 FAI_5 ( .A(A[4]), .B(B[4]), .Ci(CTMP[4]), .S(S[4]), .Co(CTMP[5]) );
  FA_891 FAI_6 ( .A(A[5]), .B(B[5]), .Ci(CTMP[5]), .S(S[5]), .Co(CTMP[6]) );
  FA_890 FAI_7 ( .A(A[6]), .B(B[6]), .Ci(CTMP[6]), .S(S[6]), .Co(CTMP[7]) );
  FA_889 FAI_8 ( .A(A[7]), .B(B[7]), .Ci(CTMP[7]), .S(S[7]), .Co(CTMP[8]) );
  FA_888 FAI_9 ( .A(A[8]), .B(B[8]), .Ci(CTMP[8]), .S(S[8]), .Co(CTMP[9]) );
  FA_887 FAI_10 ( .A(A[9]), .B(B[9]), .Ci(CTMP[9]), .S(S[9]), .Co(CTMP[10]) );
  FA_886 FAI_11 ( .A(A[10]), .B(B[10]), .Ci(CTMP[10]), .S(S[10]), .Co(CTMP[11]) );
  FA_885 FAI_12 ( .A(A[11]), .B(B[11]), .Ci(CTMP[11]), .S(S[11]), .Co(CTMP[12]) );
  FA_884 FAI_13 ( .A(A[12]), .B(B[12]), .Ci(CTMP[12]), .S(S[12]), .Co(CTMP[13]) );
  FA_883 FAI_14 ( .A(A[13]), .B(B[13]), .Ci(CTMP[13]), .S(S[13]), .Co(CTMP[14]) );
  FA_882 FAI_15 ( .A(A[14]), .B(B[14]), .Ci(CTMP[14]), .S(S[14]), .Co(CTMP[15]) );
  FA_881 FAI_16 ( .A(A[15]), .B(B[15]), .Ci(CTMP[15]), .S(S[15]), .Co(CTMP[16]) );
  FA_880 FAI_17 ( .A(A[16]), .B(B[16]), .Ci(CTMP[16]), .S(S[16]), .Co(CTMP[17]) );
  FA_879 FAI_18 ( .A(A[17]), .B(B[17]), .Ci(CTMP[17]), .S(S[17]), .Co(CTMP[18]) );
  FA_878 FAI_19 ( .A(A[18]), .B(B[18]), .Ci(CTMP[18]), .S(S[18]), .Co(CTMP[19]) );
  FA_877 FAI_20 ( .A(A[19]), .B(B[19]), .Ci(CTMP[19]), .S(S[19]), .Co(CTMP[20]) );
  FA_876 FAI_21 ( .A(A[20]), .B(B[20]), .Ci(CTMP[20]), .S(S[20]), .Co(CTMP[21]) );
  FA_875 FAI_22 ( .A(A[21]), .B(B[21]), .Ci(CTMP[21]), .S(S[21]), .Co(CTMP[22]) );
  FA_874 FAI_23 ( .A(A[22]), .B(B[22]), .Ci(CTMP[22]), .S(S[22]), .Co(CTMP[23]) );
  FA_873 FAI_24 ( .A(A[23]), .B(B[23]), .Ci(CTMP[23]), .S(S[23]), .Co(CTMP[24]) );
  FA_872 FAI_25 ( .A(A[24]), .B(B[24]), .Ci(CTMP[24]), .S(S[24]), .Co(CTMP[25]) );
  FA_871 FAI_26 ( .A(A[25]), .B(B[25]), .Ci(CTMP[25]), .S(S[25]), .Co(CTMP[26]) );
  FA_870 FAI_27 ( .A(A[26]), .B(B[26]), .Ci(CTMP[26]), .S(S[26]), .Co(CTMP[27]) );
  FA_869 FAI_28 ( .A(A[27]), .B(B[27]), .Ci(CTMP[27]), .S(S[27]), .Co(CTMP[28]) );
  FA_868 FAI_29 ( .A(A[28]), .B(B[28]), .Ci(CTMP[28]), .S(S[28]), .Co(CTMP[29]) );
  FA_867 FAI_30 ( .A(A[29]), .B(B[29]), .Ci(CTMP[29]), .S(S[29]), .Co(CTMP[30]) );
  FA_866 FAI_31 ( .A(A[30]), .B(B[30]), .Ci(CTMP[30]), .S(S[30]), .Co(CTMP[31]) );
  FA_865 FAI_32 ( .A(A[31]), .B(B[31]), .Ci(CTMP[31]), .S(S[31]), .Co(CTMP[32]) );
  FA_864 FAI_33 ( .A(A[32]), .B(B[32]), .Ci(CTMP[32]), .S(S[32]), .Co(CTMP[33]) );
  FA_863 FAI_34 ( .A(A[33]), .B(B[33]), .Ci(CTMP[33]), .S(S[33]), .Co(CTMP[34]) );
  FA_862 FAI_35 ( .A(A[34]), .B(B[34]), .Ci(CTMP[34]), .S(S[34]), .Co(CTMP[35]) );
  FA_861 FAI_36 ( .A(A[35]), .B(B[35]), .Ci(CTMP[35]), .S(S[35]), .Co(CTMP[36]) );
  FA_860 FAI_37 ( .A(A[36]), .B(B[36]), .Ci(CTMP[36]), .S(S[36]), .Co(CTMP[37]) );
  FA_859 FAI_38 ( .A(A[37]), .B(B[37]), .Ci(CTMP[37]), .S(S[37]), .Co(CTMP[38]) );
  FA_858 FAI_39 ( .A(A[38]), .B(B[38]), .Ci(CTMP[38]), .S(S[38]), .Co(CTMP[39]) );
  FA_857 FAI_40 ( .A(A[39]), .B(B[39]), .Ci(CTMP[39]), .S(S[39]), .Co(CTMP[40]) );
  FA_856 FAI_41 ( .A(A[40]), .B(B[40]), .Ci(CTMP[40]), .S(S[40]), .Co(CTMP[41]) );
  FA_855 FAI_42 ( .A(A[41]), .B(B[41]), .Ci(CTMP[41]), .S(S[41]), .Co(CTMP[42]) );
  FA_854 FAI_43 ( .A(A[42]), .B(B[42]), .Ci(CTMP[42]), .S(S[42]), .Co(CTMP[43]) );
  FA_853 FAI_44 ( .A(A[43]), .B(B[43]), .Ci(CTMP[43]), .S(S[43]), .Co(CTMP[44]) );
  FA_852 FAI_45 ( .A(A[44]), .B(B[44]), .Ci(CTMP[44]), .S(S[44]), .Co(CTMP[45]) );
  FA_851 FAI_46 ( .A(A[45]), .B(B[45]), .Ci(CTMP[45]), .S(S[45]), .Co(CTMP[46]) );
  FA_850 FAI_47 ( .A(A[46]), .B(B[46]), .Ci(CTMP[46]), .S(S[46]), .Co(CTMP[47]) );
  FA_849 FAI_48 ( .A(A[47]), .B(B[47]), .Ci(CTMP[47]), .S(S[47]), .Co(CTMP[48]) );
  FA_848 FAI_49 ( .A(A[48]), .B(B[48]), .Ci(CTMP[48]), .S(S[48]), .Co(CTMP[49]) );
  FA_847 FAI_50 ( .A(A[49]), .B(B[49]), .Ci(CTMP[49]), .S(S[49]), .Co(CTMP[50]) );
  FA_846 FAI_51 ( .A(A[50]), .B(B[50]), .Ci(CTMP[50]), .S(S[50]), .Co(CTMP[51]) );
  FA_845 FAI_52 ( .A(A[51]), .B(B[51]), .Ci(CTMP[51]), .S(S[51]), .Co(CTMP[52]) );
  FA_844 FAI_53 ( .A(A[52]), .B(B[52]), .Ci(CTMP[52]), .S(S[52]), .Co(CTMP[53]) );
  FA_843 FAI_54 ( .A(A[53]), .B(B[53]), .Ci(CTMP[53]), .S(S[53]), .Co(CTMP[54]) );
  FA_842 FAI_55 ( .A(A[54]), .B(B[54]), .Ci(CTMP[54]), .S(S[54]), .Co(CTMP[55]) );
  FA_841 FAI_56 ( .A(A[55]), .B(B[55]), .Ci(CTMP[55]), .S(S[55]), .Co(CTMP[56]) );
  FA_840 FAI_57 ( .A(A[56]), .B(B[56]), .Ci(CTMP[56]), .S(S[56]), .Co(CTMP[57]) );
  FA_839 FAI_58 ( .A(A[57]), .B(B[57]), .Ci(CTMP[57]), .S(S[57]), .Co(CTMP[58]) );
  FA_838 FAI_59 ( .A(A[58]), .B(B[58]), .Ci(CTMP[58]), .S(S[58]), .Co(CTMP[59]) );
  FA_837 FAI_60 ( .A(A[59]), .B(B[59]), .Ci(CTMP[59]), .S(S[59]), .Co(CTMP[60]) );
  FA_836 FAI_61 ( .A(A[60]), .B(B[60]), .Ci(CTMP[60]), .S(S[60]), .Co(CTMP[61]) );
  FA_835 FAI_62 ( .A(A[61]), .B(B[61]), .Ci(CTMP[61]), .S(S[61]), .Co(CTMP[62]) );
  FA_834 FAI_63 ( .A(A[62]), .B(B[62]), .Ci(CTMP[62]), .S(S[62]), .Co(CTMP[63]) );
  FA_833 FAI_64 ( .A(A[63]), .B(B[63]), .Ci(CTMP[63]), .S(S[63]), .Co(Co) );
endmodule


module booth_mul_row_N64_RADIX3_14 ( prevA, prevSum, encoderIn, nextA, nextSum
 );
  input [63:0] prevA;
  input [63:0] prevSum;
  input [2:0] encoderIn;
  output [63:0] nextA;
  output [63:0] nextSum;
  wire   n4, n5;
  wire   [2:0] encoder_to_mux;
  wire   [63:0] plus2A_s;
  wire   [63:0] minus2A_s;
  wire   [63:0] minus4A_s;
  tri   [63:0] mux_to_adder;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign nextA[51] = n4;
  assign nextA[39] = n5;
  assign nextA[0] = 1'b0;

  encoder_N64_RADIX3_14 encoder_1 ( .X(encoderIn), .Z(encoder_to_mux) );
  ShiftnCompl_N64_14 ShiftnCompl_1 ( .plusA(prevA), .plus2A_out({
        plus2A_s[63:1], SYNOPSYS_UNCONNECTED__0}), .minus2A_out(minus2A_s), 
        .plus4A_out({nextA[63:52], n4, nextA[50:40], n5, nextA[38:1], 
        SYNOPSYS_UNCONNECTED__1}), .minus4A_out(minus4A_s) );
  MUX_GENERIC_N64_RADIX3_14 mux_1 ( .plusA({plus2A_s[63:1], 1'b0}), .minusA(
        minus2A_s), .plus2A({nextA[63:52], n4, nextA[50:40], n5, nextA[38:1], 
        1'b0}), .minus2A(minus4A_s), .SEL(encoder_to_mux), .Y(mux_to_adder) );
  RCA_N64_14 rca_1 ( .A(mux_to_adder), .B(prevSum), .Ci(1'b0), .S(nextSum) );
endmodule


module encoder_N64_RADIX3_13 ( X, Z );
  input [2:0] X;
  output [2:0] Z;
  wire   n5, n7, n8;

  OAI22_X1 U1 ( .A1(n8), .A2(n5), .B1(X[2]), .B2(n7), .ZN(Z[1]) );
  INV_X1 U2 ( .A(X[2]), .ZN(n5) );
  AOI21_X1 U3 ( .B1(n8), .B2(n7), .A(X[2]), .ZN(Z[0]) );
  OAI21_X1 U4 ( .B1(X[1]), .B2(X[0]), .A(n7), .ZN(n8) );
  AND3_X1 U5 ( .A1(X[2]), .A2(n7), .A3(n8), .ZN(Z[2]) );
  NAND2_X1 U6 ( .A1(X[1]), .A2(X[0]), .ZN(n7) );
endmodule


module shifter_N64_26 ( \input , shiftLeftOnePos );
  input [63:0] \input ;
  output [63:0] shiftLeftOnePos;
  wire   \input[62] , \input[61] , \input[60] , \input[59] , \input[58] ,
         \input[57] , \input[56] , \input[55] , \input[54] , \input[53] ,
         \input[52] , \input[51] , \input[50] , \input[49] , \input[48] ,
         \input[47] , \input[46] , \input[45] , \input[44] , \input[43] ,
         \input[42] , \input[41] , \input[40] , \input[39] , \input[38] ,
         \input[37] , \input[36] , \input[35] , \input[34] , \input[33] ,
         \input[32] , \input[31] , \input[30] , \input[29] , \input[28] ,
         \input[27] , \input[26] , \input[25] , \input[24] , \input[23] ,
         \input[22] , \input[21] , \input[20] , \input[19] , \input[18] ,
         \input[17] , \input[16] , \input[15] , \input[14] , \input[13] ,
         \input[12] , \input[11] , \input[10] , \input[9] , \input[8] ,
         \input[7] , \input[6] , \input[5] , \input[4] , \input[3] ,
         \input[2] , \input[1] , \input[0] ;
  assign shiftLeftOnePos[0] = 1'b0;
  assign shiftLeftOnePos[63] = \input[62] ;
  assign \input[62]  = \input  [62];
  assign shiftLeftOnePos[62] = \input[61] ;
  assign \input[61]  = \input  [61];
  assign shiftLeftOnePos[61] = \input[60] ;
  assign \input[60]  = \input  [60];
  assign shiftLeftOnePos[60] = \input[59] ;
  assign \input[59]  = \input  [59];
  assign shiftLeftOnePos[59] = \input[58] ;
  assign \input[58]  = \input  [58];
  assign shiftLeftOnePos[58] = \input[57] ;
  assign \input[57]  = \input  [57];
  assign shiftLeftOnePos[57] = \input[56] ;
  assign \input[56]  = \input  [56];
  assign shiftLeftOnePos[56] = \input[55] ;
  assign \input[55]  = \input  [55];
  assign shiftLeftOnePos[55] = \input[54] ;
  assign \input[54]  = \input  [54];
  assign shiftLeftOnePos[54] = \input[53] ;
  assign \input[53]  = \input  [53];
  assign shiftLeftOnePos[53] = \input[52] ;
  assign \input[52]  = \input  [52];
  assign shiftLeftOnePos[52] = \input[51] ;
  assign \input[51]  = \input  [51];
  assign shiftLeftOnePos[51] = \input[50] ;
  assign \input[50]  = \input  [50];
  assign shiftLeftOnePos[50] = \input[49] ;
  assign \input[49]  = \input  [49];
  assign shiftLeftOnePos[49] = \input[48] ;
  assign \input[48]  = \input  [48];
  assign shiftLeftOnePos[48] = \input[47] ;
  assign \input[47]  = \input  [47];
  assign shiftLeftOnePos[47] = \input[46] ;
  assign \input[46]  = \input  [46];
  assign shiftLeftOnePos[46] = \input[45] ;
  assign \input[45]  = \input  [45];
  assign shiftLeftOnePos[45] = \input[44] ;
  assign \input[44]  = \input  [44];
  assign shiftLeftOnePos[44] = \input[43] ;
  assign \input[43]  = \input  [43];
  assign shiftLeftOnePos[43] = \input[42] ;
  assign \input[42]  = \input  [42];
  assign shiftLeftOnePos[42] = \input[41] ;
  assign \input[41]  = \input  [41];
  assign shiftLeftOnePos[41] = \input[40] ;
  assign \input[40]  = \input  [40];
  assign shiftLeftOnePos[40] = \input[39] ;
  assign \input[39]  = \input  [39];
  assign shiftLeftOnePos[39] = \input[38] ;
  assign \input[38]  = \input  [38];
  assign shiftLeftOnePos[38] = \input[37] ;
  assign \input[37]  = \input  [37];
  assign shiftLeftOnePos[37] = \input[36] ;
  assign \input[36]  = \input  [36];
  assign shiftLeftOnePos[36] = \input[35] ;
  assign \input[35]  = \input  [35];
  assign shiftLeftOnePos[35] = \input[34] ;
  assign \input[34]  = \input  [34];
  assign shiftLeftOnePos[34] = \input[33] ;
  assign \input[33]  = \input  [33];
  assign shiftLeftOnePos[33] = \input[32] ;
  assign \input[32]  = \input  [32];
  assign shiftLeftOnePos[32] = \input[31] ;
  assign \input[31]  = \input  [31];
  assign shiftLeftOnePos[31] = \input[30] ;
  assign \input[30]  = \input  [30];
  assign shiftLeftOnePos[30] = \input[29] ;
  assign \input[29]  = \input  [29];
  assign shiftLeftOnePos[29] = \input[28] ;
  assign \input[28]  = \input  [28];
  assign shiftLeftOnePos[28] = \input[27] ;
  assign \input[27]  = \input  [27];
  assign shiftLeftOnePos[27] = \input[26] ;
  assign \input[26]  = \input  [26];
  assign shiftLeftOnePos[26] = \input[25] ;
  assign \input[25]  = \input  [25];
  assign shiftLeftOnePos[25] = \input[24] ;
  assign \input[24]  = \input  [24];
  assign shiftLeftOnePos[24] = \input[23] ;
  assign \input[23]  = \input  [23];
  assign shiftLeftOnePos[23] = \input[22] ;
  assign \input[22]  = \input  [22];
  assign shiftLeftOnePos[22] = \input[21] ;
  assign \input[21]  = \input  [21];
  assign shiftLeftOnePos[21] = \input[20] ;
  assign \input[20]  = \input  [20];
  assign shiftLeftOnePos[20] = \input[19] ;
  assign \input[19]  = \input  [19];
  assign shiftLeftOnePos[19] = \input[18] ;
  assign \input[18]  = \input  [18];
  assign shiftLeftOnePos[18] = \input[17] ;
  assign \input[17]  = \input  [17];
  assign shiftLeftOnePos[17] = \input[16] ;
  assign \input[16]  = \input  [16];
  assign shiftLeftOnePos[16] = \input[15] ;
  assign \input[15]  = \input  [15];
  assign shiftLeftOnePos[15] = \input[14] ;
  assign \input[14]  = \input  [14];
  assign shiftLeftOnePos[14] = \input[13] ;
  assign \input[13]  = \input  [13];
  assign shiftLeftOnePos[13] = \input[12] ;
  assign \input[12]  = \input  [12];
  assign shiftLeftOnePos[12] = \input[11] ;
  assign \input[11]  = \input  [11];
  assign shiftLeftOnePos[11] = \input[10] ;
  assign \input[10]  = \input  [10];
  assign shiftLeftOnePos[10] = \input[9] ;
  assign \input[9]  = \input  [9];
  assign shiftLeftOnePos[9] = \input[8] ;
  assign \input[8]  = \input  [8];
  assign shiftLeftOnePos[8] = \input[7] ;
  assign \input[7]  = \input  [7];
  assign shiftLeftOnePos[7] = \input[6] ;
  assign \input[6]  = \input  [6];
  assign shiftLeftOnePos[6] = \input[5] ;
  assign \input[5]  = \input  [5];
  assign shiftLeftOnePos[5] = \input[4] ;
  assign \input[4]  = \input  [4];
  assign shiftLeftOnePos[4] = \input[3] ;
  assign \input[3]  = \input  [3];
  assign shiftLeftOnePos[3] = \input[2] ;
  assign \input[2]  = \input  [2];
  assign shiftLeftOnePos[2] = \input[1] ;
  assign \input[1]  = \input  [1];
  assign shiftLeftOnePos[1] = \input[0] ;
  assign \input[0]  = \input  [0];

endmodule


module shifter_N64_25 ( \input , shiftLeftOnePos );
  input [63:0] \input ;
  output [63:0] shiftLeftOnePos;
  wire   \input[62] , \input[61] , \input[60] , \input[59] , \input[58] ,
         \input[57] , \input[56] , \input[55] , \input[54] , \input[53] ,
         \input[52] , \input[51] , \input[50] , \input[49] , \input[48] ,
         \input[47] , \input[46] , \input[45] , \input[44] , \input[43] ,
         \input[42] , \input[41] , \input[40] , \input[39] , \input[38] ,
         \input[37] , \input[36] , \input[35] , \input[34] , \input[33] ,
         \input[32] , \input[31] , \input[30] , \input[29] , \input[28] ,
         \input[27] , \input[26] , \input[25] , \input[24] , \input[23] ,
         \input[22] , \input[21] , \input[20] , \input[19] , \input[18] ,
         \input[17] , \input[16] , \input[15] , \input[14] , \input[13] ,
         \input[12] , \input[11] , \input[10] , \input[9] , \input[8] ,
         \input[7] , \input[6] , \input[5] , \input[4] , \input[3] ,
         \input[2] , \input[1] , \input[0] ;
  assign shiftLeftOnePos[0] = 1'b0;
  assign shiftLeftOnePos[63] = \input[62] ;
  assign \input[62]  = \input  [62];
  assign shiftLeftOnePos[62] = \input[61] ;
  assign \input[61]  = \input  [61];
  assign shiftLeftOnePos[61] = \input[60] ;
  assign \input[60]  = \input  [60];
  assign shiftLeftOnePos[60] = \input[59] ;
  assign \input[59]  = \input  [59];
  assign shiftLeftOnePos[59] = \input[58] ;
  assign \input[58]  = \input  [58];
  assign shiftLeftOnePos[58] = \input[57] ;
  assign \input[57]  = \input  [57];
  assign shiftLeftOnePos[57] = \input[56] ;
  assign \input[56]  = \input  [56];
  assign shiftLeftOnePos[56] = \input[55] ;
  assign \input[55]  = \input  [55];
  assign shiftLeftOnePos[55] = \input[54] ;
  assign \input[54]  = \input  [54];
  assign shiftLeftOnePos[54] = \input[53] ;
  assign \input[53]  = \input  [53];
  assign shiftLeftOnePos[53] = \input[52] ;
  assign \input[52]  = \input  [52];
  assign shiftLeftOnePos[52] = \input[51] ;
  assign \input[51]  = \input  [51];
  assign shiftLeftOnePos[51] = \input[50] ;
  assign \input[50]  = \input  [50];
  assign shiftLeftOnePos[50] = \input[49] ;
  assign \input[49]  = \input  [49];
  assign shiftLeftOnePos[49] = \input[48] ;
  assign \input[48]  = \input  [48];
  assign shiftLeftOnePos[48] = \input[47] ;
  assign \input[47]  = \input  [47];
  assign shiftLeftOnePos[47] = \input[46] ;
  assign \input[46]  = \input  [46];
  assign shiftLeftOnePos[46] = \input[45] ;
  assign \input[45]  = \input  [45];
  assign shiftLeftOnePos[45] = \input[44] ;
  assign \input[44]  = \input  [44];
  assign shiftLeftOnePos[44] = \input[43] ;
  assign \input[43]  = \input  [43];
  assign shiftLeftOnePos[43] = \input[42] ;
  assign \input[42]  = \input  [42];
  assign shiftLeftOnePos[42] = \input[41] ;
  assign \input[41]  = \input  [41];
  assign shiftLeftOnePos[41] = \input[40] ;
  assign \input[40]  = \input  [40];
  assign shiftLeftOnePos[40] = \input[39] ;
  assign \input[39]  = \input  [39];
  assign shiftLeftOnePos[39] = \input[38] ;
  assign \input[38]  = \input  [38];
  assign shiftLeftOnePos[38] = \input[37] ;
  assign \input[37]  = \input  [37];
  assign shiftLeftOnePos[37] = \input[36] ;
  assign \input[36]  = \input  [36];
  assign shiftLeftOnePos[36] = \input[35] ;
  assign \input[35]  = \input  [35];
  assign shiftLeftOnePos[35] = \input[34] ;
  assign \input[34]  = \input  [34];
  assign shiftLeftOnePos[34] = \input[33] ;
  assign \input[33]  = \input  [33];
  assign shiftLeftOnePos[33] = \input[32] ;
  assign \input[32]  = \input  [32];
  assign shiftLeftOnePos[32] = \input[31] ;
  assign \input[31]  = \input  [31];
  assign shiftLeftOnePos[31] = \input[30] ;
  assign \input[30]  = \input  [30];
  assign shiftLeftOnePos[30] = \input[29] ;
  assign \input[29]  = \input  [29];
  assign shiftLeftOnePos[29] = \input[28] ;
  assign \input[28]  = \input  [28];
  assign shiftLeftOnePos[28] = \input[27] ;
  assign \input[27]  = \input  [27];
  assign shiftLeftOnePos[27] = \input[26] ;
  assign \input[26]  = \input  [26];
  assign shiftLeftOnePos[26] = \input[25] ;
  assign \input[25]  = \input  [25];
  assign shiftLeftOnePos[25] = \input[24] ;
  assign \input[24]  = \input  [24];
  assign shiftLeftOnePos[24] = \input[23] ;
  assign \input[23]  = \input  [23];
  assign shiftLeftOnePos[23] = \input[22] ;
  assign \input[22]  = \input  [22];
  assign shiftLeftOnePos[22] = \input[21] ;
  assign \input[21]  = \input  [21];
  assign shiftLeftOnePos[21] = \input[20] ;
  assign \input[20]  = \input  [20];
  assign shiftLeftOnePos[20] = \input[19] ;
  assign \input[19]  = \input  [19];
  assign shiftLeftOnePos[19] = \input[18] ;
  assign \input[18]  = \input  [18];
  assign shiftLeftOnePos[18] = \input[17] ;
  assign \input[17]  = \input  [17];
  assign shiftLeftOnePos[17] = \input[16] ;
  assign \input[16]  = \input  [16];
  assign shiftLeftOnePos[16] = \input[15] ;
  assign \input[15]  = \input  [15];
  assign shiftLeftOnePos[15] = \input[14] ;
  assign \input[14]  = \input  [14];
  assign shiftLeftOnePos[14] = \input[13] ;
  assign \input[13]  = \input  [13];
  assign shiftLeftOnePos[13] = \input[12] ;
  assign \input[12]  = \input  [12];
  assign shiftLeftOnePos[12] = \input[11] ;
  assign \input[11]  = \input  [11];
  assign shiftLeftOnePos[11] = \input[10] ;
  assign \input[10]  = \input  [10];
  assign shiftLeftOnePos[10] = \input[9] ;
  assign \input[9]  = \input  [9];
  assign shiftLeftOnePos[9] = \input[8] ;
  assign \input[8]  = \input  [8];
  assign shiftLeftOnePos[8] = \input[7] ;
  assign \input[7]  = \input  [7];
  assign shiftLeftOnePos[7] = \input[6] ;
  assign \input[6]  = \input  [6];
  assign shiftLeftOnePos[6] = \input[5] ;
  assign \input[5]  = \input  [5];
  assign shiftLeftOnePos[5] = \input[4] ;
  assign \input[4]  = \input  [4];
  assign shiftLeftOnePos[4] = \input[3] ;
  assign \input[3]  = \input  [3];
  assign shiftLeftOnePos[3] = \input[2] ;
  assign \input[2]  = \input  [2];
  assign shiftLeftOnePos[2] = \input[1] ;
  assign \input[1]  = \input  [1];
  assign shiftLeftOnePos[1] = \input[0] ;
  assign \input[0]  = \input  [0];

endmodule


module complementer_N64_26_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n190, n191, n192, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n189, n193;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U81 ( .A(n190), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U82 ( .A(n192), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U84 ( .A(n195), .B(B[63]), .Z(DIFF[63]) );
  XOR2_X1 U85 ( .A(n196), .B(B[62]), .Z(DIFF[62]) );
  XOR2_X1 U86 ( .A(n194), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U87 ( .A(n198), .B(B[59]), .Z(DIFF[59]) );
  XOR2_X1 U88 ( .A(n201), .B(B[58]), .Z(DIFF[58]) );
  XOR2_X1 U89 ( .A(n200), .B(B[57]), .Z(DIFF[57]) );
  XOR2_X1 U90 ( .A(n202), .B(B[55]), .Z(DIFF[55]) );
  XOR2_X1 U91 ( .A(n205), .B(B[54]), .Z(DIFF[54]) );
  XOR2_X1 U92 ( .A(n204), .B(B[53]), .Z(DIFF[53]) );
  XOR2_X1 U93 ( .A(n206), .B(B[51]), .Z(DIFF[51]) );
  XOR2_X1 U94 ( .A(n209), .B(B[50]), .Z(DIFF[50]) );
  XOR2_X1 U95 ( .A(n208), .B(B[49]), .Z(DIFF[49]) );
  XOR2_X1 U96 ( .A(n212), .B(B[47]), .Z(DIFF[47]) );
  XOR2_X1 U97 ( .A(n215), .B(B[46]), .Z(DIFF[46]) );
  XOR2_X1 U98 ( .A(n214), .B(B[45]), .Z(DIFF[45]) );
  XOR2_X1 U99 ( .A(n216), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U100 ( .A(n219), .B(B[42]), .Z(DIFF[42]) );
  XOR2_X1 U101 ( .A(n218), .B(B[41]), .Z(DIFF[41]) );
  XOR2_X1 U102 ( .A(n211), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U103 ( .A(n220), .B(B[39]), .Z(DIFF[39]) );
  XOR2_X1 U104 ( .A(n223), .B(B[38]), .Z(DIFF[38]) );
  XOR2_X1 U105 ( .A(n222), .B(B[37]), .Z(DIFF[37]) );
  XOR2_X1 U106 ( .A(n224), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U107 ( .A(n227), .B(B[34]), .Z(DIFF[34]) );
  XOR2_X1 U108 ( .A(n226), .B(B[33]), .Z(DIFF[33]) );
  XOR2_X1 U109 ( .A(n228), .B(B[31]), .Z(DIFF[31]) );
  XOR2_X1 U110 ( .A(n231), .B(B[30]), .Z(DIFF[30]) );
  XOR2_X1 U111 ( .A(n230), .B(B[29]), .Z(DIFF[29]) );
  XOR2_X1 U112 ( .A(n233), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U113 ( .A(n236), .B(B[26]), .Z(DIFF[26]) );
  XOR2_X1 U114 ( .A(n235), .B(B[25]), .Z(DIFF[25]) );
  XOR2_X1 U115 ( .A(n237), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U116 ( .A(n240), .B(B[22]), .Z(DIFF[22]) );
  XOR2_X1 U117 ( .A(n239), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U118 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U119 ( .A(n241), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U120 ( .A(n244), .B(B[18]), .Z(DIFF[18]) );
  XOR2_X1 U121 ( .A(n243), .B(B[17]), .Z(DIFF[17]) );
  XOR2_X1 U122 ( .A(n245), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U123 ( .A(n248), .B(B[14]), .Z(DIFF[14]) );
  XOR2_X1 U124 ( .A(n247), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U125 ( .A(n249), .B(B[11]), .Z(DIFF[11]) );
  XOR2_X1 U126 ( .A(n251), .B(B[10]), .Z(DIFF[10]) );
  NOR2_X1 U1 ( .A1(B[43]), .A2(n216), .ZN(n217) );
  NAND2_X1 U2 ( .A1(n197), .A2(n193), .ZN(n196) );
  OR3_X1 U3 ( .A1(B[53]), .A2(B[54]), .A3(n204), .ZN(n202) );
  OR3_X1 U4 ( .A1(B[43]), .A2(B[44]), .A3(n216), .ZN(n214) );
  OR2_X1 U5 ( .A1(n204), .A2(B[53]), .ZN(n205) );
  OR2_X1 U6 ( .A1(n208), .A2(B[49]), .ZN(n209) );
  NOR2_X1 U7 ( .A1(B[59]), .A2(n198), .ZN(n199) );
  NOR3_X1 U8 ( .A1(B[59]), .A2(B[60]), .A3(n198), .ZN(n197) );
  NOR2_X1 U9 ( .A1(B[47]), .A2(n212), .ZN(n213) );
  NOR2_X1 U10 ( .A1(B[55]), .A2(n202), .ZN(n203) );
  NOR2_X1 U11 ( .A1(B[51]), .A2(n206), .ZN(n207) );
  NOR2_X1 U12 ( .A1(B[39]), .A2(n220), .ZN(n221) );
  OR3_X1 U13 ( .A1(B[45]), .A2(B[46]), .A3(n214), .ZN(n212) );
  OR3_X1 U14 ( .A1(B[57]), .A2(B[58]), .A3(n200), .ZN(n198) );
  OR3_X1 U15 ( .A1(B[49]), .A2(B[50]), .A3(n208), .ZN(n206) );
  OR3_X1 U16 ( .A1(B[41]), .A2(B[42]), .A3(n218), .ZN(n216) );
  OR3_X1 U17 ( .A1(B[47]), .A2(B[48]), .A3(n212), .ZN(n208) );
  OR3_X1 U18 ( .A1(B[55]), .A2(B[56]), .A3(n202), .ZN(n200) );
  OR3_X1 U19 ( .A1(B[51]), .A2(B[52]), .A3(n206), .ZN(n204) );
  OR3_X1 U20 ( .A1(B[39]), .A2(B[40]), .A3(n220), .ZN(n218) );
  XNOR2_X1 U21 ( .A(B[44]), .B(n217), .ZN(DIFF[44]) );
  XNOR2_X1 U22 ( .A(B[56]), .B(n203), .ZN(DIFF[56]) );
  XNOR2_X1 U23 ( .A(B[52]), .B(n207), .ZN(DIFF[52]) );
  XNOR2_X1 U24 ( .A(B[48]), .B(n213), .ZN(DIFF[48]) );
  XNOR2_X1 U25 ( .A(B[40]), .B(n221), .ZN(DIFF[40]) );
  OR2_X1 U26 ( .A1(n214), .A2(B[45]), .ZN(n215) );
  OR2_X1 U27 ( .A1(n200), .A2(B[57]), .ZN(n201) );
  OR2_X1 U28 ( .A1(n218), .A2(B[41]), .ZN(n219) );
  XNOR2_X1 U29 ( .A(n197), .B(B[61]), .ZN(DIFF[61]) );
  XNOR2_X1 U30 ( .A(B[60]), .B(n199), .ZN(DIFF[60]) );
  OR2_X1 U31 ( .A1(n196), .A2(B[62]), .ZN(n195) );
  OR3_X1 U32 ( .A1(B[37]), .A2(B[38]), .A3(n222), .ZN(n220) );
  XNOR2_X1 U33 ( .A(B[36]), .B(n225), .ZN(DIFF[36]) );
  OR2_X1 U34 ( .A1(n222), .A2(B[37]), .ZN(n223) );
  NOR2_X1 U35 ( .A1(B[11]), .A2(n249), .ZN(n250) );
  NOR2_X1 U36 ( .A1(B[7]), .A2(n192), .ZN(n191) );
  OR3_X1 U37 ( .A1(B[10]), .A2(B[9]), .A3(n190), .ZN(n249) );
  OR3_X1 U38 ( .A1(B[7]), .A2(B[8]), .A3(n192), .ZN(n190) );
  XNOR2_X1 U39 ( .A(B[12]), .B(n250), .ZN(DIFF[12]) );
  XNOR2_X1 U40 ( .A(B[8]), .B(n191), .ZN(DIFF[8]) );
  NOR2_X1 U41 ( .A1(B[31]), .A2(n228), .ZN(n229) );
  NOR2_X1 U42 ( .A1(B[27]), .A2(n233), .ZN(n234) );
  NOR2_X1 U43 ( .A1(B[23]), .A2(n237), .ZN(n238) );
  NOR2_X1 U44 ( .A1(B[19]), .A2(n241), .ZN(n242) );
  NOR2_X1 U45 ( .A1(B[15]), .A2(n245), .ZN(n246) );
  OR3_X1 U46 ( .A1(B[29]), .A2(B[30]), .A3(n230), .ZN(n228) );
  OR3_X1 U47 ( .A1(B[25]), .A2(B[26]), .A3(n235), .ZN(n233) );
  OR3_X1 U48 ( .A1(B[21]), .A2(B[22]), .A3(n239), .ZN(n237) );
  OR3_X1 U49 ( .A1(B[17]), .A2(B[18]), .A3(n243), .ZN(n241) );
  OR3_X1 U50 ( .A1(B[13]), .A2(B[14]), .A3(n247), .ZN(n245) );
  OR3_X1 U51 ( .A1(B[31]), .A2(B[32]), .A3(n228), .ZN(n226) );
  OR3_X1 U52 ( .A1(B[27]), .A2(B[28]), .A3(n233), .ZN(n230) );
  OR3_X1 U53 ( .A1(B[23]), .A2(B[24]), .A3(n237), .ZN(n235) );
  OR3_X1 U54 ( .A1(B[19]), .A2(B[20]), .A3(n241), .ZN(n239) );
  OR3_X1 U55 ( .A1(B[15]), .A2(B[16]), .A3(n245), .ZN(n243) );
  OR3_X1 U56 ( .A1(B[11]), .A2(B[12]), .A3(n249), .ZN(n247) );
  XNOR2_X1 U57 ( .A(B[32]), .B(n229), .ZN(DIFF[32]) );
  XNOR2_X1 U58 ( .A(B[28]), .B(n234), .ZN(DIFF[28]) );
  XNOR2_X1 U59 ( .A(B[24]), .B(n238), .ZN(DIFF[24]) );
  XNOR2_X1 U60 ( .A(B[20]), .B(n242), .ZN(DIFF[20]) );
  XNOR2_X1 U61 ( .A(B[16]), .B(n246), .ZN(DIFF[16]) );
  OR2_X1 U62 ( .A1(n226), .A2(B[33]), .ZN(n227) );
  OR2_X1 U63 ( .A1(n230), .A2(B[29]), .ZN(n231) );
  OR2_X1 U64 ( .A1(n235), .A2(B[25]), .ZN(n236) );
  OR2_X1 U65 ( .A1(n239), .A2(B[21]), .ZN(n240) );
  OR2_X1 U66 ( .A1(n243), .A2(B[17]), .ZN(n244) );
  OR2_X1 U67 ( .A1(n247), .A2(B[13]), .ZN(n248) );
  OR2_X1 U68 ( .A1(n190), .A2(B[9]), .ZN(n251) );
  NOR2_X1 U69 ( .A1(B[35]), .A2(n224), .ZN(n225) );
  OR3_X1 U70 ( .A1(B[33]), .A2(B[34]), .A3(n226), .ZN(n224) );
  OR3_X1 U71 ( .A1(B[35]), .A2(B[36]), .A3(n224), .ZN(n222) );
  XNOR2_X1 U72 ( .A(n189), .B(B[6]), .ZN(DIFF[6]) );
  NOR2_X1 U73 ( .A1(n194), .A2(B[5]), .ZN(n189) );
  OR3_X1 U74 ( .A1(B[5]), .A2(B[6]), .A3(n194), .ZN(n192) );
  NOR2_X1 U75 ( .A1(B[3]), .A2(n211), .ZN(n210) );
  OR3_X1 U76 ( .A1(B[3]), .A2(B[4]), .A3(n211), .ZN(n194) );
  XNOR2_X1 U77 ( .A(B[4]), .B(n210), .ZN(DIFF[4]) );
  XNOR2_X1 U78 ( .A(B[2]), .B(n232), .ZN(DIFF[2]) );
  OR3_X1 U79 ( .A1(B[1]), .A2(B[2]), .A3(\B[0] ), .ZN(n211) );
  NOR2_X1 U80 ( .A1(\B[0] ), .A2(B[1]), .ZN(n232) );
  INV_X1 U83 ( .A(B[61]), .ZN(n193) );
endmodule


module complementer_N64_26 ( \input , complement2 );
  input [63:0] \input ;
  output [63:0] complement2;


  complementer_N64_26_DW01_sub_0 sub_add_31_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(\input ), .CI(1'b0), .DIFF(complement2) );
endmodule


module complementer_N64_25_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n190, n191, n192, n193, n194, n196, n197, n198, n199, n200,
         n202, n203, n204, n206, n207, n208, n210, n211, n212, n213, n214,
         n216, n217, n218, n220, n221, n222, n224, n225, n226, n228, n229,
         n230, n232, n233, n234, n235, n237, n238, n239, n241, n242, n243,
         n245, n246, n247, n249, n250, n189, n195, n201, n205, n209, n215,
         n219, n223, n227, n231, n236, n240, n244, n248, n251;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U81 ( .A(n190), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U82 ( .A(n192), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U83 ( .A(n193), .B(B[6]), .Z(DIFF[6]) );
  XOR2_X1 U85 ( .A(n196), .B(B[62]), .Z(DIFF[62]) );
  XOR2_X1 U86 ( .A(n194), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U87 ( .A(n198), .B(B[59]), .Z(DIFF[59]) );
  XOR2_X1 U89 ( .A(n200), .B(B[57]), .Z(DIFF[57]) );
  XOR2_X1 U90 ( .A(n202), .B(B[55]), .Z(DIFF[55]) );
  XOR2_X1 U92 ( .A(n204), .B(B[53]), .Z(DIFF[53]) );
  XOR2_X1 U93 ( .A(n206), .B(B[51]), .Z(DIFF[51]) );
  XOR2_X1 U95 ( .A(n208), .B(B[49]), .Z(DIFF[49]) );
  XOR2_X1 U96 ( .A(n212), .B(B[47]), .Z(DIFF[47]) );
  XOR2_X1 U98 ( .A(n214), .B(B[45]), .Z(DIFF[45]) );
  XOR2_X1 U99 ( .A(n216), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U101 ( .A(n218), .B(B[41]), .Z(DIFF[41]) );
  XOR2_X1 U102 ( .A(n211), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U103 ( .A(n220), .B(B[39]), .Z(DIFF[39]) );
  XOR2_X1 U105 ( .A(n222), .B(B[37]), .Z(DIFF[37]) );
  XOR2_X1 U106 ( .A(n224), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U108 ( .A(n226), .B(B[33]), .Z(DIFF[33]) );
  XOR2_X1 U109 ( .A(n228), .B(B[31]), .Z(DIFF[31]) );
  XOR2_X1 U111 ( .A(n230), .B(B[29]), .Z(DIFF[29]) );
  XOR2_X1 U112 ( .A(n233), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U114 ( .A(n235), .B(B[25]), .Z(DIFF[25]) );
  XOR2_X1 U115 ( .A(n237), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U117 ( .A(n239), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U118 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U119 ( .A(n241), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U121 ( .A(n243), .B(B[17]), .Z(DIFF[17]) );
  XOR2_X1 U122 ( .A(n245), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U124 ( .A(n247), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U125 ( .A(n249), .B(B[11]), .Z(DIFF[11]) );
  NOR3_X1 U1 ( .A1(B[59]), .A2(B[60]), .A3(n198), .ZN(n197) );
  XNOR2_X1 U2 ( .A(B[44]), .B(n217), .ZN(DIFF[44]) );
  NOR2_X1 U3 ( .A1(B[43]), .A2(n216), .ZN(n217) );
  NAND2_X1 U4 ( .A1(n197), .A2(n251), .ZN(n196) );
  OR3_X1 U5 ( .A1(B[53]), .A2(B[54]), .A3(n204), .ZN(n202) );
  OR3_X1 U6 ( .A1(B[49]), .A2(B[50]), .A3(n208), .ZN(n206) );
  OR3_X1 U7 ( .A1(B[43]), .A2(B[44]), .A3(n216), .ZN(n214) );
  XNOR2_X1 U8 ( .A(n189), .B(B[54]), .ZN(DIFF[54]) );
  NOR2_X1 U9 ( .A1(n204), .A2(B[53]), .ZN(n189) );
  XNOR2_X1 U10 ( .A(n195), .B(B[50]), .ZN(DIFF[50]) );
  NOR2_X1 U11 ( .A1(n208), .A2(B[49]), .ZN(n195) );
  XNOR2_X1 U12 ( .A(B[60]), .B(n199), .ZN(DIFF[60]) );
  NOR2_X1 U13 ( .A1(B[59]), .A2(n198), .ZN(n199) );
  XOR2_X1 U14 ( .A(n197), .B(n251), .Z(DIFF[61]) );
  XNOR2_X1 U15 ( .A(B[56]), .B(n203), .ZN(DIFF[56]) );
  NOR2_X1 U16 ( .A1(B[55]), .A2(n202), .ZN(n203) );
  XNOR2_X1 U17 ( .A(B[52]), .B(n207), .ZN(DIFF[52]) );
  NOR2_X1 U18 ( .A1(B[51]), .A2(n206), .ZN(n207) );
  XNOR2_X1 U19 ( .A(B[48]), .B(n213), .ZN(DIFF[48]) );
  NOR2_X1 U20 ( .A1(B[47]), .A2(n212), .ZN(n213) );
  XNOR2_X1 U21 ( .A(B[40]), .B(n221), .ZN(DIFF[40]) );
  NOR2_X1 U22 ( .A1(B[39]), .A2(n220), .ZN(n221) );
  OR3_X1 U23 ( .A1(B[45]), .A2(B[46]), .A3(n214), .ZN(n212) );
  OR3_X1 U24 ( .A1(B[57]), .A2(B[58]), .A3(n200), .ZN(n198) );
  OR3_X1 U25 ( .A1(B[41]), .A2(B[42]), .A3(n218), .ZN(n216) );
  OR3_X1 U26 ( .A1(B[47]), .A2(B[48]), .A3(n212), .ZN(n208) );
  OR3_X1 U27 ( .A1(B[55]), .A2(B[56]), .A3(n202), .ZN(n200) );
  OR3_X1 U28 ( .A1(B[51]), .A2(B[52]), .A3(n206), .ZN(n204) );
  OR3_X1 U29 ( .A1(B[39]), .A2(B[40]), .A3(n220), .ZN(n218) );
  XNOR2_X1 U30 ( .A(n201), .B(B[46]), .ZN(DIFF[46]) );
  NOR2_X1 U31 ( .A1(n214), .A2(B[45]), .ZN(n201) );
  XNOR2_X1 U32 ( .A(n205), .B(B[58]), .ZN(DIFF[58]) );
  NOR2_X1 U33 ( .A1(n200), .A2(B[57]), .ZN(n205) );
  XNOR2_X1 U34 ( .A(n209), .B(B[42]), .ZN(DIFF[42]) );
  NOR2_X1 U35 ( .A1(n218), .A2(B[41]), .ZN(n209) );
  XNOR2_X1 U36 ( .A(n215), .B(B[63]), .ZN(DIFF[63]) );
  NOR2_X1 U37 ( .A1(n196), .A2(B[62]), .ZN(n215) );
  XNOR2_X1 U38 ( .A(B[12]), .B(n250), .ZN(DIFF[12]) );
  NOR2_X1 U39 ( .A1(B[11]), .A2(n249), .ZN(n250) );
  OR3_X1 U40 ( .A1(B[10]), .A2(B[9]), .A3(n190), .ZN(n249) );
  XNOR2_X1 U41 ( .A(n219), .B(B[34]), .ZN(DIFF[34]) );
  NOR2_X1 U42 ( .A1(n226), .A2(B[33]), .ZN(n219) );
  XNOR2_X1 U43 ( .A(n223), .B(B[30]), .ZN(DIFF[30]) );
  NOR2_X1 U44 ( .A1(n230), .A2(B[29]), .ZN(n223) );
  XNOR2_X1 U45 ( .A(n227), .B(B[26]), .ZN(DIFF[26]) );
  NOR2_X1 U46 ( .A1(n235), .A2(B[25]), .ZN(n227) );
  XNOR2_X1 U47 ( .A(n231), .B(B[22]), .ZN(DIFF[22]) );
  NOR2_X1 U48 ( .A1(n239), .A2(B[21]), .ZN(n231) );
  XNOR2_X1 U49 ( .A(n236), .B(B[18]), .ZN(DIFF[18]) );
  NOR2_X1 U50 ( .A1(n243), .A2(B[17]), .ZN(n236) );
  XNOR2_X1 U51 ( .A(n240), .B(B[14]), .ZN(DIFF[14]) );
  NOR2_X1 U52 ( .A1(n247), .A2(B[13]), .ZN(n240) );
  XNOR2_X1 U53 ( .A(n244), .B(B[10]), .ZN(DIFF[10]) );
  NOR2_X1 U54 ( .A1(n190), .A2(B[9]), .ZN(n244) );
  XNOR2_X1 U55 ( .A(B[32]), .B(n229), .ZN(DIFF[32]) );
  NOR2_X1 U56 ( .A1(B[31]), .A2(n228), .ZN(n229) );
  XNOR2_X1 U57 ( .A(B[28]), .B(n234), .ZN(DIFF[28]) );
  NOR2_X1 U58 ( .A1(B[27]), .A2(n233), .ZN(n234) );
  XNOR2_X1 U59 ( .A(B[24]), .B(n238), .ZN(DIFF[24]) );
  NOR2_X1 U60 ( .A1(B[23]), .A2(n237), .ZN(n238) );
  XNOR2_X1 U61 ( .A(B[20]), .B(n242), .ZN(DIFF[20]) );
  NOR2_X1 U62 ( .A1(B[19]), .A2(n241), .ZN(n242) );
  XNOR2_X1 U63 ( .A(B[16]), .B(n246), .ZN(DIFF[16]) );
  NOR2_X1 U64 ( .A1(B[15]), .A2(n245), .ZN(n246) );
  OR3_X1 U65 ( .A1(B[13]), .A2(B[14]), .A3(n247), .ZN(n245) );
  OR3_X1 U66 ( .A1(B[17]), .A2(B[18]), .A3(n243), .ZN(n241) );
  OR3_X1 U67 ( .A1(B[21]), .A2(B[22]), .A3(n239), .ZN(n237) );
  OR3_X1 U68 ( .A1(B[25]), .A2(B[26]), .A3(n235), .ZN(n233) );
  OR3_X1 U69 ( .A1(B[29]), .A2(B[30]), .A3(n230), .ZN(n228) );
  OR3_X1 U70 ( .A1(B[11]), .A2(B[12]), .A3(n249), .ZN(n247) );
  OR3_X1 U71 ( .A1(B[15]), .A2(B[16]), .A3(n245), .ZN(n243) );
  OR3_X1 U72 ( .A1(B[19]), .A2(B[20]), .A3(n241), .ZN(n239) );
  OR3_X1 U73 ( .A1(B[23]), .A2(B[24]), .A3(n237), .ZN(n235) );
  OR3_X1 U74 ( .A1(B[27]), .A2(B[28]), .A3(n233), .ZN(n230) );
  OR3_X1 U75 ( .A1(B[31]), .A2(B[32]), .A3(n228), .ZN(n226) );
  XNOR2_X1 U76 ( .A(B[36]), .B(n225), .ZN(DIFF[36]) );
  NOR2_X1 U77 ( .A1(B[35]), .A2(n224), .ZN(n225) );
  OR3_X1 U78 ( .A1(B[33]), .A2(B[34]), .A3(n226), .ZN(n224) );
  OR3_X1 U79 ( .A1(B[37]), .A2(B[38]), .A3(n222), .ZN(n220) );
  OR3_X1 U80 ( .A1(B[35]), .A2(B[36]), .A3(n224), .ZN(n222) );
  XNOR2_X1 U84 ( .A(n248), .B(B[38]), .ZN(DIFF[38]) );
  NOR2_X1 U88 ( .A1(n222), .A2(B[37]), .ZN(n248) );
  XNOR2_X1 U91 ( .A(B[8]), .B(n191), .ZN(DIFF[8]) );
  NOR2_X1 U94 ( .A1(B[7]), .A2(n192), .ZN(n191) );
  OR3_X1 U97 ( .A1(B[7]), .A2(B[8]), .A3(n192), .ZN(n190) );
  XNOR2_X1 U100 ( .A(B[2]), .B(n232), .ZN(DIFF[2]) );
  NOR2_X1 U104 ( .A1(\B[0] ), .A2(B[1]), .ZN(n232) );
  XNOR2_X1 U107 ( .A(B[4]), .B(n210), .ZN(DIFF[4]) );
  NOR2_X1 U110 ( .A1(B[3]), .A2(n211), .ZN(n210) );
  OR3_X1 U113 ( .A1(B[5]), .A2(B[6]), .A3(n194), .ZN(n192) );
  OR3_X1 U116 ( .A1(B[3]), .A2(B[4]), .A3(n211), .ZN(n194) );
  OR2_X1 U120 ( .A1(n194), .A2(B[5]), .ZN(n193) );
  OR3_X1 U123 ( .A1(B[1]), .A2(B[2]), .A3(\B[0] ), .ZN(n211) );
  INV_X1 U126 ( .A(B[61]), .ZN(n251) );
endmodule


module complementer_N64_25 ( \input , complement2 );
  input [63:0] \input ;
  output [63:0] complement2;


  complementer_N64_25_DW01_sub_0 sub_add_31_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(\input ), .CI(1'b0), .DIFF(complement2) );
endmodule


module ShiftnCompl_N64_13 ( plusA, plus2A_out, minus2A_out, plus4A_out, 
        minus4A_out );
  input [63:0] plusA;
  output [63:0] plus2A_out;
  output [63:0] minus2A_out;
  output [63:0] plus4A_out;
  output [63:0] minus4A_out;
  wire   n46, n47, n3, n48, n49, n4, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign plus2A_out[0] = 1'b0;
  assign plus2A_out[51] = n3;
  assign plus2A_out[39] = n4;
  assign plus4A_out[0] = 1'b0;

  shifter_N64_26 shifter_1 ( .\input (plusA), .shiftLeftOnePos({
        plus2A_out[63:59], n46, plus2A_out[57:54], n47, plus2A_out[52], n3, 
        plus2A_out[50:49], n48, plus2A_out[47:44], n49, plus2A_out[42:40], n4, 
        n50, n51, n52, plus2A_out[35:1], SYNOPSYS_UNCONNECTED__0}) );
  shifter_N64_25 shifter_2 ( .\input ({plus2A_out[63:52], n3, 
        plus2A_out[50:40], n4, plus2A_out[38:1], 1'b0}), .shiftLeftOnePos({
        plus4A_out[63:59], n53, plus4A_out[57:54], n54, plus4A_out[52:49], n55, 
        plus4A_out[47:44], n56, plus4A_out[42:37], n57, n58, n59, n60, n61, 
        n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, 
        n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, plus4A_out[6:1], 
        SYNOPSYS_UNCONNECTED__1}) );
  complementer_N64_26 complementer_1 ( .\input ({plus2A_out[63:52], n3, 
        plus2A_out[50:40], n4, plus2A_out[38:1], 1'b0}), .complement2(
        minus2A_out) );
  complementer_N64_25 complementer_2 ( .\input ({plus4A_out[63:1], 1'b0}), 
        .complement2(minus4A_out) );
  BUF_X1 U1 ( .A(n50), .Z(plus2A_out[38]) );
  BUF_X1 U2 ( .A(n49), .Z(plus2A_out[43]) );
  BUF_X1 U5 ( .A(n56), .Z(plus4A_out[43]) );
  BUF_X1 U6 ( .A(n48), .Z(plus2A_out[48]) );
  BUF_X1 U7 ( .A(n55), .Z(plus4A_out[48]) );
  BUF_X1 U8 ( .A(n47), .Z(plus2A_out[53]) );
  BUF_X1 U9 ( .A(n54), .Z(plus4A_out[53]) );
  BUF_X1 U10 ( .A(n46), .Z(plus2A_out[58]) );
  BUF_X1 U11 ( .A(n53), .Z(plus4A_out[58]) );
  BUF_X1 U12 ( .A(n78), .Z(plus4A_out[15]) );
  BUF_X1 U13 ( .A(n76), .Z(plus4A_out[17]) );
  BUF_X1 U14 ( .A(n80), .Z(plus4A_out[13]) );
  BUF_X1 U15 ( .A(n82), .Z(plus4A_out[11]) );
  BUF_X1 U16 ( .A(n84), .Z(plus4A_out[9]) );
  BUF_X1 U17 ( .A(n79), .Z(plus4A_out[14]) );
  BUF_X1 U18 ( .A(n77), .Z(plus4A_out[16]) );
  BUF_X1 U19 ( .A(n81), .Z(plus4A_out[12]) );
  BUF_X1 U20 ( .A(n83), .Z(plus4A_out[10]) );
  BUF_X1 U21 ( .A(n66), .Z(plus4A_out[27]) );
  BUF_X1 U22 ( .A(n70), .Z(plus4A_out[23]) );
  BUF_X1 U23 ( .A(n74), .Z(plus4A_out[19]) );
  BUF_X1 U24 ( .A(n68), .Z(plus4A_out[25]) );
  BUF_X1 U25 ( .A(n72), .Z(plus4A_out[21]) );
  BUF_X1 U26 ( .A(n67), .Z(plus4A_out[26]) );
  BUF_X1 U27 ( .A(n71), .Z(plus4A_out[22]) );
  BUF_X1 U28 ( .A(n75), .Z(plus4A_out[18]) );
  BUF_X1 U29 ( .A(n65), .Z(plus4A_out[28]) );
  BUF_X1 U30 ( .A(n69), .Z(plus4A_out[24]) );
  BUF_X1 U31 ( .A(n73), .Z(plus4A_out[20]) );
  BUF_X1 U32 ( .A(n58), .Z(plus4A_out[35]) );
  BUF_X1 U33 ( .A(n62), .Z(plus4A_out[31]) );
  BUF_X1 U34 ( .A(n60), .Z(plus4A_out[33]) );
  BUF_X1 U35 ( .A(n64), .Z(plus4A_out[29]) );
  BUF_X1 U36 ( .A(n59), .Z(plus4A_out[34]) );
  BUF_X1 U37 ( .A(n63), .Z(plus4A_out[30]) );
  BUF_X1 U38 ( .A(n52), .Z(plus2A_out[36]) );
  BUF_X1 U39 ( .A(n57), .Z(plus4A_out[36]) );
  BUF_X1 U40 ( .A(n61), .Z(plus4A_out[32]) );
  BUF_X1 U41 ( .A(n51), .Z(plus2A_out[37]) );
  BUF_X1 U42 ( .A(n86), .Z(plus4A_out[7]) );
  BUF_X1 U43 ( .A(n85), .Z(plus4A_out[8]) );
endmodule


module MUX_GENERIC_N64_RADIX3_13 ( plusA, minusA, plus2A, minus2A, SEL, Y );
  input [63:0] plusA;
  input [63:0] minusA;
  input [63:0] plus2A;
  input [63:0] minus2A;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502;
  tri   [63:0] Y;

  TBUF_X1 \Y_tri[60]  ( .A(n441), .EN(n301), .Z(Y[60]) );
  TBUF_X1 \Y_tri[61]  ( .A(n440), .EN(n301), .Z(Y[61]) );
  TBUF_X1 \Y_tri[63]  ( .A(n438), .EN(n301), .Z(Y[63]) );
  TBUF_X1 \Y_tri[55]  ( .A(n446), .EN(n301), .Z(Y[55]) );
  TBUF_X1 \Y_tri[56]  ( .A(n445), .EN(n301), .Z(Y[56]) );
  TBUF_X1 \Y_tri[57]  ( .A(n444), .EN(n301), .Z(Y[57]) );
  TBUF_X1 \Y_tri[58]  ( .A(n443), .EN(n301), .Z(Y[58]) );
  TBUF_X1 \Y_tri[59]  ( .A(n442), .EN(n301), .Z(Y[59]) );
  TBUF_X1 \Y_tri[35]  ( .A(n466), .EN(n299), .Z(Y[35]) );
  TBUF_X1 \Y_tri[36]  ( .A(n465), .EN(n299), .Z(Y[36]) );
  TBUF_X1 \Y_tri[37]  ( .A(n464), .EN(n299), .Z(Y[37]) );
  TBUF_X1 \Y_tri[38]  ( .A(n463), .EN(n299), .Z(Y[38]) );
  TBUF_X1 \Y_tri[39]  ( .A(n462), .EN(n299), .Z(Y[39]) );
  TBUF_X1 \Y_tri[40]  ( .A(n461), .EN(n299), .Z(Y[40]) );
  TBUF_X1 \Y_tri[41]  ( .A(n460), .EN(n299), .Z(Y[41]) );
  TBUF_X1 \Y_tri[42]  ( .A(n459), .EN(n299), .Z(Y[42]) );
  TBUF_X1 \Y_tri[43]  ( .A(n458), .EN(n299), .Z(Y[43]) );
  TBUF_X1 \Y_tri[44]  ( .A(n457), .EN(n300), .Z(Y[44]) );
  TBUF_X1 \Y_tri[45]  ( .A(n456), .EN(n300), .Z(Y[45]) );
  TBUF_X1 \Y_tri[46]  ( .A(n455), .EN(n300), .Z(Y[46]) );
  TBUF_X1 \Y_tri[47]  ( .A(n454), .EN(n300), .Z(Y[47]) );
  TBUF_X1 \Y_tri[48]  ( .A(n453), .EN(n300), .Z(Y[48]) );
  TBUF_X1 \Y_tri[49]  ( .A(n452), .EN(n300), .Z(Y[49]) );
  TBUF_X1 \Y_tri[50]  ( .A(n451), .EN(n300), .Z(Y[50]) );
  TBUF_X1 \Y_tri[51]  ( .A(n450), .EN(n300), .Z(Y[51]) );
  TBUF_X1 \Y_tri[52]  ( .A(n449), .EN(n300), .Z(Y[52]) );
  TBUF_X1 \Y_tri[53]  ( .A(n448), .EN(n300), .Z(Y[53]) );
  TBUF_X1 \Y_tri[54]  ( .A(n447), .EN(n300), .Z(Y[54]) );
  TBUF_X1 \Y_tri[10]  ( .A(n491), .EN(n296), .Z(Y[10]) );
  TBUF_X1 \Y_tri[11]  ( .A(n490), .EN(n297), .Z(Y[11]) );
  TBUF_X1 \Y_tri[13]  ( .A(n488), .EN(n297), .Z(Y[13]) );
  TBUF_X1 \Y_tri[14]  ( .A(n487), .EN(n297), .Z(Y[14]) );
  TBUF_X1 \Y_tri[15]  ( .A(n486), .EN(n297), .Z(Y[15]) );
  TBUF_X1 \Y_tri[16]  ( .A(n485), .EN(n297), .Z(Y[16]) );
  TBUF_X1 \Y_tri[17]  ( .A(n484), .EN(n297), .Z(Y[17]) );
  TBUF_X1 \Y_tri[18]  ( .A(n483), .EN(n297), .Z(Y[18]) );
  TBUF_X1 \Y_tri[19]  ( .A(n482), .EN(n297), .Z(Y[19]) );
  TBUF_X1 \Y_tri[20]  ( .A(n481), .EN(n297), .Z(Y[20]) );
  TBUF_X1 \Y_tri[21]  ( .A(n480), .EN(n297), .Z(Y[21]) );
  TBUF_X1 \Y_tri[22]  ( .A(n479), .EN(n298), .Z(Y[22]) );
  TBUF_X1 \Y_tri[25]  ( .A(n476), .EN(n298), .Z(Y[25]) );
  TBUF_X1 \Y_tri[26]  ( .A(n475), .EN(n298), .Z(Y[26]) );
  TBUF_X1 \Y_tri[27]  ( .A(n474), .EN(n298), .Z(Y[27]) );
  TBUF_X1 \Y_tri[29]  ( .A(n472), .EN(n298), .Z(Y[29]) );
  TBUF_X1 \Y_tri[30]  ( .A(n471), .EN(n298), .Z(Y[30]) );
  TBUF_X1 \Y_tri[0]  ( .A(n502), .EN(n296), .Z(Y[0]) );
  TBUF_X1 \Y_tri[1]  ( .A(n501), .EN(n296), .Z(Y[1]) );
  TBUF_X1 \Y_tri[2]  ( .A(n500), .EN(n296), .Z(Y[2]) );
  TBUF_X1 \Y_tri[3]  ( .A(n499), .EN(n296), .Z(Y[3]) );
  TBUF_X1 \Y_tri[4]  ( .A(n498), .EN(n296), .Z(Y[4]) );
  TBUF_X1 \Y_tri[6]  ( .A(n496), .EN(n296), .Z(Y[6]) );
  TBUF_X1 \Y_tri[8]  ( .A(n494), .EN(n296), .Z(Y[8]) );
  TBUF_X1 \Y_tri[9]  ( .A(n492), .EN(n296), .Z(Y[9]) );
  TBUF_X1 \Y_tri[5]  ( .A(n497), .EN(n296), .Z(Y[5]) );
  TBUF_X1 \Y_tri[7]  ( .A(n495), .EN(n296), .Z(Y[7]) );
  TBUF_X1 \Y_tri[12]  ( .A(n489), .EN(n297), .Z(Y[12]) );
  TBUF_X1 \Y_tri[23]  ( .A(n478), .EN(n298), .Z(Y[23]) );
  TBUF_X1 \Y_tri[24]  ( .A(n477), .EN(n298), .Z(Y[24]) );
  TBUF_X1 \Y_tri[28]  ( .A(n473), .EN(n298), .Z(Y[28]) );
  TBUF_X1 \Y_tri[31]  ( .A(n470), .EN(n298), .Z(Y[31]) );
  TBUF_X1 \Y_tri[32]  ( .A(n469), .EN(n298), .Z(Y[32]) );
  TBUF_X1 \Y_tri[33]  ( .A(n468), .EN(n299), .Z(Y[33]) );
  TBUF_X1 \Y_tri[34]  ( .A(n467), .EN(n299), .Z(Y[34]) );
  TBUF_X1 \Y_tri[62]  ( .A(n439), .EN(n301), .Z(Y[62]) );
  NAND2_X1 U2 ( .A1(n399), .A2(n398), .ZN(n455) );
  AOI22_X1 U3 ( .A1(plusA[46]), .A2(n281), .B1(plus2A[46]), .B2(n275), .ZN(
        n399) );
  AOI22_X1 U4 ( .A1(minus2A[46]), .A2(n293), .B1(minusA[46]), .B2(n287), .ZN(
        n398) );
  NAND2_X1 U5 ( .A1(n401), .A2(n400), .ZN(n454) );
  AOI22_X1 U6 ( .A1(plusA[47]), .A2(n281), .B1(plus2A[47]), .B2(n275), .ZN(
        n401) );
  AOI22_X1 U7 ( .A1(minus2A[47]), .A2(n293), .B1(minusA[47]), .B2(n287), .ZN(
        n400) );
  NAND2_X1 U8 ( .A1(n395), .A2(n394), .ZN(n457) );
  AOI22_X1 U9 ( .A1(plusA[44]), .A2(n281), .B1(plus2A[44]), .B2(n275), .ZN(
        n395) );
  AOI22_X1 U10 ( .A1(minus2A[44]), .A2(n293), .B1(minusA[44]), .B2(n287), .ZN(
        n394) );
  NAND2_X1 U11 ( .A1(n397), .A2(n396), .ZN(n456) );
  AOI22_X1 U12 ( .A1(plusA[45]), .A2(n281), .B1(plus2A[45]), .B2(n275), .ZN(
        n397) );
  AOI22_X1 U13 ( .A1(minus2A[45]), .A2(n293), .B1(minusA[45]), .B2(n287), .ZN(
        n396) );
  NAND2_X1 U14 ( .A1(n393), .A2(n392), .ZN(n458) );
  AOI22_X1 U15 ( .A1(plusA[43]), .A2(n281), .B1(plus2A[43]), .B2(n275), .ZN(
        n393) );
  AOI22_X1 U16 ( .A1(minus2A[43]), .A2(n293), .B1(minusA[43]), .B2(n287), .ZN(
        n392) );
  NAND2_X1 U17 ( .A1(n419), .A2(n418), .ZN(n445) );
  AOI22_X1 U18 ( .A1(plusA[56]), .A2(n282), .B1(plus2A[56]), .B2(n276), .ZN(
        n419) );
  AOI22_X1 U19 ( .A1(minus2A[56]), .A2(n294), .B1(minusA[56]), .B2(n288), .ZN(
        n418) );
  NAND2_X1 U20 ( .A1(n421), .A2(n420), .ZN(n444) );
  AOI22_X1 U21 ( .A1(plusA[57]), .A2(n282), .B1(plus2A[57]), .B2(n276), .ZN(
        n421) );
  AOI22_X1 U22 ( .A1(minus2A[57]), .A2(n294), .B1(minusA[57]), .B2(n288), .ZN(
        n420) );
  NAND2_X1 U23 ( .A1(n415), .A2(n414), .ZN(n447) );
  AOI22_X1 U24 ( .A1(plusA[54]), .A2(n282), .B1(plus2A[54]), .B2(n276), .ZN(
        n415) );
  AOI22_X1 U25 ( .A1(minus2A[54]), .A2(n294), .B1(minusA[54]), .B2(n288), .ZN(
        n414) );
  NAND2_X1 U26 ( .A1(n383), .A2(n382), .ZN(n463) );
  AOI22_X1 U27 ( .A1(plusA[38]), .A2(n281), .B1(plus2A[38]), .B2(n275), .ZN(
        n383) );
  AOI22_X1 U28 ( .A1(minus2A[38]), .A2(n293), .B1(minusA[38]), .B2(n287), .ZN(
        n382) );
  NAND2_X1 U29 ( .A1(n417), .A2(n416), .ZN(n446) );
  AOI22_X1 U30 ( .A1(plusA[55]), .A2(n282), .B1(plus2A[55]), .B2(n276), .ZN(
        n417) );
  AOI22_X1 U31 ( .A1(minus2A[55]), .A2(n294), .B1(minusA[55]), .B2(n288), .ZN(
        n416) );
  NAND2_X1 U32 ( .A1(n413), .A2(n412), .ZN(n448) );
  AOI22_X1 U33 ( .A1(plusA[53]), .A2(n282), .B1(plus2A[53]), .B2(n276), .ZN(
        n413) );
  AOI22_X1 U34 ( .A1(minus2A[53]), .A2(n294), .B1(minusA[53]), .B2(n288), .ZN(
        n412) );
  NAND2_X1 U35 ( .A1(n409), .A2(n408), .ZN(n450) );
  AOI22_X1 U36 ( .A1(plusA[51]), .A2(n282), .B1(plus2A[51]), .B2(n276), .ZN(
        n409) );
  AOI22_X1 U37 ( .A1(minus2A[51]), .A2(n294), .B1(minusA[51]), .B2(n288), .ZN(
        n408) );
  NAND2_X1 U38 ( .A1(n411), .A2(n410), .ZN(n449) );
  AOI22_X1 U39 ( .A1(plusA[52]), .A2(n282), .B1(plus2A[52]), .B2(n276), .ZN(
        n411) );
  AOI22_X1 U40 ( .A1(minus2A[52]), .A2(n294), .B1(minusA[52]), .B2(n288), .ZN(
        n410) );
  NAND2_X1 U41 ( .A1(n405), .A2(n404), .ZN(n452) );
  AOI22_X1 U42 ( .A1(plusA[49]), .A2(n282), .B1(plus2A[49]), .B2(n276), .ZN(
        n405) );
  AOI22_X1 U43 ( .A1(minus2A[49]), .A2(n294), .B1(minusA[49]), .B2(n288), .ZN(
        n404) );
  NAND2_X1 U44 ( .A1(n407), .A2(n406), .ZN(n451) );
  AOI22_X1 U45 ( .A1(plusA[50]), .A2(n282), .B1(plus2A[50]), .B2(n276), .ZN(
        n407) );
  AOI22_X1 U46 ( .A1(minus2A[50]), .A2(n294), .B1(minusA[50]), .B2(n288), .ZN(
        n406) );
  NAND2_X1 U47 ( .A1(n403), .A2(n402), .ZN(n453) );
  AOI22_X1 U48 ( .A1(plusA[48]), .A2(n282), .B1(plus2A[48]), .B2(n276), .ZN(
        n403) );
  AOI22_X1 U49 ( .A1(minus2A[48]), .A2(n294), .B1(minusA[48]), .B2(n288), .ZN(
        n402) );
  NAND2_X1 U50 ( .A1(n389), .A2(n388), .ZN(n460) );
  AOI22_X1 U51 ( .A1(plusA[41]), .A2(n281), .B1(plus2A[41]), .B2(n275), .ZN(
        n389) );
  AOI22_X1 U52 ( .A1(minus2A[41]), .A2(n293), .B1(minusA[41]), .B2(n287), .ZN(
        n388) );
  NAND2_X1 U53 ( .A1(n391), .A2(n390), .ZN(n459) );
  AOI22_X1 U54 ( .A1(plusA[42]), .A2(n281), .B1(plus2A[42]), .B2(n275), .ZN(
        n391) );
  AOI22_X1 U55 ( .A1(minus2A[42]), .A2(n293), .B1(minusA[42]), .B2(n287), .ZN(
        n390) );
  NAND2_X1 U56 ( .A1(n385), .A2(n384), .ZN(n462) );
  AOI22_X1 U57 ( .A1(plusA[39]), .A2(n281), .B1(plus2A[39]), .B2(n275), .ZN(
        n385) );
  AOI22_X1 U58 ( .A1(minus2A[39]), .A2(n293), .B1(minusA[39]), .B2(n287), .ZN(
        n384) );
  NAND2_X1 U59 ( .A1(n387), .A2(n386), .ZN(n461) );
  AOI22_X1 U60 ( .A1(plusA[40]), .A2(n281), .B1(plus2A[40]), .B2(n275), .ZN(
        n387) );
  AOI22_X1 U61 ( .A1(minus2A[40]), .A2(n293), .B1(minusA[40]), .B2(n287), .ZN(
        n386) );
  NAND2_X1 U62 ( .A1(n431), .A2(n430), .ZN(n439) );
  AOI22_X1 U63 ( .A1(plusA[62]), .A2(n283), .B1(plus2A[62]), .B2(n277), .ZN(
        n431) );
  AOI22_X1 U64 ( .A1(minus2A[62]), .A2(n295), .B1(minusA[62]), .B2(n289), .ZN(
        n430) );
  NAND2_X1 U65 ( .A1(n423), .A2(n422), .ZN(n443) );
  AOI22_X1 U66 ( .A1(plusA[58]), .A2(n282), .B1(plus2A[58]), .B2(n276), .ZN(
        n423) );
  AOI22_X1 U67 ( .A1(minus2A[58]), .A2(n294), .B1(minusA[58]), .B2(n288), .ZN(
        n422) );
  NAND2_X1 U68 ( .A1(n425), .A2(n424), .ZN(n442) );
  AOI22_X1 U69 ( .A1(plusA[59]), .A2(n282), .B1(plus2A[59]), .B2(n276), .ZN(
        n425) );
  AOI22_X1 U70 ( .A1(minus2A[59]), .A2(n294), .B1(minusA[59]), .B2(n288), .ZN(
        n424) );
  NAND2_X1 U71 ( .A1(n437), .A2(n436), .ZN(n438) );
  AOI22_X1 U72 ( .A1(plusA[63]), .A2(n283), .B1(plus2A[63]), .B2(n277), .ZN(
        n437) );
  AOI22_X1 U73 ( .A1(minus2A[63]), .A2(n295), .B1(minusA[63]), .B2(n289), .ZN(
        n436) );
  NAND2_X1 U74 ( .A1(n429), .A2(n428), .ZN(n440) );
  AOI22_X1 U75 ( .A1(plusA[61]), .A2(n283), .B1(plus2A[61]), .B2(n277), .ZN(
        n429) );
  AOI22_X1 U76 ( .A1(minus2A[61]), .A2(n295), .B1(minusA[61]), .B2(n289), .ZN(
        n428) );
  NAND2_X1 U77 ( .A1(n427), .A2(n426), .ZN(n441) );
  AOI22_X1 U78 ( .A1(plusA[60]), .A2(n283), .B1(plus2A[60]), .B2(n277), .ZN(
        n427) );
  AOI22_X1 U79 ( .A1(minus2A[60]), .A2(n295), .B1(minusA[60]), .B2(n289), .ZN(
        n426) );
  BUF_X1 U80 ( .A(n433), .Z(n279) );
  BUF_X1 U81 ( .A(n433), .Z(n278) );
  BUF_X1 U82 ( .A(n435), .Z(n291) );
  BUF_X1 U83 ( .A(n435), .Z(n290) );
  BUF_X1 U84 ( .A(n434), .Z(n285) );
  BUF_X1 U85 ( .A(n432), .Z(n273) );
  BUF_X1 U86 ( .A(n434), .Z(n284) );
  BUF_X1 U87 ( .A(n432), .Z(n272) );
  BUF_X1 U88 ( .A(n493), .Z(n297) );
  BUF_X1 U89 ( .A(n493), .Z(n296) );
  BUF_X1 U90 ( .A(n433), .Z(n280) );
  BUF_X1 U91 ( .A(n434), .Z(n286) );
  BUF_X1 U92 ( .A(n432), .Z(n274) );
  BUF_X1 U93 ( .A(n493), .Z(n298) );
  BUF_X1 U94 ( .A(n435), .Z(n292) );
  BUF_X1 U95 ( .A(n493), .Z(n299) );
  NAND2_X1 U96 ( .A1(n381), .A2(n380), .ZN(n464) );
  AOI22_X1 U97 ( .A1(plusA[37]), .A2(n281), .B1(plus2A[37]), .B2(n275), .ZN(
        n381) );
  AOI22_X1 U98 ( .A1(minus2A[37]), .A2(n293), .B1(minusA[37]), .B2(n287), .ZN(
        n380) );
  NAND2_X1 U99 ( .A1(n379), .A2(n378), .ZN(n465) );
  AOI22_X1 U100 ( .A1(plusA[36]), .A2(n281), .B1(plus2A[36]), .B2(n275), .ZN(
        n379) );
  AOI22_X1 U101 ( .A1(minus2A[36]), .A2(n293), .B1(minusA[36]), .B2(n287), 
        .ZN(n378) );
  BUF_X1 U102 ( .A(n433), .Z(n281) );
  BUF_X1 U103 ( .A(n435), .Z(n293) );
  BUF_X1 U104 ( .A(n434), .Z(n287) );
  BUF_X1 U105 ( .A(n432), .Z(n275) );
  BUF_X1 U106 ( .A(n433), .Z(n282) );
  BUF_X1 U107 ( .A(n435), .Z(n294) );
  BUF_X1 U108 ( .A(n434), .Z(n288) );
  BUF_X1 U109 ( .A(n432), .Z(n276) );
  BUF_X1 U110 ( .A(n493), .Z(n300) );
  BUF_X1 U111 ( .A(n493), .Z(n301) );
  NOR3_X1 U112 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n302), .ZN(n434) );
  NOR3_X1 U113 ( .A1(n302), .A2(SEL[2]), .A3(n303), .ZN(n432) );
  NOR3_X1 U114 ( .A1(SEL[1]), .A2(SEL[2]), .A3(n303), .ZN(n433) );
  NOR2_X1 U115 ( .A1(n323), .A2(n304), .ZN(n493) );
  INV_X1 U116 ( .A(SEL[2]), .ZN(n304) );
  NOR2_X1 U117 ( .A1(SEL[1]), .A2(SEL[0]), .ZN(n323) );
  AND2_X1 U118 ( .A1(SEL[2]), .A2(n323), .ZN(n435) );
  INV_X1 U119 ( .A(SEL[1]), .ZN(n302) );
  INV_X1 U120 ( .A(SEL[0]), .ZN(n303) );
  NAND2_X1 U121 ( .A1(n320), .A2(n319), .ZN(n495) );
  AOI22_X1 U122 ( .A1(plusA[7]), .A2(n278), .B1(plus2A[7]), .B2(n272), .ZN(
        n320) );
  AOI22_X1 U123 ( .A1(minus2A[7]), .A2(n290), .B1(minusA[7]), .B2(n284), .ZN(
        n319) );
  NAND2_X1 U124 ( .A1(n325), .A2(n324), .ZN(n492) );
  AOI22_X1 U125 ( .A1(plusA[9]), .A2(n278), .B1(plus2A[9]), .B2(n272), .ZN(
        n325) );
  AOI22_X1 U126 ( .A1(minus2A[9]), .A2(n290), .B1(minusA[9]), .B2(n284), .ZN(
        n324) );
  NAND2_X1 U127 ( .A1(n331), .A2(n330), .ZN(n489) );
  AOI22_X1 U128 ( .A1(plusA[12]), .A2(n279), .B1(plus2A[12]), .B2(n273), .ZN(
        n331) );
  AOI22_X1 U129 ( .A1(minus2A[12]), .A2(n291), .B1(minusA[12]), .B2(n285), 
        .ZN(n330) );
  NAND2_X1 U130 ( .A1(n322), .A2(n321), .ZN(n494) );
  AOI22_X1 U131 ( .A1(plusA[8]), .A2(n278), .B1(plus2A[8]), .B2(n272), .ZN(
        n322) );
  AOI22_X1 U132 ( .A1(minus2A[8]), .A2(n290), .B1(minusA[8]), .B2(n284), .ZN(
        n321) );
  NAND2_X1 U133 ( .A1(n369), .A2(n368), .ZN(n470) );
  AOI22_X1 U134 ( .A1(plusA[31]), .A2(n280), .B1(plus2A[31]), .B2(n274), .ZN(
        n369) );
  AOI22_X1 U135 ( .A1(minus2A[31]), .A2(n292), .B1(minusA[31]), .B2(n286), 
        .ZN(n368) );
  NAND2_X1 U136 ( .A1(n367), .A2(n366), .ZN(n471) );
  AOI22_X1 U137 ( .A1(plusA[30]), .A2(n280), .B1(plus2A[30]), .B2(n274), .ZN(
        n367) );
  AOI22_X1 U138 ( .A1(minus2A[30]), .A2(n292), .B1(minusA[30]), .B2(n286), 
        .ZN(n366) );
  NAND2_X1 U139 ( .A1(n365), .A2(n364), .ZN(n472) );
  AOI22_X1 U140 ( .A1(plusA[29]), .A2(n280), .B1(plus2A[29]), .B2(n274), .ZN(
        n365) );
  AOI22_X1 U141 ( .A1(minus2A[29]), .A2(n292), .B1(minusA[29]), .B2(n286), 
        .ZN(n364) );
  NAND2_X1 U142 ( .A1(n361), .A2(n360), .ZN(n474) );
  AOI22_X1 U143 ( .A1(plusA[27]), .A2(n280), .B1(plus2A[27]), .B2(n274), .ZN(
        n361) );
  AOI22_X1 U144 ( .A1(minus2A[27]), .A2(n292), .B1(minusA[27]), .B2(n286), 
        .ZN(n360) );
  NAND2_X1 U145 ( .A1(n359), .A2(n358), .ZN(n475) );
  AOI22_X1 U146 ( .A1(plusA[26]), .A2(n280), .B1(plus2A[26]), .B2(n274), .ZN(
        n359) );
  AOI22_X1 U147 ( .A1(minus2A[26]), .A2(n292), .B1(minusA[26]), .B2(n286), 
        .ZN(n358) );
  NAND2_X1 U148 ( .A1(n357), .A2(n356), .ZN(n476) );
  AOI22_X1 U149 ( .A1(plusA[25]), .A2(n280), .B1(plus2A[25]), .B2(n274), .ZN(
        n357) );
  AOI22_X1 U150 ( .A1(minus2A[25]), .A2(n292), .B1(minusA[25]), .B2(n286), 
        .ZN(n356) );
  NAND2_X1 U151 ( .A1(n353), .A2(n352), .ZN(n478) );
  AOI22_X1 U152 ( .A1(plusA[23]), .A2(n279), .B1(plus2A[23]), .B2(n273), .ZN(
        n353) );
  AOI22_X1 U153 ( .A1(minus2A[23]), .A2(n291), .B1(minusA[23]), .B2(n285), 
        .ZN(n352) );
  NAND2_X1 U154 ( .A1(n351), .A2(n350), .ZN(n479) );
  AOI22_X1 U155 ( .A1(plusA[22]), .A2(n279), .B1(plus2A[22]), .B2(n273), .ZN(
        n351) );
  AOI22_X1 U156 ( .A1(minus2A[22]), .A2(n291), .B1(minusA[22]), .B2(n285), 
        .ZN(n350) );
  NAND2_X1 U157 ( .A1(n349), .A2(n348), .ZN(n480) );
  AOI22_X1 U158 ( .A1(plusA[21]), .A2(n279), .B1(plus2A[21]), .B2(n273), .ZN(
        n349) );
  AOI22_X1 U159 ( .A1(minus2A[21]), .A2(n291), .B1(minusA[21]), .B2(n285), 
        .ZN(n348) );
  NAND2_X1 U160 ( .A1(n345), .A2(n344), .ZN(n482) );
  AOI22_X1 U161 ( .A1(plusA[19]), .A2(n279), .B1(plus2A[19]), .B2(n273), .ZN(
        n345) );
  AOI22_X1 U162 ( .A1(minus2A[19]), .A2(n291), .B1(minusA[19]), .B2(n285), 
        .ZN(n344) );
  NAND2_X1 U163 ( .A1(n343), .A2(n342), .ZN(n483) );
  AOI22_X1 U164 ( .A1(plusA[18]), .A2(n279), .B1(plus2A[18]), .B2(n273), .ZN(
        n343) );
  AOI22_X1 U165 ( .A1(minus2A[18]), .A2(n291), .B1(minusA[18]), .B2(n285), 
        .ZN(n342) );
  NAND2_X1 U166 ( .A1(n341), .A2(n340), .ZN(n484) );
  AOI22_X1 U167 ( .A1(plusA[17]), .A2(n279), .B1(plus2A[17]), .B2(n273), .ZN(
        n341) );
  AOI22_X1 U168 ( .A1(minus2A[17]), .A2(n291), .B1(minusA[17]), .B2(n285), 
        .ZN(n340) );
  NAND2_X1 U169 ( .A1(n337), .A2(n336), .ZN(n486) );
  AOI22_X1 U170 ( .A1(plusA[15]), .A2(n279), .B1(plus2A[15]), .B2(n273), .ZN(
        n337) );
  AOI22_X1 U171 ( .A1(minus2A[15]), .A2(n291), .B1(minusA[15]), .B2(n285), 
        .ZN(n336) );
  NAND2_X1 U172 ( .A1(n335), .A2(n334), .ZN(n487) );
  AOI22_X1 U173 ( .A1(plusA[14]), .A2(n279), .B1(plus2A[14]), .B2(n273), .ZN(
        n335) );
  AOI22_X1 U174 ( .A1(minus2A[14]), .A2(n291), .B1(minusA[14]), .B2(n285), 
        .ZN(n334) );
  NAND2_X1 U175 ( .A1(n333), .A2(n332), .ZN(n488) );
  AOI22_X1 U176 ( .A1(plusA[13]), .A2(n279), .B1(plus2A[13]), .B2(n273), .ZN(
        n333) );
  AOI22_X1 U177 ( .A1(minus2A[13]), .A2(n291), .B1(minusA[13]), .B2(n285), 
        .ZN(n332) );
  NAND2_X1 U178 ( .A1(n329), .A2(n328), .ZN(n490) );
  AOI22_X1 U179 ( .A1(plusA[11]), .A2(n278), .B1(plus2A[11]), .B2(n272), .ZN(
        n329) );
  AOI22_X1 U180 ( .A1(minus2A[11]), .A2(n290), .B1(minusA[11]), .B2(n284), 
        .ZN(n328) );
  NAND2_X1 U181 ( .A1(n373), .A2(n372), .ZN(n468) );
  AOI22_X1 U182 ( .A1(plusA[33]), .A2(n280), .B1(plus2A[33]), .B2(n274), .ZN(
        n373) );
  AOI22_X1 U183 ( .A1(minus2A[33]), .A2(n292), .B1(minusA[33]), .B2(n286), 
        .ZN(n372) );
  NAND2_X1 U184 ( .A1(n371), .A2(n370), .ZN(n469) );
  AOI22_X1 U185 ( .A1(plusA[32]), .A2(n280), .B1(plus2A[32]), .B2(n274), .ZN(
        n371) );
  AOI22_X1 U186 ( .A1(minus2A[32]), .A2(n292), .B1(minusA[32]), .B2(n286), 
        .ZN(n370) );
  NAND2_X1 U187 ( .A1(n363), .A2(n362), .ZN(n473) );
  AOI22_X1 U188 ( .A1(plusA[28]), .A2(n280), .B1(plus2A[28]), .B2(n274), .ZN(
        n363) );
  AOI22_X1 U189 ( .A1(minus2A[28]), .A2(n292), .B1(minusA[28]), .B2(n286), 
        .ZN(n362) );
  NAND2_X1 U190 ( .A1(n355), .A2(n354), .ZN(n477) );
  AOI22_X1 U191 ( .A1(plusA[24]), .A2(n280), .B1(plus2A[24]), .B2(n274), .ZN(
        n355) );
  AOI22_X1 U192 ( .A1(minus2A[24]), .A2(n292), .B1(minusA[24]), .B2(n286), 
        .ZN(n354) );
  NAND2_X1 U193 ( .A1(n347), .A2(n346), .ZN(n481) );
  AOI22_X1 U194 ( .A1(plusA[20]), .A2(n279), .B1(plus2A[20]), .B2(n273), .ZN(
        n347) );
  AOI22_X1 U195 ( .A1(minus2A[20]), .A2(n291), .B1(minusA[20]), .B2(n285), 
        .ZN(n346) );
  NAND2_X1 U196 ( .A1(n339), .A2(n338), .ZN(n485) );
  AOI22_X1 U197 ( .A1(plusA[16]), .A2(n279), .B1(plus2A[16]), .B2(n273), .ZN(
        n339) );
  AOI22_X1 U198 ( .A1(minus2A[16]), .A2(n291), .B1(minusA[16]), .B2(n285), 
        .ZN(n338) );
  NAND2_X1 U199 ( .A1(n375), .A2(n374), .ZN(n467) );
  AOI22_X1 U200 ( .A1(plusA[34]), .A2(n280), .B1(plus2A[34]), .B2(n274), .ZN(
        n375) );
  AOI22_X1 U201 ( .A1(minus2A[34]), .A2(n292), .B1(minusA[34]), .B2(n286), 
        .ZN(n374) );
  NAND2_X1 U202 ( .A1(n327), .A2(n326), .ZN(n491) );
  AOI22_X1 U203 ( .A1(plusA[10]), .A2(n278), .B1(plus2A[10]), .B2(n272), .ZN(
        n327) );
  AOI22_X1 U204 ( .A1(minus2A[10]), .A2(n290), .B1(minusA[10]), .B2(n284), 
        .ZN(n326) );
  NAND2_X1 U205 ( .A1(n377), .A2(n376), .ZN(n466) );
  AOI22_X1 U206 ( .A1(plusA[35]), .A2(n280), .B1(plus2A[35]), .B2(n274), .ZN(
        n377) );
  AOI22_X1 U207 ( .A1(minus2A[35]), .A2(n292), .B1(minusA[35]), .B2(n286), 
        .ZN(n376) );
  NAND2_X1 U208 ( .A1(n318), .A2(n317), .ZN(n496) );
  AOI22_X1 U209 ( .A1(plusA[6]), .A2(n278), .B1(plus2A[6]), .B2(n272), .ZN(
        n318) );
  AOI22_X1 U210 ( .A1(minus2A[6]), .A2(n290), .B1(minusA[6]), .B2(n284), .ZN(
        n317) );
  NAND2_X1 U211 ( .A1(n316), .A2(n315), .ZN(n497) );
  AOI22_X1 U212 ( .A1(plusA[5]), .A2(n278), .B1(plus2A[5]), .B2(n272), .ZN(
        n316) );
  AOI22_X1 U213 ( .A1(minus2A[5]), .A2(n290), .B1(minusA[5]), .B2(n284), .ZN(
        n315) );
  NAND2_X1 U214 ( .A1(n312), .A2(n311), .ZN(n499) );
  AOI22_X1 U215 ( .A1(plusA[3]), .A2(n278), .B1(plus2A[3]), .B2(n272), .ZN(
        n312) );
  AOI22_X1 U216 ( .A1(minus2A[3]), .A2(n290), .B1(minusA[3]), .B2(n284), .ZN(
        n311) );
  NAND2_X1 U217 ( .A1(n314), .A2(n313), .ZN(n498) );
  AOI22_X1 U218 ( .A1(plusA[4]), .A2(n278), .B1(plus2A[4]), .B2(n272), .ZN(
        n314) );
  AOI22_X1 U219 ( .A1(minus2A[4]), .A2(n290), .B1(minusA[4]), .B2(n284), .ZN(
        n313) );
  NAND2_X1 U220 ( .A1(n310), .A2(n309), .ZN(n500) );
  AOI22_X1 U221 ( .A1(plusA[2]), .A2(n278), .B1(plus2A[2]), .B2(n272), .ZN(
        n310) );
  AOI22_X1 U222 ( .A1(minus2A[2]), .A2(n290), .B1(minusA[2]), .B2(n284), .ZN(
        n309) );
  NAND2_X1 U223 ( .A1(n308), .A2(n307), .ZN(n501) );
  AOI22_X1 U224 ( .A1(plusA[1]), .A2(n278), .B1(plus2A[1]), .B2(n272), .ZN(
        n308) );
  AOI22_X1 U225 ( .A1(minus2A[1]), .A2(n290), .B1(minusA[1]), .B2(n284), .ZN(
        n307) );
  NAND2_X1 U226 ( .A1(n306), .A2(n305), .ZN(n502) );
  AOI22_X1 U227 ( .A1(plusA[0]), .A2(n278), .B1(plus2A[0]), .B2(n272), .ZN(
        n306) );
  AOI22_X1 U228 ( .A1(minus2A[0]), .A2(n290), .B1(minusA[0]), .B2(n284), .ZN(
        n305) );
  CLKBUF_X1 U229 ( .A(n432), .Z(n277) );
  CLKBUF_X1 U230 ( .A(n433), .Z(n283) );
  CLKBUF_X1 U231 ( .A(n434), .Z(n289) );
  CLKBUF_X1 U232 ( .A(n435), .Z(n295) );
endmodule


module FA_832 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_831 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_830 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_829 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_828 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_827 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  AOI22_X1 U4 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
  INV_X1 U5 ( .A(n7), .ZN(Co) );
endmodule


module FA_826 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_825 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  AOI22_X1 U4 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
  INV_X1 U5 ( .A(n7), .ZN(Co) );
endmodule


module FA_824 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_823 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_822 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_821 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_820 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  AOI22_X1 U4 ( .A1(B), .A2(A), .B1(Ci), .B2(n6), .ZN(n7) );
  INV_X1 U5 ( .A(n7), .ZN(Co) );
endmodule


module FA_819 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_818 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_817 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_816 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_815 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_814 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_813 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_812 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_811 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_810 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_809 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  AOI22_X1 U4 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
  INV_X1 U5 ( .A(n7), .ZN(Co) );
endmodule


module FA_808 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_807 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_806 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_805 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_804 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  AOI22_X1 U4 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
  INV_X1 U5 ( .A(n7), .ZN(Co) );
endmodule


module FA_803 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_802 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_801 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  AOI22_X1 U4 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
  INV_X1 U5 ( .A(n7), .ZN(Co) );
endmodule


module FA_800 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_799 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  AOI22_X1 U4 ( .A1(B), .A2(A), .B1(Ci), .B2(n6), .ZN(n7) );
  INV_X1 U5 ( .A(n7), .ZN(Co) );
endmodule


module FA_798 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  AOI22_X1 U4 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
  INV_X1 U5 ( .A(n7), .ZN(Co) );
endmodule


module FA_797 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_796 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_795 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_794 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_793 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_792 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_791 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_790 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_789 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_788 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_787 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_786 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_785 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_784 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_783 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_782 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_781 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_780 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_779 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_778 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_777 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_776 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_775 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_774 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_773 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_772 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_771 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_770 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_769 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N64_13 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Ci;
  output Co;

  wire   [63:1] CTMP;
  tri   [63:0] A;

  FA_832 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_831 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_830 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_829 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(CTMP[4]) );
  FA_828 FAI_5 ( .A(A[4]), .B(B[4]), .Ci(CTMP[4]), .S(S[4]), .Co(CTMP[5]) );
  FA_827 FAI_6 ( .A(A[5]), .B(B[5]), .Ci(CTMP[5]), .S(S[5]), .Co(CTMP[6]) );
  FA_826 FAI_7 ( .A(A[6]), .B(B[6]), .Ci(CTMP[6]), .S(S[6]), .Co(CTMP[7]) );
  FA_825 FAI_8 ( .A(A[7]), .B(B[7]), .Ci(CTMP[7]), .S(S[7]), .Co(CTMP[8]) );
  FA_824 FAI_9 ( .A(A[8]), .B(B[8]), .Ci(CTMP[8]), .S(S[8]), .Co(CTMP[9]) );
  FA_823 FAI_10 ( .A(A[9]), .B(B[9]), .Ci(CTMP[9]), .S(S[9]), .Co(CTMP[10]) );
  FA_822 FAI_11 ( .A(A[10]), .B(B[10]), .Ci(CTMP[10]), .S(S[10]), .Co(CTMP[11]) );
  FA_821 FAI_12 ( .A(A[11]), .B(B[11]), .Ci(CTMP[11]), .S(S[11]), .Co(CTMP[12]) );
  FA_820 FAI_13 ( .A(A[12]), .B(B[12]), .Ci(CTMP[12]), .S(S[12]), .Co(CTMP[13]) );
  FA_819 FAI_14 ( .A(A[13]), .B(B[13]), .Ci(CTMP[13]), .S(S[13]), .Co(CTMP[14]) );
  FA_818 FAI_15 ( .A(A[14]), .B(B[14]), .Ci(CTMP[14]), .S(S[14]), .Co(CTMP[15]) );
  FA_817 FAI_16 ( .A(A[15]), .B(B[15]), .Ci(CTMP[15]), .S(S[15]), .Co(CTMP[16]) );
  FA_816 FAI_17 ( .A(A[16]), .B(B[16]), .Ci(CTMP[16]), .S(S[16]), .Co(CTMP[17]) );
  FA_815 FAI_18 ( .A(A[17]), .B(B[17]), .Ci(CTMP[17]), .S(S[17]), .Co(CTMP[18]) );
  FA_814 FAI_19 ( .A(A[18]), .B(B[18]), .Ci(CTMP[18]), .S(S[18]), .Co(CTMP[19]) );
  FA_813 FAI_20 ( .A(A[19]), .B(B[19]), .Ci(CTMP[19]), .S(S[19]), .Co(CTMP[20]) );
  FA_812 FAI_21 ( .A(A[20]), .B(B[20]), .Ci(CTMP[20]), .S(S[20]), .Co(CTMP[21]) );
  FA_811 FAI_22 ( .A(A[21]), .B(B[21]), .Ci(CTMP[21]), .S(S[21]), .Co(CTMP[22]) );
  FA_810 FAI_23 ( .A(A[22]), .B(B[22]), .Ci(CTMP[22]), .S(S[22]), .Co(CTMP[23]) );
  FA_809 FAI_24 ( .A(A[23]), .B(B[23]), .Ci(CTMP[23]), .S(S[23]), .Co(CTMP[24]) );
  FA_808 FAI_25 ( .A(A[24]), .B(B[24]), .Ci(CTMP[24]), .S(S[24]), .Co(CTMP[25]) );
  FA_807 FAI_26 ( .A(A[25]), .B(B[25]), .Ci(CTMP[25]), .S(S[25]), .Co(CTMP[26]) );
  FA_806 FAI_27 ( .A(A[26]), .B(B[26]), .Ci(CTMP[26]), .S(S[26]), .Co(CTMP[27]) );
  FA_805 FAI_28 ( .A(A[27]), .B(B[27]), .Ci(CTMP[27]), .S(S[27]), .Co(CTMP[28]) );
  FA_804 FAI_29 ( .A(A[28]), .B(B[28]), .Ci(CTMP[28]), .S(S[28]), .Co(CTMP[29]) );
  FA_803 FAI_30 ( .A(A[29]), .B(B[29]), .Ci(CTMP[29]), .S(S[29]), .Co(CTMP[30]) );
  FA_802 FAI_31 ( .A(A[30]), .B(B[30]), .Ci(CTMP[30]), .S(S[30]), .Co(CTMP[31]) );
  FA_801 FAI_32 ( .A(A[31]), .B(B[31]), .Ci(CTMP[31]), .S(S[31]), .Co(CTMP[32]) );
  FA_800 FAI_33 ( .A(A[32]), .B(B[32]), .Ci(CTMP[32]), .S(S[32]), .Co(CTMP[33]) );
  FA_799 FAI_34 ( .A(A[33]), .B(B[33]), .Ci(CTMP[33]), .S(S[33]), .Co(CTMP[34]) );
  FA_798 FAI_35 ( .A(A[34]), .B(B[34]), .Ci(CTMP[34]), .S(S[34]), .Co(CTMP[35]) );
  FA_797 FAI_36 ( .A(A[35]), .B(B[35]), .Ci(CTMP[35]), .S(S[35]), .Co(CTMP[36]) );
  FA_796 FAI_37 ( .A(A[36]), .B(B[36]), .Ci(CTMP[36]), .S(S[36]), .Co(CTMP[37]) );
  FA_795 FAI_38 ( .A(A[37]), .B(B[37]), .Ci(CTMP[37]), .S(S[37]), .Co(CTMP[38]) );
  FA_794 FAI_39 ( .A(A[38]), .B(B[38]), .Ci(CTMP[38]), .S(S[38]), .Co(CTMP[39]) );
  FA_793 FAI_40 ( .A(A[39]), .B(B[39]), .Ci(CTMP[39]), .S(S[39]), .Co(CTMP[40]) );
  FA_792 FAI_41 ( .A(A[40]), .B(B[40]), .Ci(CTMP[40]), .S(S[40]), .Co(CTMP[41]) );
  FA_791 FAI_42 ( .A(A[41]), .B(B[41]), .Ci(CTMP[41]), .S(S[41]), .Co(CTMP[42]) );
  FA_790 FAI_43 ( .A(A[42]), .B(B[42]), .Ci(CTMP[42]), .S(S[42]), .Co(CTMP[43]) );
  FA_789 FAI_44 ( .A(A[43]), .B(B[43]), .Ci(CTMP[43]), .S(S[43]), .Co(CTMP[44]) );
  FA_788 FAI_45 ( .A(A[44]), .B(B[44]), .Ci(CTMP[44]), .S(S[44]), .Co(CTMP[45]) );
  FA_787 FAI_46 ( .A(A[45]), .B(B[45]), .Ci(CTMP[45]), .S(S[45]), .Co(CTMP[46]) );
  FA_786 FAI_47 ( .A(A[46]), .B(B[46]), .Ci(CTMP[46]), .S(S[46]), .Co(CTMP[47]) );
  FA_785 FAI_48 ( .A(A[47]), .B(B[47]), .Ci(CTMP[47]), .S(S[47]), .Co(CTMP[48]) );
  FA_784 FAI_49 ( .A(A[48]), .B(B[48]), .Ci(CTMP[48]), .S(S[48]), .Co(CTMP[49]) );
  FA_783 FAI_50 ( .A(A[49]), .B(B[49]), .Ci(CTMP[49]), .S(S[49]), .Co(CTMP[50]) );
  FA_782 FAI_51 ( .A(A[50]), .B(B[50]), .Ci(CTMP[50]), .S(S[50]), .Co(CTMP[51]) );
  FA_781 FAI_52 ( .A(A[51]), .B(B[51]), .Ci(CTMP[51]), .S(S[51]), .Co(CTMP[52]) );
  FA_780 FAI_53 ( .A(A[52]), .B(B[52]), .Ci(CTMP[52]), .S(S[52]), .Co(CTMP[53]) );
  FA_779 FAI_54 ( .A(A[53]), .B(B[53]), .Ci(CTMP[53]), .S(S[53]), .Co(CTMP[54]) );
  FA_778 FAI_55 ( .A(A[54]), .B(B[54]), .Ci(CTMP[54]), .S(S[54]), .Co(CTMP[55]) );
  FA_777 FAI_56 ( .A(A[55]), .B(B[55]), .Ci(CTMP[55]), .S(S[55]), .Co(CTMP[56]) );
  FA_776 FAI_57 ( .A(A[56]), .B(B[56]), .Ci(CTMP[56]), .S(S[56]), .Co(CTMP[57]) );
  FA_775 FAI_58 ( .A(A[57]), .B(B[57]), .Ci(CTMP[57]), .S(S[57]), .Co(CTMP[58]) );
  FA_774 FAI_59 ( .A(A[58]), .B(B[58]), .Ci(CTMP[58]), .S(S[58]), .Co(CTMP[59]) );
  FA_773 FAI_60 ( .A(A[59]), .B(B[59]), .Ci(CTMP[59]), .S(S[59]), .Co(CTMP[60]) );
  FA_772 FAI_61 ( .A(A[60]), .B(B[60]), .Ci(CTMP[60]), .S(S[60]), .Co(CTMP[61]) );
  FA_771 FAI_62 ( .A(A[61]), .B(B[61]), .Ci(CTMP[61]), .S(S[61]), .Co(CTMP[62]) );
  FA_770 FAI_63 ( .A(A[62]), .B(B[62]), .Ci(CTMP[62]), .S(S[62]), .Co(CTMP[63]) );
  FA_769 FAI_64 ( .A(A[63]), .B(B[63]), .Ci(CTMP[63]), .S(S[63]), .Co(Co) );
endmodule


module booth_mul_row_N64_RADIX3_13 ( prevA, prevSum, encoderIn, nextA, nextSum
 );
  input [63:0] prevA;
  input [63:0] prevSum;
  input [2:0] encoderIn;
  output [63:0] nextA;
  output [63:0] nextSum;
  wire   n5, n6, n7;
  wire   [2:0] encoder_to_mux;
  wire   [63:0] plus2A_s;
  wire   [63:0] minus2A_s;
  wire   [63:0] minus4A_s;
  tri   [63:0] mux_to_adder;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign nextA[51] = n5;
  assign nextA[39] = n6;
  assign nextA[38] = n7;
  assign nextA[0] = 1'b0;

  encoder_N64_RADIX3_13 encoder_1 ( .X(encoderIn), .Z(encoder_to_mux) );
  ShiftnCompl_N64_13 ShiftnCompl_1 ( .plusA(prevA), .plus2A_out({
        plus2A_s[63:1], SYNOPSYS_UNCONNECTED__0}), .minus2A_out(minus2A_s), 
        .plus4A_out({nextA[63:52], n5, nextA[50:40], n6, n7, nextA[37:1], 
        SYNOPSYS_UNCONNECTED__1}), .minus4A_out(minus4A_s) );
  MUX_GENERIC_N64_RADIX3_13 mux_1 ( .plusA({plus2A_s[63:1], 1'b0}), .minusA(
        minus2A_s), .plus2A({nextA[63:52], n5, nextA[50:40], n6, n7, 
        nextA[37:1], 1'b0}), .minus2A(minus4A_s), .SEL(encoder_to_mux), .Y(
        mux_to_adder) );
  RCA_N64_13 rca_1 ( .A(mux_to_adder), .B(prevSum), .Ci(1'b0), .S(nextSum) );
endmodule


module encoder_N64_RADIX3_12 ( X, Z );
  input [2:0] X;
  output [2:0] Z;
  wire   n5, n7, n8;

  OAI22_X1 U1 ( .A1(n8), .A2(n5), .B1(X[2]), .B2(n7), .ZN(Z[1]) );
  INV_X1 U2 ( .A(X[2]), .ZN(n5) );
  AOI21_X1 U3 ( .B1(n8), .B2(n7), .A(X[2]), .ZN(Z[0]) );
  OAI21_X1 U4 ( .B1(X[1]), .B2(X[0]), .A(n7), .ZN(n8) );
  AND3_X1 U5 ( .A1(X[2]), .A2(n7), .A3(n8), .ZN(Z[2]) );
  NAND2_X1 U6 ( .A1(X[1]), .A2(X[0]), .ZN(n7) );
endmodule


module shifter_N64_24 ( \input , shiftLeftOnePos );
  input [63:0] \input ;
  output [63:0] shiftLeftOnePos;
  wire   \input[62] , \input[61] , \input[60] , \input[59] , \input[58] ,
         \input[57] , \input[56] , \input[55] , \input[54] , \input[53] ,
         \input[52] , \input[51] , \input[50] , \input[49] , \input[48] ,
         \input[47] , \input[46] , \input[45] , \input[44] , \input[43] ,
         \input[42] , \input[41] , \input[40] , \input[39] , \input[38] ,
         \input[37] , \input[36] , \input[35] , \input[34] , \input[33] ,
         \input[32] , \input[31] , \input[30] , \input[29] , \input[28] ,
         \input[27] , \input[26] , \input[25] , \input[24] , \input[23] ,
         \input[22] , \input[21] , \input[20] , \input[19] , \input[18] ,
         \input[17] , \input[16] , \input[15] , \input[14] , \input[13] ,
         \input[12] , \input[11] , \input[10] , \input[9] , \input[8] ,
         \input[7] , \input[6] , \input[5] , \input[4] , \input[3] ,
         \input[2] , \input[1] , \input[0] ;
  assign shiftLeftOnePos[0] = 1'b0;
  assign shiftLeftOnePos[63] = \input[62] ;
  assign \input[62]  = \input  [62];
  assign shiftLeftOnePos[62] = \input[61] ;
  assign \input[61]  = \input  [61];
  assign shiftLeftOnePos[61] = \input[60] ;
  assign \input[60]  = \input  [60];
  assign shiftLeftOnePos[60] = \input[59] ;
  assign \input[59]  = \input  [59];
  assign shiftLeftOnePos[59] = \input[58] ;
  assign \input[58]  = \input  [58];
  assign shiftLeftOnePos[58] = \input[57] ;
  assign \input[57]  = \input  [57];
  assign shiftLeftOnePos[57] = \input[56] ;
  assign \input[56]  = \input  [56];
  assign shiftLeftOnePos[56] = \input[55] ;
  assign \input[55]  = \input  [55];
  assign shiftLeftOnePos[55] = \input[54] ;
  assign \input[54]  = \input  [54];
  assign shiftLeftOnePos[54] = \input[53] ;
  assign \input[53]  = \input  [53];
  assign shiftLeftOnePos[53] = \input[52] ;
  assign \input[52]  = \input  [52];
  assign shiftLeftOnePos[52] = \input[51] ;
  assign \input[51]  = \input  [51];
  assign shiftLeftOnePos[51] = \input[50] ;
  assign \input[50]  = \input  [50];
  assign shiftLeftOnePos[50] = \input[49] ;
  assign \input[49]  = \input  [49];
  assign shiftLeftOnePos[49] = \input[48] ;
  assign \input[48]  = \input  [48];
  assign shiftLeftOnePos[48] = \input[47] ;
  assign \input[47]  = \input  [47];
  assign shiftLeftOnePos[47] = \input[46] ;
  assign \input[46]  = \input  [46];
  assign shiftLeftOnePos[46] = \input[45] ;
  assign \input[45]  = \input  [45];
  assign shiftLeftOnePos[45] = \input[44] ;
  assign \input[44]  = \input  [44];
  assign shiftLeftOnePos[44] = \input[43] ;
  assign \input[43]  = \input  [43];
  assign shiftLeftOnePos[43] = \input[42] ;
  assign \input[42]  = \input  [42];
  assign shiftLeftOnePos[42] = \input[41] ;
  assign \input[41]  = \input  [41];
  assign shiftLeftOnePos[41] = \input[40] ;
  assign \input[40]  = \input  [40];
  assign shiftLeftOnePos[40] = \input[39] ;
  assign \input[39]  = \input  [39];
  assign shiftLeftOnePos[39] = \input[38] ;
  assign \input[38]  = \input  [38];
  assign shiftLeftOnePos[38] = \input[37] ;
  assign \input[37]  = \input  [37];
  assign shiftLeftOnePos[37] = \input[36] ;
  assign \input[36]  = \input  [36];
  assign shiftLeftOnePos[36] = \input[35] ;
  assign \input[35]  = \input  [35];
  assign shiftLeftOnePos[35] = \input[34] ;
  assign \input[34]  = \input  [34];
  assign shiftLeftOnePos[34] = \input[33] ;
  assign \input[33]  = \input  [33];
  assign shiftLeftOnePos[33] = \input[32] ;
  assign \input[32]  = \input  [32];
  assign shiftLeftOnePos[32] = \input[31] ;
  assign \input[31]  = \input  [31];
  assign shiftLeftOnePos[31] = \input[30] ;
  assign \input[30]  = \input  [30];
  assign shiftLeftOnePos[30] = \input[29] ;
  assign \input[29]  = \input  [29];
  assign shiftLeftOnePos[29] = \input[28] ;
  assign \input[28]  = \input  [28];
  assign shiftLeftOnePos[28] = \input[27] ;
  assign \input[27]  = \input  [27];
  assign shiftLeftOnePos[27] = \input[26] ;
  assign \input[26]  = \input  [26];
  assign shiftLeftOnePos[26] = \input[25] ;
  assign \input[25]  = \input  [25];
  assign shiftLeftOnePos[25] = \input[24] ;
  assign \input[24]  = \input  [24];
  assign shiftLeftOnePos[24] = \input[23] ;
  assign \input[23]  = \input  [23];
  assign shiftLeftOnePos[23] = \input[22] ;
  assign \input[22]  = \input  [22];
  assign shiftLeftOnePos[22] = \input[21] ;
  assign \input[21]  = \input  [21];
  assign shiftLeftOnePos[21] = \input[20] ;
  assign \input[20]  = \input  [20];
  assign shiftLeftOnePos[20] = \input[19] ;
  assign \input[19]  = \input  [19];
  assign shiftLeftOnePos[19] = \input[18] ;
  assign \input[18]  = \input  [18];
  assign shiftLeftOnePos[18] = \input[17] ;
  assign \input[17]  = \input  [17];
  assign shiftLeftOnePos[17] = \input[16] ;
  assign \input[16]  = \input  [16];
  assign shiftLeftOnePos[16] = \input[15] ;
  assign \input[15]  = \input  [15];
  assign shiftLeftOnePos[15] = \input[14] ;
  assign \input[14]  = \input  [14];
  assign shiftLeftOnePos[14] = \input[13] ;
  assign \input[13]  = \input  [13];
  assign shiftLeftOnePos[13] = \input[12] ;
  assign \input[12]  = \input  [12];
  assign shiftLeftOnePos[12] = \input[11] ;
  assign \input[11]  = \input  [11];
  assign shiftLeftOnePos[11] = \input[10] ;
  assign \input[10]  = \input  [10];
  assign shiftLeftOnePos[10] = \input[9] ;
  assign \input[9]  = \input  [9];
  assign shiftLeftOnePos[9] = \input[8] ;
  assign \input[8]  = \input  [8];
  assign shiftLeftOnePos[8] = \input[7] ;
  assign \input[7]  = \input  [7];
  assign shiftLeftOnePos[7] = \input[6] ;
  assign \input[6]  = \input  [6];
  assign shiftLeftOnePos[6] = \input[5] ;
  assign \input[5]  = \input  [5];
  assign shiftLeftOnePos[5] = \input[4] ;
  assign \input[4]  = \input  [4];
  assign shiftLeftOnePos[4] = \input[3] ;
  assign \input[3]  = \input  [3];
  assign shiftLeftOnePos[3] = \input[2] ;
  assign \input[2]  = \input  [2];
  assign shiftLeftOnePos[2] = \input[1] ;
  assign \input[1]  = \input  [1];
  assign shiftLeftOnePos[1] = \input[0] ;
  assign \input[0]  = \input  [0];

endmodule


module shifter_N64_23 ( \input , shiftLeftOnePos );
  input [63:0] \input ;
  output [63:0] shiftLeftOnePos;
  wire   \input[62] , \input[61] , \input[60] , \input[59] , \input[58] ,
         \input[57] , \input[56] , \input[55] , \input[54] , \input[53] ,
         \input[52] , \input[51] , \input[50] , \input[49] , \input[48] ,
         \input[47] , \input[46] , \input[45] , \input[44] , \input[43] ,
         \input[42] , \input[41] , \input[40] , \input[39] , \input[38] ,
         \input[37] , \input[36] , \input[35] , \input[34] , \input[33] ,
         \input[32] , \input[31] , \input[30] , \input[29] , \input[28] ,
         \input[27] , \input[26] , \input[25] , \input[24] , \input[23] ,
         \input[22] , \input[21] , \input[20] , \input[19] , \input[18] ,
         \input[17] , \input[16] , \input[15] , \input[14] , \input[13] ,
         \input[12] , \input[11] , \input[10] , \input[9] , \input[8] ,
         \input[7] , \input[6] , \input[5] , \input[4] , \input[3] ,
         \input[2] , \input[1] , \input[0] ;
  assign shiftLeftOnePos[0] = 1'b0;
  assign shiftLeftOnePos[63] = \input[62] ;
  assign \input[62]  = \input  [62];
  assign shiftLeftOnePos[62] = \input[61] ;
  assign \input[61]  = \input  [61];
  assign shiftLeftOnePos[61] = \input[60] ;
  assign \input[60]  = \input  [60];
  assign shiftLeftOnePos[60] = \input[59] ;
  assign \input[59]  = \input  [59];
  assign shiftLeftOnePos[59] = \input[58] ;
  assign \input[58]  = \input  [58];
  assign shiftLeftOnePos[58] = \input[57] ;
  assign \input[57]  = \input  [57];
  assign shiftLeftOnePos[57] = \input[56] ;
  assign \input[56]  = \input  [56];
  assign shiftLeftOnePos[56] = \input[55] ;
  assign \input[55]  = \input  [55];
  assign shiftLeftOnePos[55] = \input[54] ;
  assign \input[54]  = \input  [54];
  assign shiftLeftOnePos[54] = \input[53] ;
  assign \input[53]  = \input  [53];
  assign shiftLeftOnePos[53] = \input[52] ;
  assign \input[52]  = \input  [52];
  assign shiftLeftOnePos[52] = \input[51] ;
  assign \input[51]  = \input  [51];
  assign shiftLeftOnePos[51] = \input[50] ;
  assign \input[50]  = \input  [50];
  assign shiftLeftOnePos[50] = \input[49] ;
  assign \input[49]  = \input  [49];
  assign shiftLeftOnePos[49] = \input[48] ;
  assign \input[48]  = \input  [48];
  assign shiftLeftOnePos[48] = \input[47] ;
  assign \input[47]  = \input  [47];
  assign shiftLeftOnePos[47] = \input[46] ;
  assign \input[46]  = \input  [46];
  assign shiftLeftOnePos[46] = \input[45] ;
  assign \input[45]  = \input  [45];
  assign shiftLeftOnePos[45] = \input[44] ;
  assign \input[44]  = \input  [44];
  assign shiftLeftOnePos[44] = \input[43] ;
  assign \input[43]  = \input  [43];
  assign shiftLeftOnePos[43] = \input[42] ;
  assign \input[42]  = \input  [42];
  assign shiftLeftOnePos[42] = \input[41] ;
  assign \input[41]  = \input  [41];
  assign shiftLeftOnePos[41] = \input[40] ;
  assign \input[40]  = \input  [40];
  assign shiftLeftOnePos[40] = \input[39] ;
  assign \input[39]  = \input  [39];
  assign shiftLeftOnePos[39] = \input[38] ;
  assign \input[38]  = \input  [38];
  assign shiftLeftOnePos[38] = \input[37] ;
  assign \input[37]  = \input  [37];
  assign shiftLeftOnePos[37] = \input[36] ;
  assign \input[36]  = \input  [36];
  assign shiftLeftOnePos[36] = \input[35] ;
  assign \input[35]  = \input  [35];
  assign shiftLeftOnePos[35] = \input[34] ;
  assign \input[34]  = \input  [34];
  assign shiftLeftOnePos[34] = \input[33] ;
  assign \input[33]  = \input  [33];
  assign shiftLeftOnePos[33] = \input[32] ;
  assign \input[32]  = \input  [32];
  assign shiftLeftOnePos[32] = \input[31] ;
  assign \input[31]  = \input  [31];
  assign shiftLeftOnePos[31] = \input[30] ;
  assign \input[30]  = \input  [30];
  assign shiftLeftOnePos[30] = \input[29] ;
  assign \input[29]  = \input  [29];
  assign shiftLeftOnePos[29] = \input[28] ;
  assign \input[28]  = \input  [28];
  assign shiftLeftOnePos[28] = \input[27] ;
  assign \input[27]  = \input  [27];
  assign shiftLeftOnePos[27] = \input[26] ;
  assign \input[26]  = \input  [26];
  assign shiftLeftOnePos[26] = \input[25] ;
  assign \input[25]  = \input  [25];
  assign shiftLeftOnePos[25] = \input[24] ;
  assign \input[24]  = \input  [24];
  assign shiftLeftOnePos[24] = \input[23] ;
  assign \input[23]  = \input  [23];
  assign shiftLeftOnePos[23] = \input[22] ;
  assign \input[22]  = \input  [22];
  assign shiftLeftOnePos[22] = \input[21] ;
  assign \input[21]  = \input  [21];
  assign shiftLeftOnePos[21] = \input[20] ;
  assign \input[20]  = \input  [20];
  assign shiftLeftOnePos[20] = \input[19] ;
  assign \input[19]  = \input  [19];
  assign shiftLeftOnePos[19] = \input[18] ;
  assign \input[18]  = \input  [18];
  assign shiftLeftOnePos[18] = \input[17] ;
  assign \input[17]  = \input  [17];
  assign shiftLeftOnePos[17] = \input[16] ;
  assign \input[16]  = \input  [16];
  assign shiftLeftOnePos[16] = \input[15] ;
  assign \input[15]  = \input  [15];
  assign shiftLeftOnePos[15] = \input[14] ;
  assign \input[14]  = \input  [14];
  assign shiftLeftOnePos[14] = \input[13] ;
  assign \input[13]  = \input  [13];
  assign shiftLeftOnePos[13] = \input[12] ;
  assign \input[12]  = \input  [12];
  assign shiftLeftOnePos[12] = \input[11] ;
  assign \input[11]  = \input  [11];
  assign shiftLeftOnePos[11] = \input[10] ;
  assign \input[10]  = \input  [10];
  assign shiftLeftOnePos[10] = \input[9] ;
  assign \input[9]  = \input  [9];
  assign shiftLeftOnePos[9] = \input[8] ;
  assign \input[8]  = \input  [8];
  assign shiftLeftOnePos[8] = \input[7] ;
  assign \input[7]  = \input  [7];
  assign shiftLeftOnePos[7] = \input[6] ;
  assign \input[6]  = \input  [6];
  assign shiftLeftOnePos[6] = \input[5] ;
  assign \input[5]  = \input  [5];
  assign shiftLeftOnePos[5] = \input[4] ;
  assign \input[4]  = \input  [4];
  assign shiftLeftOnePos[4] = \input[3] ;
  assign \input[3]  = \input  [3];
  assign shiftLeftOnePos[3] = \input[2] ;
  assign \input[2]  = \input  [2];
  assign shiftLeftOnePos[2] = \input[1] ;
  assign \input[1]  = \input  [1];
  assign shiftLeftOnePos[1] = \input[0] ;
  assign \input[0]  = \input  [0];

endmodule


module complementer_N64_24_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n190, n191, n192, n193, n194, n196, n197, n198, n199, n200,
         n202, n203, n204, n206, n207, n208, n210, n211, n212, n213, n214,
         n216, n217, n218, n220, n221, n222, n224, n225, n226, n228, n229,
         n230, n232, n233, n234, n235, n237, n238, n239, n241, n242, n243,
         n245, n246, n247, n249, n250, n189, n195, n201, n205, n209, n215,
         n219, n223, n227, n231, n236, n240, n244, n248, n251;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U81 ( .A(n190), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U82 ( .A(n192), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U83 ( .A(n193), .B(B[6]), .Z(DIFF[6]) );
  XOR2_X1 U85 ( .A(n196), .B(B[62]), .Z(DIFF[62]) );
  XOR2_X1 U86 ( .A(n194), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U87 ( .A(n198), .B(B[59]), .Z(DIFF[59]) );
  XOR2_X1 U89 ( .A(n200), .B(B[57]), .Z(DIFF[57]) );
  XOR2_X1 U90 ( .A(n202), .B(B[55]), .Z(DIFF[55]) );
  XOR2_X1 U92 ( .A(n204), .B(B[53]), .Z(DIFF[53]) );
  XOR2_X1 U93 ( .A(n206), .B(B[51]), .Z(DIFF[51]) );
  XOR2_X1 U95 ( .A(n208), .B(B[49]), .Z(DIFF[49]) );
  XOR2_X1 U96 ( .A(n212), .B(B[47]), .Z(DIFF[47]) );
  XOR2_X1 U98 ( .A(n214), .B(B[45]), .Z(DIFF[45]) );
  XOR2_X1 U99 ( .A(n216), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U101 ( .A(n218), .B(B[41]), .Z(DIFF[41]) );
  XOR2_X1 U102 ( .A(n211), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U103 ( .A(n220), .B(B[39]), .Z(DIFF[39]) );
  XOR2_X1 U105 ( .A(n222), .B(B[37]), .Z(DIFF[37]) );
  XOR2_X1 U106 ( .A(n224), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U108 ( .A(n226), .B(B[33]), .Z(DIFF[33]) );
  XOR2_X1 U109 ( .A(n228), .B(B[31]), .Z(DIFF[31]) );
  XOR2_X1 U111 ( .A(n230), .B(B[29]), .Z(DIFF[29]) );
  XOR2_X1 U112 ( .A(n233), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U114 ( .A(n235), .B(B[25]), .Z(DIFF[25]) );
  XOR2_X1 U115 ( .A(n237), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U117 ( .A(n239), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U118 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U119 ( .A(n241), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U121 ( .A(n243), .B(B[17]), .Z(DIFF[17]) );
  XOR2_X1 U122 ( .A(n245), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U124 ( .A(n247), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U125 ( .A(n249), .B(B[11]), .Z(DIFF[11]) );
  XOR2_X1 U1 ( .A(n197), .B(n251), .Z(DIFF[61]) );
  NAND2_X1 U2 ( .A1(n197), .A2(n251), .ZN(n196) );
  XNOR2_X1 U3 ( .A(B[44]), .B(n217), .ZN(DIFF[44]) );
  NOR2_X1 U4 ( .A1(B[43]), .A2(n216), .ZN(n217) );
  OR3_X1 U5 ( .A1(B[45]), .A2(B[46]), .A3(n214), .ZN(n212) );
  OR3_X1 U6 ( .A1(B[53]), .A2(B[54]), .A3(n204), .ZN(n202) );
  OR3_X1 U7 ( .A1(B[49]), .A2(B[50]), .A3(n208), .ZN(n206) );
  OR3_X1 U8 ( .A1(B[43]), .A2(B[44]), .A3(n216), .ZN(n214) );
  OR3_X1 U9 ( .A1(B[55]), .A2(B[56]), .A3(n202), .ZN(n200) );
  XNOR2_X1 U10 ( .A(n189), .B(B[46]), .ZN(DIFF[46]) );
  NOR2_X1 U11 ( .A1(n214), .A2(B[45]), .ZN(n189) );
  XNOR2_X1 U12 ( .A(n195), .B(B[54]), .ZN(DIFF[54]) );
  NOR2_X1 U13 ( .A1(n204), .A2(B[53]), .ZN(n195) );
  XNOR2_X1 U14 ( .A(n201), .B(B[50]), .ZN(DIFF[50]) );
  NOR2_X1 U15 ( .A1(n208), .A2(B[49]), .ZN(n201) );
  NOR3_X1 U16 ( .A1(B[59]), .A2(B[60]), .A3(n198), .ZN(n197) );
  XNOR2_X1 U17 ( .A(B[56]), .B(n203), .ZN(DIFF[56]) );
  NOR2_X1 U18 ( .A1(B[55]), .A2(n202), .ZN(n203) );
  XNOR2_X1 U19 ( .A(B[60]), .B(n199), .ZN(DIFF[60]) );
  NOR2_X1 U20 ( .A1(B[59]), .A2(n198), .ZN(n199) );
  XNOR2_X1 U21 ( .A(B[52]), .B(n207), .ZN(DIFF[52]) );
  NOR2_X1 U22 ( .A1(B[51]), .A2(n206), .ZN(n207) );
  XNOR2_X1 U23 ( .A(B[48]), .B(n213), .ZN(DIFF[48]) );
  NOR2_X1 U24 ( .A1(B[47]), .A2(n212), .ZN(n213) );
  XNOR2_X1 U25 ( .A(B[40]), .B(n221), .ZN(DIFF[40]) );
  NOR2_X1 U26 ( .A1(B[39]), .A2(n220), .ZN(n221) );
  OR3_X1 U27 ( .A1(B[57]), .A2(B[58]), .A3(n200), .ZN(n198) );
  OR3_X1 U28 ( .A1(B[41]), .A2(B[42]), .A3(n218), .ZN(n216) );
  OR3_X1 U29 ( .A1(B[47]), .A2(B[48]), .A3(n212), .ZN(n208) );
  OR3_X1 U30 ( .A1(B[39]), .A2(B[40]), .A3(n220), .ZN(n218) );
  OR3_X1 U31 ( .A1(B[51]), .A2(B[52]), .A3(n206), .ZN(n204) );
  XNOR2_X1 U32 ( .A(n205), .B(B[42]), .ZN(DIFF[42]) );
  NOR2_X1 U33 ( .A1(n218), .A2(B[41]), .ZN(n205) );
  XNOR2_X1 U34 ( .A(n209), .B(B[58]), .ZN(DIFF[58]) );
  NOR2_X1 U35 ( .A1(n200), .A2(B[57]), .ZN(n209) );
  XNOR2_X1 U36 ( .A(n215), .B(B[63]), .ZN(DIFF[63]) );
  NOR2_X1 U37 ( .A1(n196), .A2(B[62]), .ZN(n215) );
  XNOR2_X1 U38 ( .A(n219), .B(B[30]), .ZN(DIFF[30]) );
  NOR2_X1 U39 ( .A1(n230), .A2(B[29]), .ZN(n219) );
  XNOR2_X1 U40 ( .A(n223), .B(B[26]), .ZN(DIFF[26]) );
  NOR2_X1 U41 ( .A1(n235), .A2(B[25]), .ZN(n223) );
  XNOR2_X1 U42 ( .A(n227), .B(B[22]), .ZN(DIFF[22]) );
  NOR2_X1 U43 ( .A1(n239), .A2(B[21]), .ZN(n227) );
  XNOR2_X1 U44 ( .A(n231), .B(B[18]), .ZN(DIFF[18]) );
  NOR2_X1 U45 ( .A1(n243), .A2(B[17]), .ZN(n231) );
  XNOR2_X1 U46 ( .A(n236), .B(B[14]), .ZN(DIFF[14]) );
  NOR2_X1 U47 ( .A1(n247), .A2(B[13]), .ZN(n236) );
  XNOR2_X1 U48 ( .A(B[28]), .B(n234), .ZN(DIFF[28]) );
  NOR2_X1 U49 ( .A1(B[27]), .A2(n233), .ZN(n234) );
  XNOR2_X1 U50 ( .A(B[24]), .B(n238), .ZN(DIFF[24]) );
  NOR2_X1 U51 ( .A1(B[23]), .A2(n237), .ZN(n238) );
  XNOR2_X1 U52 ( .A(B[20]), .B(n242), .ZN(DIFF[20]) );
  NOR2_X1 U53 ( .A1(B[19]), .A2(n241), .ZN(n242) );
  XNOR2_X1 U54 ( .A(B[16]), .B(n246), .ZN(DIFF[16]) );
  NOR2_X1 U55 ( .A1(B[15]), .A2(n245), .ZN(n246) );
  XNOR2_X1 U56 ( .A(B[12]), .B(n250), .ZN(DIFF[12]) );
  NOR2_X1 U57 ( .A1(B[11]), .A2(n249), .ZN(n250) );
  OR3_X1 U58 ( .A1(B[13]), .A2(B[14]), .A3(n247), .ZN(n245) );
  OR3_X1 U59 ( .A1(B[17]), .A2(B[18]), .A3(n243), .ZN(n241) );
  OR3_X1 U60 ( .A1(B[21]), .A2(B[22]), .A3(n239), .ZN(n237) );
  OR3_X1 U61 ( .A1(B[25]), .A2(B[26]), .A3(n235), .ZN(n233) );
  OR3_X1 U62 ( .A1(B[11]), .A2(B[12]), .A3(n249), .ZN(n247) );
  OR3_X1 U63 ( .A1(B[15]), .A2(B[16]), .A3(n245), .ZN(n243) );
  OR3_X1 U64 ( .A1(B[19]), .A2(B[20]), .A3(n241), .ZN(n239) );
  OR3_X1 U65 ( .A1(B[23]), .A2(B[24]), .A3(n237), .ZN(n235) );
  OR3_X1 U66 ( .A1(B[27]), .A2(B[28]), .A3(n233), .ZN(n230) );
  XNOR2_X1 U67 ( .A(B[36]), .B(n225), .ZN(DIFF[36]) );
  NOR2_X1 U68 ( .A1(B[35]), .A2(n224), .ZN(n225) );
  XNOR2_X1 U69 ( .A(B[32]), .B(n229), .ZN(DIFF[32]) );
  NOR2_X1 U70 ( .A1(B[31]), .A2(n228), .ZN(n229) );
  OR3_X1 U71 ( .A1(B[29]), .A2(B[30]), .A3(n230), .ZN(n228) );
  OR3_X1 U72 ( .A1(B[33]), .A2(B[34]), .A3(n226), .ZN(n224) );
  OR3_X1 U73 ( .A1(B[37]), .A2(B[38]), .A3(n222), .ZN(n220) );
  OR3_X1 U74 ( .A1(B[31]), .A2(B[32]), .A3(n228), .ZN(n226) );
  OR3_X1 U75 ( .A1(B[35]), .A2(B[36]), .A3(n224), .ZN(n222) );
  XNOR2_X1 U76 ( .A(n240), .B(B[38]), .ZN(DIFF[38]) );
  NOR2_X1 U77 ( .A1(n222), .A2(B[37]), .ZN(n240) );
  XNOR2_X1 U78 ( .A(n244), .B(B[34]), .ZN(DIFF[34]) );
  NOR2_X1 U79 ( .A1(n226), .A2(B[33]), .ZN(n244) );
  XNOR2_X1 U80 ( .A(n248), .B(B[10]), .ZN(DIFF[10]) );
  NOR2_X1 U84 ( .A1(n190), .A2(B[9]), .ZN(n248) );
  OR3_X1 U88 ( .A1(B[10]), .A2(B[9]), .A3(n190), .ZN(n249) );
  OR3_X1 U91 ( .A1(B[7]), .A2(B[8]), .A3(n192), .ZN(n190) );
  XNOR2_X1 U94 ( .A(B[8]), .B(n191), .ZN(DIFF[8]) );
  NOR2_X1 U97 ( .A1(B[7]), .A2(n192), .ZN(n191) );
  NOR2_X1 U100 ( .A1(B[3]), .A2(n211), .ZN(n210) );
  OR3_X1 U104 ( .A1(B[5]), .A2(B[6]), .A3(n194), .ZN(n192) );
  OR3_X1 U107 ( .A1(B[3]), .A2(B[4]), .A3(n211), .ZN(n194) );
  XNOR2_X1 U110 ( .A(B[4]), .B(n210), .ZN(DIFF[4]) );
  XNOR2_X1 U113 ( .A(B[2]), .B(n232), .ZN(DIFF[2]) );
  OR2_X1 U116 ( .A1(n194), .A2(B[5]), .ZN(n193) );
  OR3_X1 U120 ( .A1(B[1]), .A2(B[2]), .A3(\B[0] ), .ZN(n211) );
  NOR2_X1 U123 ( .A1(\B[0] ), .A2(B[1]), .ZN(n232) );
  INV_X1 U126 ( .A(B[61]), .ZN(n251) );
endmodule


module complementer_N64_24 ( \input , complement2 );
  input [63:0] \input ;
  output [63:0] complement2;


  complementer_N64_24_DW01_sub_0 sub_add_31_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(\input ), .CI(1'b0), .DIFF(complement2) );
endmodule


module complementer_N64_23_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n190, n191, n192, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n189, n193;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U81 ( .A(n190), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U82 ( .A(n192), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U84 ( .A(n195), .B(B[63]), .Z(DIFF[63]) );
  XOR2_X1 U85 ( .A(n196), .B(B[62]), .Z(DIFF[62]) );
  XOR2_X1 U86 ( .A(n194), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U87 ( .A(n198), .B(B[59]), .Z(DIFF[59]) );
  XOR2_X1 U88 ( .A(n201), .B(B[58]), .Z(DIFF[58]) );
  XOR2_X1 U89 ( .A(n200), .B(B[57]), .Z(DIFF[57]) );
  XOR2_X1 U90 ( .A(n202), .B(B[55]), .Z(DIFF[55]) );
  XOR2_X1 U91 ( .A(n205), .B(B[54]), .Z(DIFF[54]) );
  XOR2_X1 U92 ( .A(n204), .B(B[53]), .Z(DIFF[53]) );
  XOR2_X1 U93 ( .A(n206), .B(B[51]), .Z(DIFF[51]) );
  XOR2_X1 U94 ( .A(n209), .B(B[50]), .Z(DIFF[50]) );
  XOR2_X1 U95 ( .A(n208), .B(B[49]), .Z(DIFF[49]) );
  XOR2_X1 U96 ( .A(n212), .B(B[47]), .Z(DIFF[47]) );
  XOR2_X1 U97 ( .A(n215), .B(B[46]), .Z(DIFF[46]) );
  XOR2_X1 U98 ( .A(n214), .B(B[45]), .Z(DIFF[45]) );
  XOR2_X1 U99 ( .A(n216), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U100 ( .A(n219), .B(B[42]), .Z(DIFF[42]) );
  XOR2_X1 U101 ( .A(n218), .B(B[41]), .Z(DIFF[41]) );
  XOR2_X1 U102 ( .A(n211), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U103 ( .A(n220), .B(B[39]), .Z(DIFF[39]) );
  XOR2_X1 U104 ( .A(n223), .B(B[38]), .Z(DIFF[38]) );
  XOR2_X1 U105 ( .A(n222), .B(B[37]), .Z(DIFF[37]) );
  XOR2_X1 U106 ( .A(n224), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U107 ( .A(n227), .B(B[34]), .Z(DIFF[34]) );
  XOR2_X1 U108 ( .A(n226), .B(B[33]), .Z(DIFF[33]) );
  XOR2_X1 U109 ( .A(n228), .B(B[31]), .Z(DIFF[31]) );
  XOR2_X1 U110 ( .A(n231), .B(B[30]), .Z(DIFF[30]) );
  XOR2_X1 U111 ( .A(n230), .B(B[29]), .Z(DIFF[29]) );
  XOR2_X1 U112 ( .A(n233), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U113 ( .A(n236), .B(B[26]), .Z(DIFF[26]) );
  XOR2_X1 U114 ( .A(n235), .B(B[25]), .Z(DIFF[25]) );
  XOR2_X1 U115 ( .A(n237), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U116 ( .A(n240), .B(B[22]), .Z(DIFF[22]) );
  XOR2_X1 U117 ( .A(n239), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U118 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U119 ( .A(n241), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U120 ( .A(n244), .B(B[18]), .Z(DIFF[18]) );
  XOR2_X1 U121 ( .A(n243), .B(B[17]), .Z(DIFF[17]) );
  XOR2_X1 U122 ( .A(n245), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U123 ( .A(n248), .B(B[14]), .Z(DIFF[14]) );
  XOR2_X1 U124 ( .A(n247), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U125 ( .A(n249), .B(B[11]), .Z(DIFF[11]) );
  XOR2_X1 U126 ( .A(n251), .B(B[10]), .Z(DIFF[10]) );
  NAND2_X1 U1 ( .A1(n197), .A2(n193), .ZN(n196) );
  NOR2_X1 U2 ( .A1(B[43]), .A2(n216), .ZN(n217) );
  NOR2_X1 U3 ( .A1(B[47]), .A2(n212), .ZN(n213) );
  NOR2_X1 U4 ( .A1(B[51]), .A2(n206), .ZN(n207) );
  OR3_X1 U5 ( .A1(B[45]), .A2(B[46]), .A3(n214), .ZN(n212) );
  OR3_X1 U6 ( .A1(B[57]), .A2(B[58]), .A3(n200), .ZN(n198) );
  OR3_X1 U7 ( .A1(B[53]), .A2(B[54]), .A3(n204), .ZN(n202) );
  OR3_X1 U8 ( .A1(B[49]), .A2(B[50]), .A3(n208), .ZN(n206) );
  OR3_X1 U9 ( .A1(B[47]), .A2(B[48]), .A3(n212), .ZN(n208) );
  OR3_X1 U10 ( .A1(B[43]), .A2(B[44]), .A3(n216), .ZN(n214) );
  OR3_X1 U11 ( .A1(B[55]), .A2(B[56]), .A3(n202), .ZN(n200) );
  OR3_X1 U12 ( .A1(B[51]), .A2(B[52]), .A3(n206), .ZN(n204) );
  OR2_X1 U13 ( .A1(n214), .A2(B[45]), .ZN(n215) );
  OR2_X1 U14 ( .A1(n208), .A2(B[49]), .ZN(n209) );
  NOR3_X1 U15 ( .A1(B[59]), .A2(B[60]), .A3(n198), .ZN(n197) );
  NOR2_X1 U16 ( .A1(B[55]), .A2(n202), .ZN(n203) );
  NOR2_X1 U17 ( .A1(B[59]), .A2(n198), .ZN(n199) );
  OR2_X1 U18 ( .A1(n200), .A2(B[57]), .ZN(n201) );
  OR2_X1 U19 ( .A1(n204), .A2(B[53]), .ZN(n205) );
  OR2_X1 U20 ( .A1(n196), .A2(B[62]), .ZN(n195) );
  OR3_X1 U21 ( .A1(B[41]), .A2(B[42]), .A3(n218), .ZN(n216) );
  XNOR2_X1 U22 ( .A(B[44]), .B(n217), .ZN(DIFF[44]) );
  XNOR2_X1 U23 ( .A(B[40]), .B(n221), .ZN(DIFF[40]) );
  XNOR2_X1 U24 ( .A(B[52]), .B(n207), .ZN(DIFF[52]) );
  XNOR2_X1 U25 ( .A(B[48]), .B(n213), .ZN(DIFF[48]) );
  OR2_X1 U26 ( .A1(n218), .A2(B[41]), .ZN(n219) );
  XNOR2_X1 U27 ( .A(B[56]), .B(n203), .ZN(DIFF[56]) );
  XNOR2_X1 U28 ( .A(B[60]), .B(n199), .ZN(DIFF[60]) );
  XNOR2_X1 U29 ( .A(n197), .B(B[61]), .ZN(DIFF[61]) );
  XNOR2_X1 U30 ( .A(B[28]), .B(n234), .ZN(DIFF[28]) );
  XNOR2_X1 U31 ( .A(B[24]), .B(n238), .ZN(DIFF[24]) );
  XNOR2_X1 U32 ( .A(B[20]), .B(n242), .ZN(DIFF[20]) );
  NOR2_X1 U33 ( .A1(B[23]), .A2(n237), .ZN(n238) );
  NOR2_X1 U34 ( .A1(B[19]), .A2(n241), .ZN(n242) );
  NOR2_X1 U35 ( .A1(B[15]), .A2(n245), .ZN(n246) );
  NOR2_X1 U36 ( .A1(B[11]), .A2(n249), .ZN(n250) );
  OR3_X1 U37 ( .A1(B[25]), .A2(B[26]), .A3(n235), .ZN(n233) );
  OR3_X1 U38 ( .A1(B[21]), .A2(B[22]), .A3(n239), .ZN(n237) );
  OR3_X1 U39 ( .A1(B[17]), .A2(B[18]), .A3(n243), .ZN(n241) );
  OR3_X1 U40 ( .A1(B[13]), .A2(B[14]), .A3(n247), .ZN(n245) );
  OR3_X1 U41 ( .A1(B[27]), .A2(B[28]), .A3(n233), .ZN(n230) );
  OR3_X1 U42 ( .A1(B[23]), .A2(B[24]), .A3(n237), .ZN(n235) );
  OR3_X1 U43 ( .A1(B[19]), .A2(B[20]), .A3(n241), .ZN(n239) );
  OR3_X1 U44 ( .A1(B[15]), .A2(B[16]), .A3(n245), .ZN(n243) );
  OR3_X1 U45 ( .A1(B[11]), .A2(B[12]), .A3(n249), .ZN(n247) );
  XNOR2_X1 U46 ( .A(B[16]), .B(n246), .ZN(DIFF[16]) );
  XNOR2_X1 U47 ( .A(B[12]), .B(n250), .ZN(DIFF[12]) );
  OR2_X1 U48 ( .A1(n230), .A2(B[29]), .ZN(n231) );
  OR2_X1 U49 ( .A1(n235), .A2(B[25]), .ZN(n236) );
  OR2_X1 U50 ( .A1(n239), .A2(B[21]), .ZN(n240) );
  OR2_X1 U51 ( .A1(n243), .A2(B[17]), .ZN(n244) );
  OR2_X1 U52 ( .A1(n247), .A2(B[13]), .ZN(n248) );
  NOR2_X1 U53 ( .A1(B[35]), .A2(n224), .ZN(n225) );
  NOR2_X1 U54 ( .A1(B[31]), .A2(n228), .ZN(n229) );
  NOR2_X1 U55 ( .A1(B[27]), .A2(n233), .ZN(n234) );
  NOR2_X1 U56 ( .A1(B[39]), .A2(n220), .ZN(n221) );
  OR3_X1 U57 ( .A1(B[37]), .A2(B[38]), .A3(n222), .ZN(n220) );
  OR3_X1 U58 ( .A1(B[33]), .A2(B[34]), .A3(n226), .ZN(n224) );
  OR3_X1 U59 ( .A1(B[29]), .A2(B[30]), .A3(n230), .ZN(n228) );
  OR3_X1 U60 ( .A1(B[35]), .A2(B[36]), .A3(n224), .ZN(n222) );
  OR3_X1 U61 ( .A1(B[31]), .A2(B[32]), .A3(n228), .ZN(n226) );
  OR3_X1 U62 ( .A1(B[39]), .A2(B[40]), .A3(n220), .ZN(n218) );
  XNOR2_X1 U63 ( .A(B[36]), .B(n225), .ZN(DIFF[36]) );
  XNOR2_X1 U64 ( .A(B[32]), .B(n229), .ZN(DIFF[32]) );
  OR2_X1 U65 ( .A1(n222), .A2(B[37]), .ZN(n223) );
  OR2_X1 U66 ( .A1(n226), .A2(B[33]), .ZN(n227) );
  OR2_X1 U67 ( .A1(n190), .A2(B[9]), .ZN(n251) );
  OR3_X1 U68 ( .A1(B[10]), .A2(B[9]), .A3(n190), .ZN(n249) );
  XNOR2_X1 U69 ( .A(B[8]), .B(n191), .ZN(DIFF[8]) );
  XNOR2_X1 U70 ( .A(n189), .B(B[6]), .ZN(DIFF[6]) );
  NOR2_X1 U71 ( .A1(n194), .A2(B[5]), .ZN(n189) );
  NOR2_X1 U72 ( .A1(B[7]), .A2(n192), .ZN(n191) );
  XNOR2_X1 U73 ( .A(B[2]), .B(n232), .ZN(DIFF[2]) );
  NOR2_X1 U74 ( .A1(\B[0] ), .A2(B[1]), .ZN(n232) );
  XNOR2_X1 U75 ( .A(B[4]), .B(n210), .ZN(DIFF[4]) );
  NOR2_X1 U76 ( .A1(B[3]), .A2(n211), .ZN(n210) );
  OR3_X1 U77 ( .A1(B[5]), .A2(B[6]), .A3(n194), .ZN(n192) );
  OR3_X1 U78 ( .A1(B[7]), .A2(B[8]), .A3(n192), .ZN(n190) );
  OR3_X1 U79 ( .A1(B[3]), .A2(B[4]), .A3(n211), .ZN(n194) );
  OR3_X1 U80 ( .A1(B[1]), .A2(B[2]), .A3(\B[0] ), .ZN(n211) );
  INV_X1 U83 ( .A(B[61]), .ZN(n193) );
endmodule


module complementer_N64_23 ( \input , complement2 );
  input [63:0] \input ;
  output [63:0] complement2;


  complementer_N64_23_DW01_sub_0 sub_add_31_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(\input ), .CI(1'b0), .DIFF(complement2) );
endmodule


module ShiftnCompl_N64_12 ( plusA, plus2A_out, minus2A_out, plus4A_out, 
        minus4A_out );
  input [63:0] plusA;
  output [63:0] plus2A_out;
  output [63:0] minus2A_out;
  output [63:0] plus4A_out;
  output [63:0] minus4A_out;
  wire   n11, n12, n2, n13, n14, n15, n16, n17, n18;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign plus2A_out[0] = 1'b0;
  assign plus2A_out[51] = n2;
  assign plus4A_out[0] = 1'b0;

  shifter_N64_24 shifter_1 ( .\input (plusA), .shiftLeftOnePos({
        plus2A_out[63:59], n11, plus2A_out[57:54], n12, plus2A_out[52], n2, 
        plus2A_out[50:49], n13, plus2A_out[47:44], n14, plus2A_out[42:1], 
        SYNOPSYS_UNCONNECTED__0}) );
  shifter_N64_23 shifter_2 ( .\input ({plus2A_out[63:52], n2, plus2A_out[50:1], 
        1'b0}), .shiftLeftOnePos({plus4A_out[63:59], n15, plus4A_out[57:54], 
        n16, plus4A_out[52:49], n17, plus4A_out[47:44], n18, plus4A_out[42:1], 
        SYNOPSYS_UNCONNECTED__1}) );
  complementer_N64_24 complementer_1 ( .\input ({plus2A_out[63:52], n2, 
        plus2A_out[50:1], 1'b0}), .complement2(minus2A_out) );
  complementer_N64_23 complementer_2 ( .\input ({plus4A_out[63:1], 1'b0}), 
        .complement2(minus4A_out) );
  BUF_X1 U1 ( .A(n14), .Z(plus2A_out[43]) );
  BUF_X1 U4 ( .A(n18), .Z(plus4A_out[43]) );
  BUF_X1 U5 ( .A(n17), .Z(plus4A_out[48]) );
  BUF_X1 U6 ( .A(n13), .Z(plus2A_out[48]) );
  BUF_X1 U7 ( .A(n12), .Z(plus2A_out[53]) );
  BUF_X1 U8 ( .A(n11), .Z(plus2A_out[58]) );
  BUF_X1 U9 ( .A(n16), .Z(plus4A_out[53]) );
  BUF_X1 U10 ( .A(n15), .Z(plus4A_out[58]) );
endmodule


module MUX_GENERIC_N64_RADIX3_12 ( plusA, minusA, plus2A, minus2A, SEL, Y );
  input [63:0] plusA;
  input [63:0] minusA;
  input [63:0] plus2A;
  input [63:0] minus2A;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502;
  tri   [63:0] Y;

  TBUF_X1 \Y_tri[56]  ( .A(n445), .EN(n301), .Z(Y[56]) );
  TBUF_X1 \Y_tri[57]  ( .A(n444), .EN(n301), .Z(Y[57]) );
  TBUF_X1 \Y_tri[58]  ( .A(n443), .EN(n301), .Z(Y[58]) );
  TBUF_X1 \Y_tri[60]  ( .A(n441), .EN(n301), .Z(Y[60]) );
  TBUF_X1 \Y_tri[61]  ( .A(n440), .EN(n301), .Z(Y[61]) );
  TBUF_X1 \Y_tri[62]  ( .A(n439), .EN(n301), .Z(Y[62]) );
  TBUF_X1 \Y_tri[63]  ( .A(n438), .EN(n301), .Z(Y[63]) );
  TBUF_X1 \Y_tri[55]  ( .A(n446), .EN(n301), .Z(Y[55]) );
  TBUF_X1 \Y_tri[31]  ( .A(n470), .EN(n298), .Z(Y[31]) );
  TBUF_X1 \Y_tri[32]  ( .A(n469), .EN(n298), .Z(Y[32]) );
  TBUF_X1 \Y_tri[33]  ( .A(n468), .EN(n299), .Z(Y[33]) );
  TBUF_X1 \Y_tri[34]  ( .A(n467), .EN(n299), .Z(Y[34]) );
  TBUF_X1 \Y_tri[35]  ( .A(n466), .EN(n299), .Z(Y[35]) );
  TBUF_X1 \Y_tri[36]  ( .A(n465), .EN(n299), .Z(Y[36]) );
  TBUF_X1 \Y_tri[37]  ( .A(n464), .EN(n299), .Z(Y[37]) );
  TBUF_X1 \Y_tri[38]  ( .A(n463), .EN(n299), .Z(Y[38]) );
  TBUF_X1 \Y_tri[39]  ( .A(n462), .EN(n299), .Z(Y[39]) );
  TBUF_X1 \Y_tri[40]  ( .A(n461), .EN(n299), .Z(Y[40]) );
  TBUF_X1 \Y_tri[41]  ( .A(n460), .EN(n299), .Z(Y[41]) );
  TBUF_X1 \Y_tri[42]  ( .A(n459), .EN(n299), .Z(Y[42]) );
  TBUF_X1 \Y_tri[43]  ( .A(n458), .EN(n299), .Z(Y[43]) );
  TBUF_X1 \Y_tri[44]  ( .A(n457), .EN(n300), .Z(Y[44]) );
  TBUF_X1 \Y_tri[45]  ( .A(n456), .EN(n300), .Z(Y[45]) );
  TBUF_X1 \Y_tri[46]  ( .A(n455), .EN(n300), .Z(Y[46]) );
  TBUF_X1 \Y_tri[47]  ( .A(n454), .EN(n300), .Z(Y[47]) );
  TBUF_X1 \Y_tri[48]  ( .A(n453), .EN(n300), .Z(Y[48]) );
  TBUF_X1 \Y_tri[49]  ( .A(n452), .EN(n300), .Z(Y[49]) );
  TBUF_X1 \Y_tri[50]  ( .A(n451), .EN(n300), .Z(Y[50]) );
  TBUF_X1 \Y_tri[51]  ( .A(n450), .EN(n300), .Z(Y[51]) );
  TBUF_X1 \Y_tri[52]  ( .A(n449), .EN(n300), .Z(Y[52]) );
  TBUF_X1 \Y_tri[53]  ( .A(n448), .EN(n300), .Z(Y[53]) );
  TBUF_X1 \Y_tri[54]  ( .A(n447), .EN(n300), .Z(Y[54]) );
  TBUF_X1 \Y_tri[9]  ( .A(n492), .EN(n296), .Z(Y[9]) );
  TBUF_X1 \Y_tri[11]  ( .A(n490), .EN(n297), .Z(Y[11]) );
  TBUF_X1 \Y_tri[12]  ( .A(n489), .EN(n297), .Z(Y[12]) );
  TBUF_X1 \Y_tri[13]  ( .A(n488), .EN(n297), .Z(Y[13]) );
  TBUF_X1 \Y_tri[14]  ( .A(n487), .EN(n297), .Z(Y[14]) );
  TBUF_X1 \Y_tri[15]  ( .A(n486), .EN(n297), .Z(Y[15]) );
  TBUF_X1 \Y_tri[16]  ( .A(n485), .EN(n297), .Z(Y[16]) );
  TBUF_X1 \Y_tri[17]  ( .A(n484), .EN(n297), .Z(Y[17]) );
  TBUF_X1 \Y_tri[18]  ( .A(n483), .EN(n297), .Z(Y[18]) );
  TBUF_X1 \Y_tri[19]  ( .A(n482), .EN(n297), .Z(Y[19]) );
  TBUF_X1 \Y_tri[20]  ( .A(n481), .EN(n297), .Z(Y[20]) );
  TBUF_X1 \Y_tri[21]  ( .A(n480), .EN(n297), .Z(Y[21]) );
  TBUF_X1 \Y_tri[22]  ( .A(n479), .EN(n298), .Z(Y[22]) );
  TBUF_X1 \Y_tri[23]  ( .A(n478), .EN(n298), .Z(Y[23]) );
  TBUF_X1 \Y_tri[24]  ( .A(n477), .EN(n298), .Z(Y[24]) );
  TBUF_X1 \Y_tri[25]  ( .A(n476), .EN(n298), .Z(Y[25]) );
  TBUF_X1 \Y_tri[26]  ( .A(n475), .EN(n298), .Z(Y[26]) );
  TBUF_X1 \Y_tri[27]  ( .A(n474), .EN(n298), .Z(Y[27]) );
  TBUF_X1 \Y_tri[28]  ( .A(n473), .EN(n298), .Z(Y[28]) );
  TBUF_X1 \Y_tri[29]  ( .A(n472), .EN(n298), .Z(Y[29]) );
  TBUF_X1 \Y_tri[0]  ( .A(n502), .EN(n296), .Z(Y[0]) );
  TBUF_X1 \Y_tri[1]  ( .A(n501), .EN(n296), .Z(Y[1]) );
  TBUF_X1 \Y_tri[3]  ( .A(n499), .EN(n296), .Z(Y[3]) );
  TBUF_X1 \Y_tri[4]  ( .A(n498), .EN(n296), .Z(Y[4]) );
  TBUF_X1 \Y_tri[5]  ( .A(n497), .EN(n296), .Z(Y[5]) );
  TBUF_X1 \Y_tri[6]  ( .A(n496), .EN(n296), .Z(Y[6]) );
  TBUF_X1 \Y_tri[2]  ( .A(n500), .EN(n296), .Z(Y[2]) );
  TBUF_X1 \Y_tri[7]  ( .A(n495), .EN(n296), .Z(Y[7]) );
  TBUF_X1 \Y_tri[8]  ( .A(n494), .EN(n296), .Z(Y[8]) );
  TBUF_X1 \Y_tri[10]  ( .A(n491), .EN(n296), .Z(Y[10]) );
  TBUF_X1 \Y_tri[30]  ( .A(n471), .EN(n298), .Z(Y[30]) );
  TBUF_X1 \Y_tri[59]  ( .A(n442), .EN(n301), .Z(Y[59]) );
  NAND2_X1 U2 ( .A1(n399), .A2(n398), .ZN(n455) );
  AOI22_X1 U3 ( .A1(plusA[46]), .A2(n281), .B1(plus2A[46]), .B2(n275), .ZN(
        n399) );
  AOI22_X1 U4 ( .A1(minus2A[46]), .A2(n293), .B1(minusA[46]), .B2(n287), .ZN(
        n398) );
  NAND2_X1 U5 ( .A1(n395), .A2(n394), .ZN(n457) );
  AOI22_X1 U6 ( .A1(plusA[44]), .A2(n281), .B1(plus2A[44]), .B2(n275), .ZN(
        n395) );
  AOI22_X1 U7 ( .A1(minus2A[44]), .A2(n293), .B1(minusA[44]), .B2(n287), .ZN(
        n394) );
  NAND2_X1 U8 ( .A1(n401), .A2(n400), .ZN(n454) );
  AOI22_X1 U9 ( .A1(plusA[47]), .A2(n281), .B1(plus2A[47]), .B2(n275), .ZN(
        n401) );
  AOI22_X1 U10 ( .A1(minus2A[47]), .A2(n293), .B1(minusA[47]), .B2(n287), .ZN(
        n400) );
  NAND2_X1 U11 ( .A1(n397), .A2(n396), .ZN(n456) );
  AOI22_X1 U12 ( .A1(plusA[45]), .A2(n281), .B1(plus2A[45]), .B2(n275), .ZN(
        n397) );
  AOI22_X1 U13 ( .A1(minus2A[45]), .A2(n293), .B1(minusA[45]), .B2(n287), .ZN(
        n396) );
  NAND2_X1 U14 ( .A1(n393), .A2(n392), .ZN(n458) );
  AOI22_X1 U15 ( .A1(plusA[43]), .A2(n281), .B1(plus2A[43]), .B2(n275), .ZN(
        n393) );
  AOI22_X1 U16 ( .A1(minus2A[43]), .A2(n293), .B1(minusA[43]), .B2(n287), .ZN(
        n392) );
  NAND2_X1 U17 ( .A1(n415), .A2(n414), .ZN(n447) );
  AOI22_X1 U18 ( .A1(plusA[54]), .A2(n282), .B1(plus2A[54]), .B2(n276), .ZN(
        n415) );
  AOI22_X1 U19 ( .A1(minus2A[54]), .A2(n294), .B1(minusA[54]), .B2(n288), .ZN(
        n414) );
  NAND2_X1 U20 ( .A1(n387), .A2(n386), .ZN(n461) );
  AOI22_X1 U21 ( .A1(plusA[40]), .A2(n281), .B1(plus2A[40]), .B2(n275), .ZN(
        n387) );
  AOI22_X1 U22 ( .A1(minus2A[40]), .A2(n293), .B1(minusA[40]), .B2(n287), .ZN(
        n386) );
  NAND2_X1 U23 ( .A1(n417), .A2(n416), .ZN(n446) );
  AOI22_X1 U24 ( .A1(plusA[55]), .A2(n282), .B1(plus2A[55]), .B2(n276), .ZN(
        n417) );
  AOI22_X1 U25 ( .A1(minus2A[55]), .A2(n294), .B1(minusA[55]), .B2(n288), .ZN(
        n416) );
  NAND2_X1 U26 ( .A1(n413), .A2(n412), .ZN(n448) );
  AOI22_X1 U27 ( .A1(plusA[53]), .A2(n282), .B1(plus2A[53]), .B2(n276), .ZN(
        n413) );
  AOI22_X1 U28 ( .A1(minus2A[53]), .A2(n294), .B1(minusA[53]), .B2(n288), .ZN(
        n412) );
  NAND2_X1 U29 ( .A1(n409), .A2(n408), .ZN(n450) );
  AOI22_X1 U30 ( .A1(plusA[51]), .A2(n282), .B1(plus2A[51]), .B2(n276), .ZN(
        n409) );
  AOI22_X1 U31 ( .A1(minus2A[51]), .A2(n294), .B1(minusA[51]), .B2(n288), .ZN(
        n408) );
  NAND2_X1 U32 ( .A1(n405), .A2(n404), .ZN(n452) );
  AOI22_X1 U33 ( .A1(plusA[49]), .A2(n282), .B1(plus2A[49]), .B2(n276), .ZN(
        n405) );
  AOI22_X1 U34 ( .A1(minus2A[49]), .A2(n294), .B1(minusA[49]), .B2(n288), .ZN(
        n404) );
  NAND2_X1 U35 ( .A1(n411), .A2(n410), .ZN(n449) );
  AOI22_X1 U36 ( .A1(plusA[52]), .A2(n282), .B1(plus2A[52]), .B2(n276), .ZN(
        n411) );
  AOI22_X1 U37 ( .A1(minus2A[52]), .A2(n294), .B1(minusA[52]), .B2(n288), .ZN(
        n410) );
  NAND2_X1 U38 ( .A1(n407), .A2(n406), .ZN(n451) );
  AOI22_X1 U39 ( .A1(plusA[50]), .A2(n282), .B1(plus2A[50]), .B2(n276), .ZN(
        n407) );
  AOI22_X1 U40 ( .A1(minus2A[50]), .A2(n294), .B1(minusA[50]), .B2(n288), .ZN(
        n406) );
  NAND2_X1 U41 ( .A1(n403), .A2(n402), .ZN(n453) );
  AOI22_X1 U42 ( .A1(plusA[48]), .A2(n282), .B1(plus2A[48]), .B2(n276), .ZN(
        n403) );
  AOI22_X1 U43 ( .A1(minus2A[48]), .A2(n294), .B1(minusA[48]), .B2(n288), .ZN(
        n402) );
  NAND2_X1 U44 ( .A1(n389), .A2(n388), .ZN(n460) );
  AOI22_X1 U45 ( .A1(plusA[41]), .A2(n281), .B1(plus2A[41]), .B2(n275), .ZN(
        n389) );
  AOI22_X1 U46 ( .A1(minus2A[41]), .A2(n293), .B1(minusA[41]), .B2(n287), .ZN(
        n388) );
  NAND2_X1 U47 ( .A1(n391), .A2(n390), .ZN(n459) );
  AOI22_X1 U48 ( .A1(plusA[42]), .A2(n281), .B1(plus2A[42]), .B2(n275), .ZN(
        n391) );
  AOI22_X1 U49 ( .A1(minus2A[42]), .A2(n293), .B1(minusA[42]), .B2(n287), .ZN(
        n390) );
  NAND2_X1 U50 ( .A1(n425), .A2(n424), .ZN(n442) );
  AOI22_X1 U51 ( .A1(plusA[59]), .A2(n282), .B1(plus2A[59]), .B2(n276), .ZN(
        n425) );
  AOI22_X1 U52 ( .A1(minus2A[59]), .A2(n294), .B1(minusA[59]), .B2(n288), .ZN(
        n424) );
  NAND2_X1 U53 ( .A1(n419), .A2(n418), .ZN(n445) );
  AOI22_X1 U54 ( .A1(plusA[56]), .A2(n282), .B1(plus2A[56]), .B2(n276), .ZN(
        n419) );
  AOI22_X1 U55 ( .A1(minus2A[56]), .A2(n294), .B1(minusA[56]), .B2(n288), .ZN(
        n418) );
  NAND2_X1 U56 ( .A1(n421), .A2(n420), .ZN(n444) );
  AOI22_X1 U57 ( .A1(plusA[57]), .A2(n282), .B1(plus2A[57]), .B2(n276), .ZN(
        n421) );
  AOI22_X1 U58 ( .A1(minus2A[57]), .A2(n294), .B1(minusA[57]), .B2(n288), .ZN(
        n420) );
  NAND2_X1 U59 ( .A1(n437), .A2(n436), .ZN(n438) );
  AOI22_X1 U60 ( .A1(plusA[63]), .A2(n283), .B1(plus2A[63]), .B2(n277), .ZN(
        n437) );
  AOI22_X1 U61 ( .A1(minus2A[63]), .A2(n295), .B1(minusA[63]), .B2(n289), .ZN(
        n436) );
  NAND2_X1 U62 ( .A1(n431), .A2(n430), .ZN(n439) );
  AOI22_X1 U63 ( .A1(plusA[62]), .A2(n283), .B1(plus2A[62]), .B2(n277), .ZN(
        n431) );
  AOI22_X1 U64 ( .A1(minus2A[62]), .A2(n295), .B1(minusA[62]), .B2(n289), .ZN(
        n430) );
  NAND2_X1 U65 ( .A1(n427), .A2(n426), .ZN(n441) );
  AOI22_X1 U66 ( .A1(plusA[60]), .A2(n283), .B1(plus2A[60]), .B2(n277), .ZN(
        n427) );
  AOI22_X1 U67 ( .A1(minus2A[60]), .A2(n295), .B1(minusA[60]), .B2(n289), .ZN(
        n426) );
  NAND2_X1 U68 ( .A1(n423), .A2(n422), .ZN(n443) );
  AOI22_X1 U69 ( .A1(plusA[58]), .A2(n282), .B1(plus2A[58]), .B2(n276), .ZN(
        n423) );
  AOI22_X1 U70 ( .A1(minus2A[58]), .A2(n294), .B1(minusA[58]), .B2(n288), .ZN(
        n422) );
  NAND2_X1 U71 ( .A1(n429), .A2(n428), .ZN(n440) );
  AOI22_X1 U72 ( .A1(plusA[61]), .A2(n283), .B1(plus2A[61]), .B2(n277), .ZN(
        n429) );
  AOI22_X1 U73 ( .A1(minus2A[61]), .A2(n295), .B1(minusA[61]), .B2(n289), .ZN(
        n428) );
  BUF_X1 U74 ( .A(n433), .Z(n278) );
  BUF_X1 U75 ( .A(n435), .Z(n290) );
  BUF_X1 U76 ( .A(n434), .Z(n284) );
  BUF_X1 U77 ( .A(n432), .Z(n272) );
  BUF_X1 U78 ( .A(n493), .Z(n296) );
  NAND2_X1 U79 ( .A1(n327), .A2(n326), .ZN(n491) );
  AOI22_X1 U80 ( .A1(plusA[10]), .A2(n278), .B1(plus2A[10]), .B2(n272), .ZN(
        n327) );
  AOI22_X1 U81 ( .A1(minus2A[10]), .A2(n290), .B1(minusA[10]), .B2(n284), .ZN(
        n326) );
  BUF_X1 U82 ( .A(n433), .Z(n279) );
  BUF_X1 U83 ( .A(n435), .Z(n291) );
  BUF_X1 U84 ( .A(n434), .Z(n285) );
  BUF_X1 U85 ( .A(n432), .Z(n273) );
  BUF_X1 U86 ( .A(n493), .Z(n297) );
  NAND2_X1 U87 ( .A1(n367), .A2(n366), .ZN(n471) );
  AOI22_X1 U88 ( .A1(plusA[30]), .A2(n280), .B1(plus2A[30]), .B2(n274), .ZN(
        n367) );
  AOI22_X1 U89 ( .A1(minus2A[30]), .A2(n292), .B1(minusA[30]), .B2(n286), .ZN(
        n366) );
  NAND2_X1 U90 ( .A1(n365), .A2(n364), .ZN(n472) );
  AOI22_X1 U91 ( .A1(plusA[29]), .A2(n280), .B1(plus2A[29]), .B2(n274), .ZN(
        n365) );
  AOI22_X1 U92 ( .A1(minus2A[29]), .A2(n292), .B1(minusA[29]), .B2(n286), .ZN(
        n364) );
  NAND2_X1 U93 ( .A1(n363), .A2(n362), .ZN(n473) );
  AOI22_X1 U94 ( .A1(plusA[28]), .A2(n280), .B1(plus2A[28]), .B2(n274), .ZN(
        n363) );
  AOI22_X1 U95 ( .A1(minus2A[28]), .A2(n292), .B1(minusA[28]), .B2(n286), .ZN(
        n362) );
  NAND2_X1 U96 ( .A1(n361), .A2(n360), .ZN(n474) );
  AOI22_X1 U97 ( .A1(plusA[27]), .A2(n280), .B1(plus2A[27]), .B2(n274), .ZN(
        n361) );
  AOI22_X1 U98 ( .A1(minus2A[27]), .A2(n292), .B1(minusA[27]), .B2(n286), .ZN(
        n360) );
  NAND2_X1 U99 ( .A1(n359), .A2(n358), .ZN(n475) );
  AOI22_X1 U100 ( .A1(plusA[26]), .A2(n280), .B1(plus2A[26]), .B2(n274), .ZN(
        n359) );
  AOI22_X1 U101 ( .A1(minus2A[26]), .A2(n292), .B1(minusA[26]), .B2(n286), 
        .ZN(n358) );
  NAND2_X1 U102 ( .A1(n357), .A2(n356), .ZN(n476) );
  AOI22_X1 U103 ( .A1(plusA[25]), .A2(n280), .B1(plus2A[25]), .B2(n274), .ZN(
        n357) );
  AOI22_X1 U104 ( .A1(minus2A[25]), .A2(n292), .B1(minusA[25]), .B2(n286), 
        .ZN(n356) );
  NAND2_X1 U105 ( .A1(n355), .A2(n354), .ZN(n477) );
  AOI22_X1 U106 ( .A1(plusA[24]), .A2(n280), .B1(plus2A[24]), .B2(n274), .ZN(
        n355) );
  AOI22_X1 U107 ( .A1(minus2A[24]), .A2(n292), .B1(minusA[24]), .B2(n286), 
        .ZN(n354) );
  NAND2_X1 U108 ( .A1(n353), .A2(n352), .ZN(n478) );
  AOI22_X1 U109 ( .A1(plusA[23]), .A2(n279), .B1(plus2A[23]), .B2(n273), .ZN(
        n353) );
  AOI22_X1 U110 ( .A1(minus2A[23]), .A2(n291), .B1(minusA[23]), .B2(n285), 
        .ZN(n352) );
  NAND2_X1 U111 ( .A1(n351), .A2(n350), .ZN(n479) );
  AOI22_X1 U112 ( .A1(plusA[22]), .A2(n279), .B1(plus2A[22]), .B2(n273), .ZN(
        n351) );
  AOI22_X1 U113 ( .A1(minus2A[22]), .A2(n291), .B1(minusA[22]), .B2(n285), 
        .ZN(n350) );
  NAND2_X1 U114 ( .A1(n349), .A2(n348), .ZN(n480) );
  AOI22_X1 U115 ( .A1(plusA[21]), .A2(n279), .B1(plus2A[21]), .B2(n273), .ZN(
        n349) );
  AOI22_X1 U116 ( .A1(minus2A[21]), .A2(n291), .B1(minusA[21]), .B2(n285), 
        .ZN(n348) );
  NAND2_X1 U117 ( .A1(n347), .A2(n346), .ZN(n481) );
  AOI22_X1 U118 ( .A1(plusA[20]), .A2(n279), .B1(plus2A[20]), .B2(n273), .ZN(
        n347) );
  AOI22_X1 U119 ( .A1(minus2A[20]), .A2(n291), .B1(minusA[20]), .B2(n285), 
        .ZN(n346) );
  NAND2_X1 U120 ( .A1(n345), .A2(n344), .ZN(n482) );
  AOI22_X1 U121 ( .A1(plusA[19]), .A2(n279), .B1(plus2A[19]), .B2(n273), .ZN(
        n345) );
  AOI22_X1 U122 ( .A1(minus2A[19]), .A2(n291), .B1(minusA[19]), .B2(n285), 
        .ZN(n344) );
  NAND2_X1 U123 ( .A1(n343), .A2(n342), .ZN(n483) );
  AOI22_X1 U124 ( .A1(plusA[18]), .A2(n279), .B1(plus2A[18]), .B2(n273), .ZN(
        n343) );
  AOI22_X1 U125 ( .A1(minus2A[18]), .A2(n291), .B1(minusA[18]), .B2(n285), 
        .ZN(n342) );
  NAND2_X1 U126 ( .A1(n341), .A2(n340), .ZN(n484) );
  AOI22_X1 U127 ( .A1(plusA[17]), .A2(n279), .B1(plus2A[17]), .B2(n273), .ZN(
        n341) );
  AOI22_X1 U128 ( .A1(minus2A[17]), .A2(n291), .B1(minusA[17]), .B2(n285), 
        .ZN(n340) );
  NAND2_X1 U129 ( .A1(n337), .A2(n336), .ZN(n486) );
  AOI22_X1 U130 ( .A1(plusA[15]), .A2(n279), .B1(plus2A[15]), .B2(n273), .ZN(
        n337) );
  AOI22_X1 U131 ( .A1(minus2A[15]), .A2(n291), .B1(minusA[15]), .B2(n285), 
        .ZN(n336) );
  NAND2_X1 U132 ( .A1(n335), .A2(n334), .ZN(n487) );
  AOI22_X1 U133 ( .A1(plusA[14]), .A2(n279), .B1(plus2A[14]), .B2(n273), .ZN(
        n335) );
  AOI22_X1 U134 ( .A1(minus2A[14]), .A2(n291), .B1(minusA[14]), .B2(n285), 
        .ZN(n334) );
  NAND2_X1 U135 ( .A1(n333), .A2(n332), .ZN(n488) );
  AOI22_X1 U136 ( .A1(plusA[13]), .A2(n279), .B1(plus2A[13]), .B2(n273), .ZN(
        n333) );
  AOI22_X1 U137 ( .A1(minus2A[13]), .A2(n291), .B1(minusA[13]), .B2(n285), 
        .ZN(n332) );
  NAND2_X1 U138 ( .A1(n329), .A2(n328), .ZN(n490) );
  AOI22_X1 U139 ( .A1(plusA[11]), .A2(n278), .B1(plus2A[11]), .B2(n272), .ZN(
        n329) );
  AOI22_X1 U140 ( .A1(minus2A[11]), .A2(n290), .B1(minusA[11]), .B2(n284), 
        .ZN(n328) );
  NAND2_X1 U141 ( .A1(n339), .A2(n338), .ZN(n485) );
  AOI22_X1 U142 ( .A1(plusA[16]), .A2(n279), .B1(plus2A[16]), .B2(n273), .ZN(
        n339) );
  AOI22_X1 U143 ( .A1(minus2A[16]), .A2(n291), .B1(minusA[16]), .B2(n285), 
        .ZN(n338) );
  NAND2_X1 U144 ( .A1(n331), .A2(n330), .ZN(n489) );
  AOI22_X1 U145 ( .A1(plusA[12]), .A2(n279), .B1(plus2A[12]), .B2(n273), .ZN(
        n331) );
  AOI22_X1 U146 ( .A1(minus2A[12]), .A2(n291), .B1(minusA[12]), .B2(n285), 
        .ZN(n330) );
  BUF_X1 U147 ( .A(n433), .Z(n280) );
  BUF_X1 U148 ( .A(n435), .Z(n292) );
  BUF_X1 U149 ( .A(n434), .Z(n286) );
  BUF_X1 U150 ( .A(n432), .Z(n274) );
  BUF_X1 U151 ( .A(n493), .Z(n298) );
  NAND2_X1 U152 ( .A1(n369), .A2(n368), .ZN(n470) );
  AOI22_X1 U153 ( .A1(plusA[31]), .A2(n280), .B1(plus2A[31]), .B2(n274), .ZN(
        n369) );
  AOI22_X1 U154 ( .A1(minus2A[31]), .A2(n292), .B1(minusA[31]), .B2(n286), 
        .ZN(n368) );
  NAND2_X1 U155 ( .A1(n381), .A2(n380), .ZN(n464) );
  AOI22_X1 U156 ( .A1(plusA[37]), .A2(n281), .B1(plus2A[37]), .B2(n275), .ZN(
        n381) );
  AOI22_X1 U157 ( .A1(minus2A[37]), .A2(n293), .B1(minusA[37]), .B2(n287), 
        .ZN(n380) );
  NAND2_X1 U158 ( .A1(n373), .A2(n372), .ZN(n468) );
  AOI22_X1 U159 ( .A1(plusA[33]), .A2(n280), .B1(plus2A[33]), .B2(n274), .ZN(
        n373) );
  AOI22_X1 U160 ( .A1(minus2A[33]), .A2(n292), .B1(minusA[33]), .B2(n286), 
        .ZN(n372) );
  NAND2_X1 U161 ( .A1(n377), .A2(n376), .ZN(n466) );
  AOI22_X1 U162 ( .A1(plusA[35]), .A2(n280), .B1(plus2A[35]), .B2(n274), .ZN(
        n377) );
  AOI22_X1 U163 ( .A1(minus2A[35]), .A2(n292), .B1(minusA[35]), .B2(n286), 
        .ZN(n376) );
  NAND2_X1 U164 ( .A1(n385), .A2(n384), .ZN(n462) );
  AOI22_X1 U165 ( .A1(plusA[39]), .A2(n281), .B1(plus2A[39]), .B2(n275), .ZN(
        n385) );
  AOI22_X1 U166 ( .A1(minus2A[39]), .A2(n293), .B1(minusA[39]), .B2(n287), 
        .ZN(n384) );
  NAND2_X1 U167 ( .A1(n383), .A2(n382), .ZN(n463) );
  AOI22_X1 U168 ( .A1(plusA[38]), .A2(n281), .B1(plus2A[38]), .B2(n275), .ZN(
        n383) );
  AOI22_X1 U169 ( .A1(minus2A[38]), .A2(n293), .B1(minusA[38]), .B2(n287), 
        .ZN(n382) );
  NAND2_X1 U170 ( .A1(n375), .A2(n374), .ZN(n467) );
  AOI22_X1 U171 ( .A1(plusA[34]), .A2(n280), .B1(plus2A[34]), .B2(n274), .ZN(
        n375) );
  AOI22_X1 U172 ( .A1(minus2A[34]), .A2(n292), .B1(minusA[34]), .B2(n286), 
        .ZN(n374) );
  NAND2_X1 U173 ( .A1(n379), .A2(n378), .ZN(n465) );
  AOI22_X1 U174 ( .A1(plusA[36]), .A2(n281), .B1(plus2A[36]), .B2(n275), .ZN(
        n379) );
  AOI22_X1 U175 ( .A1(minus2A[36]), .A2(n293), .B1(minusA[36]), .B2(n287), 
        .ZN(n378) );
  NAND2_X1 U176 ( .A1(n371), .A2(n370), .ZN(n469) );
  AOI22_X1 U177 ( .A1(plusA[32]), .A2(n280), .B1(plus2A[32]), .B2(n274), .ZN(
        n371) );
  AOI22_X1 U178 ( .A1(minus2A[32]), .A2(n292), .B1(minusA[32]), .B2(n286), 
        .ZN(n370) );
  BUF_X1 U179 ( .A(n433), .Z(n281) );
  BUF_X1 U180 ( .A(n435), .Z(n293) );
  BUF_X1 U181 ( .A(n434), .Z(n287) );
  BUF_X1 U182 ( .A(n432), .Z(n275) );
  BUF_X1 U183 ( .A(n493), .Z(n299) );
  BUF_X1 U184 ( .A(n433), .Z(n282) );
  BUF_X1 U185 ( .A(n435), .Z(n294) );
  BUF_X1 U186 ( .A(n434), .Z(n288) );
  BUF_X1 U187 ( .A(n432), .Z(n276) );
  BUF_X1 U188 ( .A(n493), .Z(n300) );
  BUF_X1 U189 ( .A(n493), .Z(n301) );
  NOR3_X1 U190 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n302), .ZN(n434) );
  NOR3_X1 U191 ( .A1(SEL[1]), .A2(SEL[2]), .A3(n303), .ZN(n433) );
  NOR3_X1 U192 ( .A1(n302), .A2(SEL[2]), .A3(n303), .ZN(n432) );
  NOR2_X1 U193 ( .A1(n323), .A2(n304), .ZN(n493) );
  INV_X1 U194 ( .A(SEL[2]), .ZN(n304) );
  NOR2_X1 U195 ( .A1(SEL[1]), .A2(SEL[0]), .ZN(n323) );
  AND2_X1 U196 ( .A1(SEL[2]), .A2(n323), .ZN(n435) );
  INV_X1 U197 ( .A(SEL[1]), .ZN(n302) );
  INV_X1 U198 ( .A(SEL[0]), .ZN(n303) );
  NAND2_X1 U199 ( .A1(n325), .A2(n324), .ZN(n492) );
  AOI22_X1 U200 ( .A1(plusA[9]), .A2(n278), .B1(plus2A[9]), .B2(n272), .ZN(
        n325) );
  AOI22_X1 U201 ( .A1(minus2A[9]), .A2(n290), .B1(minusA[9]), .B2(n284), .ZN(
        n324) );
  NAND2_X1 U202 ( .A1(n322), .A2(n321), .ZN(n494) );
  AOI22_X1 U203 ( .A1(plusA[8]), .A2(n278), .B1(plus2A[8]), .B2(n272), .ZN(
        n322) );
  AOI22_X1 U204 ( .A1(minus2A[8]), .A2(n290), .B1(minusA[8]), .B2(n284), .ZN(
        n321) );
  NAND2_X1 U205 ( .A1(n320), .A2(n319), .ZN(n495) );
  AOI22_X1 U206 ( .A1(plusA[7]), .A2(n278), .B1(plus2A[7]), .B2(n272), .ZN(
        n320) );
  AOI22_X1 U207 ( .A1(minus2A[7]), .A2(n290), .B1(minusA[7]), .B2(n284), .ZN(
        n319) );
  NAND2_X1 U208 ( .A1(n318), .A2(n317), .ZN(n496) );
  AOI22_X1 U209 ( .A1(plusA[6]), .A2(n278), .B1(plus2A[6]), .B2(n272), .ZN(
        n318) );
  AOI22_X1 U210 ( .A1(minus2A[6]), .A2(n290), .B1(minusA[6]), .B2(n284), .ZN(
        n317) );
  NAND2_X1 U211 ( .A1(n316), .A2(n315), .ZN(n497) );
  AOI22_X1 U212 ( .A1(plusA[5]), .A2(n278), .B1(plus2A[5]), .B2(n272), .ZN(
        n316) );
  AOI22_X1 U213 ( .A1(minus2A[5]), .A2(n290), .B1(minusA[5]), .B2(n284), .ZN(
        n315) );
  NAND2_X1 U214 ( .A1(n312), .A2(n311), .ZN(n499) );
  AOI22_X1 U215 ( .A1(plusA[3]), .A2(n278), .B1(plus2A[3]), .B2(n272), .ZN(
        n312) );
  AOI22_X1 U216 ( .A1(minus2A[3]), .A2(n290), .B1(minusA[3]), .B2(n284), .ZN(
        n311) );
  NAND2_X1 U217 ( .A1(n314), .A2(n313), .ZN(n498) );
  AOI22_X1 U218 ( .A1(plusA[4]), .A2(n278), .B1(plus2A[4]), .B2(n272), .ZN(
        n314) );
  AOI22_X1 U219 ( .A1(minus2A[4]), .A2(n290), .B1(minusA[4]), .B2(n284), .ZN(
        n313) );
  NAND2_X1 U220 ( .A1(n310), .A2(n309), .ZN(n500) );
  AOI22_X1 U221 ( .A1(plusA[2]), .A2(n278), .B1(plus2A[2]), .B2(n272), .ZN(
        n310) );
  AOI22_X1 U222 ( .A1(minus2A[2]), .A2(n290), .B1(minusA[2]), .B2(n284), .ZN(
        n309) );
  NAND2_X1 U223 ( .A1(n308), .A2(n307), .ZN(n501) );
  AOI22_X1 U224 ( .A1(plusA[1]), .A2(n278), .B1(plus2A[1]), .B2(n272), .ZN(
        n308) );
  AOI22_X1 U225 ( .A1(minus2A[1]), .A2(n290), .B1(minusA[1]), .B2(n284), .ZN(
        n307) );
  NAND2_X1 U226 ( .A1(n306), .A2(n305), .ZN(n502) );
  AOI22_X1 U227 ( .A1(plusA[0]), .A2(n278), .B1(plus2A[0]), .B2(n272), .ZN(
        n306) );
  AOI22_X1 U228 ( .A1(minus2A[0]), .A2(n290), .B1(minusA[0]), .B2(n284), .ZN(
        n305) );
  CLKBUF_X1 U229 ( .A(n432), .Z(n277) );
  CLKBUF_X1 U230 ( .A(n433), .Z(n283) );
  CLKBUF_X1 U231 ( .A(n434), .Z(n289) );
  CLKBUF_X1 U232 ( .A(n435), .Z(n295) );
endmodule


module FA_768 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_767 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_766 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_765 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_764 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_763 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_762 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_761 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  AOI22_X1 U4 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
  INV_X1 U5 ( .A(n7), .ZN(Co) );
endmodule


module FA_760 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  AOI22_X1 U4 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
  INV_X1 U5 ( .A(n7), .ZN(Co) );
endmodule


module FA_759 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_758 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  AOI22_X1 U4 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
  INV_X1 U5 ( .A(n7), .ZN(Co) );
endmodule


module FA_757 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_756 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_755 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_754 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_753 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_752 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_751 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_750 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_749 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_748 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_747 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_746 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_745 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_744 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_743 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_742 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_741 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_740 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_739 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_738 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_737 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_736 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_735 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_734 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_733 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_732 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_731 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_730 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_729 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_728 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_727 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_726 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_725 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_724 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_723 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_722 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_721 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_720 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_719 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_718 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_717 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_716 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_715 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_714 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_713 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_712 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_711 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_710 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_709 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  AOI22_X1 U4 ( .A1(B), .A2(A), .B1(Ci), .B2(n6), .ZN(n7) );
  INV_X1 U5 ( .A(n7), .ZN(Co) );
endmodule


module FA_708 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_707 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_706 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_705 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N64_12 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Ci;
  output Co;

  wire   [63:1] CTMP;
  tri   [63:0] A;

  FA_768 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_767 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_766 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_765 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(CTMP[4]) );
  FA_764 FAI_5 ( .A(A[4]), .B(B[4]), .Ci(CTMP[4]), .S(S[4]), .Co(CTMP[5]) );
  FA_763 FAI_6 ( .A(A[5]), .B(B[5]), .Ci(CTMP[5]), .S(S[5]), .Co(CTMP[6]) );
  FA_762 FAI_7 ( .A(A[6]), .B(B[6]), .Ci(CTMP[6]), .S(S[6]), .Co(CTMP[7]) );
  FA_761 FAI_8 ( .A(A[7]), .B(B[7]), .Ci(CTMP[7]), .S(S[7]), .Co(CTMP[8]) );
  FA_760 FAI_9 ( .A(A[8]), .B(B[8]), .Ci(CTMP[8]), .S(S[8]), .Co(CTMP[9]) );
  FA_759 FAI_10 ( .A(A[9]), .B(B[9]), .Ci(CTMP[9]), .S(S[9]), .Co(CTMP[10]) );
  FA_758 FAI_11 ( .A(A[10]), .B(B[10]), .Ci(CTMP[10]), .S(S[10]), .Co(CTMP[11]) );
  FA_757 FAI_12 ( .A(A[11]), .B(B[11]), .Ci(CTMP[11]), .S(S[11]), .Co(CTMP[12]) );
  FA_756 FAI_13 ( .A(A[12]), .B(B[12]), .Ci(CTMP[12]), .S(S[12]), .Co(CTMP[13]) );
  FA_755 FAI_14 ( .A(A[13]), .B(B[13]), .Ci(CTMP[13]), .S(S[13]), .Co(CTMP[14]) );
  FA_754 FAI_15 ( .A(A[14]), .B(B[14]), .Ci(CTMP[14]), .S(S[14]), .Co(CTMP[15]) );
  FA_753 FAI_16 ( .A(A[15]), .B(B[15]), .Ci(CTMP[15]), .S(S[15]), .Co(CTMP[16]) );
  FA_752 FAI_17 ( .A(A[16]), .B(B[16]), .Ci(CTMP[16]), .S(S[16]), .Co(CTMP[17]) );
  FA_751 FAI_18 ( .A(A[17]), .B(B[17]), .Ci(CTMP[17]), .S(S[17]), .Co(CTMP[18]) );
  FA_750 FAI_19 ( .A(A[18]), .B(B[18]), .Ci(CTMP[18]), .S(S[18]), .Co(CTMP[19]) );
  FA_749 FAI_20 ( .A(A[19]), .B(B[19]), .Ci(CTMP[19]), .S(S[19]), .Co(CTMP[20]) );
  FA_748 FAI_21 ( .A(A[20]), .B(B[20]), .Ci(CTMP[20]), .S(S[20]), .Co(CTMP[21]) );
  FA_747 FAI_22 ( .A(A[21]), .B(B[21]), .Ci(CTMP[21]), .S(S[21]), .Co(CTMP[22]) );
  FA_746 FAI_23 ( .A(A[22]), .B(B[22]), .Ci(CTMP[22]), .S(S[22]), .Co(CTMP[23]) );
  FA_745 FAI_24 ( .A(A[23]), .B(B[23]), .Ci(CTMP[23]), .S(S[23]), .Co(CTMP[24]) );
  FA_744 FAI_25 ( .A(A[24]), .B(B[24]), .Ci(CTMP[24]), .S(S[24]), .Co(CTMP[25]) );
  FA_743 FAI_26 ( .A(A[25]), .B(B[25]), .Ci(CTMP[25]), .S(S[25]), .Co(CTMP[26]) );
  FA_742 FAI_27 ( .A(A[26]), .B(B[26]), .Ci(CTMP[26]), .S(S[26]), .Co(CTMP[27]) );
  FA_741 FAI_28 ( .A(A[27]), .B(B[27]), .Ci(CTMP[27]), .S(S[27]), .Co(CTMP[28]) );
  FA_740 FAI_29 ( .A(A[28]), .B(B[28]), .Ci(CTMP[28]), .S(S[28]), .Co(CTMP[29]) );
  FA_739 FAI_30 ( .A(A[29]), .B(B[29]), .Ci(CTMP[29]), .S(S[29]), .Co(CTMP[30]) );
  FA_738 FAI_31 ( .A(A[30]), .B(B[30]), .Ci(CTMP[30]), .S(S[30]), .Co(CTMP[31]) );
  FA_737 FAI_32 ( .A(A[31]), .B(B[31]), .Ci(CTMP[31]), .S(S[31]), .Co(CTMP[32]) );
  FA_736 FAI_33 ( .A(A[32]), .B(B[32]), .Ci(CTMP[32]), .S(S[32]), .Co(CTMP[33]) );
  FA_735 FAI_34 ( .A(A[33]), .B(B[33]), .Ci(CTMP[33]), .S(S[33]), .Co(CTMP[34]) );
  FA_734 FAI_35 ( .A(A[34]), .B(B[34]), .Ci(CTMP[34]), .S(S[34]), .Co(CTMP[35]) );
  FA_733 FAI_36 ( .A(A[35]), .B(B[35]), .Ci(CTMP[35]), .S(S[35]), .Co(CTMP[36]) );
  FA_732 FAI_37 ( .A(A[36]), .B(B[36]), .Ci(CTMP[36]), .S(S[36]), .Co(CTMP[37]) );
  FA_731 FAI_38 ( .A(A[37]), .B(B[37]), .Ci(CTMP[37]), .S(S[37]), .Co(CTMP[38]) );
  FA_730 FAI_39 ( .A(A[38]), .B(B[38]), .Ci(CTMP[38]), .S(S[38]), .Co(CTMP[39]) );
  FA_729 FAI_40 ( .A(A[39]), .B(B[39]), .Ci(CTMP[39]), .S(S[39]), .Co(CTMP[40]) );
  FA_728 FAI_41 ( .A(A[40]), .B(B[40]), .Ci(CTMP[40]), .S(S[40]), .Co(CTMP[41]) );
  FA_727 FAI_42 ( .A(A[41]), .B(B[41]), .Ci(CTMP[41]), .S(S[41]), .Co(CTMP[42]) );
  FA_726 FAI_43 ( .A(A[42]), .B(B[42]), .Ci(CTMP[42]), .S(S[42]), .Co(CTMP[43]) );
  FA_725 FAI_44 ( .A(A[43]), .B(B[43]), .Ci(CTMP[43]), .S(S[43]), .Co(CTMP[44]) );
  FA_724 FAI_45 ( .A(A[44]), .B(B[44]), .Ci(CTMP[44]), .S(S[44]), .Co(CTMP[45]) );
  FA_723 FAI_46 ( .A(A[45]), .B(B[45]), .Ci(CTMP[45]), .S(S[45]), .Co(CTMP[46]) );
  FA_722 FAI_47 ( .A(A[46]), .B(B[46]), .Ci(CTMP[46]), .S(S[46]), .Co(CTMP[47]) );
  FA_721 FAI_48 ( .A(A[47]), .B(B[47]), .Ci(CTMP[47]), .S(S[47]), .Co(CTMP[48]) );
  FA_720 FAI_49 ( .A(A[48]), .B(B[48]), .Ci(CTMP[48]), .S(S[48]), .Co(CTMP[49]) );
  FA_719 FAI_50 ( .A(A[49]), .B(B[49]), .Ci(CTMP[49]), .S(S[49]), .Co(CTMP[50]) );
  FA_718 FAI_51 ( .A(A[50]), .B(B[50]), .Ci(CTMP[50]), .S(S[50]), .Co(CTMP[51]) );
  FA_717 FAI_52 ( .A(A[51]), .B(B[51]), .Ci(CTMP[51]), .S(S[51]), .Co(CTMP[52]) );
  FA_716 FAI_53 ( .A(A[52]), .B(B[52]), .Ci(CTMP[52]), .S(S[52]), .Co(CTMP[53]) );
  FA_715 FAI_54 ( .A(A[53]), .B(B[53]), .Ci(CTMP[53]), .S(S[53]), .Co(CTMP[54]) );
  FA_714 FAI_55 ( .A(A[54]), .B(B[54]), .Ci(CTMP[54]), .S(S[54]), .Co(CTMP[55]) );
  FA_713 FAI_56 ( .A(A[55]), .B(B[55]), .Ci(CTMP[55]), .S(S[55]), .Co(CTMP[56]) );
  FA_712 FAI_57 ( .A(A[56]), .B(B[56]), .Ci(CTMP[56]), .S(S[56]), .Co(CTMP[57]) );
  FA_711 FAI_58 ( .A(A[57]), .B(B[57]), .Ci(CTMP[57]), .S(S[57]), .Co(CTMP[58]) );
  FA_710 FAI_59 ( .A(A[58]), .B(B[58]), .Ci(CTMP[58]), .S(S[58]), .Co(CTMP[59]) );
  FA_709 FAI_60 ( .A(A[59]), .B(B[59]), .Ci(CTMP[59]), .S(S[59]), .Co(CTMP[60]) );
  FA_708 FAI_61 ( .A(A[60]), .B(B[60]), .Ci(CTMP[60]), .S(S[60]), .Co(CTMP[61]) );
  FA_707 FAI_62 ( .A(A[61]), .B(B[61]), .Ci(CTMP[61]), .S(S[61]), .Co(CTMP[62]) );
  FA_706 FAI_63 ( .A(A[62]), .B(B[62]), .Ci(CTMP[62]), .S(S[62]), .Co(CTMP[63]) );
  FA_705 FAI_64 ( .A(A[63]), .B(B[63]), .Ci(CTMP[63]), .S(S[63]), .Co(Co) );
endmodule


module booth_mul_row_N64_RADIX3_12 ( prevA, prevSum, encoderIn, nextA, nextSum
 );
  input [63:0] prevA;
  input [63:0] prevSum;
  input [2:0] encoderIn;
  output [63:0] nextA;
  output [63:0] nextSum;
  wire   n3;
  wire   [2:0] encoder_to_mux;
  wire   [63:0] plus2A_s;
  wire   [63:0] minus2A_s;
  wire   [63:0] minus4A_s;
  tri   [63:0] mux_to_adder;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign nextA[51] = n3;
  assign nextA[0] = 1'b0;

  encoder_N64_RADIX3_12 encoder_1 ( .X(encoderIn), .Z(encoder_to_mux) );
  ShiftnCompl_N64_12 ShiftnCompl_1 ( .plusA(prevA), .plus2A_out({
        plus2A_s[63:1], SYNOPSYS_UNCONNECTED__0}), .minus2A_out(minus2A_s), 
        .plus4A_out({nextA[63:52], n3, nextA[50:1], SYNOPSYS_UNCONNECTED__1}), 
        .minus4A_out(minus4A_s) );
  MUX_GENERIC_N64_RADIX3_12 mux_1 ( .plusA({plus2A_s[63:1], 1'b0}), .minusA(
        minus2A_s), .plus2A({nextA[63:52], n3, nextA[50:1], 1'b0}), .minus2A(
        minus4A_s), .SEL(encoder_to_mux), .Y(mux_to_adder) );
  RCA_N64_12 rca_1 ( .A(mux_to_adder), .B(prevSum), .Ci(1'b0), .S(nextSum) );
endmodule


module encoder_N64_RADIX3_11 ( X, Z );
  input [2:0] X;
  output [2:0] Z;
  wire   n5, n7, n8;

  OAI22_X1 U1 ( .A1(n8), .A2(n5), .B1(X[2]), .B2(n7), .ZN(Z[1]) );
  INV_X1 U2 ( .A(X[2]), .ZN(n5) );
  AOI21_X1 U3 ( .B1(n8), .B2(n7), .A(X[2]), .ZN(Z[0]) );
  OAI21_X1 U4 ( .B1(X[1]), .B2(X[0]), .A(n7), .ZN(n8) );
  AND3_X1 U5 ( .A1(X[2]), .A2(n7), .A3(n8), .ZN(Z[2]) );
  NAND2_X1 U6 ( .A1(X[1]), .A2(X[0]), .ZN(n7) );
endmodule


module shifter_N64_22 ( \input , shiftLeftOnePos );
  input [63:0] \input ;
  output [63:0] shiftLeftOnePos;
  wire   \input[62] , \input[61] , \input[60] , \input[59] , \input[58] ,
         \input[57] , \input[56] , \input[55] , \input[54] , \input[53] ,
         \input[52] , \input[51] , \input[50] , \input[49] , \input[48] ,
         \input[47] , \input[46] , \input[45] , \input[44] , \input[43] ,
         \input[42] , \input[41] , \input[40] , \input[39] , \input[38] ,
         \input[37] , \input[36] , \input[35] , \input[34] , \input[33] ,
         \input[32] , \input[31] , \input[30] , \input[29] , \input[28] ,
         \input[27] , \input[26] , \input[25] , \input[24] , \input[23] ,
         \input[22] , \input[21] , \input[20] , \input[19] , \input[18] ,
         \input[17] , \input[16] , \input[15] , \input[14] , \input[13] ,
         \input[12] , \input[11] , \input[10] , \input[9] , \input[8] ,
         \input[7] , \input[6] , \input[5] , \input[4] , \input[3] ,
         \input[2] , \input[1] , \input[0] ;
  assign shiftLeftOnePos[0] = 1'b0;
  assign shiftLeftOnePos[63] = \input[62] ;
  assign \input[62]  = \input  [62];
  assign shiftLeftOnePos[62] = \input[61] ;
  assign \input[61]  = \input  [61];
  assign shiftLeftOnePos[61] = \input[60] ;
  assign \input[60]  = \input  [60];
  assign shiftLeftOnePos[60] = \input[59] ;
  assign \input[59]  = \input  [59];
  assign shiftLeftOnePos[59] = \input[58] ;
  assign \input[58]  = \input  [58];
  assign shiftLeftOnePos[58] = \input[57] ;
  assign \input[57]  = \input  [57];
  assign shiftLeftOnePos[57] = \input[56] ;
  assign \input[56]  = \input  [56];
  assign shiftLeftOnePos[56] = \input[55] ;
  assign \input[55]  = \input  [55];
  assign shiftLeftOnePos[55] = \input[54] ;
  assign \input[54]  = \input  [54];
  assign shiftLeftOnePos[54] = \input[53] ;
  assign \input[53]  = \input  [53];
  assign shiftLeftOnePos[53] = \input[52] ;
  assign \input[52]  = \input  [52];
  assign shiftLeftOnePos[52] = \input[51] ;
  assign \input[51]  = \input  [51];
  assign shiftLeftOnePos[51] = \input[50] ;
  assign \input[50]  = \input  [50];
  assign shiftLeftOnePos[50] = \input[49] ;
  assign \input[49]  = \input  [49];
  assign shiftLeftOnePos[49] = \input[48] ;
  assign \input[48]  = \input  [48];
  assign shiftLeftOnePos[48] = \input[47] ;
  assign \input[47]  = \input  [47];
  assign shiftLeftOnePos[47] = \input[46] ;
  assign \input[46]  = \input  [46];
  assign shiftLeftOnePos[46] = \input[45] ;
  assign \input[45]  = \input  [45];
  assign shiftLeftOnePos[45] = \input[44] ;
  assign \input[44]  = \input  [44];
  assign shiftLeftOnePos[44] = \input[43] ;
  assign \input[43]  = \input  [43];
  assign shiftLeftOnePos[43] = \input[42] ;
  assign \input[42]  = \input  [42];
  assign shiftLeftOnePos[42] = \input[41] ;
  assign \input[41]  = \input  [41];
  assign shiftLeftOnePos[41] = \input[40] ;
  assign \input[40]  = \input  [40];
  assign shiftLeftOnePos[40] = \input[39] ;
  assign \input[39]  = \input  [39];
  assign shiftLeftOnePos[39] = \input[38] ;
  assign \input[38]  = \input  [38];
  assign shiftLeftOnePos[38] = \input[37] ;
  assign \input[37]  = \input  [37];
  assign shiftLeftOnePos[37] = \input[36] ;
  assign \input[36]  = \input  [36];
  assign shiftLeftOnePos[36] = \input[35] ;
  assign \input[35]  = \input  [35];
  assign shiftLeftOnePos[35] = \input[34] ;
  assign \input[34]  = \input  [34];
  assign shiftLeftOnePos[34] = \input[33] ;
  assign \input[33]  = \input  [33];
  assign shiftLeftOnePos[33] = \input[32] ;
  assign \input[32]  = \input  [32];
  assign shiftLeftOnePos[32] = \input[31] ;
  assign \input[31]  = \input  [31];
  assign shiftLeftOnePos[31] = \input[30] ;
  assign \input[30]  = \input  [30];
  assign shiftLeftOnePos[30] = \input[29] ;
  assign \input[29]  = \input  [29];
  assign shiftLeftOnePos[29] = \input[28] ;
  assign \input[28]  = \input  [28];
  assign shiftLeftOnePos[28] = \input[27] ;
  assign \input[27]  = \input  [27];
  assign shiftLeftOnePos[27] = \input[26] ;
  assign \input[26]  = \input  [26];
  assign shiftLeftOnePos[26] = \input[25] ;
  assign \input[25]  = \input  [25];
  assign shiftLeftOnePos[25] = \input[24] ;
  assign \input[24]  = \input  [24];
  assign shiftLeftOnePos[24] = \input[23] ;
  assign \input[23]  = \input  [23];
  assign shiftLeftOnePos[23] = \input[22] ;
  assign \input[22]  = \input  [22];
  assign shiftLeftOnePos[22] = \input[21] ;
  assign \input[21]  = \input  [21];
  assign shiftLeftOnePos[21] = \input[20] ;
  assign \input[20]  = \input  [20];
  assign shiftLeftOnePos[20] = \input[19] ;
  assign \input[19]  = \input  [19];
  assign shiftLeftOnePos[19] = \input[18] ;
  assign \input[18]  = \input  [18];
  assign shiftLeftOnePos[18] = \input[17] ;
  assign \input[17]  = \input  [17];
  assign shiftLeftOnePos[17] = \input[16] ;
  assign \input[16]  = \input  [16];
  assign shiftLeftOnePos[16] = \input[15] ;
  assign \input[15]  = \input  [15];
  assign shiftLeftOnePos[15] = \input[14] ;
  assign \input[14]  = \input  [14];
  assign shiftLeftOnePos[14] = \input[13] ;
  assign \input[13]  = \input  [13];
  assign shiftLeftOnePos[13] = \input[12] ;
  assign \input[12]  = \input  [12];
  assign shiftLeftOnePos[12] = \input[11] ;
  assign \input[11]  = \input  [11];
  assign shiftLeftOnePos[11] = \input[10] ;
  assign \input[10]  = \input  [10];
  assign shiftLeftOnePos[10] = \input[9] ;
  assign \input[9]  = \input  [9];
  assign shiftLeftOnePos[9] = \input[8] ;
  assign \input[8]  = \input  [8];
  assign shiftLeftOnePos[8] = \input[7] ;
  assign \input[7]  = \input  [7];
  assign shiftLeftOnePos[7] = \input[6] ;
  assign \input[6]  = \input  [6];
  assign shiftLeftOnePos[6] = \input[5] ;
  assign \input[5]  = \input  [5];
  assign shiftLeftOnePos[5] = \input[4] ;
  assign \input[4]  = \input  [4];
  assign shiftLeftOnePos[4] = \input[3] ;
  assign \input[3]  = \input  [3];
  assign shiftLeftOnePos[3] = \input[2] ;
  assign \input[2]  = \input  [2];
  assign shiftLeftOnePos[2] = \input[1] ;
  assign \input[1]  = \input  [1];
  assign shiftLeftOnePos[1] = \input[0] ;
  assign \input[0]  = \input  [0];

endmodule


module shifter_N64_21 ( \input , shiftLeftOnePos );
  input [63:0] \input ;
  output [63:0] shiftLeftOnePos;
  wire   \input[62] , \input[61] , \input[60] , \input[59] , \input[58] ,
         \input[57] , \input[56] , \input[55] , \input[54] , \input[53] ,
         \input[52] , \input[51] , \input[50] , \input[49] , \input[48] ,
         \input[47] , \input[46] , \input[45] , \input[44] , \input[43] ,
         \input[42] , \input[41] , \input[40] , \input[39] , \input[38] ,
         \input[37] , \input[36] , \input[35] , \input[34] , \input[33] ,
         \input[32] , \input[31] , \input[30] , \input[29] , \input[28] ,
         \input[27] , \input[26] , \input[25] , \input[24] , \input[23] ,
         \input[22] , \input[21] , \input[20] , \input[19] , \input[18] ,
         \input[17] , \input[16] , \input[15] , \input[14] , \input[13] ,
         \input[12] , \input[11] , \input[10] , \input[9] , \input[8] ,
         \input[7] , \input[6] , \input[5] , \input[4] , \input[3] ,
         \input[2] , \input[1] , \input[0] ;
  assign shiftLeftOnePos[0] = 1'b0;
  assign shiftLeftOnePos[63] = \input[62] ;
  assign \input[62]  = \input  [62];
  assign shiftLeftOnePos[62] = \input[61] ;
  assign \input[61]  = \input  [61];
  assign shiftLeftOnePos[61] = \input[60] ;
  assign \input[60]  = \input  [60];
  assign shiftLeftOnePos[60] = \input[59] ;
  assign \input[59]  = \input  [59];
  assign shiftLeftOnePos[59] = \input[58] ;
  assign \input[58]  = \input  [58];
  assign shiftLeftOnePos[58] = \input[57] ;
  assign \input[57]  = \input  [57];
  assign shiftLeftOnePos[57] = \input[56] ;
  assign \input[56]  = \input  [56];
  assign shiftLeftOnePos[56] = \input[55] ;
  assign \input[55]  = \input  [55];
  assign shiftLeftOnePos[55] = \input[54] ;
  assign \input[54]  = \input  [54];
  assign shiftLeftOnePos[54] = \input[53] ;
  assign \input[53]  = \input  [53];
  assign shiftLeftOnePos[53] = \input[52] ;
  assign \input[52]  = \input  [52];
  assign shiftLeftOnePos[52] = \input[51] ;
  assign \input[51]  = \input  [51];
  assign shiftLeftOnePos[51] = \input[50] ;
  assign \input[50]  = \input  [50];
  assign shiftLeftOnePos[50] = \input[49] ;
  assign \input[49]  = \input  [49];
  assign shiftLeftOnePos[49] = \input[48] ;
  assign \input[48]  = \input  [48];
  assign shiftLeftOnePos[48] = \input[47] ;
  assign \input[47]  = \input  [47];
  assign shiftLeftOnePos[47] = \input[46] ;
  assign \input[46]  = \input  [46];
  assign shiftLeftOnePos[46] = \input[45] ;
  assign \input[45]  = \input  [45];
  assign shiftLeftOnePos[45] = \input[44] ;
  assign \input[44]  = \input  [44];
  assign shiftLeftOnePos[44] = \input[43] ;
  assign \input[43]  = \input  [43];
  assign shiftLeftOnePos[43] = \input[42] ;
  assign \input[42]  = \input  [42];
  assign shiftLeftOnePos[42] = \input[41] ;
  assign \input[41]  = \input  [41];
  assign shiftLeftOnePos[41] = \input[40] ;
  assign \input[40]  = \input  [40];
  assign shiftLeftOnePos[40] = \input[39] ;
  assign \input[39]  = \input  [39];
  assign shiftLeftOnePos[39] = \input[38] ;
  assign \input[38]  = \input  [38];
  assign shiftLeftOnePos[38] = \input[37] ;
  assign \input[37]  = \input  [37];
  assign shiftLeftOnePos[37] = \input[36] ;
  assign \input[36]  = \input  [36];
  assign shiftLeftOnePos[36] = \input[35] ;
  assign \input[35]  = \input  [35];
  assign shiftLeftOnePos[35] = \input[34] ;
  assign \input[34]  = \input  [34];
  assign shiftLeftOnePos[34] = \input[33] ;
  assign \input[33]  = \input  [33];
  assign shiftLeftOnePos[33] = \input[32] ;
  assign \input[32]  = \input  [32];
  assign shiftLeftOnePos[32] = \input[31] ;
  assign \input[31]  = \input  [31];
  assign shiftLeftOnePos[31] = \input[30] ;
  assign \input[30]  = \input  [30];
  assign shiftLeftOnePos[30] = \input[29] ;
  assign \input[29]  = \input  [29];
  assign shiftLeftOnePos[29] = \input[28] ;
  assign \input[28]  = \input  [28];
  assign shiftLeftOnePos[28] = \input[27] ;
  assign \input[27]  = \input  [27];
  assign shiftLeftOnePos[27] = \input[26] ;
  assign \input[26]  = \input  [26];
  assign shiftLeftOnePos[26] = \input[25] ;
  assign \input[25]  = \input  [25];
  assign shiftLeftOnePos[25] = \input[24] ;
  assign \input[24]  = \input  [24];
  assign shiftLeftOnePos[24] = \input[23] ;
  assign \input[23]  = \input  [23];
  assign shiftLeftOnePos[23] = \input[22] ;
  assign \input[22]  = \input  [22];
  assign shiftLeftOnePos[22] = \input[21] ;
  assign \input[21]  = \input  [21];
  assign shiftLeftOnePos[21] = \input[20] ;
  assign \input[20]  = \input  [20];
  assign shiftLeftOnePos[20] = \input[19] ;
  assign \input[19]  = \input  [19];
  assign shiftLeftOnePos[19] = \input[18] ;
  assign \input[18]  = \input  [18];
  assign shiftLeftOnePos[18] = \input[17] ;
  assign \input[17]  = \input  [17];
  assign shiftLeftOnePos[17] = \input[16] ;
  assign \input[16]  = \input  [16];
  assign shiftLeftOnePos[16] = \input[15] ;
  assign \input[15]  = \input  [15];
  assign shiftLeftOnePos[15] = \input[14] ;
  assign \input[14]  = \input  [14];
  assign shiftLeftOnePos[14] = \input[13] ;
  assign \input[13]  = \input  [13];
  assign shiftLeftOnePos[13] = \input[12] ;
  assign \input[12]  = \input  [12];
  assign shiftLeftOnePos[12] = \input[11] ;
  assign \input[11]  = \input  [11];
  assign shiftLeftOnePos[11] = \input[10] ;
  assign \input[10]  = \input  [10];
  assign shiftLeftOnePos[10] = \input[9] ;
  assign \input[9]  = \input  [9];
  assign shiftLeftOnePos[9] = \input[8] ;
  assign \input[8]  = \input  [8];
  assign shiftLeftOnePos[8] = \input[7] ;
  assign \input[7]  = \input  [7];
  assign shiftLeftOnePos[7] = \input[6] ;
  assign \input[6]  = \input  [6];
  assign shiftLeftOnePos[6] = \input[5] ;
  assign \input[5]  = \input  [5];
  assign shiftLeftOnePos[5] = \input[4] ;
  assign \input[4]  = \input  [4];
  assign shiftLeftOnePos[4] = \input[3] ;
  assign \input[3]  = \input  [3];
  assign shiftLeftOnePos[3] = \input[2] ;
  assign \input[2]  = \input  [2];
  assign shiftLeftOnePos[2] = \input[1] ;
  assign \input[1]  = \input  [1];
  assign shiftLeftOnePos[1] = \input[0] ;
  assign \input[0]  = \input  [0];

endmodule


module complementer_N64_22_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n190, n191, n192, n193, n194, n196, n197, n198, n199, n200,
         n202, n203, n204, n206, n207, n208, n210, n211, n212, n213, n214,
         n216, n217, n218, n220, n221, n222, n224, n225, n226, n228, n229,
         n230, n232, n233, n234, n235, n237, n238, n239, n241, n242, n243,
         n245, n246, n247, n249, n250, n189, n195, n201, n205, n209, n215,
         n219, n223, n227, n231, n236, n240, n244, n248, n251;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U81 ( .A(n190), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U82 ( .A(n192), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U83 ( .A(n193), .B(B[6]), .Z(DIFF[6]) );
  XOR2_X1 U85 ( .A(n196), .B(B[62]), .Z(DIFF[62]) );
  XOR2_X1 U86 ( .A(n194), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U87 ( .A(n198), .B(B[59]), .Z(DIFF[59]) );
  XOR2_X1 U89 ( .A(n200), .B(B[57]), .Z(DIFF[57]) );
  XOR2_X1 U90 ( .A(n202), .B(B[55]), .Z(DIFF[55]) );
  XOR2_X1 U92 ( .A(n204), .B(B[53]), .Z(DIFF[53]) );
  XOR2_X1 U93 ( .A(n206), .B(B[51]), .Z(DIFF[51]) );
  XOR2_X1 U95 ( .A(n208), .B(B[49]), .Z(DIFF[49]) );
  XOR2_X1 U96 ( .A(n212), .B(B[47]), .Z(DIFF[47]) );
  XOR2_X1 U98 ( .A(n214), .B(B[45]), .Z(DIFF[45]) );
  XOR2_X1 U99 ( .A(n216), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U101 ( .A(n218), .B(B[41]), .Z(DIFF[41]) );
  XOR2_X1 U102 ( .A(n211), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U103 ( .A(n220), .B(B[39]), .Z(DIFF[39]) );
  XOR2_X1 U105 ( .A(n222), .B(B[37]), .Z(DIFF[37]) );
  XOR2_X1 U106 ( .A(n224), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U108 ( .A(n226), .B(B[33]), .Z(DIFF[33]) );
  XOR2_X1 U109 ( .A(n228), .B(B[31]), .Z(DIFF[31]) );
  XOR2_X1 U111 ( .A(n230), .B(B[29]), .Z(DIFF[29]) );
  XOR2_X1 U112 ( .A(n233), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U114 ( .A(n235), .B(B[25]), .Z(DIFF[25]) );
  XOR2_X1 U115 ( .A(n237), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U117 ( .A(n239), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U118 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U119 ( .A(n241), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U121 ( .A(n243), .B(B[17]), .Z(DIFF[17]) );
  XOR2_X1 U122 ( .A(n245), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U124 ( .A(n247), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U125 ( .A(n249), .B(B[11]), .Z(DIFF[11]) );
  XOR2_X1 U1 ( .A(n197), .B(n251), .Z(DIFF[61]) );
  NAND2_X1 U2 ( .A1(n197), .A2(n251), .ZN(n196) );
  XNOR2_X1 U3 ( .A(B[44]), .B(n217), .ZN(DIFF[44]) );
  NOR2_X1 U4 ( .A1(B[43]), .A2(n216), .ZN(n217) );
  XNOR2_X1 U5 ( .A(B[48]), .B(n213), .ZN(DIFF[48]) );
  NOR2_X1 U6 ( .A1(B[47]), .A2(n212), .ZN(n213) );
  OR3_X1 U7 ( .A1(B[45]), .A2(B[46]), .A3(n214), .ZN(n212) );
  OR3_X1 U8 ( .A1(B[43]), .A2(B[44]), .A3(n216), .ZN(n214) );
  XNOR2_X1 U9 ( .A(n189), .B(B[46]), .ZN(DIFF[46]) );
  NOR2_X1 U10 ( .A1(n214), .A2(B[45]), .ZN(n189) );
  NOR3_X1 U11 ( .A1(B[59]), .A2(B[60]), .A3(n198), .ZN(n197) );
  XNOR2_X1 U12 ( .A(n195), .B(B[63]), .ZN(DIFF[63]) );
  NOR2_X1 U13 ( .A1(n196), .A2(B[62]), .ZN(n195) );
  XNOR2_X1 U14 ( .A(B[52]), .B(n207), .ZN(DIFF[52]) );
  NOR2_X1 U15 ( .A1(B[51]), .A2(n206), .ZN(n207) );
  XNOR2_X1 U16 ( .A(B[56]), .B(n203), .ZN(DIFF[56]) );
  NOR2_X1 U17 ( .A1(B[55]), .A2(n202), .ZN(n203) );
  XNOR2_X1 U18 ( .A(B[60]), .B(n199), .ZN(DIFF[60]) );
  NOR2_X1 U19 ( .A1(B[59]), .A2(n198), .ZN(n199) );
  OR3_X1 U20 ( .A1(B[57]), .A2(B[58]), .A3(n200), .ZN(n198) );
  OR3_X1 U21 ( .A1(B[53]), .A2(B[54]), .A3(n204), .ZN(n202) );
  OR3_X1 U22 ( .A1(B[49]), .A2(B[50]), .A3(n208), .ZN(n206) );
  OR3_X1 U23 ( .A1(B[47]), .A2(B[48]), .A3(n212), .ZN(n208) );
  OR3_X1 U24 ( .A1(B[55]), .A2(B[56]), .A3(n202), .ZN(n200) );
  OR3_X1 U25 ( .A1(B[51]), .A2(B[52]), .A3(n206), .ZN(n204) );
  XNOR2_X1 U26 ( .A(n201), .B(B[58]), .ZN(DIFF[58]) );
  NOR2_X1 U27 ( .A1(n200), .A2(B[57]), .ZN(n201) );
  XNOR2_X1 U28 ( .A(n205), .B(B[54]), .ZN(DIFF[54]) );
  NOR2_X1 U29 ( .A1(n204), .A2(B[53]), .ZN(n205) );
  XNOR2_X1 U30 ( .A(n209), .B(B[50]), .ZN(DIFF[50]) );
  NOR2_X1 U31 ( .A1(n208), .A2(B[49]), .ZN(n209) );
  OR3_X1 U32 ( .A1(B[41]), .A2(B[42]), .A3(n218), .ZN(n216) );
  XNOR2_X1 U33 ( .A(n215), .B(B[42]), .ZN(DIFF[42]) );
  NOR2_X1 U34 ( .A1(n218), .A2(B[41]), .ZN(n215) );
  XNOR2_X1 U35 ( .A(n219), .B(B[26]), .ZN(DIFF[26]) );
  NOR2_X1 U36 ( .A1(n235), .A2(B[25]), .ZN(n219) );
  XNOR2_X1 U37 ( .A(n223), .B(B[22]), .ZN(DIFF[22]) );
  NOR2_X1 U38 ( .A1(n239), .A2(B[21]), .ZN(n223) );
  XNOR2_X1 U39 ( .A(n227), .B(B[18]), .ZN(DIFF[18]) );
  NOR2_X1 U40 ( .A1(n243), .A2(B[17]), .ZN(n227) );
  XNOR2_X1 U41 ( .A(n231), .B(B[14]), .ZN(DIFF[14]) );
  NOR2_X1 U42 ( .A1(n247), .A2(B[13]), .ZN(n231) );
  XNOR2_X1 U43 ( .A(B[24]), .B(n238), .ZN(DIFF[24]) );
  NOR2_X1 U44 ( .A1(B[23]), .A2(n237), .ZN(n238) );
  XNOR2_X1 U45 ( .A(B[20]), .B(n242), .ZN(DIFF[20]) );
  NOR2_X1 U46 ( .A1(B[19]), .A2(n241), .ZN(n242) );
  XNOR2_X1 U47 ( .A(B[16]), .B(n246), .ZN(DIFF[16]) );
  NOR2_X1 U48 ( .A1(B[15]), .A2(n245), .ZN(n246) );
  OR3_X1 U49 ( .A1(B[13]), .A2(B[14]), .A3(n247), .ZN(n245) );
  OR3_X1 U50 ( .A1(B[17]), .A2(B[18]), .A3(n243), .ZN(n241) );
  OR3_X1 U51 ( .A1(B[21]), .A2(B[22]), .A3(n239), .ZN(n237) );
  OR3_X1 U52 ( .A1(B[25]), .A2(B[26]), .A3(n235), .ZN(n233) );
  OR3_X1 U53 ( .A1(B[29]), .A2(B[30]), .A3(n230), .ZN(n228) );
  OR3_X1 U54 ( .A1(B[15]), .A2(B[16]), .A3(n245), .ZN(n243) );
  OR3_X1 U55 ( .A1(B[19]), .A2(B[20]), .A3(n241), .ZN(n239) );
  OR3_X1 U56 ( .A1(B[23]), .A2(B[24]), .A3(n237), .ZN(n235) );
  OR3_X1 U57 ( .A1(B[27]), .A2(B[28]), .A3(n233), .ZN(n230) );
  OR3_X1 U58 ( .A1(B[31]), .A2(B[32]), .A3(n228), .ZN(n226) );
  XNOR2_X1 U59 ( .A(n236), .B(B[34]), .ZN(DIFF[34]) );
  NOR2_X1 U60 ( .A1(n226), .A2(B[33]), .ZN(n236) );
  XNOR2_X1 U61 ( .A(n240), .B(B[30]), .ZN(DIFF[30]) );
  NOR2_X1 U62 ( .A1(n230), .A2(B[29]), .ZN(n240) );
  XNOR2_X1 U63 ( .A(B[36]), .B(n225), .ZN(DIFF[36]) );
  NOR2_X1 U64 ( .A1(B[35]), .A2(n224), .ZN(n225) );
  XNOR2_X1 U65 ( .A(B[32]), .B(n229), .ZN(DIFF[32]) );
  NOR2_X1 U66 ( .A1(B[31]), .A2(n228), .ZN(n229) );
  XNOR2_X1 U67 ( .A(B[28]), .B(n234), .ZN(DIFF[28]) );
  NOR2_X1 U68 ( .A1(B[27]), .A2(n233), .ZN(n234) );
  XNOR2_X1 U69 ( .A(B[40]), .B(n221), .ZN(DIFF[40]) );
  NOR2_X1 U70 ( .A1(B[39]), .A2(n220), .ZN(n221) );
  OR3_X1 U71 ( .A1(B[33]), .A2(B[34]), .A3(n226), .ZN(n224) );
  OR3_X1 U72 ( .A1(B[37]), .A2(B[38]), .A3(n222), .ZN(n220) );
  OR3_X1 U73 ( .A1(B[35]), .A2(B[36]), .A3(n224), .ZN(n222) );
  OR3_X1 U74 ( .A1(B[39]), .A2(B[40]), .A3(n220), .ZN(n218) );
  XNOR2_X1 U75 ( .A(n244), .B(B[38]), .ZN(DIFF[38]) );
  NOR2_X1 U76 ( .A1(n222), .A2(B[37]), .ZN(n244) );
  XNOR2_X1 U77 ( .A(B[12]), .B(n250), .ZN(DIFF[12]) );
  NOR2_X1 U78 ( .A1(B[11]), .A2(n249), .ZN(n250) );
  OR3_X1 U79 ( .A1(B[11]), .A2(B[12]), .A3(n249), .ZN(n247) );
  XNOR2_X1 U80 ( .A(n248), .B(B[10]), .ZN(DIFF[10]) );
  NOR2_X1 U84 ( .A1(n190), .A2(B[9]), .ZN(n248) );
  OR3_X1 U88 ( .A1(B[10]), .A2(B[9]), .A3(n190), .ZN(n249) );
  NOR2_X1 U91 ( .A1(B[7]), .A2(n192), .ZN(n191) );
  NOR2_X1 U94 ( .A1(B[3]), .A2(n211), .ZN(n210) );
  OR3_X1 U97 ( .A1(B[5]), .A2(B[6]), .A3(n194), .ZN(n192) );
  OR3_X1 U100 ( .A1(B[7]), .A2(B[8]), .A3(n192), .ZN(n190) );
  OR3_X1 U104 ( .A1(B[3]), .A2(B[4]), .A3(n211), .ZN(n194) );
  XNOR2_X1 U107 ( .A(B[8]), .B(n191), .ZN(DIFF[8]) );
  XNOR2_X1 U110 ( .A(B[4]), .B(n210), .ZN(DIFF[4]) );
  XNOR2_X1 U113 ( .A(B[2]), .B(n232), .ZN(DIFF[2]) );
  OR2_X1 U116 ( .A1(n194), .A2(B[5]), .ZN(n193) );
  OR3_X1 U120 ( .A1(B[1]), .A2(B[2]), .A3(\B[0] ), .ZN(n211) );
  NOR2_X1 U123 ( .A1(\B[0] ), .A2(B[1]), .ZN(n232) );
  INV_X1 U126 ( .A(B[61]), .ZN(n251) );
endmodule


module complementer_N64_22 ( \input , complement2 );
  input [63:0] \input ;
  output [63:0] complement2;


  complementer_N64_22_DW01_sub_0 sub_add_31_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(\input ), .CI(1'b0), .DIFF(complement2) );
endmodule


module complementer_N64_21_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n190, n191, n192, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n189, n193;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U81 ( .A(n190), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U82 ( .A(n192), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U84 ( .A(n195), .B(B[63]), .Z(DIFF[63]) );
  XOR2_X1 U85 ( .A(n196), .B(B[62]), .Z(DIFF[62]) );
  XOR2_X1 U86 ( .A(n194), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U87 ( .A(n198), .B(B[59]), .Z(DIFF[59]) );
  XOR2_X1 U88 ( .A(n201), .B(B[58]), .Z(DIFF[58]) );
  XOR2_X1 U89 ( .A(n200), .B(B[57]), .Z(DIFF[57]) );
  XOR2_X1 U90 ( .A(n202), .B(B[55]), .Z(DIFF[55]) );
  XOR2_X1 U91 ( .A(n205), .B(B[54]), .Z(DIFF[54]) );
  XOR2_X1 U92 ( .A(n204), .B(B[53]), .Z(DIFF[53]) );
  XOR2_X1 U93 ( .A(n206), .B(B[51]), .Z(DIFF[51]) );
  XOR2_X1 U94 ( .A(n209), .B(B[50]), .Z(DIFF[50]) );
  XOR2_X1 U95 ( .A(n208), .B(B[49]), .Z(DIFF[49]) );
  XOR2_X1 U96 ( .A(n212), .B(B[47]), .Z(DIFF[47]) );
  XOR2_X1 U97 ( .A(n215), .B(B[46]), .Z(DIFF[46]) );
  XOR2_X1 U98 ( .A(n214), .B(B[45]), .Z(DIFF[45]) );
  XOR2_X1 U99 ( .A(n216), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U100 ( .A(n219), .B(B[42]), .Z(DIFF[42]) );
  XOR2_X1 U101 ( .A(n218), .B(B[41]), .Z(DIFF[41]) );
  XOR2_X1 U102 ( .A(n211), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U103 ( .A(n220), .B(B[39]), .Z(DIFF[39]) );
  XOR2_X1 U104 ( .A(n223), .B(B[38]), .Z(DIFF[38]) );
  XOR2_X1 U105 ( .A(n222), .B(B[37]), .Z(DIFF[37]) );
  XOR2_X1 U106 ( .A(n224), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U107 ( .A(n227), .B(B[34]), .Z(DIFF[34]) );
  XOR2_X1 U108 ( .A(n226), .B(B[33]), .Z(DIFF[33]) );
  XOR2_X1 U109 ( .A(n228), .B(B[31]), .Z(DIFF[31]) );
  XOR2_X1 U110 ( .A(n231), .B(B[30]), .Z(DIFF[30]) );
  XOR2_X1 U111 ( .A(n230), .B(B[29]), .Z(DIFF[29]) );
  XOR2_X1 U112 ( .A(n233), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U113 ( .A(n236), .B(B[26]), .Z(DIFF[26]) );
  XOR2_X1 U114 ( .A(n235), .B(B[25]), .Z(DIFF[25]) );
  XOR2_X1 U115 ( .A(n237), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U116 ( .A(n240), .B(B[22]), .Z(DIFF[22]) );
  XOR2_X1 U117 ( .A(n239), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U118 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U119 ( .A(n241), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U120 ( .A(n244), .B(B[18]), .Z(DIFF[18]) );
  XOR2_X1 U121 ( .A(n243), .B(B[17]), .Z(DIFF[17]) );
  XOR2_X1 U122 ( .A(n245), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U123 ( .A(n248), .B(B[14]), .Z(DIFF[14]) );
  XOR2_X1 U124 ( .A(n247), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U125 ( .A(n249), .B(B[11]), .Z(DIFF[11]) );
  XOR2_X1 U126 ( .A(n251), .B(B[10]), .Z(DIFF[10]) );
  NOR2_X1 U1 ( .A1(B[59]), .A2(n198), .ZN(n199) );
  NAND2_X1 U2 ( .A1(n197), .A2(n193), .ZN(n196) );
  OR3_X1 U3 ( .A1(B[53]), .A2(B[54]), .A3(n204), .ZN(n202) );
  OR2_X1 U4 ( .A1(n204), .A2(B[53]), .ZN(n205) );
  OR2_X1 U5 ( .A1(n208), .A2(B[49]), .ZN(n209) );
  NOR2_X1 U6 ( .A1(B[43]), .A2(n216), .ZN(n217) );
  OR3_X1 U7 ( .A1(B[43]), .A2(B[44]), .A3(n216), .ZN(n214) );
  NOR3_X1 U8 ( .A1(B[59]), .A2(B[60]), .A3(n198), .ZN(n197) );
  NOR2_X1 U9 ( .A1(B[47]), .A2(n212), .ZN(n213) );
  NOR2_X1 U10 ( .A1(B[55]), .A2(n202), .ZN(n203) );
  NOR2_X1 U11 ( .A1(B[51]), .A2(n206), .ZN(n207) );
  OR3_X1 U12 ( .A1(B[45]), .A2(B[46]), .A3(n214), .ZN(n212) );
  OR3_X1 U13 ( .A1(B[57]), .A2(B[58]), .A3(n200), .ZN(n198) );
  OR3_X1 U14 ( .A1(B[49]), .A2(B[50]), .A3(n208), .ZN(n206) );
  OR3_X1 U15 ( .A1(B[47]), .A2(B[48]), .A3(n212), .ZN(n208) );
  OR3_X1 U16 ( .A1(B[55]), .A2(B[56]), .A3(n202), .ZN(n200) );
  OR3_X1 U17 ( .A1(B[51]), .A2(B[52]), .A3(n206), .ZN(n204) );
  OR2_X1 U18 ( .A1(n214), .A2(B[45]), .ZN(n215) );
  OR2_X1 U19 ( .A1(n200), .A2(B[57]), .ZN(n201) );
  OR2_X1 U20 ( .A1(n196), .A2(B[62]), .ZN(n195) );
  OR3_X1 U21 ( .A1(B[41]), .A2(B[42]), .A3(n218), .ZN(n216) );
  XNOR2_X1 U22 ( .A(B[44]), .B(n217), .ZN(DIFF[44]) );
  XNOR2_X1 U23 ( .A(B[48]), .B(n213), .ZN(DIFF[48]) );
  OR2_X1 U24 ( .A1(n218), .A2(B[41]), .ZN(n219) );
  XNOR2_X1 U25 ( .A(B[56]), .B(n203), .ZN(DIFF[56]) );
  XNOR2_X1 U26 ( .A(B[52]), .B(n207), .ZN(DIFF[52]) );
  XNOR2_X1 U27 ( .A(n197), .B(B[61]), .ZN(DIFF[61]) );
  XNOR2_X1 U28 ( .A(B[60]), .B(n199), .ZN(DIFF[60]) );
  XNOR2_X1 U29 ( .A(B[20]), .B(n242), .ZN(DIFF[20]) );
  XNOR2_X1 U30 ( .A(B[12]), .B(n250), .ZN(DIFF[12]) );
  NOR2_X1 U31 ( .A1(B[23]), .A2(n237), .ZN(n238) );
  NOR2_X1 U32 ( .A1(B[19]), .A2(n241), .ZN(n242) );
  NOR2_X1 U33 ( .A1(B[15]), .A2(n245), .ZN(n246) );
  OR3_X1 U34 ( .A1(B[21]), .A2(B[22]), .A3(n239), .ZN(n237) );
  OR3_X1 U35 ( .A1(B[17]), .A2(B[18]), .A3(n243), .ZN(n241) );
  OR3_X1 U36 ( .A1(B[13]), .A2(B[14]), .A3(n247), .ZN(n245) );
  OR3_X1 U37 ( .A1(B[23]), .A2(B[24]), .A3(n237), .ZN(n235) );
  OR3_X1 U38 ( .A1(B[19]), .A2(B[20]), .A3(n241), .ZN(n239) );
  OR3_X1 U39 ( .A1(B[15]), .A2(B[16]), .A3(n245), .ZN(n243) );
  XNOR2_X1 U40 ( .A(B[24]), .B(n238), .ZN(DIFF[24]) );
  XNOR2_X1 U41 ( .A(B[16]), .B(n246), .ZN(DIFF[16]) );
  OR2_X1 U42 ( .A1(n235), .A2(B[25]), .ZN(n236) );
  OR2_X1 U43 ( .A1(n243), .A2(B[17]), .ZN(n244) );
  OR2_X1 U44 ( .A1(n247), .A2(B[13]), .ZN(n248) );
  NOR2_X1 U45 ( .A1(B[39]), .A2(n220), .ZN(n221) );
  NOR2_X1 U46 ( .A1(B[35]), .A2(n224), .ZN(n225) );
  NOR2_X1 U47 ( .A1(B[31]), .A2(n228), .ZN(n229) );
  NOR2_X1 U48 ( .A1(B[27]), .A2(n233), .ZN(n234) );
  OR3_X1 U49 ( .A1(B[37]), .A2(B[38]), .A3(n222), .ZN(n220) );
  OR3_X1 U50 ( .A1(B[33]), .A2(B[34]), .A3(n226), .ZN(n224) );
  OR3_X1 U51 ( .A1(B[29]), .A2(B[30]), .A3(n230), .ZN(n228) );
  OR3_X1 U52 ( .A1(B[25]), .A2(B[26]), .A3(n235), .ZN(n233) );
  OR3_X1 U53 ( .A1(B[39]), .A2(B[40]), .A3(n220), .ZN(n218) );
  OR3_X1 U54 ( .A1(B[35]), .A2(B[36]), .A3(n224), .ZN(n222) );
  OR3_X1 U55 ( .A1(B[31]), .A2(B[32]), .A3(n228), .ZN(n226) );
  OR3_X1 U56 ( .A1(B[27]), .A2(B[28]), .A3(n233), .ZN(n230) );
  XNOR2_X1 U57 ( .A(B[40]), .B(n221), .ZN(DIFF[40]) );
  XNOR2_X1 U58 ( .A(B[36]), .B(n225), .ZN(DIFF[36]) );
  XNOR2_X1 U59 ( .A(B[32]), .B(n229), .ZN(DIFF[32]) );
  XNOR2_X1 U60 ( .A(B[28]), .B(n234), .ZN(DIFF[28]) );
  OR2_X1 U61 ( .A1(n222), .A2(B[37]), .ZN(n223) );
  OR2_X1 U62 ( .A1(n226), .A2(B[33]), .ZN(n227) );
  OR2_X1 U63 ( .A1(n230), .A2(B[29]), .ZN(n231) );
  OR2_X1 U64 ( .A1(n239), .A2(B[21]), .ZN(n240) );
  NOR2_X1 U65 ( .A1(B[11]), .A2(n249), .ZN(n250) );
  OR3_X1 U66 ( .A1(B[11]), .A2(B[12]), .A3(n249), .ZN(n247) );
  XNOR2_X1 U67 ( .A(n189), .B(B[6]), .ZN(DIFF[6]) );
  NOR2_X1 U68 ( .A1(n194), .A2(B[5]), .ZN(n189) );
  XNOR2_X1 U69 ( .A(B[8]), .B(n191), .ZN(DIFF[8]) );
  NOR2_X1 U70 ( .A1(B[7]), .A2(n192), .ZN(n191) );
  XNOR2_X1 U71 ( .A(B[2]), .B(n232), .ZN(DIFF[2]) );
  NOR2_X1 U72 ( .A1(\B[0] ), .A2(B[1]), .ZN(n232) );
  XNOR2_X1 U73 ( .A(B[4]), .B(n210), .ZN(DIFF[4]) );
  NOR2_X1 U74 ( .A1(B[3]), .A2(n211), .ZN(n210) );
  OR3_X1 U75 ( .A1(B[5]), .A2(B[6]), .A3(n194), .ZN(n192) );
  OR3_X1 U76 ( .A1(B[10]), .A2(B[9]), .A3(n190), .ZN(n249) );
  OR3_X1 U77 ( .A1(B[7]), .A2(B[8]), .A3(n192), .ZN(n190) );
  OR3_X1 U78 ( .A1(B[3]), .A2(B[4]), .A3(n211), .ZN(n194) );
  OR2_X1 U79 ( .A1(n190), .A2(B[9]), .ZN(n251) );
  OR3_X1 U80 ( .A1(B[1]), .A2(B[2]), .A3(\B[0] ), .ZN(n211) );
  INV_X1 U83 ( .A(B[61]), .ZN(n193) );
endmodule


module complementer_N64_21 ( \input , complement2 );
  input [63:0] \input ;
  output [63:0] complement2;


  complementer_N64_21_DW01_sub_0 sub_add_31_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(\input ), .CI(1'b0), .DIFF(complement2) );
endmodule


module ShiftnCompl_N64_11 ( plusA, plus2A_out, minus2A_out, plus4A_out, 
        minus4A_out );
  input [63:0] plusA;
  output [63:0] plus2A_out;
  output [63:0] minus2A_out;
  output [63:0] plus4A_out;
  output [63:0] minus4A_out;
  wire   n13, n14, n2, n15, n16, n17, n18, n19, n20, n21, n22;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign plus2A_out[0] = 1'b0;
  assign plus2A_out[51] = n2;
  assign plus4A_out[0] = 1'b0;

  shifter_N64_22 shifter_1 ( .\input (plusA), .shiftLeftOnePos({
        plus2A_out[63:59], n13, plus2A_out[57:54], n14, plus2A_out[52], n2, 
        plus2A_out[50:49], n15, plus2A_out[47:44], n16, plus2A_out[42:1], 
        SYNOPSYS_UNCONNECTED__0}) );
  shifter_N64_21 shifter_2 ( .\input ({plus2A_out[63:52], n2, plus2A_out[50:1], 
        1'b0}), .shiftLeftOnePos({plus4A_out[63:59], n17, plus4A_out[57:54], 
        n18, plus4A_out[52:49], n19, plus4A_out[47:44], n20, n21, n22, 
        plus4A_out[40:1], SYNOPSYS_UNCONNECTED__1}) );
  complementer_N64_22 complementer_1 ( .\input ({plus2A_out[63:52], n2, 
        plus2A_out[50:1], 1'b0}), .complement2(minus2A_out) );
  complementer_N64_21 complementer_2 ( .\input ({plus4A_out[63:1], 1'b0}), 
        .complement2(minus4A_out) );
  BUF_X1 U1 ( .A(n16), .Z(plus2A_out[43]) );
  BUF_X1 U4 ( .A(n20), .Z(plus4A_out[43]) );
  BUF_X1 U5 ( .A(n18), .Z(plus4A_out[53]) );
  BUF_X1 U6 ( .A(n22), .Z(plus4A_out[41]) );
  BUF_X1 U7 ( .A(n15), .Z(plus2A_out[48]) );
  BUF_X1 U8 ( .A(n19), .Z(plus4A_out[48]) );
  BUF_X1 U9 ( .A(n21), .Z(plus4A_out[42]) );
  BUF_X1 U10 ( .A(n14), .Z(plus2A_out[53]) );
  BUF_X1 U11 ( .A(n17), .Z(plus4A_out[58]) );
  BUF_X1 U12 ( .A(n13), .Z(plus2A_out[58]) );
endmodule


module MUX_GENERIC_N64_RADIX3_11 ( plusA, minusA, plus2A, minus2A, SEL, Y );
  input [63:0] plusA;
  input [63:0] minusA;
  input [63:0] plus2A;
  input [63:0] minus2A;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502;
  tri   [63:0] Y;

  TBUF_X1 \Y_tri[55]  ( .A(n446), .EN(n301), .Z(Y[55]) );
  TBUF_X1 \Y_tri[56]  ( .A(n445), .EN(n301), .Z(Y[56]) );
  TBUF_X1 \Y_tri[57]  ( .A(n444), .EN(n301), .Z(Y[57]) );
  TBUF_X1 \Y_tri[58]  ( .A(n443), .EN(n301), .Z(Y[58]) );
  TBUF_X1 \Y_tri[59]  ( .A(n442), .EN(n301), .Z(Y[59]) );
  TBUF_X1 \Y_tri[60]  ( .A(n441), .EN(n301), .Z(Y[60]) );
  TBUF_X1 \Y_tri[61]  ( .A(n440), .EN(n301), .Z(Y[61]) );
  TBUF_X1 \Y_tri[63]  ( .A(n438), .EN(n301), .Z(Y[63]) );
  TBUF_X1 \Y_tri[49]  ( .A(n452), .EN(n300), .Z(Y[49]) );
  TBUF_X1 \Y_tri[50]  ( .A(n451), .EN(n300), .Z(Y[50]) );
  TBUF_X1 \Y_tri[51]  ( .A(n450), .EN(n300), .Z(Y[51]) );
  TBUF_X1 \Y_tri[52]  ( .A(n449), .EN(n300), .Z(Y[52]) );
  TBUF_X1 \Y_tri[53]  ( .A(n448), .EN(n300), .Z(Y[53]) );
  TBUF_X1 \Y_tri[54]  ( .A(n447), .EN(n300), .Z(Y[54]) );
  TBUF_X1 \Y_tri[25]  ( .A(n476), .EN(n298), .Z(Y[25]) );
  TBUF_X1 \Y_tri[27]  ( .A(n474), .EN(n298), .Z(Y[27]) );
  TBUF_X1 \Y_tri[28]  ( .A(n473), .EN(n298), .Z(Y[28]) );
  TBUF_X1 \Y_tri[30]  ( .A(n471), .EN(n298), .Z(Y[30]) );
  TBUF_X1 \Y_tri[31]  ( .A(n470), .EN(n298), .Z(Y[31]) );
  TBUF_X1 \Y_tri[32]  ( .A(n469), .EN(n298), .Z(Y[32]) );
  TBUF_X1 \Y_tri[35]  ( .A(n466), .EN(n299), .Z(Y[35]) );
  TBUF_X1 \Y_tri[36]  ( .A(n465), .EN(n299), .Z(Y[36]) );
  TBUF_X1 \Y_tri[37]  ( .A(n464), .EN(n299), .Z(Y[37]) );
  TBUF_X1 \Y_tri[38]  ( .A(n463), .EN(n299), .Z(Y[38]) );
  TBUF_X1 \Y_tri[39]  ( .A(n462), .EN(n299), .Z(Y[39]) );
  TBUF_X1 \Y_tri[40]  ( .A(n461), .EN(n299), .Z(Y[40]) );
  TBUF_X1 \Y_tri[41]  ( .A(n460), .EN(n299), .Z(Y[41]) );
  TBUF_X1 \Y_tri[42]  ( .A(n459), .EN(n299), .Z(Y[42]) );
  TBUF_X1 \Y_tri[43]  ( .A(n458), .EN(n299), .Z(Y[43]) );
  TBUF_X1 \Y_tri[44]  ( .A(n457), .EN(n300), .Z(Y[44]) );
  TBUF_X1 \Y_tri[45]  ( .A(n456), .EN(n300), .Z(Y[45]) );
  TBUF_X1 \Y_tri[46]  ( .A(n455), .EN(n300), .Z(Y[46]) );
  TBUF_X1 \Y_tri[47]  ( .A(n454), .EN(n300), .Z(Y[47]) );
  TBUF_X1 \Y_tri[48]  ( .A(n453), .EN(n300), .Z(Y[48]) );
  TBUF_X1 \Y_tri[29]  ( .A(n472), .EN(n298), .Z(Y[29]) );
  TBUF_X1 \Y_tri[6]  ( .A(n496), .EN(n296), .Z(Y[6]) );
  TBUF_X1 \Y_tri[7]  ( .A(n495), .EN(n296), .Z(Y[7]) );
  TBUF_X1 \Y_tri[8]  ( .A(n494), .EN(n296), .Z(Y[8]) );
  TBUF_X1 \Y_tri[9]  ( .A(n492), .EN(n296), .Z(Y[9]) );
  TBUF_X1 \Y_tri[10]  ( .A(n491), .EN(n296), .Z(Y[10]) );
  TBUF_X1 \Y_tri[11]  ( .A(n490), .EN(n297), .Z(Y[11]) );
  TBUF_X1 \Y_tri[12]  ( .A(n489), .EN(n297), .Z(Y[12]) );
  TBUF_X1 \Y_tri[13]  ( .A(n488), .EN(n297), .Z(Y[13]) );
  TBUF_X1 \Y_tri[14]  ( .A(n487), .EN(n297), .Z(Y[14]) );
  TBUF_X1 \Y_tri[15]  ( .A(n486), .EN(n297), .Z(Y[15]) );
  TBUF_X1 \Y_tri[17]  ( .A(n484), .EN(n297), .Z(Y[17]) );
  TBUF_X1 \Y_tri[18]  ( .A(n483), .EN(n297), .Z(Y[18]) );
  TBUF_X1 \Y_tri[19]  ( .A(n482), .EN(n297), .Z(Y[19]) );
  TBUF_X1 \Y_tri[20]  ( .A(n481), .EN(n297), .Z(Y[20]) );
  TBUF_X1 \Y_tri[21]  ( .A(n480), .EN(n297), .Z(Y[21]) );
  TBUF_X1 \Y_tri[22]  ( .A(n479), .EN(n298), .Z(Y[22]) );
  TBUF_X1 \Y_tri[23]  ( .A(n478), .EN(n298), .Z(Y[23]) );
  TBUF_X1 \Y_tri[0]  ( .A(n502), .EN(n296), .Z(Y[0]) );
  TBUF_X1 \Y_tri[2]  ( .A(n500), .EN(n296), .Z(Y[2]) );
  TBUF_X1 \Y_tri[3]  ( .A(n499), .EN(n296), .Z(Y[3]) );
  TBUF_X1 \Y_tri[5]  ( .A(n497), .EN(n296), .Z(Y[5]) );
  TBUF_X1 \Y_tri[1]  ( .A(n501), .EN(n296), .Z(Y[1]) );
  TBUF_X1 \Y_tri[4]  ( .A(n498), .EN(n296), .Z(Y[4]) );
  TBUF_X1 \Y_tri[16]  ( .A(n485), .EN(n297), .Z(Y[16]) );
  TBUF_X1 \Y_tri[24]  ( .A(n477), .EN(n298), .Z(Y[24]) );
  TBUF_X1 \Y_tri[26]  ( .A(n475), .EN(n298), .Z(Y[26]) );
  TBUF_X1 \Y_tri[33]  ( .A(n468), .EN(n299), .Z(Y[33]) );
  TBUF_X1 \Y_tri[34]  ( .A(n467), .EN(n299), .Z(Y[34]) );
  TBUF_X1 \Y_tri[62]  ( .A(n439), .EN(n301), .Z(Y[62]) );
  NAND2_X1 U2 ( .A1(n399), .A2(n398), .ZN(n455) );
  AOI22_X1 U3 ( .A1(plusA[46]), .A2(n281), .B1(plus2A[46]), .B2(n275), .ZN(
        n399) );
  AOI22_X1 U4 ( .A1(minus2A[46]), .A2(n293), .B1(minusA[46]), .B2(n287), .ZN(
        n398) );
  NAND2_X1 U5 ( .A1(n395), .A2(n394), .ZN(n457) );
  AOI22_X1 U6 ( .A1(plusA[44]), .A2(n281), .B1(plus2A[44]), .B2(n275), .ZN(
        n395) );
  AOI22_X1 U7 ( .A1(minus2A[44]), .A2(n293), .B1(minusA[44]), .B2(n287), .ZN(
        n394) );
  NAND2_X1 U8 ( .A1(n401), .A2(n400), .ZN(n454) );
  AOI22_X1 U9 ( .A1(plusA[47]), .A2(n281), .B1(plus2A[47]), .B2(n275), .ZN(
        n401) );
  AOI22_X1 U10 ( .A1(minus2A[47]), .A2(n293), .B1(minusA[47]), .B2(n287), .ZN(
        n400) );
  NAND2_X1 U11 ( .A1(n397), .A2(n396), .ZN(n456) );
  AOI22_X1 U12 ( .A1(plusA[45]), .A2(n281), .B1(plus2A[45]), .B2(n275), .ZN(
        n397) );
  AOI22_X1 U13 ( .A1(minus2A[45]), .A2(n293), .B1(minusA[45]), .B2(n287), .ZN(
        n396) );
  NAND2_X1 U14 ( .A1(n393), .A2(n392), .ZN(n458) );
  AOI22_X1 U15 ( .A1(plusA[43]), .A2(n281), .B1(plus2A[43]), .B2(n275), .ZN(
        n393) );
  AOI22_X1 U16 ( .A1(minus2A[43]), .A2(n293), .B1(minusA[43]), .B2(n287), .ZN(
        n392) );
  NAND2_X1 U17 ( .A1(n389), .A2(n388), .ZN(n460) );
  AOI22_X1 U18 ( .A1(plusA[41]), .A2(n281), .B1(plus2A[41]), .B2(n275), .ZN(
        n389) );
  AOI22_X1 U19 ( .A1(minus2A[41]), .A2(n293), .B1(minusA[41]), .B2(n287), .ZN(
        n388) );
  NAND2_X1 U20 ( .A1(n403), .A2(n402), .ZN(n453) );
  AOI22_X1 U21 ( .A1(plusA[48]), .A2(n282), .B1(plus2A[48]), .B2(n276), .ZN(
        n403) );
  AOI22_X1 U22 ( .A1(minus2A[48]), .A2(n294), .B1(minusA[48]), .B2(n288), .ZN(
        n402) );
  NAND2_X1 U23 ( .A1(n391), .A2(n390), .ZN(n459) );
  AOI22_X1 U24 ( .A1(plusA[42]), .A2(n281), .B1(plus2A[42]), .B2(n275), .ZN(
        n391) );
  AOI22_X1 U25 ( .A1(minus2A[42]), .A2(n293), .B1(minusA[42]), .B2(n287), .ZN(
        n390) );
  NAND2_X1 U26 ( .A1(n419), .A2(n418), .ZN(n445) );
  AOI22_X1 U27 ( .A1(plusA[56]), .A2(n282), .B1(plus2A[56]), .B2(n276), .ZN(
        n419) );
  AOI22_X1 U28 ( .A1(minus2A[56]), .A2(n294), .B1(minusA[56]), .B2(n288), .ZN(
        n418) );
  NAND2_X1 U29 ( .A1(n415), .A2(n414), .ZN(n447) );
  AOI22_X1 U30 ( .A1(plusA[54]), .A2(n282), .B1(plus2A[54]), .B2(n276), .ZN(
        n415) );
  AOI22_X1 U31 ( .A1(minus2A[54]), .A2(n294), .B1(minusA[54]), .B2(n288), .ZN(
        n414) );
  NAND2_X1 U32 ( .A1(n421), .A2(n420), .ZN(n444) );
  AOI22_X1 U33 ( .A1(plusA[57]), .A2(n282), .B1(plus2A[57]), .B2(n276), .ZN(
        n421) );
  AOI22_X1 U34 ( .A1(minus2A[57]), .A2(n294), .B1(minusA[57]), .B2(n288), .ZN(
        n420) );
  NAND2_X1 U35 ( .A1(n417), .A2(n416), .ZN(n446) );
  AOI22_X1 U36 ( .A1(plusA[55]), .A2(n282), .B1(plus2A[55]), .B2(n276), .ZN(
        n417) );
  AOI22_X1 U37 ( .A1(minus2A[55]), .A2(n294), .B1(minusA[55]), .B2(n288), .ZN(
        n416) );
  NAND2_X1 U38 ( .A1(n413), .A2(n412), .ZN(n448) );
  AOI22_X1 U39 ( .A1(plusA[53]), .A2(n282), .B1(plus2A[53]), .B2(n276), .ZN(
        n413) );
  AOI22_X1 U40 ( .A1(minus2A[53]), .A2(n294), .B1(minusA[53]), .B2(n288), .ZN(
        n412) );
  NAND2_X1 U41 ( .A1(n409), .A2(n408), .ZN(n450) );
  AOI22_X1 U42 ( .A1(plusA[51]), .A2(n282), .B1(plus2A[51]), .B2(n276), .ZN(
        n409) );
  AOI22_X1 U43 ( .A1(minus2A[51]), .A2(n294), .B1(minusA[51]), .B2(n288), .ZN(
        n408) );
  NAND2_X1 U44 ( .A1(n405), .A2(n404), .ZN(n452) );
  AOI22_X1 U45 ( .A1(plusA[49]), .A2(n282), .B1(plus2A[49]), .B2(n276), .ZN(
        n405) );
  AOI22_X1 U46 ( .A1(minus2A[49]), .A2(n294), .B1(minusA[49]), .B2(n288), .ZN(
        n404) );
  NAND2_X1 U47 ( .A1(n411), .A2(n410), .ZN(n449) );
  AOI22_X1 U48 ( .A1(plusA[52]), .A2(n282), .B1(plus2A[52]), .B2(n276), .ZN(
        n411) );
  AOI22_X1 U49 ( .A1(minus2A[52]), .A2(n294), .B1(minusA[52]), .B2(n288), .ZN(
        n410) );
  NAND2_X1 U50 ( .A1(n407), .A2(n406), .ZN(n451) );
  AOI22_X1 U51 ( .A1(plusA[50]), .A2(n282), .B1(plus2A[50]), .B2(n276), .ZN(
        n407) );
  AOI22_X1 U52 ( .A1(minus2A[50]), .A2(n294), .B1(minusA[50]), .B2(n288), .ZN(
        n406) );
  NAND2_X1 U53 ( .A1(n431), .A2(n430), .ZN(n439) );
  AOI22_X1 U54 ( .A1(plusA[62]), .A2(n283), .B1(plus2A[62]), .B2(n277), .ZN(
        n431) );
  AOI22_X1 U55 ( .A1(minus2A[62]), .A2(n295), .B1(minusA[62]), .B2(n289), .ZN(
        n430) );
  NAND2_X1 U56 ( .A1(n437), .A2(n436), .ZN(n438) );
  AOI22_X1 U57 ( .A1(plusA[63]), .A2(n283), .B1(plus2A[63]), .B2(n277), .ZN(
        n437) );
  AOI22_X1 U58 ( .A1(minus2A[63]), .A2(n295), .B1(minusA[63]), .B2(n289), .ZN(
        n436) );
  NAND2_X1 U59 ( .A1(n429), .A2(n428), .ZN(n440) );
  AOI22_X1 U60 ( .A1(plusA[61]), .A2(n283), .B1(plus2A[61]), .B2(n277), .ZN(
        n429) );
  AOI22_X1 U61 ( .A1(minus2A[61]), .A2(n295), .B1(minusA[61]), .B2(n289), .ZN(
        n428) );
  NAND2_X1 U62 ( .A1(n427), .A2(n426), .ZN(n441) );
  AOI22_X1 U63 ( .A1(plusA[60]), .A2(n283), .B1(plus2A[60]), .B2(n277), .ZN(
        n427) );
  AOI22_X1 U64 ( .A1(minus2A[60]), .A2(n295), .B1(minusA[60]), .B2(n289), .ZN(
        n426) );
  NAND2_X1 U65 ( .A1(n425), .A2(n424), .ZN(n442) );
  AOI22_X1 U66 ( .A1(plusA[59]), .A2(n282), .B1(plus2A[59]), .B2(n276), .ZN(
        n425) );
  AOI22_X1 U67 ( .A1(minus2A[59]), .A2(n294), .B1(minusA[59]), .B2(n288), .ZN(
        n424) );
  NAND2_X1 U68 ( .A1(n423), .A2(n422), .ZN(n443) );
  AOI22_X1 U69 ( .A1(plusA[58]), .A2(n282), .B1(plus2A[58]), .B2(n276), .ZN(
        n423) );
  AOI22_X1 U70 ( .A1(minus2A[58]), .A2(n294), .B1(minusA[58]), .B2(n288), .ZN(
        n422) );
  BUF_X1 U71 ( .A(n493), .Z(n296) );
  BUF_X1 U72 ( .A(n433), .Z(n279) );
  BUF_X1 U73 ( .A(n433), .Z(n278) );
  BUF_X1 U74 ( .A(n435), .Z(n291) );
  BUF_X1 U75 ( .A(n435), .Z(n290) );
  BUF_X1 U76 ( .A(n434), .Z(n285) );
  BUF_X1 U77 ( .A(n432), .Z(n273) );
  BUF_X1 U78 ( .A(n434), .Z(n284) );
  BUF_X1 U79 ( .A(n432), .Z(n272) );
  BUF_X1 U80 ( .A(n493), .Z(n297) );
  NAND2_X1 U81 ( .A1(n373), .A2(n372), .ZN(n468) );
  AOI22_X1 U82 ( .A1(plusA[33]), .A2(n280), .B1(plus2A[33]), .B2(n274), .ZN(
        n373) );
  AOI22_X1 U83 ( .A1(minus2A[33]), .A2(n292), .B1(minusA[33]), .B2(n286), .ZN(
        n372) );
  NAND2_X1 U84 ( .A1(n359), .A2(n358), .ZN(n475) );
  AOI22_X1 U85 ( .A1(plusA[26]), .A2(n280), .B1(plus2A[26]), .B2(n274), .ZN(
        n359) );
  AOI22_X1 U86 ( .A1(minus2A[26]), .A2(n292), .B1(minusA[26]), .B2(n286), .ZN(
        n358) );
  NAND2_X1 U87 ( .A1(n353), .A2(n352), .ZN(n478) );
  AOI22_X1 U88 ( .A1(plusA[23]), .A2(n279), .B1(plus2A[23]), .B2(n273), .ZN(
        n353) );
  AOI22_X1 U89 ( .A1(minus2A[23]), .A2(n291), .B1(minusA[23]), .B2(n285), .ZN(
        n352) );
  NAND2_X1 U90 ( .A1(n351), .A2(n350), .ZN(n479) );
  AOI22_X1 U91 ( .A1(plusA[22]), .A2(n279), .B1(plus2A[22]), .B2(n273), .ZN(
        n351) );
  AOI22_X1 U92 ( .A1(minus2A[22]), .A2(n291), .B1(minusA[22]), .B2(n285), .ZN(
        n350) );
  NAND2_X1 U93 ( .A1(n349), .A2(n348), .ZN(n480) );
  AOI22_X1 U94 ( .A1(plusA[21]), .A2(n279), .B1(plus2A[21]), .B2(n273), .ZN(
        n349) );
  AOI22_X1 U95 ( .A1(minus2A[21]), .A2(n291), .B1(minusA[21]), .B2(n285), .ZN(
        n348) );
  NAND2_X1 U96 ( .A1(n347), .A2(n346), .ZN(n481) );
  AOI22_X1 U97 ( .A1(plusA[20]), .A2(n279), .B1(plus2A[20]), .B2(n273), .ZN(
        n347) );
  AOI22_X1 U98 ( .A1(minus2A[20]), .A2(n291), .B1(minusA[20]), .B2(n285), .ZN(
        n346) );
  NAND2_X1 U99 ( .A1(n345), .A2(n344), .ZN(n482) );
  AOI22_X1 U100 ( .A1(plusA[19]), .A2(n279), .B1(plus2A[19]), .B2(n273), .ZN(
        n345) );
  AOI22_X1 U101 ( .A1(minus2A[19]), .A2(n291), .B1(minusA[19]), .B2(n285), 
        .ZN(n344) );
  NAND2_X1 U102 ( .A1(n343), .A2(n342), .ZN(n483) );
  AOI22_X1 U103 ( .A1(plusA[18]), .A2(n279), .B1(plus2A[18]), .B2(n273), .ZN(
        n343) );
  AOI22_X1 U104 ( .A1(minus2A[18]), .A2(n291), .B1(minusA[18]), .B2(n285), 
        .ZN(n342) );
  NAND2_X1 U105 ( .A1(n341), .A2(n340), .ZN(n484) );
  AOI22_X1 U106 ( .A1(plusA[17]), .A2(n279), .B1(plus2A[17]), .B2(n273), .ZN(
        n341) );
  AOI22_X1 U107 ( .A1(minus2A[17]), .A2(n291), .B1(minusA[17]), .B2(n285), 
        .ZN(n340) );
  NAND2_X1 U108 ( .A1(n337), .A2(n336), .ZN(n486) );
  AOI22_X1 U109 ( .A1(plusA[15]), .A2(n279), .B1(plus2A[15]), .B2(n273), .ZN(
        n337) );
  AOI22_X1 U110 ( .A1(minus2A[15]), .A2(n291), .B1(minusA[15]), .B2(n285), 
        .ZN(n336) );
  NAND2_X1 U111 ( .A1(n335), .A2(n334), .ZN(n487) );
  AOI22_X1 U112 ( .A1(plusA[14]), .A2(n279), .B1(plus2A[14]), .B2(n273), .ZN(
        n335) );
  AOI22_X1 U113 ( .A1(minus2A[14]), .A2(n291), .B1(minusA[14]), .B2(n285), 
        .ZN(n334) );
  NAND2_X1 U114 ( .A1(n333), .A2(n332), .ZN(n488) );
  AOI22_X1 U115 ( .A1(plusA[13]), .A2(n279), .B1(plus2A[13]), .B2(n273), .ZN(
        n333) );
  AOI22_X1 U116 ( .A1(minus2A[13]), .A2(n291), .B1(minusA[13]), .B2(n285), 
        .ZN(n332) );
  NAND2_X1 U117 ( .A1(n331), .A2(n330), .ZN(n489) );
  AOI22_X1 U118 ( .A1(plusA[12]), .A2(n279), .B1(plus2A[12]), .B2(n273), .ZN(
        n331) );
  AOI22_X1 U119 ( .A1(minus2A[12]), .A2(n291), .B1(minusA[12]), .B2(n285), 
        .ZN(n330) );
  NAND2_X1 U120 ( .A1(n355), .A2(n354), .ZN(n477) );
  AOI22_X1 U121 ( .A1(plusA[24]), .A2(n280), .B1(plus2A[24]), .B2(n274), .ZN(
        n355) );
  AOI22_X1 U122 ( .A1(minus2A[24]), .A2(n292), .B1(minusA[24]), .B2(n286), 
        .ZN(n354) );
  NAND2_X1 U123 ( .A1(n339), .A2(n338), .ZN(n485) );
  AOI22_X1 U124 ( .A1(plusA[16]), .A2(n279), .B1(plus2A[16]), .B2(n273), .ZN(
        n339) );
  AOI22_X1 U125 ( .A1(minus2A[16]), .A2(n291), .B1(minusA[16]), .B2(n285), 
        .ZN(n338) );
  BUF_X1 U126 ( .A(n433), .Z(n280) );
  BUF_X1 U127 ( .A(n435), .Z(n292) );
  BUF_X1 U128 ( .A(n434), .Z(n286) );
  BUF_X1 U129 ( .A(n432), .Z(n274) );
  BUF_X1 U130 ( .A(n493), .Z(n298) );
  NAND2_X1 U131 ( .A1(n375), .A2(n374), .ZN(n467) );
  AOI22_X1 U132 ( .A1(plusA[34]), .A2(n280), .B1(plus2A[34]), .B2(n274), .ZN(
        n375) );
  AOI22_X1 U133 ( .A1(minus2A[34]), .A2(n292), .B1(minusA[34]), .B2(n286), 
        .ZN(n374) );
  NAND2_X1 U134 ( .A1(n367), .A2(n366), .ZN(n471) );
  AOI22_X1 U135 ( .A1(plusA[30]), .A2(n280), .B1(plus2A[30]), .B2(n274), .ZN(
        n367) );
  AOI22_X1 U136 ( .A1(minus2A[30]), .A2(n292), .B1(minusA[30]), .B2(n286), 
        .ZN(n366) );
  NAND2_X1 U137 ( .A1(n365), .A2(n364), .ZN(n472) );
  AOI22_X1 U138 ( .A1(plusA[29]), .A2(n280), .B1(plus2A[29]), .B2(n274), .ZN(
        n365) );
  AOI22_X1 U139 ( .A1(minus2A[29]), .A2(n292), .B1(minusA[29]), .B2(n286), 
        .ZN(n364) );
  NAND2_X1 U140 ( .A1(n361), .A2(n360), .ZN(n474) );
  AOI22_X1 U141 ( .A1(plusA[27]), .A2(n280), .B1(plus2A[27]), .B2(n274), .ZN(
        n361) );
  AOI22_X1 U142 ( .A1(minus2A[27]), .A2(n292), .B1(minusA[27]), .B2(n286), 
        .ZN(n360) );
  NAND2_X1 U143 ( .A1(n357), .A2(n356), .ZN(n476) );
  AOI22_X1 U144 ( .A1(plusA[25]), .A2(n280), .B1(plus2A[25]), .B2(n274), .ZN(
        n357) );
  AOI22_X1 U145 ( .A1(minus2A[25]), .A2(n292), .B1(minusA[25]), .B2(n286), 
        .ZN(n356) );
  NAND2_X1 U146 ( .A1(n385), .A2(n384), .ZN(n462) );
  AOI22_X1 U147 ( .A1(plusA[39]), .A2(n281), .B1(plus2A[39]), .B2(n275), .ZN(
        n385) );
  AOI22_X1 U148 ( .A1(minus2A[39]), .A2(n293), .B1(minusA[39]), .B2(n287), 
        .ZN(n384) );
  NAND2_X1 U149 ( .A1(n377), .A2(n376), .ZN(n466) );
  AOI22_X1 U150 ( .A1(plusA[35]), .A2(n280), .B1(plus2A[35]), .B2(n274), .ZN(
        n377) );
  AOI22_X1 U151 ( .A1(minus2A[35]), .A2(n292), .B1(minusA[35]), .B2(n286), 
        .ZN(n376) );
  NAND2_X1 U152 ( .A1(n369), .A2(n368), .ZN(n470) );
  AOI22_X1 U153 ( .A1(plusA[31]), .A2(n280), .B1(plus2A[31]), .B2(n274), .ZN(
        n369) );
  AOI22_X1 U154 ( .A1(minus2A[31]), .A2(n292), .B1(minusA[31]), .B2(n286), 
        .ZN(n368) );
  NAND2_X1 U155 ( .A1(n381), .A2(n380), .ZN(n464) );
  AOI22_X1 U156 ( .A1(plusA[37]), .A2(n281), .B1(plus2A[37]), .B2(n275), .ZN(
        n381) );
  AOI22_X1 U157 ( .A1(minus2A[37]), .A2(n293), .B1(minusA[37]), .B2(n287), 
        .ZN(n380) );
  NAND2_X1 U158 ( .A1(n387), .A2(n386), .ZN(n461) );
  AOI22_X1 U159 ( .A1(plusA[40]), .A2(n281), .B1(plus2A[40]), .B2(n275), .ZN(
        n387) );
  AOI22_X1 U160 ( .A1(minus2A[40]), .A2(n293), .B1(minusA[40]), .B2(n287), 
        .ZN(n386) );
  NAND2_X1 U161 ( .A1(n379), .A2(n378), .ZN(n465) );
  AOI22_X1 U162 ( .A1(plusA[36]), .A2(n281), .B1(plus2A[36]), .B2(n275), .ZN(
        n379) );
  AOI22_X1 U163 ( .A1(minus2A[36]), .A2(n293), .B1(minusA[36]), .B2(n287), 
        .ZN(n378) );
  NAND2_X1 U164 ( .A1(n371), .A2(n370), .ZN(n469) );
  AOI22_X1 U165 ( .A1(plusA[32]), .A2(n280), .B1(plus2A[32]), .B2(n274), .ZN(
        n371) );
  AOI22_X1 U166 ( .A1(minus2A[32]), .A2(n292), .B1(minusA[32]), .B2(n286), 
        .ZN(n370) );
  NAND2_X1 U167 ( .A1(n363), .A2(n362), .ZN(n473) );
  AOI22_X1 U168 ( .A1(plusA[28]), .A2(n280), .B1(plus2A[28]), .B2(n274), .ZN(
        n363) );
  AOI22_X1 U169 ( .A1(minus2A[28]), .A2(n292), .B1(minusA[28]), .B2(n286), 
        .ZN(n362) );
  NAND2_X1 U170 ( .A1(n383), .A2(n382), .ZN(n463) );
  AOI22_X1 U171 ( .A1(plusA[38]), .A2(n281), .B1(plus2A[38]), .B2(n275), .ZN(
        n383) );
  AOI22_X1 U172 ( .A1(minus2A[38]), .A2(n293), .B1(minusA[38]), .B2(n287), 
        .ZN(n382) );
  BUF_X1 U173 ( .A(n433), .Z(n281) );
  BUF_X1 U174 ( .A(n435), .Z(n293) );
  BUF_X1 U175 ( .A(n434), .Z(n287) );
  BUF_X1 U176 ( .A(n432), .Z(n275) );
  BUF_X1 U177 ( .A(n493), .Z(n299) );
  BUF_X1 U178 ( .A(n493), .Z(n300) );
  BUF_X1 U179 ( .A(n433), .Z(n282) );
  BUF_X1 U180 ( .A(n435), .Z(n294) );
  BUF_X1 U181 ( .A(n434), .Z(n288) );
  BUF_X1 U182 ( .A(n432), .Z(n276) );
  BUF_X1 U183 ( .A(n493), .Z(n301) );
  NOR2_X1 U184 ( .A1(n323), .A2(n304), .ZN(n493) );
  INV_X1 U185 ( .A(SEL[2]), .ZN(n304) );
  NOR2_X1 U186 ( .A1(SEL[1]), .A2(SEL[0]), .ZN(n323) );
  NOR3_X1 U187 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n302), .ZN(n434) );
  NOR3_X1 U188 ( .A1(SEL[1]), .A2(SEL[2]), .A3(n303), .ZN(n433) );
  NOR3_X1 U189 ( .A1(n302), .A2(SEL[2]), .A3(n303), .ZN(n432) );
  NAND2_X1 U190 ( .A1(n329), .A2(n328), .ZN(n490) );
  AOI22_X1 U191 ( .A1(plusA[11]), .A2(n278), .B1(plus2A[11]), .B2(n272), .ZN(
        n329) );
  AOI22_X1 U192 ( .A1(minus2A[11]), .A2(n290), .B1(minusA[11]), .B2(n284), 
        .ZN(n328) );
  AND2_X1 U193 ( .A1(SEL[2]), .A2(n323), .ZN(n435) );
  INV_X1 U194 ( .A(SEL[1]), .ZN(n302) );
  INV_X1 U195 ( .A(SEL[0]), .ZN(n303) );
  NAND2_X1 U196 ( .A1(n327), .A2(n326), .ZN(n491) );
  AOI22_X1 U197 ( .A1(plusA[10]), .A2(n278), .B1(plus2A[10]), .B2(n272), .ZN(
        n327) );
  AOI22_X1 U198 ( .A1(minus2A[10]), .A2(n290), .B1(minusA[10]), .B2(n284), 
        .ZN(n326) );
  NAND2_X1 U199 ( .A1(n325), .A2(n324), .ZN(n492) );
  AOI22_X1 U200 ( .A1(plusA[9]), .A2(n278), .B1(plus2A[9]), .B2(n272), .ZN(
        n325) );
  AOI22_X1 U201 ( .A1(minus2A[9]), .A2(n290), .B1(minusA[9]), .B2(n284), .ZN(
        n324) );
  NAND2_X1 U202 ( .A1(n320), .A2(n319), .ZN(n495) );
  AOI22_X1 U203 ( .A1(plusA[7]), .A2(n278), .B1(plus2A[7]), .B2(n272), .ZN(
        n320) );
  AOI22_X1 U204 ( .A1(minus2A[7]), .A2(n290), .B1(minusA[7]), .B2(n284), .ZN(
        n319) );
  NAND2_X1 U205 ( .A1(n318), .A2(n317), .ZN(n496) );
  AOI22_X1 U206 ( .A1(plusA[6]), .A2(n278), .B1(plus2A[6]), .B2(n272), .ZN(
        n318) );
  AOI22_X1 U207 ( .A1(minus2A[6]), .A2(n290), .B1(minusA[6]), .B2(n284), .ZN(
        n317) );
  NAND2_X1 U208 ( .A1(n316), .A2(n315), .ZN(n497) );
  AOI22_X1 U209 ( .A1(plusA[5]), .A2(n278), .B1(plus2A[5]), .B2(n272), .ZN(
        n316) );
  AOI22_X1 U210 ( .A1(minus2A[5]), .A2(n290), .B1(minusA[5]), .B2(n284), .ZN(
        n315) );
  NAND2_X1 U211 ( .A1(n312), .A2(n311), .ZN(n499) );
  AOI22_X1 U212 ( .A1(plusA[3]), .A2(n278), .B1(plus2A[3]), .B2(n272), .ZN(
        n312) );
  AOI22_X1 U213 ( .A1(minus2A[3]), .A2(n290), .B1(minusA[3]), .B2(n284), .ZN(
        n311) );
  NAND2_X1 U214 ( .A1(n322), .A2(n321), .ZN(n494) );
  AOI22_X1 U215 ( .A1(plusA[8]), .A2(n278), .B1(plus2A[8]), .B2(n272), .ZN(
        n322) );
  AOI22_X1 U216 ( .A1(minus2A[8]), .A2(n290), .B1(minusA[8]), .B2(n284), .ZN(
        n321) );
  NAND2_X1 U217 ( .A1(n314), .A2(n313), .ZN(n498) );
  AOI22_X1 U218 ( .A1(plusA[4]), .A2(n278), .B1(plus2A[4]), .B2(n272), .ZN(
        n314) );
  AOI22_X1 U219 ( .A1(minus2A[4]), .A2(n290), .B1(minusA[4]), .B2(n284), .ZN(
        n313) );
  NAND2_X1 U220 ( .A1(n310), .A2(n309), .ZN(n500) );
  AOI22_X1 U221 ( .A1(plusA[2]), .A2(n278), .B1(plus2A[2]), .B2(n272), .ZN(
        n310) );
  AOI22_X1 U222 ( .A1(minus2A[2]), .A2(n290), .B1(minusA[2]), .B2(n284), .ZN(
        n309) );
  NAND2_X1 U223 ( .A1(n308), .A2(n307), .ZN(n501) );
  AOI22_X1 U224 ( .A1(plusA[1]), .A2(n278), .B1(plus2A[1]), .B2(n272), .ZN(
        n308) );
  AOI22_X1 U225 ( .A1(minus2A[1]), .A2(n290), .B1(minusA[1]), .B2(n284), .ZN(
        n307) );
  NAND2_X1 U226 ( .A1(n306), .A2(n305), .ZN(n502) );
  AOI22_X1 U227 ( .A1(plusA[0]), .A2(n278), .B1(plus2A[0]), .B2(n272), .ZN(
        n306) );
  AOI22_X1 U228 ( .A1(minus2A[0]), .A2(n290), .B1(minusA[0]), .B2(n284), .ZN(
        n305) );
  CLKBUF_X1 U229 ( .A(n432), .Z(n277) );
  CLKBUF_X1 U230 ( .A(n433), .Z(n283) );
  CLKBUF_X1 U231 ( .A(n434), .Z(n289) );
  CLKBUF_X1 U232 ( .A(n435), .Z(n295) );
endmodule


module FA_704 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_703 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_702 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_701 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_700 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  XNOR2_X1 U4 ( .A(n4), .B(B), .ZN(n6) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_699 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_698 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_697 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_696 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_695 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_694 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_693 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_692 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_691 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_690 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_689 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_688 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  AOI22_X1 U4 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
  INV_X1 U5 ( .A(n7), .ZN(Co) );
endmodule


module FA_687 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_686 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_685 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_684 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_683 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_682 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_681 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_680 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  AOI22_X1 U4 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
  INV_X1 U5 ( .A(n7), .ZN(Co) );
endmodule


module FA_679 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_678 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  AOI22_X1 U4 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
  INV_X1 U5 ( .A(n7), .ZN(Co) );
endmodule


module FA_677 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_676 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_675 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_674 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_673 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_672 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_671 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_670 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  AOI22_X1 U4 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
  INV_X1 U5 ( .A(n7), .ZN(Co) );
endmodule


module FA_669 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_668 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_667 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_666 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_665 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_664 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_663 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_662 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_661 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_660 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_659 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_658 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_657 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_656 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_655 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_654 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_653 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_652 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_651 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_650 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_649 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_648 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_647 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_646 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_645 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_644 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_643 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_642 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  XNOR2_X1 U4 ( .A(n4), .B(B), .ZN(n6) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_641 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N64_11 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Ci;
  output Co;

  wire   [63:1] CTMP;
  tri   [63:0] A;

  FA_704 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_703 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_702 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_701 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(CTMP[4]) );
  FA_700 FAI_5 ( .A(A[4]), .B(B[4]), .Ci(CTMP[4]), .S(S[4]), .Co(CTMP[5]) );
  FA_699 FAI_6 ( .A(A[5]), .B(B[5]), .Ci(CTMP[5]), .S(S[5]), .Co(CTMP[6]) );
  FA_698 FAI_7 ( .A(A[6]), .B(B[6]), .Ci(CTMP[6]), .S(S[6]), .Co(CTMP[7]) );
  FA_697 FAI_8 ( .A(A[7]), .B(B[7]), .Ci(CTMP[7]), .S(S[7]), .Co(CTMP[8]) );
  FA_696 FAI_9 ( .A(A[8]), .B(B[8]), .Ci(CTMP[8]), .S(S[8]), .Co(CTMP[9]) );
  FA_695 FAI_10 ( .A(A[9]), .B(B[9]), .Ci(CTMP[9]), .S(S[9]), .Co(CTMP[10]) );
  FA_694 FAI_11 ( .A(A[10]), .B(B[10]), .Ci(CTMP[10]), .S(S[10]), .Co(CTMP[11]) );
  FA_693 FAI_12 ( .A(A[11]), .B(B[11]), .Ci(CTMP[11]), .S(S[11]), .Co(CTMP[12]) );
  FA_692 FAI_13 ( .A(A[12]), .B(B[12]), .Ci(CTMP[12]), .S(S[12]), .Co(CTMP[13]) );
  FA_691 FAI_14 ( .A(A[13]), .B(B[13]), .Ci(CTMP[13]), .S(S[13]), .Co(CTMP[14]) );
  FA_690 FAI_15 ( .A(A[14]), .B(B[14]), .Ci(CTMP[14]), .S(S[14]), .Co(CTMP[15]) );
  FA_689 FAI_16 ( .A(A[15]), .B(B[15]), .Ci(CTMP[15]), .S(S[15]), .Co(CTMP[16]) );
  FA_688 FAI_17 ( .A(A[16]), .B(B[16]), .Ci(CTMP[16]), .S(S[16]), .Co(CTMP[17]) );
  FA_687 FAI_18 ( .A(A[17]), .B(B[17]), .Ci(CTMP[17]), .S(S[17]), .Co(CTMP[18]) );
  FA_686 FAI_19 ( .A(A[18]), .B(B[18]), .Ci(CTMP[18]), .S(S[18]), .Co(CTMP[19]) );
  FA_685 FAI_20 ( .A(A[19]), .B(B[19]), .Ci(CTMP[19]), .S(S[19]), .Co(CTMP[20]) );
  FA_684 FAI_21 ( .A(A[20]), .B(B[20]), .Ci(CTMP[20]), .S(S[20]), .Co(CTMP[21]) );
  FA_683 FAI_22 ( .A(A[21]), .B(B[21]), .Ci(CTMP[21]), .S(S[21]), .Co(CTMP[22]) );
  FA_682 FAI_23 ( .A(A[22]), .B(B[22]), .Ci(CTMP[22]), .S(S[22]), .Co(CTMP[23]) );
  FA_681 FAI_24 ( .A(A[23]), .B(B[23]), .Ci(CTMP[23]), .S(S[23]), .Co(CTMP[24]) );
  FA_680 FAI_25 ( .A(A[24]), .B(B[24]), .Ci(CTMP[24]), .S(S[24]), .Co(CTMP[25]) );
  FA_679 FAI_26 ( .A(A[25]), .B(B[25]), .Ci(CTMP[25]), .S(S[25]), .Co(CTMP[26]) );
  FA_678 FAI_27 ( .A(A[26]), .B(B[26]), .Ci(CTMP[26]), .S(S[26]), .Co(CTMP[27]) );
  FA_677 FAI_28 ( .A(A[27]), .B(B[27]), .Ci(CTMP[27]), .S(S[27]), .Co(CTMP[28]) );
  FA_676 FAI_29 ( .A(A[28]), .B(B[28]), .Ci(CTMP[28]), .S(S[28]), .Co(CTMP[29]) );
  FA_675 FAI_30 ( .A(A[29]), .B(B[29]), .Ci(CTMP[29]), .S(S[29]), .Co(CTMP[30]) );
  FA_674 FAI_31 ( .A(A[30]), .B(B[30]), .Ci(CTMP[30]), .S(S[30]), .Co(CTMP[31]) );
  FA_673 FAI_32 ( .A(A[31]), .B(B[31]), .Ci(CTMP[31]), .S(S[31]), .Co(CTMP[32]) );
  FA_672 FAI_33 ( .A(A[32]), .B(B[32]), .Ci(CTMP[32]), .S(S[32]), .Co(CTMP[33]) );
  FA_671 FAI_34 ( .A(A[33]), .B(B[33]), .Ci(CTMP[33]), .S(S[33]), .Co(CTMP[34]) );
  FA_670 FAI_35 ( .A(A[34]), .B(B[34]), .Ci(CTMP[34]), .S(S[34]), .Co(CTMP[35]) );
  FA_669 FAI_36 ( .A(A[35]), .B(B[35]), .Ci(CTMP[35]), .S(S[35]), .Co(CTMP[36]) );
  FA_668 FAI_37 ( .A(A[36]), .B(B[36]), .Ci(CTMP[36]), .S(S[36]), .Co(CTMP[37]) );
  FA_667 FAI_38 ( .A(A[37]), .B(B[37]), .Ci(CTMP[37]), .S(S[37]), .Co(CTMP[38]) );
  FA_666 FAI_39 ( .A(A[38]), .B(B[38]), .Ci(CTMP[38]), .S(S[38]), .Co(CTMP[39]) );
  FA_665 FAI_40 ( .A(A[39]), .B(B[39]), .Ci(CTMP[39]), .S(S[39]), .Co(CTMP[40]) );
  FA_664 FAI_41 ( .A(A[40]), .B(B[40]), .Ci(CTMP[40]), .S(S[40]), .Co(CTMP[41]) );
  FA_663 FAI_42 ( .A(A[41]), .B(B[41]), .Ci(CTMP[41]), .S(S[41]), .Co(CTMP[42]) );
  FA_662 FAI_43 ( .A(A[42]), .B(B[42]), .Ci(CTMP[42]), .S(S[42]), .Co(CTMP[43]) );
  FA_661 FAI_44 ( .A(A[43]), .B(B[43]), .Ci(CTMP[43]), .S(S[43]), .Co(CTMP[44]) );
  FA_660 FAI_45 ( .A(A[44]), .B(B[44]), .Ci(CTMP[44]), .S(S[44]), .Co(CTMP[45]) );
  FA_659 FAI_46 ( .A(A[45]), .B(B[45]), .Ci(CTMP[45]), .S(S[45]), .Co(CTMP[46]) );
  FA_658 FAI_47 ( .A(A[46]), .B(B[46]), .Ci(CTMP[46]), .S(S[46]), .Co(CTMP[47]) );
  FA_657 FAI_48 ( .A(A[47]), .B(B[47]), .Ci(CTMP[47]), .S(S[47]), .Co(CTMP[48]) );
  FA_656 FAI_49 ( .A(A[48]), .B(B[48]), .Ci(CTMP[48]), .S(S[48]), .Co(CTMP[49]) );
  FA_655 FAI_50 ( .A(A[49]), .B(B[49]), .Ci(CTMP[49]), .S(S[49]), .Co(CTMP[50]) );
  FA_654 FAI_51 ( .A(A[50]), .B(B[50]), .Ci(CTMP[50]), .S(S[50]), .Co(CTMP[51]) );
  FA_653 FAI_52 ( .A(A[51]), .B(B[51]), .Ci(CTMP[51]), .S(S[51]), .Co(CTMP[52]) );
  FA_652 FAI_53 ( .A(A[52]), .B(B[52]), .Ci(CTMP[52]), .S(S[52]), .Co(CTMP[53]) );
  FA_651 FAI_54 ( .A(A[53]), .B(B[53]), .Ci(CTMP[53]), .S(S[53]), .Co(CTMP[54]) );
  FA_650 FAI_55 ( .A(A[54]), .B(B[54]), .Ci(CTMP[54]), .S(S[54]), .Co(CTMP[55]) );
  FA_649 FAI_56 ( .A(A[55]), .B(B[55]), .Ci(CTMP[55]), .S(S[55]), .Co(CTMP[56]) );
  FA_648 FAI_57 ( .A(A[56]), .B(B[56]), .Ci(CTMP[56]), .S(S[56]), .Co(CTMP[57]) );
  FA_647 FAI_58 ( .A(A[57]), .B(B[57]), .Ci(CTMP[57]), .S(S[57]), .Co(CTMP[58]) );
  FA_646 FAI_59 ( .A(A[58]), .B(B[58]), .Ci(CTMP[58]), .S(S[58]), .Co(CTMP[59]) );
  FA_645 FAI_60 ( .A(A[59]), .B(B[59]), .Ci(CTMP[59]), .S(S[59]), .Co(CTMP[60]) );
  FA_644 FAI_61 ( .A(A[60]), .B(B[60]), .Ci(CTMP[60]), .S(S[60]), .Co(CTMP[61]) );
  FA_643 FAI_62 ( .A(A[61]), .B(B[61]), .Ci(CTMP[61]), .S(S[61]), .Co(CTMP[62]) );
  FA_642 FAI_63 ( .A(A[62]), .B(B[62]), .Ci(CTMP[62]), .S(S[62]), .Co(CTMP[63]) );
  FA_641 FAI_64 ( .A(A[63]), .B(B[63]), .Ci(CTMP[63]), .S(S[63]), .Co(Co) );
endmodule


module booth_mul_row_N64_RADIX3_11 ( prevA, prevSum, encoderIn, nextA, nextSum
 );
  input [63:0] prevA;
  input [63:0] prevSum;
  input [2:0] encoderIn;
  output [63:0] nextA;
  output [63:0] nextSum;
  wire   n3;
  wire   [2:0] encoder_to_mux;
  wire   [63:0] plus2A_s;
  wire   [63:0] minus2A_s;
  wire   [63:0] minus4A_s;
  tri   [63:0] mux_to_adder;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign nextA[51] = n3;
  assign nextA[0] = 1'b0;

  encoder_N64_RADIX3_11 encoder_1 ( .X(encoderIn), .Z(encoder_to_mux) );
  ShiftnCompl_N64_11 ShiftnCompl_1 ( .plusA(prevA), .plus2A_out({
        plus2A_s[63:1], SYNOPSYS_UNCONNECTED__0}), .minus2A_out(minus2A_s), 
        .plus4A_out({nextA[63:52], n3, nextA[50:1], SYNOPSYS_UNCONNECTED__1}), 
        .minus4A_out(minus4A_s) );
  MUX_GENERIC_N64_RADIX3_11 mux_1 ( .plusA({plus2A_s[63:1], 1'b0}), .minusA(
        minus2A_s), .plus2A({nextA[63:52], n3, nextA[50:1], 1'b0}), .minus2A(
        minus4A_s), .SEL(encoder_to_mux), .Y(mux_to_adder) );
  RCA_N64_11 rca_1 ( .A(mux_to_adder), .B(prevSum), .Ci(1'b0), .S(nextSum) );
endmodule


module encoder_N64_RADIX3_10 ( X, Z );
  input [2:0] X;
  output [2:0] Z;
  wire   n5, n7, n8;

  OAI22_X1 U1 ( .A1(n8), .A2(n5), .B1(X[2]), .B2(n7), .ZN(Z[1]) );
  INV_X1 U2 ( .A(X[2]), .ZN(n5) );
  AOI21_X1 U3 ( .B1(n8), .B2(n7), .A(X[2]), .ZN(Z[0]) );
  OAI21_X1 U4 ( .B1(X[1]), .B2(X[0]), .A(n7), .ZN(n8) );
  AND3_X1 U5 ( .A1(X[2]), .A2(n7), .A3(n8), .ZN(Z[2]) );
  NAND2_X1 U6 ( .A1(X[1]), .A2(X[0]), .ZN(n7) );
endmodule


module shifter_N64_20 ( \input , shiftLeftOnePos );
  input [63:0] \input ;
  output [63:0] shiftLeftOnePos;
  wire   \input[62] , \input[61] , \input[60] , \input[59] , \input[58] ,
         \input[57] , \input[56] , \input[55] , \input[54] , \input[53] ,
         \input[52] , \input[51] , \input[50] , \input[49] , \input[48] ,
         \input[47] , \input[46] , \input[45] , \input[44] , \input[43] ,
         \input[42] , \input[41] , \input[40] , \input[39] , \input[38] ,
         \input[37] , \input[36] , \input[35] , \input[34] , \input[33] ,
         \input[32] , \input[31] , \input[30] , \input[29] , \input[28] ,
         \input[27] , \input[26] , \input[25] , \input[24] , \input[23] ,
         \input[22] , \input[21] , \input[20] , \input[19] , \input[18] ,
         \input[17] , \input[16] , \input[15] , \input[14] , \input[13] ,
         \input[12] , \input[11] , \input[10] , \input[9] , \input[8] ,
         \input[7] , \input[6] , \input[5] , \input[4] , \input[3] ,
         \input[2] , \input[1] , \input[0] ;
  assign shiftLeftOnePos[0] = 1'b0;
  assign shiftLeftOnePos[63] = \input[62] ;
  assign \input[62]  = \input  [62];
  assign shiftLeftOnePos[62] = \input[61] ;
  assign \input[61]  = \input  [61];
  assign shiftLeftOnePos[61] = \input[60] ;
  assign \input[60]  = \input  [60];
  assign shiftLeftOnePos[60] = \input[59] ;
  assign \input[59]  = \input  [59];
  assign shiftLeftOnePos[59] = \input[58] ;
  assign \input[58]  = \input  [58];
  assign shiftLeftOnePos[58] = \input[57] ;
  assign \input[57]  = \input  [57];
  assign shiftLeftOnePos[57] = \input[56] ;
  assign \input[56]  = \input  [56];
  assign shiftLeftOnePos[56] = \input[55] ;
  assign \input[55]  = \input  [55];
  assign shiftLeftOnePos[55] = \input[54] ;
  assign \input[54]  = \input  [54];
  assign shiftLeftOnePos[54] = \input[53] ;
  assign \input[53]  = \input  [53];
  assign shiftLeftOnePos[53] = \input[52] ;
  assign \input[52]  = \input  [52];
  assign shiftLeftOnePos[52] = \input[51] ;
  assign \input[51]  = \input  [51];
  assign shiftLeftOnePos[51] = \input[50] ;
  assign \input[50]  = \input  [50];
  assign shiftLeftOnePos[50] = \input[49] ;
  assign \input[49]  = \input  [49];
  assign shiftLeftOnePos[49] = \input[48] ;
  assign \input[48]  = \input  [48];
  assign shiftLeftOnePos[48] = \input[47] ;
  assign \input[47]  = \input  [47];
  assign shiftLeftOnePos[47] = \input[46] ;
  assign \input[46]  = \input  [46];
  assign shiftLeftOnePos[46] = \input[45] ;
  assign \input[45]  = \input  [45];
  assign shiftLeftOnePos[45] = \input[44] ;
  assign \input[44]  = \input  [44];
  assign shiftLeftOnePos[44] = \input[43] ;
  assign \input[43]  = \input  [43];
  assign shiftLeftOnePos[43] = \input[42] ;
  assign \input[42]  = \input  [42];
  assign shiftLeftOnePos[42] = \input[41] ;
  assign \input[41]  = \input  [41];
  assign shiftLeftOnePos[41] = \input[40] ;
  assign \input[40]  = \input  [40];
  assign shiftLeftOnePos[40] = \input[39] ;
  assign \input[39]  = \input  [39];
  assign shiftLeftOnePos[39] = \input[38] ;
  assign \input[38]  = \input  [38];
  assign shiftLeftOnePos[38] = \input[37] ;
  assign \input[37]  = \input  [37];
  assign shiftLeftOnePos[37] = \input[36] ;
  assign \input[36]  = \input  [36];
  assign shiftLeftOnePos[36] = \input[35] ;
  assign \input[35]  = \input  [35];
  assign shiftLeftOnePos[35] = \input[34] ;
  assign \input[34]  = \input  [34];
  assign shiftLeftOnePos[34] = \input[33] ;
  assign \input[33]  = \input  [33];
  assign shiftLeftOnePos[33] = \input[32] ;
  assign \input[32]  = \input  [32];
  assign shiftLeftOnePos[32] = \input[31] ;
  assign \input[31]  = \input  [31];
  assign shiftLeftOnePos[31] = \input[30] ;
  assign \input[30]  = \input  [30];
  assign shiftLeftOnePos[30] = \input[29] ;
  assign \input[29]  = \input  [29];
  assign shiftLeftOnePos[29] = \input[28] ;
  assign \input[28]  = \input  [28];
  assign shiftLeftOnePos[28] = \input[27] ;
  assign \input[27]  = \input  [27];
  assign shiftLeftOnePos[27] = \input[26] ;
  assign \input[26]  = \input  [26];
  assign shiftLeftOnePos[26] = \input[25] ;
  assign \input[25]  = \input  [25];
  assign shiftLeftOnePos[25] = \input[24] ;
  assign \input[24]  = \input  [24];
  assign shiftLeftOnePos[24] = \input[23] ;
  assign \input[23]  = \input  [23];
  assign shiftLeftOnePos[23] = \input[22] ;
  assign \input[22]  = \input  [22];
  assign shiftLeftOnePos[22] = \input[21] ;
  assign \input[21]  = \input  [21];
  assign shiftLeftOnePos[21] = \input[20] ;
  assign \input[20]  = \input  [20];
  assign shiftLeftOnePos[20] = \input[19] ;
  assign \input[19]  = \input  [19];
  assign shiftLeftOnePos[19] = \input[18] ;
  assign \input[18]  = \input  [18];
  assign shiftLeftOnePos[18] = \input[17] ;
  assign \input[17]  = \input  [17];
  assign shiftLeftOnePos[17] = \input[16] ;
  assign \input[16]  = \input  [16];
  assign shiftLeftOnePos[16] = \input[15] ;
  assign \input[15]  = \input  [15];
  assign shiftLeftOnePos[15] = \input[14] ;
  assign \input[14]  = \input  [14];
  assign shiftLeftOnePos[14] = \input[13] ;
  assign \input[13]  = \input  [13];
  assign shiftLeftOnePos[13] = \input[12] ;
  assign \input[12]  = \input  [12];
  assign shiftLeftOnePos[12] = \input[11] ;
  assign \input[11]  = \input  [11];
  assign shiftLeftOnePos[11] = \input[10] ;
  assign \input[10]  = \input  [10];
  assign shiftLeftOnePos[10] = \input[9] ;
  assign \input[9]  = \input  [9];
  assign shiftLeftOnePos[9] = \input[8] ;
  assign \input[8]  = \input  [8];
  assign shiftLeftOnePos[8] = \input[7] ;
  assign \input[7]  = \input  [7];
  assign shiftLeftOnePos[7] = \input[6] ;
  assign \input[6]  = \input  [6];
  assign shiftLeftOnePos[6] = \input[5] ;
  assign \input[5]  = \input  [5];
  assign shiftLeftOnePos[5] = \input[4] ;
  assign \input[4]  = \input  [4];
  assign shiftLeftOnePos[4] = \input[3] ;
  assign \input[3]  = \input  [3];
  assign shiftLeftOnePos[3] = \input[2] ;
  assign \input[2]  = \input  [2];
  assign shiftLeftOnePos[2] = \input[1] ;
  assign \input[1]  = \input  [1];
  assign shiftLeftOnePos[1] = \input[0] ;
  assign \input[0]  = \input  [0];

endmodule


module shifter_N64_19 ( \input , shiftLeftOnePos );
  input [63:0] \input ;
  output [63:0] shiftLeftOnePos;
  wire   \input[62] , \input[61] , \input[60] , \input[59] , \input[58] ,
         \input[57] , \input[56] , \input[55] , \input[54] , \input[53] ,
         \input[52] , \input[51] , \input[50] , \input[49] , \input[48] ,
         \input[47] , \input[46] , \input[45] , \input[44] , \input[43] ,
         \input[42] , \input[41] , \input[40] , \input[39] , \input[38] ,
         \input[37] , \input[36] , \input[35] , \input[34] , \input[33] ,
         \input[32] , \input[31] , \input[30] , \input[29] , \input[28] ,
         \input[27] , \input[26] , \input[25] , \input[24] , \input[23] ,
         \input[22] , \input[21] , \input[20] , \input[19] , \input[18] ,
         \input[17] , \input[16] , \input[15] , \input[14] , \input[13] ,
         \input[12] , \input[11] , \input[10] , \input[9] , \input[8] ,
         \input[7] , \input[6] , \input[5] , \input[4] , \input[3] ,
         \input[2] , \input[1] , \input[0] ;
  assign shiftLeftOnePos[0] = 1'b0;
  assign shiftLeftOnePos[63] = \input[62] ;
  assign \input[62]  = \input  [62];
  assign shiftLeftOnePos[62] = \input[61] ;
  assign \input[61]  = \input  [61];
  assign shiftLeftOnePos[61] = \input[60] ;
  assign \input[60]  = \input  [60];
  assign shiftLeftOnePos[60] = \input[59] ;
  assign \input[59]  = \input  [59];
  assign shiftLeftOnePos[59] = \input[58] ;
  assign \input[58]  = \input  [58];
  assign shiftLeftOnePos[58] = \input[57] ;
  assign \input[57]  = \input  [57];
  assign shiftLeftOnePos[57] = \input[56] ;
  assign \input[56]  = \input  [56];
  assign shiftLeftOnePos[56] = \input[55] ;
  assign \input[55]  = \input  [55];
  assign shiftLeftOnePos[55] = \input[54] ;
  assign \input[54]  = \input  [54];
  assign shiftLeftOnePos[54] = \input[53] ;
  assign \input[53]  = \input  [53];
  assign shiftLeftOnePos[53] = \input[52] ;
  assign \input[52]  = \input  [52];
  assign shiftLeftOnePos[52] = \input[51] ;
  assign \input[51]  = \input  [51];
  assign shiftLeftOnePos[51] = \input[50] ;
  assign \input[50]  = \input  [50];
  assign shiftLeftOnePos[50] = \input[49] ;
  assign \input[49]  = \input  [49];
  assign shiftLeftOnePos[49] = \input[48] ;
  assign \input[48]  = \input  [48];
  assign shiftLeftOnePos[48] = \input[47] ;
  assign \input[47]  = \input  [47];
  assign shiftLeftOnePos[47] = \input[46] ;
  assign \input[46]  = \input  [46];
  assign shiftLeftOnePos[46] = \input[45] ;
  assign \input[45]  = \input  [45];
  assign shiftLeftOnePos[45] = \input[44] ;
  assign \input[44]  = \input  [44];
  assign shiftLeftOnePos[44] = \input[43] ;
  assign \input[43]  = \input  [43];
  assign shiftLeftOnePos[43] = \input[42] ;
  assign \input[42]  = \input  [42];
  assign shiftLeftOnePos[42] = \input[41] ;
  assign \input[41]  = \input  [41];
  assign shiftLeftOnePos[41] = \input[40] ;
  assign \input[40]  = \input  [40];
  assign shiftLeftOnePos[40] = \input[39] ;
  assign \input[39]  = \input  [39];
  assign shiftLeftOnePos[39] = \input[38] ;
  assign \input[38]  = \input  [38];
  assign shiftLeftOnePos[38] = \input[37] ;
  assign \input[37]  = \input  [37];
  assign shiftLeftOnePos[37] = \input[36] ;
  assign \input[36]  = \input  [36];
  assign shiftLeftOnePos[36] = \input[35] ;
  assign \input[35]  = \input  [35];
  assign shiftLeftOnePos[35] = \input[34] ;
  assign \input[34]  = \input  [34];
  assign shiftLeftOnePos[34] = \input[33] ;
  assign \input[33]  = \input  [33];
  assign shiftLeftOnePos[33] = \input[32] ;
  assign \input[32]  = \input  [32];
  assign shiftLeftOnePos[32] = \input[31] ;
  assign \input[31]  = \input  [31];
  assign shiftLeftOnePos[31] = \input[30] ;
  assign \input[30]  = \input  [30];
  assign shiftLeftOnePos[30] = \input[29] ;
  assign \input[29]  = \input  [29];
  assign shiftLeftOnePos[29] = \input[28] ;
  assign \input[28]  = \input  [28];
  assign shiftLeftOnePos[28] = \input[27] ;
  assign \input[27]  = \input  [27];
  assign shiftLeftOnePos[27] = \input[26] ;
  assign \input[26]  = \input  [26];
  assign shiftLeftOnePos[26] = \input[25] ;
  assign \input[25]  = \input  [25];
  assign shiftLeftOnePos[25] = \input[24] ;
  assign \input[24]  = \input  [24];
  assign shiftLeftOnePos[24] = \input[23] ;
  assign \input[23]  = \input  [23];
  assign shiftLeftOnePos[23] = \input[22] ;
  assign \input[22]  = \input  [22];
  assign shiftLeftOnePos[22] = \input[21] ;
  assign \input[21]  = \input  [21];
  assign shiftLeftOnePos[21] = \input[20] ;
  assign \input[20]  = \input  [20];
  assign shiftLeftOnePos[20] = \input[19] ;
  assign \input[19]  = \input  [19];
  assign shiftLeftOnePos[19] = \input[18] ;
  assign \input[18]  = \input  [18];
  assign shiftLeftOnePos[18] = \input[17] ;
  assign \input[17]  = \input  [17];
  assign shiftLeftOnePos[17] = \input[16] ;
  assign \input[16]  = \input  [16];
  assign shiftLeftOnePos[16] = \input[15] ;
  assign \input[15]  = \input  [15];
  assign shiftLeftOnePos[15] = \input[14] ;
  assign \input[14]  = \input  [14];
  assign shiftLeftOnePos[14] = \input[13] ;
  assign \input[13]  = \input  [13];
  assign shiftLeftOnePos[13] = \input[12] ;
  assign \input[12]  = \input  [12];
  assign shiftLeftOnePos[12] = \input[11] ;
  assign \input[11]  = \input  [11];
  assign shiftLeftOnePos[11] = \input[10] ;
  assign \input[10]  = \input  [10];
  assign shiftLeftOnePos[10] = \input[9] ;
  assign \input[9]  = \input  [9];
  assign shiftLeftOnePos[9] = \input[8] ;
  assign \input[8]  = \input  [8];
  assign shiftLeftOnePos[8] = \input[7] ;
  assign \input[7]  = \input  [7];
  assign shiftLeftOnePos[7] = \input[6] ;
  assign \input[6]  = \input  [6];
  assign shiftLeftOnePos[6] = \input[5] ;
  assign \input[5]  = \input  [5];
  assign shiftLeftOnePos[5] = \input[4] ;
  assign \input[4]  = \input  [4];
  assign shiftLeftOnePos[4] = \input[3] ;
  assign \input[3]  = \input  [3];
  assign shiftLeftOnePos[3] = \input[2] ;
  assign \input[2]  = \input  [2];
  assign shiftLeftOnePos[2] = \input[1] ;
  assign \input[1]  = \input  [1];
  assign shiftLeftOnePos[1] = \input[0] ;
  assign \input[0]  = \input  [0];

endmodule


module complementer_N64_20_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n190, n191, n192, n193, n194, n196, n197, n198, n199, n200,
         n202, n203, n204, n206, n207, n208, n210, n211, n212, n213, n214,
         n216, n217, n218, n220, n221, n222, n224, n225, n226, n228, n229,
         n230, n232, n233, n234, n235, n237, n238, n239, n241, n242, n243,
         n245, n246, n247, n249, n250, n251, n189, n195, n201, n205, n209,
         n215, n219, n223, n227, n231, n236, n240, n244, n248;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U81 ( .A(n190), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U82 ( .A(n192), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U83 ( .A(n193), .B(B[6]), .Z(DIFF[6]) );
  XOR2_X1 U85 ( .A(n196), .B(B[62]), .Z(DIFF[62]) );
  XOR2_X1 U86 ( .A(n194), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U87 ( .A(n198), .B(B[59]), .Z(DIFF[59]) );
  XOR2_X1 U89 ( .A(n200), .B(B[57]), .Z(DIFF[57]) );
  XOR2_X1 U90 ( .A(n202), .B(B[55]), .Z(DIFF[55]) );
  XOR2_X1 U92 ( .A(n204), .B(B[53]), .Z(DIFF[53]) );
  XOR2_X1 U93 ( .A(n206), .B(B[51]), .Z(DIFF[51]) );
  XOR2_X1 U95 ( .A(n208), .B(B[49]), .Z(DIFF[49]) );
  XOR2_X1 U96 ( .A(n212), .B(B[47]), .Z(DIFF[47]) );
  XOR2_X1 U98 ( .A(n214), .B(B[45]), .Z(DIFF[45]) );
  XOR2_X1 U99 ( .A(n216), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U101 ( .A(n218), .B(B[41]), .Z(DIFF[41]) );
  XOR2_X1 U102 ( .A(n211), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U103 ( .A(n220), .B(B[39]), .Z(DIFF[39]) );
  XOR2_X1 U105 ( .A(n222), .B(B[37]), .Z(DIFF[37]) );
  XOR2_X1 U106 ( .A(n224), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U108 ( .A(n226), .B(B[33]), .Z(DIFF[33]) );
  XOR2_X1 U109 ( .A(n228), .B(B[31]), .Z(DIFF[31]) );
  XOR2_X1 U111 ( .A(n230), .B(B[29]), .Z(DIFF[29]) );
  XOR2_X1 U112 ( .A(n233), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U114 ( .A(n235), .B(B[25]), .Z(DIFF[25]) );
  XOR2_X1 U115 ( .A(n237), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U117 ( .A(n239), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U118 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U119 ( .A(n241), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U121 ( .A(n243), .B(B[17]), .Z(DIFF[17]) );
  XOR2_X1 U122 ( .A(n245), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U124 ( .A(n247), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U125 ( .A(n249), .B(B[11]), .Z(DIFF[11]) );
  XOR2_X1 U126 ( .A(n251), .B(B[10]), .Z(DIFF[10]) );
  NOR3_X1 U1 ( .A1(B[59]), .A2(B[60]), .A3(n198), .ZN(n197) );
  XNOR2_X1 U2 ( .A(B[60]), .B(n199), .ZN(DIFF[60]) );
  NOR2_X1 U3 ( .A1(B[59]), .A2(n198), .ZN(n199) );
  XOR2_X1 U4 ( .A(n197), .B(n248), .Z(DIFF[61]) );
  NAND2_X1 U5 ( .A1(n197), .A2(n248), .ZN(n196) );
  OR3_X1 U6 ( .A1(B[53]), .A2(B[54]), .A3(n204), .ZN(n202) );
  OR3_X1 U7 ( .A1(B[49]), .A2(B[50]), .A3(n208), .ZN(n206) );
  XNOR2_X1 U8 ( .A(n189), .B(B[54]), .ZN(DIFF[54]) );
  NOR2_X1 U9 ( .A1(n204), .A2(B[53]), .ZN(n189) );
  XNOR2_X1 U10 ( .A(n195), .B(B[50]), .ZN(DIFF[50]) );
  NOR2_X1 U11 ( .A1(n208), .A2(B[49]), .ZN(n195) );
  XNOR2_X1 U12 ( .A(B[44]), .B(n217), .ZN(DIFF[44]) );
  NOR2_X1 U13 ( .A1(B[43]), .A2(n216), .ZN(n217) );
  OR3_X1 U14 ( .A1(B[43]), .A2(B[44]), .A3(n216), .ZN(n214) );
  XNOR2_X1 U15 ( .A(B[56]), .B(n203), .ZN(DIFF[56]) );
  NOR2_X1 U16 ( .A1(B[55]), .A2(n202), .ZN(n203) );
  XNOR2_X1 U17 ( .A(B[52]), .B(n207), .ZN(DIFF[52]) );
  NOR2_X1 U18 ( .A1(B[51]), .A2(n206), .ZN(n207) );
  XNOR2_X1 U19 ( .A(B[48]), .B(n213), .ZN(DIFF[48]) );
  NOR2_X1 U20 ( .A1(B[47]), .A2(n212), .ZN(n213) );
  OR3_X1 U21 ( .A1(B[45]), .A2(B[46]), .A3(n214), .ZN(n212) );
  OR3_X1 U22 ( .A1(B[57]), .A2(B[58]), .A3(n200), .ZN(n198) );
  OR3_X1 U23 ( .A1(B[47]), .A2(B[48]), .A3(n212), .ZN(n208) );
  OR3_X1 U24 ( .A1(B[55]), .A2(B[56]), .A3(n202), .ZN(n200) );
  OR3_X1 U25 ( .A1(B[51]), .A2(B[52]), .A3(n206), .ZN(n204) );
  XNOR2_X1 U26 ( .A(n201), .B(B[46]), .ZN(DIFF[46]) );
  NOR2_X1 U27 ( .A1(n214), .A2(B[45]), .ZN(n201) );
  XNOR2_X1 U28 ( .A(n205), .B(B[58]), .ZN(DIFF[58]) );
  NOR2_X1 U29 ( .A1(n200), .A2(B[57]), .ZN(n205) );
  XNOR2_X1 U30 ( .A(n209), .B(B[63]), .ZN(DIFF[63]) );
  NOR2_X1 U31 ( .A1(n196), .A2(B[62]), .ZN(n209) );
  XNOR2_X1 U32 ( .A(n215), .B(B[26]), .ZN(DIFF[26]) );
  NOR2_X1 U33 ( .A1(n235), .A2(B[25]), .ZN(n215) );
  XNOR2_X1 U34 ( .A(n219), .B(B[18]), .ZN(DIFF[18]) );
  NOR2_X1 U35 ( .A1(n243), .A2(B[17]), .ZN(n219) );
  XNOR2_X1 U36 ( .A(B[20]), .B(n242), .ZN(DIFF[20]) );
  NOR2_X1 U37 ( .A1(B[19]), .A2(n241), .ZN(n242) );
  XNOR2_X1 U38 ( .A(B[24]), .B(n238), .ZN(DIFF[24]) );
  NOR2_X1 U39 ( .A1(B[23]), .A2(n237), .ZN(n238) );
  OR3_X1 U40 ( .A1(B[17]), .A2(B[18]), .A3(n243), .ZN(n241) );
  OR3_X1 U41 ( .A1(B[21]), .A2(B[22]), .A3(n239), .ZN(n237) );
  OR3_X1 U42 ( .A1(B[25]), .A2(B[26]), .A3(n235), .ZN(n233) );
  OR3_X1 U43 ( .A1(B[19]), .A2(B[20]), .A3(n241), .ZN(n239) );
  OR3_X1 U44 ( .A1(B[23]), .A2(B[24]), .A3(n237), .ZN(n235) );
  XNOR2_X1 U45 ( .A(n223), .B(B[22]), .ZN(DIFF[22]) );
  NOR2_X1 U46 ( .A1(n239), .A2(B[21]), .ZN(n223) );
  XNOR2_X1 U47 ( .A(B[28]), .B(n234), .ZN(DIFF[28]) );
  NOR2_X1 U48 ( .A1(B[27]), .A2(n233), .ZN(n234) );
  XNOR2_X1 U49 ( .A(B[40]), .B(n221), .ZN(DIFF[40]) );
  NOR2_X1 U50 ( .A1(B[39]), .A2(n220), .ZN(n221) );
  XNOR2_X1 U51 ( .A(B[36]), .B(n225), .ZN(DIFF[36]) );
  NOR2_X1 U52 ( .A1(B[35]), .A2(n224), .ZN(n225) );
  XNOR2_X1 U53 ( .A(B[32]), .B(n229), .ZN(DIFF[32]) );
  NOR2_X1 U54 ( .A1(B[31]), .A2(n228), .ZN(n229) );
  OR3_X1 U55 ( .A1(B[29]), .A2(B[30]), .A3(n230), .ZN(n228) );
  OR3_X1 U56 ( .A1(B[33]), .A2(B[34]), .A3(n226), .ZN(n224) );
  OR3_X1 U57 ( .A1(B[37]), .A2(B[38]), .A3(n222), .ZN(n220) );
  OR3_X1 U58 ( .A1(B[41]), .A2(B[42]), .A3(n218), .ZN(n216) );
  OR3_X1 U59 ( .A1(B[27]), .A2(B[28]), .A3(n233), .ZN(n230) );
  OR3_X1 U60 ( .A1(B[31]), .A2(B[32]), .A3(n228), .ZN(n226) );
  OR3_X1 U61 ( .A1(B[35]), .A2(B[36]), .A3(n224), .ZN(n222) );
  OR3_X1 U62 ( .A1(B[39]), .A2(B[40]), .A3(n220), .ZN(n218) );
  XNOR2_X1 U63 ( .A(n227), .B(B[42]), .ZN(DIFF[42]) );
  NOR2_X1 U64 ( .A1(n218), .A2(B[41]), .ZN(n227) );
  XNOR2_X1 U65 ( .A(n231), .B(B[38]), .ZN(DIFF[38]) );
  NOR2_X1 U66 ( .A1(n222), .A2(B[37]), .ZN(n231) );
  XNOR2_X1 U67 ( .A(n236), .B(B[34]), .ZN(DIFF[34]) );
  NOR2_X1 U68 ( .A1(n226), .A2(B[33]), .ZN(n236) );
  XNOR2_X1 U69 ( .A(n240), .B(B[30]), .ZN(DIFF[30]) );
  NOR2_X1 U70 ( .A1(n230), .A2(B[29]), .ZN(n240) );
  XNOR2_X1 U71 ( .A(B[16]), .B(n246), .ZN(DIFF[16]) );
  NOR2_X1 U72 ( .A1(B[15]), .A2(n245), .ZN(n246) );
  OR3_X1 U73 ( .A1(B[15]), .A2(B[16]), .A3(n245), .ZN(n243) );
  XNOR2_X1 U74 ( .A(n244), .B(B[14]), .ZN(DIFF[14]) );
  NOR2_X1 U75 ( .A1(n247), .A2(B[13]), .ZN(n244) );
  OR3_X1 U76 ( .A1(B[13]), .A2(B[14]), .A3(n247), .ZN(n245) );
  OR3_X1 U77 ( .A1(B[11]), .A2(B[12]), .A3(n249), .ZN(n247) );
  XNOR2_X1 U78 ( .A(B[12]), .B(n250), .ZN(DIFF[12]) );
  NOR2_X1 U79 ( .A1(B[11]), .A2(n249), .ZN(n250) );
  NOR2_X1 U80 ( .A1(B[7]), .A2(n192), .ZN(n191) );
  NOR2_X1 U84 ( .A1(B[3]), .A2(n211), .ZN(n210) );
  OR3_X1 U88 ( .A1(B[10]), .A2(B[9]), .A3(n190), .ZN(n249) );
  OR3_X1 U91 ( .A1(B[5]), .A2(B[6]), .A3(n194), .ZN(n192) );
  OR3_X1 U94 ( .A1(B[7]), .A2(B[8]), .A3(n192), .ZN(n190) );
  OR3_X1 U97 ( .A1(B[3]), .A2(B[4]), .A3(n211), .ZN(n194) );
  XNOR2_X1 U100 ( .A(B[8]), .B(n191), .ZN(DIFF[8]) );
  XNOR2_X1 U104 ( .A(B[4]), .B(n210), .ZN(DIFF[4]) );
  XNOR2_X1 U107 ( .A(B[2]), .B(n232), .ZN(DIFF[2]) );
  OR2_X1 U110 ( .A1(n190), .A2(B[9]), .ZN(n251) );
  OR2_X1 U113 ( .A1(n194), .A2(B[5]), .ZN(n193) );
  OR3_X1 U116 ( .A1(B[1]), .A2(B[2]), .A3(\B[0] ), .ZN(n211) );
  NOR2_X1 U120 ( .A1(\B[0] ), .A2(B[1]), .ZN(n232) );
  INV_X1 U123 ( .A(B[61]), .ZN(n248) );
endmodule


module complementer_N64_20 ( \input , complement2 );
  input [63:0] \input ;
  output [63:0] complement2;


  complementer_N64_20_DW01_sub_0 sub_add_31_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(\input ), .CI(1'b0), .DIFF(complement2) );
endmodule


module complementer_N64_19_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n190, n191, n192, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n189, n193, n251;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U81 ( .A(n190), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U82 ( .A(n192), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U84 ( .A(n195), .B(B[63]), .Z(DIFF[63]) );
  XOR2_X1 U85 ( .A(n196), .B(B[62]), .Z(DIFF[62]) );
  XOR2_X1 U86 ( .A(n194), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U87 ( .A(n198), .B(B[59]), .Z(DIFF[59]) );
  XOR2_X1 U88 ( .A(n201), .B(B[58]), .Z(DIFF[58]) );
  XOR2_X1 U89 ( .A(n200), .B(B[57]), .Z(DIFF[57]) );
  XOR2_X1 U90 ( .A(n202), .B(B[55]), .Z(DIFF[55]) );
  XOR2_X1 U91 ( .A(n205), .B(B[54]), .Z(DIFF[54]) );
  XOR2_X1 U92 ( .A(n204), .B(B[53]), .Z(DIFF[53]) );
  XOR2_X1 U93 ( .A(n206), .B(B[51]), .Z(DIFF[51]) );
  XOR2_X1 U94 ( .A(n209), .B(B[50]), .Z(DIFF[50]) );
  XOR2_X1 U95 ( .A(n208), .B(B[49]), .Z(DIFF[49]) );
  XOR2_X1 U96 ( .A(n212), .B(B[47]), .Z(DIFF[47]) );
  XOR2_X1 U97 ( .A(n215), .B(B[46]), .Z(DIFF[46]) );
  XOR2_X1 U98 ( .A(n214), .B(B[45]), .Z(DIFF[45]) );
  XOR2_X1 U99 ( .A(n216), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U100 ( .A(n219), .B(B[42]), .Z(DIFF[42]) );
  XOR2_X1 U101 ( .A(n218), .B(B[41]), .Z(DIFF[41]) );
  XOR2_X1 U102 ( .A(n211), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U103 ( .A(n220), .B(B[39]), .Z(DIFF[39]) );
  XOR2_X1 U104 ( .A(n223), .B(B[38]), .Z(DIFF[38]) );
  XOR2_X1 U105 ( .A(n222), .B(B[37]), .Z(DIFF[37]) );
  XOR2_X1 U106 ( .A(n224), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U107 ( .A(n227), .B(B[34]), .Z(DIFF[34]) );
  XOR2_X1 U108 ( .A(n226), .B(B[33]), .Z(DIFF[33]) );
  XOR2_X1 U109 ( .A(n228), .B(B[31]), .Z(DIFF[31]) );
  XOR2_X1 U110 ( .A(n231), .B(B[30]), .Z(DIFF[30]) );
  XOR2_X1 U111 ( .A(n230), .B(B[29]), .Z(DIFF[29]) );
  XOR2_X1 U112 ( .A(n233), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U113 ( .A(n236), .B(B[26]), .Z(DIFF[26]) );
  XOR2_X1 U114 ( .A(n235), .B(B[25]), .Z(DIFF[25]) );
  XOR2_X1 U115 ( .A(n237), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U116 ( .A(n240), .B(B[22]), .Z(DIFF[22]) );
  XOR2_X1 U117 ( .A(n239), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U118 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U119 ( .A(n241), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U120 ( .A(n244), .B(B[18]), .Z(DIFF[18]) );
  XOR2_X1 U121 ( .A(n243), .B(B[17]), .Z(DIFF[17]) );
  XOR2_X1 U122 ( .A(n245), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U123 ( .A(n248), .B(B[14]), .Z(DIFF[14]) );
  XOR2_X1 U124 ( .A(n247), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U125 ( .A(n249), .B(B[11]), .Z(DIFF[11]) );
  NAND2_X1 U1 ( .A1(n197), .A2(n251), .ZN(n196) );
  NOR3_X1 U2 ( .A1(B[59]), .A2(B[60]), .A3(n198), .ZN(n197) );
  NOR2_X1 U3 ( .A1(B[55]), .A2(n202), .ZN(n203) );
  NOR2_X1 U4 ( .A1(B[51]), .A2(n206), .ZN(n207) );
  NOR2_X1 U5 ( .A1(B[59]), .A2(n198), .ZN(n199) );
  OR3_X1 U6 ( .A1(B[53]), .A2(B[54]), .A3(n204), .ZN(n202) );
  OR3_X1 U7 ( .A1(B[49]), .A2(B[50]), .A3(n208), .ZN(n206) );
  OR3_X1 U8 ( .A1(B[55]), .A2(B[56]), .A3(n202), .ZN(n200) );
  OR2_X1 U9 ( .A1(n204), .A2(B[53]), .ZN(n205) );
  OR2_X1 U10 ( .A1(n208), .A2(B[49]), .ZN(n209) );
  NOR2_X1 U11 ( .A1(B[47]), .A2(n212), .ZN(n213) );
  OR3_X1 U12 ( .A1(B[45]), .A2(B[46]), .A3(n214), .ZN(n212) );
  OR3_X1 U13 ( .A1(B[57]), .A2(B[58]), .A3(n200), .ZN(n198) );
  OR3_X1 U14 ( .A1(B[47]), .A2(B[48]), .A3(n212), .ZN(n208) );
  OR3_X1 U15 ( .A1(B[51]), .A2(B[52]), .A3(n206), .ZN(n204) );
  OR2_X1 U16 ( .A1(n214), .A2(B[45]), .ZN(n215) );
  OR2_X1 U17 ( .A1(n200), .A2(B[57]), .ZN(n201) );
  OR2_X1 U18 ( .A1(n196), .A2(B[62]), .ZN(n195) );
  XNOR2_X1 U19 ( .A(B[20]), .B(n242), .ZN(DIFF[20]) );
  XNOR2_X1 U20 ( .A(B[16]), .B(n246), .ZN(DIFF[16]) );
  NOR2_X1 U21 ( .A1(B[23]), .A2(n237), .ZN(n238) );
  OR3_X1 U22 ( .A1(B[25]), .A2(B[26]), .A3(n235), .ZN(n233) );
  OR3_X1 U23 ( .A1(B[21]), .A2(B[22]), .A3(n239), .ZN(n237) );
  OR3_X1 U24 ( .A1(B[17]), .A2(B[18]), .A3(n243), .ZN(n241) );
  OR3_X1 U25 ( .A1(B[23]), .A2(B[24]), .A3(n237), .ZN(n235) );
  OR3_X1 U26 ( .A1(B[19]), .A2(B[20]), .A3(n241), .ZN(n239) );
  XNOR2_X1 U27 ( .A(B[24]), .B(n238), .ZN(DIFF[24]) );
  OR2_X1 U28 ( .A1(n235), .A2(B[25]), .ZN(n236) );
  XNOR2_X1 U29 ( .A(B[28]), .B(n234), .ZN(DIFF[28]) );
  NOR2_X1 U30 ( .A1(B[39]), .A2(n220), .ZN(n221) );
  NOR2_X1 U31 ( .A1(B[35]), .A2(n224), .ZN(n225) );
  NOR2_X1 U32 ( .A1(B[31]), .A2(n228), .ZN(n229) );
  NOR2_X1 U33 ( .A1(B[27]), .A2(n233), .ZN(n234) );
  NOR2_X1 U34 ( .A1(B[19]), .A2(n241), .ZN(n242) );
  OR3_X1 U35 ( .A1(B[41]), .A2(B[42]), .A3(n218), .ZN(n216) );
  OR3_X1 U36 ( .A1(B[37]), .A2(B[38]), .A3(n222), .ZN(n220) );
  OR3_X1 U37 ( .A1(B[33]), .A2(B[34]), .A3(n226), .ZN(n224) );
  OR3_X1 U38 ( .A1(B[29]), .A2(B[30]), .A3(n230), .ZN(n228) );
  OR3_X1 U39 ( .A1(B[39]), .A2(B[40]), .A3(n220), .ZN(n218) );
  OR3_X1 U40 ( .A1(B[35]), .A2(B[36]), .A3(n224), .ZN(n222) );
  OR3_X1 U41 ( .A1(B[31]), .A2(B[32]), .A3(n228), .ZN(n226) );
  OR3_X1 U42 ( .A1(B[27]), .A2(B[28]), .A3(n233), .ZN(n230) );
  OR3_X1 U43 ( .A1(B[43]), .A2(B[44]), .A3(n216), .ZN(n214) );
  XNOR2_X1 U44 ( .A(B[40]), .B(n221), .ZN(DIFF[40]) );
  XNOR2_X1 U45 ( .A(B[36]), .B(n225), .ZN(DIFF[36]) );
  XNOR2_X1 U46 ( .A(B[32]), .B(n229), .ZN(DIFF[32]) );
  XNOR2_X1 U47 ( .A(B[44]), .B(n217), .ZN(DIFF[44]) );
  OR2_X1 U48 ( .A1(n218), .A2(B[41]), .ZN(n219) );
  OR2_X1 U49 ( .A1(n222), .A2(B[37]), .ZN(n223) );
  OR2_X1 U50 ( .A1(n226), .A2(B[33]), .ZN(n227) );
  OR2_X1 U51 ( .A1(n230), .A2(B[29]), .ZN(n231) );
  OR2_X1 U52 ( .A1(n239), .A2(B[21]), .ZN(n240) );
  OR2_X1 U53 ( .A1(n243), .A2(B[17]), .ZN(n244) );
  NOR2_X1 U54 ( .A1(B[43]), .A2(n216), .ZN(n217) );
  XNOR2_X1 U55 ( .A(B[56]), .B(n203), .ZN(DIFF[56]) );
  XNOR2_X1 U56 ( .A(B[52]), .B(n207), .ZN(DIFF[52]) );
  XNOR2_X1 U57 ( .A(B[48]), .B(n213), .ZN(DIFF[48]) );
  XNOR2_X1 U58 ( .A(n197), .B(B[61]), .ZN(DIFF[61]) );
  XNOR2_X1 U59 ( .A(B[60]), .B(n199), .ZN(DIFF[60]) );
  NOR2_X1 U60 ( .A1(B[15]), .A2(n245), .ZN(n246) );
  OR3_X1 U61 ( .A1(B[15]), .A2(B[16]), .A3(n245), .ZN(n243) );
  OR3_X1 U62 ( .A1(B[13]), .A2(B[14]), .A3(n247), .ZN(n245) );
  OR2_X1 U63 ( .A1(n247), .A2(B[13]), .ZN(n248) );
  XNOR2_X1 U64 ( .A(B[12]), .B(n250), .ZN(DIFF[12]) );
  XNOR2_X1 U65 ( .A(n189), .B(B[6]), .ZN(DIFF[6]) );
  NOR2_X1 U66 ( .A1(n194), .A2(B[5]), .ZN(n189) );
  XNOR2_X1 U67 ( .A(n193), .B(B[10]), .ZN(DIFF[10]) );
  NOR2_X1 U68 ( .A1(n190), .A2(B[9]), .ZN(n193) );
  NOR2_X1 U69 ( .A1(B[11]), .A2(n249), .ZN(n250) );
  XNOR2_X1 U70 ( .A(B[8]), .B(n191), .ZN(DIFF[8]) );
  NOR2_X1 U71 ( .A1(B[7]), .A2(n192), .ZN(n191) );
  XNOR2_X1 U72 ( .A(B[2]), .B(n232), .ZN(DIFF[2]) );
  NOR2_X1 U73 ( .A1(\B[0] ), .A2(B[1]), .ZN(n232) );
  XNOR2_X1 U74 ( .A(B[4]), .B(n210), .ZN(DIFF[4]) );
  NOR2_X1 U75 ( .A1(B[3]), .A2(n211), .ZN(n210) );
  OR3_X1 U76 ( .A1(B[5]), .A2(B[6]), .A3(n194), .ZN(n192) );
  OR3_X1 U77 ( .A1(B[10]), .A2(B[9]), .A3(n190), .ZN(n249) );
  OR3_X1 U78 ( .A1(B[7]), .A2(B[8]), .A3(n192), .ZN(n190) );
  OR3_X1 U79 ( .A1(B[11]), .A2(B[12]), .A3(n249), .ZN(n247) );
  OR3_X1 U80 ( .A1(B[3]), .A2(B[4]), .A3(n211), .ZN(n194) );
  OR3_X1 U83 ( .A1(B[1]), .A2(B[2]), .A3(\B[0] ), .ZN(n211) );
  INV_X1 U126 ( .A(B[61]), .ZN(n251) );
endmodule


module complementer_N64_19 ( \input , complement2 );
  input [63:0] \input ;
  output [63:0] complement2;


  complementer_N64_19_DW01_sub_0 sub_add_31_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(\input ), .CI(1'b0), .DIFF(complement2) );
endmodule


module ShiftnCompl_N64_10 ( plusA, plus2A_out, minus2A_out, plus4A_out, 
        minus4A_out );
  input [63:0] plusA;
  output [63:0] plus2A_out;
  output [63:0] minus2A_out;
  output [63:0] plus4A_out;
  output [63:0] minus4A_out;
  wire   n39, n40, n2, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign plus2A_out[0] = 1'b0;
  assign plus2A_out[51] = n2;
  assign plus4A_out[0] = 1'b0;

  shifter_N64_20 shifter_1 ( .\input (plusA), .shiftLeftOnePos({
        plus2A_out[63:59], n39, plus2A_out[57:54], n40, plus2A_out[52], n2, 
        plus2A_out[50:49], n41, plus2A_out[47:42], n42, n43, n44, n45, n46, 
        n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, 
        n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, 
        plus2A_out[11:1], SYNOPSYS_UNCONNECTED__0}) );
  shifter_N64_19 shifter_2 ( .\input ({plus2A_out[63:52], n2, plus2A_out[50:1], 
        1'b0}), .shiftLeftOnePos({plus4A_out[63:59], n72, plus4A_out[57:54], 
        n73, plus4A_out[52:49], n74, plus4A_out[47:1], SYNOPSYS_UNCONNECTED__1}) );
  complementer_N64_20 complementer_1 ( .\input ({plus2A_out[63:52], n2, 
        plus2A_out[50:1], 1'b0}), .complement2(minus2A_out) );
  complementer_N64_19 complementer_2 ( .\input ({plus4A_out[63:1], 1'b0}), 
        .complement2(minus4A_out) );
  BUF_X1 U1 ( .A(n64), .Z(plus2A_out[19]) );
  BUF_X1 U4 ( .A(n60), .Z(plus2A_out[23]) );
  BUF_X1 U5 ( .A(n62), .Z(plus2A_out[21]) );
  BUF_X1 U6 ( .A(n66), .Z(plus2A_out[17]) );
  BUF_X1 U7 ( .A(n61), .Z(plus2A_out[22]) );
  BUF_X1 U8 ( .A(n63), .Z(plus2A_out[20]) );
  BUF_X1 U9 ( .A(n65), .Z(plus2A_out[18]) );
  BUF_X1 U10 ( .A(n52), .Z(plus2A_out[31]) );
  BUF_X1 U11 ( .A(n50), .Z(plus2A_out[33]) );
  BUF_X1 U12 ( .A(n54), .Z(plus2A_out[29]) );
  BUF_X1 U13 ( .A(n56), .Z(plus2A_out[27]) );
  BUF_X1 U14 ( .A(n58), .Z(plus2A_out[25]) );
  BUF_X1 U15 ( .A(n49), .Z(plus2A_out[34]) );
  BUF_X1 U16 ( .A(n53), .Z(plus2A_out[30]) );
  BUF_X1 U17 ( .A(n57), .Z(plus2A_out[26]) );
  BUF_X1 U18 ( .A(n51), .Z(plus2A_out[32]) );
  BUF_X1 U19 ( .A(n55), .Z(plus2A_out[28]) );
  BUF_X1 U20 ( .A(n59), .Z(plus2A_out[24]) );
  BUF_X1 U21 ( .A(n44), .Z(plus2A_out[39]) );
  BUF_X1 U22 ( .A(n48), .Z(plus2A_out[35]) );
  BUF_X1 U23 ( .A(n42), .Z(plus2A_out[41]) );
  BUF_X1 U24 ( .A(n46), .Z(plus2A_out[37]) );
  BUF_X1 U25 ( .A(n45), .Z(plus2A_out[38]) );
  BUF_X1 U26 ( .A(n43), .Z(plus2A_out[40]) );
  BUF_X1 U27 ( .A(n47), .Z(plus2A_out[36]) );
  BUF_X1 U28 ( .A(n41), .Z(plus2A_out[48]) );
  BUF_X1 U29 ( .A(n74), .Z(plus4A_out[48]) );
  BUF_X1 U30 ( .A(n40), .Z(plus2A_out[53]) );
  BUF_X1 U31 ( .A(n73), .Z(plus4A_out[53]) );
  BUF_X1 U32 ( .A(n72), .Z(plus4A_out[58]) );
  BUF_X1 U33 ( .A(n39), .Z(plus2A_out[58]) );
  BUF_X1 U34 ( .A(n68), .Z(plus2A_out[15]) );
  BUF_X1 U35 ( .A(n70), .Z(plus2A_out[13]) );
  BUF_X1 U36 ( .A(n67), .Z(plus2A_out[16]) );
  BUF_X1 U37 ( .A(n71), .Z(plus2A_out[12]) );
  BUF_X1 U38 ( .A(n69), .Z(plus2A_out[14]) );
endmodule


module MUX_GENERIC_N64_RADIX3_10 ( plusA, minusA, plus2A, minus2A, SEL, Y );
  input [63:0] plusA;
  input [63:0] minusA;
  input [63:0] plus2A;
  input [63:0] minus2A;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502;
  tri   [63:0] Y;

  TBUF_X1 \Y_tri[55]  ( .A(n446), .EN(n301), .Z(Y[55]) );
  TBUF_X1 \Y_tri[56]  ( .A(n445), .EN(n301), .Z(Y[56]) );
  TBUF_X1 \Y_tri[57]  ( .A(n444), .EN(n301), .Z(Y[57]) );
  TBUF_X1 \Y_tri[58]  ( .A(n443), .EN(n301), .Z(Y[58]) );
  TBUF_X1 \Y_tri[59]  ( .A(n442), .EN(n301), .Z(Y[59]) );
  TBUF_X1 \Y_tri[60]  ( .A(n441), .EN(n301), .Z(Y[60]) );
  TBUF_X1 \Y_tri[61]  ( .A(n440), .EN(n301), .Z(Y[61]) );
  TBUF_X1 \Y_tri[62]  ( .A(n439), .EN(n301), .Z(Y[62]) );
  TBUF_X1 \Y_tri[63]  ( .A(n438), .EN(n301), .Z(Y[63]) );
  TBUF_X1 \Y_tri[47]  ( .A(n454), .EN(n300), .Z(Y[47]) );
  TBUF_X1 \Y_tri[48]  ( .A(n453), .EN(n300), .Z(Y[48]) );
  TBUF_X1 \Y_tri[49]  ( .A(n452), .EN(n300), .Z(Y[49]) );
  TBUF_X1 \Y_tri[50]  ( .A(n451), .EN(n300), .Z(Y[50]) );
  TBUF_X1 \Y_tri[51]  ( .A(n450), .EN(n300), .Z(Y[51]) );
  TBUF_X1 \Y_tri[53]  ( .A(n448), .EN(n300), .Z(Y[53]) );
  TBUF_X1 \Y_tri[54]  ( .A(n447), .EN(n300), .Z(Y[54]) );
  TBUF_X1 \Y_tri[46]  ( .A(n455), .EN(n300), .Z(Y[46]) );
  TBUF_X1 \Y_tri[52]  ( .A(n449), .EN(n300), .Z(Y[52]) );
  TBUF_X1 \Y_tri[21]  ( .A(n480), .EN(n297), .Z(Y[21]) );
  TBUF_X1 \Y_tri[22]  ( .A(n479), .EN(n298), .Z(Y[22]) );
  TBUF_X1 \Y_tri[28]  ( .A(n473), .EN(n298), .Z(Y[28]) );
  TBUF_X1 \Y_tri[29]  ( .A(n472), .EN(n298), .Z(Y[29]) );
  TBUF_X1 \Y_tri[30]  ( .A(n471), .EN(n298), .Z(Y[30]) );
  TBUF_X1 \Y_tri[31]  ( .A(n470), .EN(n298), .Z(Y[31]) );
  TBUF_X1 \Y_tri[32]  ( .A(n469), .EN(n298), .Z(Y[32]) );
  TBUF_X1 \Y_tri[33]  ( .A(n468), .EN(n299), .Z(Y[33]) );
  TBUF_X1 \Y_tri[34]  ( .A(n467), .EN(n299), .Z(Y[34]) );
  TBUF_X1 \Y_tri[35]  ( .A(n466), .EN(n299), .Z(Y[35]) );
  TBUF_X1 \Y_tri[36]  ( .A(n465), .EN(n299), .Z(Y[36]) );
  TBUF_X1 \Y_tri[37]  ( .A(n464), .EN(n299), .Z(Y[37]) );
  TBUF_X1 \Y_tri[38]  ( .A(n463), .EN(n299), .Z(Y[38]) );
  TBUF_X1 \Y_tri[39]  ( .A(n462), .EN(n299), .Z(Y[39]) );
  TBUF_X1 \Y_tri[40]  ( .A(n461), .EN(n299), .Z(Y[40]) );
  TBUF_X1 \Y_tri[41]  ( .A(n460), .EN(n299), .Z(Y[41]) );
  TBUF_X1 \Y_tri[42]  ( .A(n459), .EN(n299), .Z(Y[42]) );
  TBUF_X1 \Y_tri[43]  ( .A(n458), .EN(n299), .Z(Y[43]) );
  TBUF_X1 \Y_tri[44]  ( .A(n457), .EN(n300), .Z(Y[44]) );
  TBUF_X1 \Y_tri[25]  ( .A(n476), .EN(n298), .Z(Y[25]) );
  TBUF_X1 \Y_tri[4]  ( .A(n498), .EN(n296), .Z(Y[4]) );
  TBUF_X1 \Y_tri[5]  ( .A(n497), .EN(n296), .Z(Y[5]) );
  TBUF_X1 \Y_tri[7]  ( .A(n495), .EN(n296), .Z(Y[7]) );
  TBUF_X1 \Y_tri[8]  ( .A(n494), .EN(n296), .Z(Y[8]) );
  TBUF_X1 \Y_tri[10]  ( .A(n491), .EN(n296), .Z(Y[10]) );
  TBUF_X1 \Y_tri[11]  ( .A(n490), .EN(n297), .Z(Y[11]) );
  TBUF_X1 \Y_tri[12]  ( .A(n489), .EN(n297), .Z(Y[12]) );
  TBUF_X1 \Y_tri[14]  ( .A(n487), .EN(n297), .Z(Y[14]) );
  TBUF_X1 \Y_tri[15]  ( .A(n486), .EN(n297), .Z(Y[15]) );
  TBUF_X1 \Y_tri[16]  ( .A(n485), .EN(n297), .Z(Y[16]) );
  TBUF_X1 \Y_tri[17]  ( .A(n484), .EN(n297), .Z(Y[17]) );
  TBUF_X1 \Y_tri[18]  ( .A(n483), .EN(n297), .Z(Y[18]) );
  TBUF_X1 \Y_tri[19]  ( .A(n482), .EN(n297), .Z(Y[19]) );
  TBUF_X1 \Y_tri[20]  ( .A(n481), .EN(n297), .Z(Y[20]) );
  TBUF_X1 \Y_tri[9]  ( .A(n492), .EN(n296), .Z(Y[9]) );
  TBUF_X1 \Y_tri[0]  ( .A(n502), .EN(n296), .Z(Y[0]) );
  TBUF_X1 \Y_tri[2]  ( .A(n500), .EN(n296), .Z(Y[2]) );
  TBUF_X1 \Y_tri[3]  ( .A(n499), .EN(n296), .Z(Y[3]) );
  TBUF_X1 \Y_tri[1]  ( .A(n501), .EN(n296), .Z(Y[1]) );
  TBUF_X1 \Y_tri[6]  ( .A(n496), .EN(n296), .Z(Y[6]) );
  TBUF_X1 \Y_tri[13]  ( .A(n488), .EN(n297), .Z(Y[13]) );
  TBUF_X1 \Y_tri[23]  ( .A(n478), .EN(n298), .Z(Y[23]) );
  TBUF_X1 \Y_tri[24]  ( .A(n477), .EN(n298), .Z(Y[24]) );
  TBUF_X1 \Y_tri[26]  ( .A(n475), .EN(n298), .Z(Y[26]) );
  TBUF_X1 \Y_tri[27]  ( .A(n474), .EN(n298), .Z(Y[27]) );
  TBUF_X1 \Y_tri[45]  ( .A(n456), .EN(n300), .Z(Y[45]) );
  NAND2_X1 U2 ( .A1(n361), .A2(n360), .ZN(n474) );
  AOI22_X1 U3 ( .A1(plusA[27]), .A2(n280), .B1(plus2A[27]), .B2(n274), .ZN(
        n361) );
  AOI22_X1 U4 ( .A1(minus2A[27]), .A2(n292), .B1(minusA[27]), .B2(n286), .ZN(
        n360) );
  NAND2_X1 U5 ( .A1(n359), .A2(n358), .ZN(n475) );
  AOI22_X1 U6 ( .A1(plusA[26]), .A2(n280), .B1(plus2A[26]), .B2(n274), .ZN(
        n359) );
  AOI22_X1 U7 ( .A1(minus2A[26]), .A2(n292), .B1(minusA[26]), .B2(n286), .ZN(
        n358) );
  NAND2_X1 U8 ( .A1(n353), .A2(n352), .ZN(n478) );
  AOI22_X1 U9 ( .A1(plusA[23]), .A2(n279), .B1(plus2A[23]), .B2(n273), .ZN(
        n353) );
  AOI22_X1 U10 ( .A1(minus2A[23]), .A2(n291), .B1(minusA[23]), .B2(n285), .ZN(
        n352) );
  NAND2_X1 U11 ( .A1(n347), .A2(n346), .ZN(n481) );
  AOI22_X1 U12 ( .A1(plusA[20]), .A2(n279), .B1(plus2A[20]), .B2(n273), .ZN(
        n347) );
  AOI22_X1 U13 ( .A1(minus2A[20]), .A2(n291), .B1(minusA[20]), .B2(n285), .ZN(
        n346) );
  NAND2_X1 U14 ( .A1(n345), .A2(n344), .ZN(n482) );
  AOI22_X1 U15 ( .A1(plusA[19]), .A2(n279), .B1(plus2A[19]), .B2(n273), .ZN(
        n345) );
  AOI22_X1 U16 ( .A1(minus2A[19]), .A2(n291), .B1(minusA[19]), .B2(n285), .ZN(
        n344) );
  NAND2_X1 U17 ( .A1(n343), .A2(n342), .ZN(n483) );
  AOI22_X1 U18 ( .A1(plusA[18]), .A2(n279), .B1(plus2A[18]), .B2(n273), .ZN(
        n343) );
  AOI22_X1 U19 ( .A1(minus2A[18]), .A2(n291), .B1(minusA[18]), .B2(n285), .ZN(
        n342) );
  NAND2_X1 U20 ( .A1(n341), .A2(n340), .ZN(n484) );
  AOI22_X1 U21 ( .A1(plusA[17]), .A2(n279), .B1(plus2A[17]), .B2(n273), .ZN(
        n341) );
  AOI22_X1 U22 ( .A1(minus2A[17]), .A2(n291), .B1(minusA[17]), .B2(n285), .ZN(
        n340) );
  NAND2_X1 U23 ( .A1(n339), .A2(n338), .ZN(n485) );
  AOI22_X1 U24 ( .A1(plusA[16]), .A2(n279), .B1(plus2A[16]), .B2(n273), .ZN(
        n339) );
  AOI22_X1 U25 ( .A1(minus2A[16]), .A2(n291), .B1(minusA[16]), .B2(n285), .ZN(
        n338) );
  NAND2_X1 U26 ( .A1(n355), .A2(n354), .ZN(n477) );
  AOI22_X1 U27 ( .A1(plusA[24]), .A2(n280), .B1(plus2A[24]), .B2(n274), .ZN(
        n355) );
  AOI22_X1 U28 ( .A1(minus2A[24]), .A2(n292), .B1(minusA[24]), .B2(n286), .ZN(
        n354) );
  NAND2_X1 U29 ( .A1(n363), .A2(n362), .ZN(n473) );
  AOI22_X1 U30 ( .A1(plusA[28]), .A2(n280), .B1(plus2A[28]), .B2(n274), .ZN(
        n363) );
  AOI22_X1 U31 ( .A1(minus2A[28]), .A2(n292), .B1(minusA[28]), .B2(n286), .ZN(
        n362) );
  NAND2_X1 U32 ( .A1(n357), .A2(n356), .ZN(n476) );
  AOI22_X1 U33 ( .A1(plusA[25]), .A2(n280), .B1(plus2A[25]), .B2(n274), .ZN(
        n357) );
  AOI22_X1 U34 ( .A1(minus2A[25]), .A2(n292), .B1(minusA[25]), .B2(n286), .ZN(
        n356) );
  NAND2_X1 U35 ( .A1(n351), .A2(n350), .ZN(n479) );
  AOI22_X1 U36 ( .A1(plusA[22]), .A2(n279), .B1(plus2A[22]), .B2(n273), .ZN(
        n351) );
  AOI22_X1 U37 ( .A1(minus2A[22]), .A2(n291), .B1(minusA[22]), .B2(n285), .ZN(
        n350) );
  NAND2_X1 U38 ( .A1(n349), .A2(n348), .ZN(n480) );
  AOI22_X1 U39 ( .A1(plusA[21]), .A2(n279), .B1(plus2A[21]), .B2(n273), .ZN(
        n349) );
  AOI22_X1 U40 ( .A1(minus2A[21]), .A2(n291), .B1(minusA[21]), .B2(n285), .ZN(
        n348) );
  NAND2_X1 U41 ( .A1(n387), .A2(n386), .ZN(n461) );
  AOI22_X1 U42 ( .A1(plusA[40]), .A2(n281), .B1(plus2A[40]), .B2(n275), .ZN(
        n387) );
  AOI22_X1 U43 ( .A1(minus2A[40]), .A2(n293), .B1(minusA[40]), .B2(n287), .ZN(
        n386) );
  NAND2_X1 U44 ( .A1(n379), .A2(n378), .ZN(n465) );
  AOI22_X1 U45 ( .A1(plusA[36]), .A2(n281), .B1(plus2A[36]), .B2(n275), .ZN(
        n379) );
  AOI22_X1 U46 ( .A1(minus2A[36]), .A2(n293), .B1(minusA[36]), .B2(n287), .ZN(
        n378) );
  NAND2_X1 U47 ( .A1(n371), .A2(n370), .ZN(n469) );
  AOI22_X1 U48 ( .A1(plusA[32]), .A2(n280), .B1(plus2A[32]), .B2(n274), .ZN(
        n371) );
  AOI22_X1 U49 ( .A1(minus2A[32]), .A2(n292), .B1(minusA[32]), .B2(n286), .ZN(
        n370) );
  NAND2_X1 U50 ( .A1(n397), .A2(n396), .ZN(n456) );
  AOI22_X1 U51 ( .A1(plusA[45]), .A2(n281), .B1(plus2A[45]), .B2(n275), .ZN(
        n397) );
  AOI22_X1 U52 ( .A1(minus2A[45]), .A2(n293), .B1(minusA[45]), .B2(n287), .ZN(
        n396) );
  NAND2_X1 U53 ( .A1(n391), .A2(n390), .ZN(n459) );
  AOI22_X1 U54 ( .A1(plusA[42]), .A2(n281), .B1(plus2A[42]), .B2(n275), .ZN(
        n391) );
  AOI22_X1 U55 ( .A1(minus2A[42]), .A2(n293), .B1(minusA[42]), .B2(n287), .ZN(
        n390) );
  NAND2_X1 U56 ( .A1(n383), .A2(n382), .ZN(n463) );
  AOI22_X1 U57 ( .A1(plusA[38]), .A2(n281), .B1(plus2A[38]), .B2(n275), .ZN(
        n383) );
  AOI22_X1 U58 ( .A1(minus2A[38]), .A2(n293), .B1(minusA[38]), .B2(n287), .ZN(
        n382) );
  NAND2_X1 U59 ( .A1(n375), .A2(n374), .ZN(n467) );
  AOI22_X1 U60 ( .A1(plusA[34]), .A2(n280), .B1(plus2A[34]), .B2(n274), .ZN(
        n375) );
  AOI22_X1 U61 ( .A1(minus2A[34]), .A2(n292), .B1(minusA[34]), .B2(n286), .ZN(
        n374) );
  NAND2_X1 U62 ( .A1(n367), .A2(n366), .ZN(n471) );
  AOI22_X1 U63 ( .A1(plusA[30]), .A2(n280), .B1(plus2A[30]), .B2(n274), .ZN(
        n367) );
  AOI22_X1 U64 ( .A1(minus2A[30]), .A2(n292), .B1(minusA[30]), .B2(n286), .ZN(
        n366) );
  NAND2_X1 U65 ( .A1(n393), .A2(n392), .ZN(n458) );
  AOI22_X1 U66 ( .A1(plusA[43]), .A2(n281), .B1(plus2A[43]), .B2(n275), .ZN(
        n393) );
  AOI22_X1 U67 ( .A1(minus2A[43]), .A2(n293), .B1(minusA[43]), .B2(n287), .ZN(
        n392) );
  NAND2_X1 U68 ( .A1(n389), .A2(n388), .ZN(n460) );
  AOI22_X1 U69 ( .A1(plusA[41]), .A2(n281), .B1(plus2A[41]), .B2(n275), .ZN(
        n389) );
  AOI22_X1 U70 ( .A1(minus2A[41]), .A2(n293), .B1(minusA[41]), .B2(n287), .ZN(
        n388) );
  NAND2_X1 U71 ( .A1(n381), .A2(n380), .ZN(n464) );
  AOI22_X1 U72 ( .A1(plusA[37]), .A2(n281), .B1(plus2A[37]), .B2(n275), .ZN(
        n381) );
  AOI22_X1 U73 ( .A1(minus2A[37]), .A2(n293), .B1(minusA[37]), .B2(n287), .ZN(
        n380) );
  NAND2_X1 U74 ( .A1(n373), .A2(n372), .ZN(n468) );
  AOI22_X1 U75 ( .A1(plusA[33]), .A2(n280), .B1(plus2A[33]), .B2(n274), .ZN(
        n373) );
  AOI22_X1 U76 ( .A1(minus2A[33]), .A2(n292), .B1(minusA[33]), .B2(n286), .ZN(
        n372) );
  NAND2_X1 U77 ( .A1(n365), .A2(n364), .ZN(n472) );
  AOI22_X1 U78 ( .A1(plusA[29]), .A2(n280), .B1(plus2A[29]), .B2(n274), .ZN(
        n365) );
  AOI22_X1 U79 ( .A1(minus2A[29]), .A2(n292), .B1(minusA[29]), .B2(n286), .ZN(
        n364) );
  NAND2_X1 U80 ( .A1(n385), .A2(n384), .ZN(n462) );
  AOI22_X1 U81 ( .A1(plusA[39]), .A2(n281), .B1(plus2A[39]), .B2(n275), .ZN(
        n385) );
  AOI22_X1 U82 ( .A1(minus2A[39]), .A2(n293), .B1(minusA[39]), .B2(n287), .ZN(
        n384) );
  NAND2_X1 U83 ( .A1(n377), .A2(n376), .ZN(n466) );
  AOI22_X1 U84 ( .A1(plusA[35]), .A2(n280), .B1(plus2A[35]), .B2(n274), .ZN(
        n377) );
  AOI22_X1 U85 ( .A1(minus2A[35]), .A2(n292), .B1(minusA[35]), .B2(n286), .ZN(
        n376) );
  NAND2_X1 U86 ( .A1(n369), .A2(n368), .ZN(n470) );
  AOI22_X1 U87 ( .A1(plusA[31]), .A2(n280), .B1(plus2A[31]), .B2(n274), .ZN(
        n369) );
  AOI22_X1 U88 ( .A1(minus2A[31]), .A2(n292), .B1(minusA[31]), .B2(n286), .ZN(
        n368) );
  NAND2_X1 U89 ( .A1(n395), .A2(n394), .ZN(n457) );
  AOI22_X1 U90 ( .A1(plusA[44]), .A2(n281), .B1(plus2A[44]), .B2(n275), .ZN(
        n395) );
  AOI22_X1 U91 ( .A1(minus2A[44]), .A2(n293), .B1(minusA[44]), .B2(n287), .ZN(
        n394) );
  NAND2_X1 U92 ( .A1(n399), .A2(n398), .ZN(n455) );
  AOI22_X1 U93 ( .A1(plusA[46]), .A2(n281), .B1(plus2A[46]), .B2(n275), .ZN(
        n399) );
  AOI22_X1 U94 ( .A1(minus2A[46]), .A2(n293), .B1(minusA[46]), .B2(n287), .ZN(
        n398) );
  NAND2_X1 U95 ( .A1(n401), .A2(n400), .ZN(n454) );
  AOI22_X1 U96 ( .A1(plusA[47]), .A2(n281), .B1(plus2A[47]), .B2(n275), .ZN(
        n401) );
  AOI22_X1 U97 ( .A1(minus2A[47]), .A2(n293), .B1(minusA[47]), .B2(n287), .ZN(
        n400) );
  NAND2_X1 U98 ( .A1(n419), .A2(n418), .ZN(n445) );
  AOI22_X1 U99 ( .A1(plusA[56]), .A2(n282), .B1(plus2A[56]), .B2(n276), .ZN(
        n419) );
  AOI22_X1 U100 ( .A1(minus2A[56]), .A2(n294), .B1(minusA[56]), .B2(n288), 
        .ZN(n418) );
  NAND2_X1 U101 ( .A1(n415), .A2(n414), .ZN(n447) );
  AOI22_X1 U102 ( .A1(plusA[54]), .A2(n282), .B1(plus2A[54]), .B2(n276), .ZN(
        n415) );
  AOI22_X1 U103 ( .A1(minus2A[54]), .A2(n294), .B1(minusA[54]), .B2(n288), 
        .ZN(n414) );
  NAND2_X1 U104 ( .A1(n421), .A2(n420), .ZN(n444) );
  AOI22_X1 U105 ( .A1(plusA[57]), .A2(n282), .B1(plus2A[57]), .B2(n276), .ZN(
        n421) );
  AOI22_X1 U106 ( .A1(minus2A[57]), .A2(n294), .B1(minusA[57]), .B2(n288), 
        .ZN(n420) );
  NAND2_X1 U107 ( .A1(n417), .A2(n416), .ZN(n446) );
  AOI22_X1 U108 ( .A1(plusA[55]), .A2(n282), .B1(plus2A[55]), .B2(n276), .ZN(
        n417) );
  AOI22_X1 U109 ( .A1(minus2A[55]), .A2(n294), .B1(minusA[55]), .B2(n288), 
        .ZN(n416) );
  NAND2_X1 U110 ( .A1(n413), .A2(n412), .ZN(n448) );
  AOI22_X1 U111 ( .A1(plusA[53]), .A2(n282), .B1(plus2A[53]), .B2(n276), .ZN(
        n413) );
  AOI22_X1 U112 ( .A1(minus2A[53]), .A2(n294), .B1(minusA[53]), .B2(n288), 
        .ZN(n412) );
  NAND2_X1 U113 ( .A1(n409), .A2(n408), .ZN(n450) );
  AOI22_X1 U114 ( .A1(plusA[51]), .A2(n282), .B1(plus2A[51]), .B2(n276), .ZN(
        n409) );
  AOI22_X1 U115 ( .A1(minus2A[51]), .A2(n294), .B1(minusA[51]), .B2(n288), 
        .ZN(n408) );
  NAND2_X1 U116 ( .A1(n405), .A2(n404), .ZN(n452) );
  AOI22_X1 U117 ( .A1(plusA[49]), .A2(n282), .B1(plus2A[49]), .B2(n276), .ZN(
        n405) );
  AOI22_X1 U118 ( .A1(minus2A[49]), .A2(n294), .B1(minusA[49]), .B2(n288), 
        .ZN(n404) );
  NAND2_X1 U119 ( .A1(n411), .A2(n410), .ZN(n449) );
  AOI22_X1 U120 ( .A1(plusA[52]), .A2(n282), .B1(plus2A[52]), .B2(n276), .ZN(
        n411) );
  AOI22_X1 U121 ( .A1(minus2A[52]), .A2(n294), .B1(minusA[52]), .B2(n288), 
        .ZN(n410) );
  NAND2_X1 U122 ( .A1(n407), .A2(n406), .ZN(n451) );
  AOI22_X1 U123 ( .A1(plusA[50]), .A2(n282), .B1(plus2A[50]), .B2(n276), .ZN(
        n407) );
  AOI22_X1 U124 ( .A1(minus2A[50]), .A2(n294), .B1(minusA[50]), .B2(n288), 
        .ZN(n406) );
  NAND2_X1 U125 ( .A1(n403), .A2(n402), .ZN(n453) );
  AOI22_X1 U126 ( .A1(plusA[48]), .A2(n282), .B1(plus2A[48]), .B2(n276), .ZN(
        n403) );
  AOI22_X1 U127 ( .A1(minus2A[48]), .A2(n294), .B1(minusA[48]), .B2(n288), 
        .ZN(n402) );
  NAND2_X1 U128 ( .A1(n437), .A2(n436), .ZN(n438) );
  AOI22_X1 U129 ( .A1(plusA[63]), .A2(n283), .B1(plus2A[63]), .B2(n277), .ZN(
        n437) );
  AOI22_X1 U130 ( .A1(minus2A[63]), .A2(n295), .B1(minusA[63]), .B2(n289), 
        .ZN(n436) );
  NAND2_X1 U131 ( .A1(n431), .A2(n430), .ZN(n439) );
  AOI22_X1 U132 ( .A1(plusA[62]), .A2(n283), .B1(plus2A[62]), .B2(n277), .ZN(
        n431) );
  AOI22_X1 U133 ( .A1(minus2A[62]), .A2(n295), .B1(minusA[62]), .B2(n289), 
        .ZN(n430) );
  NAND2_X1 U134 ( .A1(n429), .A2(n428), .ZN(n440) );
  AOI22_X1 U135 ( .A1(plusA[61]), .A2(n283), .B1(plus2A[61]), .B2(n277), .ZN(
        n429) );
  AOI22_X1 U136 ( .A1(minus2A[61]), .A2(n295), .B1(minusA[61]), .B2(n289), 
        .ZN(n428) );
  NAND2_X1 U137 ( .A1(n427), .A2(n426), .ZN(n441) );
  AOI22_X1 U138 ( .A1(plusA[60]), .A2(n283), .B1(plus2A[60]), .B2(n277), .ZN(
        n427) );
  AOI22_X1 U139 ( .A1(minus2A[60]), .A2(n295), .B1(minusA[60]), .B2(n289), 
        .ZN(n426) );
  NAND2_X1 U140 ( .A1(n425), .A2(n424), .ZN(n442) );
  AOI22_X1 U141 ( .A1(plusA[59]), .A2(n282), .B1(plus2A[59]), .B2(n276), .ZN(
        n425) );
  AOI22_X1 U142 ( .A1(minus2A[59]), .A2(n294), .B1(minusA[59]), .B2(n288), 
        .ZN(n424) );
  NAND2_X1 U143 ( .A1(n423), .A2(n422), .ZN(n443) );
  AOI22_X1 U144 ( .A1(plusA[58]), .A2(n282), .B1(plus2A[58]), .B2(n276), .ZN(
        n423) );
  AOI22_X1 U145 ( .A1(minus2A[58]), .A2(n294), .B1(minusA[58]), .B2(n288), 
        .ZN(n422) );
  BUF_X1 U146 ( .A(n493), .Z(n296) );
  BUF_X1 U147 ( .A(n433), .Z(n279) );
  BUF_X1 U148 ( .A(n435), .Z(n291) );
  BUF_X1 U149 ( .A(n434), .Z(n285) );
  BUF_X1 U150 ( .A(n432), .Z(n273) );
  BUF_X1 U151 ( .A(n493), .Z(n297) );
  NAND2_X1 U152 ( .A1(n337), .A2(n336), .ZN(n486) );
  AOI22_X1 U153 ( .A1(plusA[15]), .A2(n279), .B1(plus2A[15]), .B2(n273), .ZN(
        n337) );
  AOI22_X1 U154 ( .A1(minus2A[15]), .A2(n291), .B1(minusA[15]), .B2(n285), 
        .ZN(n336) );
  NAND2_X1 U155 ( .A1(n335), .A2(n334), .ZN(n487) );
  AOI22_X1 U156 ( .A1(plusA[14]), .A2(n279), .B1(plus2A[14]), .B2(n273), .ZN(
        n335) );
  AOI22_X1 U157 ( .A1(minus2A[14]), .A2(n291), .B1(minusA[14]), .B2(n285), 
        .ZN(n334) );
  BUF_X1 U158 ( .A(n433), .Z(n280) );
  BUF_X1 U159 ( .A(n435), .Z(n292) );
  BUF_X1 U160 ( .A(n434), .Z(n286) );
  BUF_X1 U161 ( .A(n432), .Z(n274) );
  BUF_X1 U162 ( .A(n493), .Z(n298) );
  BUF_X1 U163 ( .A(n493), .Z(n299) );
  BUF_X1 U164 ( .A(n433), .Z(n281) );
  BUF_X1 U165 ( .A(n435), .Z(n293) );
  BUF_X1 U166 ( .A(n434), .Z(n287) );
  BUF_X1 U167 ( .A(n432), .Z(n275) );
  BUF_X1 U168 ( .A(n493), .Z(n300) );
  BUF_X1 U169 ( .A(n433), .Z(n282) );
  BUF_X1 U170 ( .A(n435), .Z(n294) );
  BUF_X1 U171 ( .A(n434), .Z(n288) );
  BUF_X1 U172 ( .A(n432), .Z(n276) );
  BUF_X1 U173 ( .A(n493), .Z(n301) );
  BUF_X1 U174 ( .A(n433), .Z(n278) );
  BUF_X1 U175 ( .A(n435), .Z(n290) );
  BUF_X1 U176 ( .A(n434), .Z(n284) );
  BUF_X1 U177 ( .A(n432), .Z(n272) );
  NOR2_X1 U178 ( .A1(n323), .A2(n304), .ZN(n493) );
  INV_X1 U179 ( .A(SEL[2]), .ZN(n304) );
  NOR2_X1 U180 ( .A1(SEL[1]), .A2(SEL[0]), .ZN(n323) );
  NOR3_X1 U181 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n302), .ZN(n434) );
  NOR3_X1 U182 ( .A1(SEL[1]), .A2(SEL[2]), .A3(n303), .ZN(n433) );
  NOR3_X1 U183 ( .A1(n302), .A2(SEL[2]), .A3(n303), .ZN(n432) );
  NAND2_X1 U184 ( .A1(n333), .A2(n332), .ZN(n488) );
  AOI22_X1 U185 ( .A1(plusA[13]), .A2(n279), .B1(plus2A[13]), .B2(n273), .ZN(
        n333) );
  AOI22_X1 U186 ( .A1(minus2A[13]), .A2(n291), .B1(minusA[13]), .B2(n285), 
        .ZN(n332) );
  AND2_X1 U187 ( .A1(SEL[2]), .A2(n323), .ZN(n435) );
  INV_X1 U188 ( .A(SEL[1]), .ZN(n302) );
  INV_X1 U189 ( .A(SEL[0]), .ZN(n303) );
  NAND2_X1 U190 ( .A1(n331), .A2(n330), .ZN(n489) );
  AOI22_X1 U191 ( .A1(plusA[12]), .A2(n279), .B1(plus2A[12]), .B2(n273), .ZN(
        n331) );
  AOI22_X1 U192 ( .A1(minus2A[12]), .A2(n291), .B1(minusA[12]), .B2(n285), 
        .ZN(n330) );
  NAND2_X1 U193 ( .A1(n329), .A2(n328), .ZN(n490) );
  AOI22_X1 U194 ( .A1(plusA[11]), .A2(n278), .B1(plus2A[11]), .B2(n272), .ZN(
        n329) );
  AOI22_X1 U195 ( .A1(minus2A[11]), .A2(n290), .B1(minusA[11]), .B2(n284), 
        .ZN(n328) );
  NAND2_X1 U196 ( .A1(n327), .A2(n326), .ZN(n491) );
  AOI22_X1 U197 ( .A1(plusA[10]), .A2(n278), .B1(plus2A[10]), .B2(n272), .ZN(
        n327) );
  AOI22_X1 U198 ( .A1(minus2A[10]), .A2(n290), .B1(minusA[10]), .B2(n284), 
        .ZN(n326) );
  NAND2_X1 U199 ( .A1(n325), .A2(n324), .ZN(n492) );
  AOI22_X1 U200 ( .A1(plusA[9]), .A2(n278), .B1(plus2A[9]), .B2(n272), .ZN(
        n325) );
  AOI22_X1 U201 ( .A1(minus2A[9]), .A2(n290), .B1(minusA[9]), .B2(n284), .ZN(
        n324) );
  NAND2_X1 U202 ( .A1(n320), .A2(n319), .ZN(n495) );
  AOI22_X1 U203 ( .A1(plusA[7]), .A2(n278), .B1(plus2A[7]), .B2(n272), .ZN(
        n320) );
  AOI22_X1 U204 ( .A1(minus2A[7]), .A2(n290), .B1(minusA[7]), .B2(n284), .ZN(
        n319) );
  NAND2_X1 U205 ( .A1(n318), .A2(n317), .ZN(n496) );
  AOI22_X1 U206 ( .A1(plusA[6]), .A2(n278), .B1(plus2A[6]), .B2(n272), .ZN(
        n318) );
  AOI22_X1 U207 ( .A1(minus2A[6]), .A2(n290), .B1(minusA[6]), .B2(n284), .ZN(
        n317) );
  NAND2_X1 U208 ( .A1(n316), .A2(n315), .ZN(n497) );
  AOI22_X1 U209 ( .A1(plusA[5]), .A2(n278), .B1(plus2A[5]), .B2(n272), .ZN(
        n316) );
  AOI22_X1 U210 ( .A1(minus2A[5]), .A2(n290), .B1(minusA[5]), .B2(n284), .ZN(
        n315) );
  NAND2_X1 U211 ( .A1(n312), .A2(n311), .ZN(n499) );
  AOI22_X1 U212 ( .A1(plusA[3]), .A2(n278), .B1(plus2A[3]), .B2(n272), .ZN(
        n312) );
  AOI22_X1 U213 ( .A1(minus2A[3]), .A2(n290), .B1(minusA[3]), .B2(n284), .ZN(
        n311) );
  NAND2_X1 U214 ( .A1(n322), .A2(n321), .ZN(n494) );
  AOI22_X1 U215 ( .A1(plusA[8]), .A2(n278), .B1(plus2A[8]), .B2(n272), .ZN(
        n322) );
  AOI22_X1 U216 ( .A1(minus2A[8]), .A2(n290), .B1(minusA[8]), .B2(n284), .ZN(
        n321) );
  NAND2_X1 U217 ( .A1(n314), .A2(n313), .ZN(n498) );
  AOI22_X1 U218 ( .A1(plusA[4]), .A2(n278), .B1(plus2A[4]), .B2(n272), .ZN(
        n314) );
  AOI22_X1 U219 ( .A1(minus2A[4]), .A2(n290), .B1(minusA[4]), .B2(n284), .ZN(
        n313) );
  NAND2_X1 U220 ( .A1(n310), .A2(n309), .ZN(n500) );
  AOI22_X1 U221 ( .A1(plusA[2]), .A2(n278), .B1(plus2A[2]), .B2(n272), .ZN(
        n310) );
  AOI22_X1 U222 ( .A1(minus2A[2]), .A2(n290), .B1(minusA[2]), .B2(n284), .ZN(
        n309) );
  NAND2_X1 U223 ( .A1(n308), .A2(n307), .ZN(n501) );
  AOI22_X1 U224 ( .A1(plusA[1]), .A2(n278), .B1(plus2A[1]), .B2(n272), .ZN(
        n308) );
  AOI22_X1 U225 ( .A1(minus2A[1]), .A2(n290), .B1(minusA[1]), .B2(n284), .ZN(
        n307) );
  NAND2_X1 U226 ( .A1(n306), .A2(n305), .ZN(n502) );
  AOI22_X1 U227 ( .A1(plusA[0]), .A2(n278), .B1(plus2A[0]), .B2(n272), .ZN(
        n306) );
  AOI22_X1 U228 ( .A1(minus2A[0]), .A2(n290), .B1(minusA[0]), .B2(n284), .ZN(
        n305) );
  CLKBUF_X1 U229 ( .A(n432), .Z(n277) );
  CLKBUF_X1 U230 ( .A(n433), .Z(n283) );
  CLKBUF_X1 U231 ( .A(n434), .Z(n289) );
  CLKBUF_X1 U232 ( .A(n435), .Z(n295) );
endmodule


module FA_640 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_639 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;
  tri   A;

  XOR2_X1 U3 ( .A(n6), .B(Ci), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  XNOR2_X1 U4 ( .A(n4), .B(B), .ZN(n6) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_638 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_637 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_636 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_635 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_634 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_633 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_632 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_631 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_630 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_629 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_628 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_627 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  AOI22_X1 U4 ( .A1(B), .A2(A), .B1(Ci), .B2(n6), .ZN(n7) );
  INV_X1 U5 ( .A(n7), .ZN(Co) );
endmodule


module FA_626 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_625 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_624 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_623 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  XOR2_X1 U1 ( .A(Ci), .B(n5), .Z(S) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_622 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(n5), .B(Ci), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_621 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_620 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_619 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_618 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_617 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  AOI22_X1 U4 ( .A1(B), .A2(A), .B1(Ci), .B2(n6), .ZN(n7) );
  INV_X1 U5 ( .A(n7), .ZN(Co) );
endmodule


module FA_616 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_615 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_614 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  AOI22_X1 U4 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
  INV_X1 U5 ( .A(n7), .ZN(Co) );
endmodule


module FA_613 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  AOI22_X1 U4 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
  INV_X1 U5 ( .A(n7), .ZN(Co) );
endmodule


module FA_612 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_611 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_610 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_609 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_608 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_607 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_606 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_605 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_604 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_603 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_602 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_601 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_600 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_599 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_598 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_597 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_596 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_595 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  AOI22_X1 U4 ( .A1(B), .A2(A), .B1(Ci), .B2(n6), .ZN(n7) );
  INV_X1 U5 ( .A(n7), .ZN(Co) );
endmodule


module FA_594 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_593 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_592 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_591 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_590 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_589 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_588 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_587 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_586 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_585 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_584 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_583 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_582 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_581 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_580 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_579 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_578 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_577 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N64_10 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Ci;
  output Co;

  wire   [63:1] CTMP;
  tri   [63:0] A;

  FA_640 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_639 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_638 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_637 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(CTMP[4]) );
  FA_636 FAI_5 ( .A(A[4]), .B(B[4]), .Ci(CTMP[4]), .S(S[4]), .Co(CTMP[5]) );
  FA_635 FAI_6 ( .A(A[5]), .B(B[5]), .Ci(CTMP[5]), .S(S[5]), .Co(CTMP[6]) );
  FA_634 FAI_7 ( .A(A[6]), .B(B[6]), .Ci(CTMP[6]), .S(S[6]), .Co(CTMP[7]) );
  FA_633 FAI_8 ( .A(A[7]), .B(B[7]), .Ci(CTMP[7]), .S(S[7]), .Co(CTMP[8]) );
  FA_632 FAI_9 ( .A(A[8]), .B(B[8]), .Ci(CTMP[8]), .S(S[8]), .Co(CTMP[9]) );
  FA_631 FAI_10 ( .A(A[9]), .B(B[9]), .Ci(CTMP[9]), .S(S[9]), .Co(CTMP[10]) );
  FA_630 FAI_11 ( .A(A[10]), .B(B[10]), .Ci(CTMP[10]), .S(S[10]), .Co(CTMP[11]) );
  FA_629 FAI_12 ( .A(A[11]), .B(B[11]), .Ci(CTMP[11]), .S(S[11]), .Co(CTMP[12]) );
  FA_628 FAI_13 ( .A(A[12]), .B(B[12]), .Ci(CTMP[12]), .S(S[12]), .Co(CTMP[13]) );
  FA_627 FAI_14 ( .A(A[13]), .B(B[13]), .Ci(CTMP[13]), .S(S[13]), .Co(CTMP[14]) );
  FA_626 FAI_15 ( .A(A[14]), .B(B[14]), .Ci(CTMP[14]), .S(S[14]), .Co(CTMP[15]) );
  FA_625 FAI_16 ( .A(A[15]), .B(B[15]), .Ci(CTMP[15]), .S(S[15]), .Co(CTMP[16]) );
  FA_624 FAI_17 ( .A(A[16]), .B(B[16]), .Ci(CTMP[16]), .S(S[16]), .Co(CTMP[17]) );
  FA_623 FAI_18 ( .A(A[17]), .B(B[17]), .Ci(CTMP[17]), .S(S[17]), .Co(CTMP[18]) );
  FA_622 FAI_19 ( .A(A[18]), .B(B[18]), .Ci(CTMP[18]), .S(S[18]), .Co(CTMP[19]) );
  FA_621 FAI_20 ( .A(A[19]), .B(B[19]), .Ci(CTMP[19]), .S(S[19]), .Co(CTMP[20]) );
  FA_620 FAI_21 ( .A(A[20]), .B(B[20]), .Ci(CTMP[20]), .S(S[20]), .Co(CTMP[21]) );
  FA_619 FAI_22 ( .A(A[21]), .B(B[21]), .Ci(CTMP[21]), .S(S[21]), .Co(CTMP[22]) );
  FA_618 FAI_23 ( .A(A[22]), .B(B[22]), .Ci(CTMP[22]), .S(S[22]), .Co(CTMP[23]) );
  FA_617 FAI_24 ( .A(A[23]), .B(B[23]), .Ci(CTMP[23]), .S(S[23]), .Co(CTMP[24]) );
  FA_616 FAI_25 ( .A(A[24]), .B(B[24]), .Ci(CTMP[24]), .S(S[24]), .Co(CTMP[25]) );
  FA_615 FAI_26 ( .A(A[25]), .B(B[25]), .Ci(CTMP[25]), .S(S[25]), .Co(CTMP[26]) );
  FA_614 FAI_27 ( .A(A[26]), .B(B[26]), .Ci(CTMP[26]), .S(S[26]), .Co(CTMP[27]) );
  FA_613 FAI_28 ( .A(A[27]), .B(B[27]), .Ci(CTMP[27]), .S(S[27]), .Co(CTMP[28]) );
  FA_612 FAI_29 ( .A(A[28]), .B(B[28]), .Ci(CTMP[28]), .S(S[28]), .Co(CTMP[29]) );
  FA_611 FAI_30 ( .A(A[29]), .B(B[29]), .Ci(CTMP[29]), .S(S[29]), .Co(CTMP[30]) );
  FA_610 FAI_31 ( .A(A[30]), .B(B[30]), .Ci(CTMP[30]), .S(S[30]), .Co(CTMP[31]) );
  FA_609 FAI_32 ( .A(A[31]), .B(B[31]), .Ci(CTMP[31]), .S(S[31]), .Co(CTMP[32]) );
  FA_608 FAI_33 ( .A(A[32]), .B(B[32]), .Ci(CTMP[32]), .S(S[32]), .Co(CTMP[33]) );
  FA_607 FAI_34 ( .A(A[33]), .B(B[33]), .Ci(CTMP[33]), .S(S[33]), .Co(CTMP[34]) );
  FA_606 FAI_35 ( .A(A[34]), .B(B[34]), .Ci(CTMP[34]), .S(S[34]), .Co(CTMP[35]) );
  FA_605 FAI_36 ( .A(A[35]), .B(B[35]), .Ci(CTMP[35]), .S(S[35]), .Co(CTMP[36]) );
  FA_604 FAI_37 ( .A(A[36]), .B(B[36]), .Ci(CTMP[36]), .S(S[36]), .Co(CTMP[37]) );
  FA_603 FAI_38 ( .A(A[37]), .B(B[37]), .Ci(CTMP[37]), .S(S[37]), .Co(CTMP[38]) );
  FA_602 FAI_39 ( .A(A[38]), .B(B[38]), .Ci(CTMP[38]), .S(S[38]), .Co(CTMP[39]) );
  FA_601 FAI_40 ( .A(A[39]), .B(B[39]), .Ci(CTMP[39]), .S(S[39]), .Co(CTMP[40]) );
  FA_600 FAI_41 ( .A(A[40]), .B(B[40]), .Ci(CTMP[40]), .S(S[40]), .Co(CTMP[41]) );
  FA_599 FAI_42 ( .A(A[41]), .B(B[41]), .Ci(CTMP[41]), .S(S[41]), .Co(CTMP[42]) );
  FA_598 FAI_43 ( .A(A[42]), .B(B[42]), .Ci(CTMP[42]), .S(S[42]), .Co(CTMP[43]) );
  FA_597 FAI_44 ( .A(A[43]), .B(B[43]), .Ci(CTMP[43]), .S(S[43]), .Co(CTMP[44]) );
  FA_596 FAI_45 ( .A(A[44]), .B(B[44]), .Ci(CTMP[44]), .S(S[44]), .Co(CTMP[45]) );
  FA_595 FAI_46 ( .A(A[45]), .B(B[45]), .Ci(CTMP[45]), .S(S[45]), .Co(CTMP[46]) );
  FA_594 FAI_47 ( .A(A[46]), .B(B[46]), .Ci(CTMP[46]), .S(S[46]), .Co(CTMP[47]) );
  FA_593 FAI_48 ( .A(A[47]), .B(B[47]), .Ci(CTMP[47]), .S(S[47]), .Co(CTMP[48]) );
  FA_592 FAI_49 ( .A(A[48]), .B(B[48]), .Ci(CTMP[48]), .S(S[48]), .Co(CTMP[49]) );
  FA_591 FAI_50 ( .A(A[49]), .B(B[49]), .Ci(CTMP[49]), .S(S[49]), .Co(CTMP[50]) );
  FA_590 FAI_51 ( .A(A[50]), .B(B[50]), .Ci(CTMP[50]), .S(S[50]), .Co(CTMP[51]) );
  FA_589 FAI_52 ( .A(A[51]), .B(B[51]), .Ci(CTMP[51]), .S(S[51]), .Co(CTMP[52]) );
  FA_588 FAI_53 ( .A(A[52]), .B(B[52]), .Ci(CTMP[52]), .S(S[52]), .Co(CTMP[53]) );
  FA_587 FAI_54 ( .A(A[53]), .B(B[53]), .Ci(CTMP[53]), .S(S[53]), .Co(CTMP[54]) );
  FA_586 FAI_55 ( .A(A[54]), .B(B[54]), .Ci(CTMP[54]), .S(S[54]), .Co(CTMP[55]) );
  FA_585 FAI_56 ( .A(A[55]), .B(B[55]), .Ci(CTMP[55]), .S(S[55]), .Co(CTMP[56]) );
  FA_584 FAI_57 ( .A(A[56]), .B(B[56]), .Ci(CTMP[56]), .S(S[56]), .Co(CTMP[57]) );
  FA_583 FAI_58 ( .A(A[57]), .B(B[57]), .Ci(CTMP[57]), .S(S[57]), .Co(CTMP[58]) );
  FA_582 FAI_59 ( .A(A[58]), .B(B[58]), .Ci(CTMP[58]), .S(S[58]), .Co(CTMP[59]) );
  FA_581 FAI_60 ( .A(A[59]), .B(B[59]), .Ci(CTMP[59]), .S(S[59]), .Co(CTMP[60]) );
  FA_580 FAI_61 ( .A(A[60]), .B(B[60]), .Ci(CTMP[60]), .S(S[60]), .Co(CTMP[61]) );
  FA_579 FAI_62 ( .A(A[61]), .B(B[61]), .Ci(CTMP[61]), .S(S[61]), .Co(CTMP[62]) );
  FA_578 FAI_63 ( .A(A[62]), .B(B[62]), .Ci(CTMP[62]), .S(S[62]), .Co(CTMP[63]) );
  FA_577 FAI_64 ( .A(A[63]), .B(B[63]), .Ci(CTMP[63]), .S(S[63]), .Co(Co) );
endmodule


module booth_mul_row_N64_RADIX3_10 ( prevA, prevSum, encoderIn, nextA, nextSum
 );
  input [63:0] prevA;
  input [63:0] prevSum;
  input [2:0] encoderIn;
  output [63:0] nextA;
  output [63:0] nextSum;
  wire   n3;
  wire   [2:0] encoder_to_mux;
  wire   [63:0] plus2A_s;
  wire   [63:0] minus2A_s;
  wire   [63:0] minus4A_s;
  tri   [63:0] mux_to_adder;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign nextA[51] = n3;
  assign nextA[0] = 1'b0;

  encoder_N64_RADIX3_10 encoder_1 ( .X(encoderIn), .Z(encoder_to_mux) );
  ShiftnCompl_N64_10 ShiftnCompl_1 ( .plusA(prevA), .plus2A_out({
        plus2A_s[63:1], SYNOPSYS_UNCONNECTED__0}), .minus2A_out(minus2A_s), 
        .plus4A_out({nextA[63:52], n3, nextA[50:1], SYNOPSYS_UNCONNECTED__1}), 
        .minus4A_out(minus4A_s) );
  MUX_GENERIC_N64_RADIX3_10 mux_1 ( .plusA({plus2A_s[63:1], 1'b0}), .minusA(
        minus2A_s), .plus2A({nextA[63:52], n3, nextA[50:1], 1'b0}), .minus2A(
        minus4A_s), .SEL(encoder_to_mux), .Y(mux_to_adder) );
  RCA_N64_10 rca_1 ( .A(mux_to_adder), .B(prevSum), .Ci(1'b0), .S(nextSum) );
endmodule


module encoder_N64_RADIX3_9 ( X, Z );
  input [2:0] X;
  output [2:0] Z;
  wire   n5, n7, n8;

  OAI22_X1 U1 ( .A1(n8), .A2(n5), .B1(X[2]), .B2(n7), .ZN(Z[1]) );
  INV_X1 U2 ( .A(X[2]), .ZN(n5) );
  AOI21_X1 U3 ( .B1(n8), .B2(n7), .A(X[2]), .ZN(Z[0]) );
  OAI21_X1 U4 ( .B1(X[1]), .B2(X[0]), .A(n7), .ZN(n8) );
  AND3_X1 U5 ( .A1(X[2]), .A2(n7), .A3(n8), .ZN(Z[2]) );
  NAND2_X1 U6 ( .A1(X[1]), .A2(X[0]), .ZN(n7) );
endmodule


module shifter_N64_18 ( \input , shiftLeftOnePos );
  input [63:0] \input ;
  output [63:0] shiftLeftOnePos;
  wire   \input[62] , \input[61] , \input[60] , \input[59] , \input[58] ,
         \input[57] , \input[56] , \input[55] , \input[54] , \input[53] ,
         \input[52] , \input[51] , \input[50] , \input[49] , \input[48] ,
         \input[47] , \input[46] , \input[45] , \input[44] , \input[43] ,
         \input[42] , \input[41] , \input[40] , \input[39] , \input[38] ,
         \input[37] , \input[36] , \input[35] , \input[34] , \input[33] ,
         \input[32] , \input[31] , \input[30] , \input[29] , \input[28] ,
         \input[27] , \input[26] , \input[25] , \input[24] , \input[23] ,
         \input[22] , \input[21] , \input[20] , \input[19] , \input[18] ,
         \input[17] , \input[16] , \input[15] , \input[14] , \input[13] ,
         \input[12] , \input[11] , \input[10] , \input[9] , \input[8] ,
         \input[7] , \input[6] , \input[5] , \input[4] , \input[3] ,
         \input[2] , \input[1] , \input[0] ;
  assign shiftLeftOnePos[0] = 1'b0;
  assign shiftLeftOnePos[63] = \input[62] ;
  assign \input[62]  = \input  [62];
  assign shiftLeftOnePos[62] = \input[61] ;
  assign \input[61]  = \input  [61];
  assign shiftLeftOnePos[61] = \input[60] ;
  assign \input[60]  = \input  [60];
  assign shiftLeftOnePos[60] = \input[59] ;
  assign \input[59]  = \input  [59];
  assign shiftLeftOnePos[59] = \input[58] ;
  assign \input[58]  = \input  [58];
  assign shiftLeftOnePos[58] = \input[57] ;
  assign \input[57]  = \input  [57];
  assign shiftLeftOnePos[57] = \input[56] ;
  assign \input[56]  = \input  [56];
  assign shiftLeftOnePos[56] = \input[55] ;
  assign \input[55]  = \input  [55];
  assign shiftLeftOnePos[55] = \input[54] ;
  assign \input[54]  = \input  [54];
  assign shiftLeftOnePos[54] = \input[53] ;
  assign \input[53]  = \input  [53];
  assign shiftLeftOnePos[53] = \input[52] ;
  assign \input[52]  = \input  [52];
  assign shiftLeftOnePos[52] = \input[51] ;
  assign \input[51]  = \input  [51];
  assign shiftLeftOnePos[51] = \input[50] ;
  assign \input[50]  = \input  [50];
  assign shiftLeftOnePos[50] = \input[49] ;
  assign \input[49]  = \input  [49];
  assign shiftLeftOnePos[49] = \input[48] ;
  assign \input[48]  = \input  [48];
  assign shiftLeftOnePos[48] = \input[47] ;
  assign \input[47]  = \input  [47];
  assign shiftLeftOnePos[47] = \input[46] ;
  assign \input[46]  = \input  [46];
  assign shiftLeftOnePos[46] = \input[45] ;
  assign \input[45]  = \input  [45];
  assign shiftLeftOnePos[45] = \input[44] ;
  assign \input[44]  = \input  [44];
  assign shiftLeftOnePos[44] = \input[43] ;
  assign \input[43]  = \input  [43];
  assign shiftLeftOnePos[43] = \input[42] ;
  assign \input[42]  = \input  [42];
  assign shiftLeftOnePos[42] = \input[41] ;
  assign \input[41]  = \input  [41];
  assign shiftLeftOnePos[41] = \input[40] ;
  assign \input[40]  = \input  [40];
  assign shiftLeftOnePos[40] = \input[39] ;
  assign \input[39]  = \input  [39];
  assign shiftLeftOnePos[39] = \input[38] ;
  assign \input[38]  = \input  [38];
  assign shiftLeftOnePos[38] = \input[37] ;
  assign \input[37]  = \input  [37];
  assign shiftLeftOnePos[37] = \input[36] ;
  assign \input[36]  = \input  [36];
  assign shiftLeftOnePos[36] = \input[35] ;
  assign \input[35]  = \input  [35];
  assign shiftLeftOnePos[35] = \input[34] ;
  assign \input[34]  = \input  [34];
  assign shiftLeftOnePos[34] = \input[33] ;
  assign \input[33]  = \input  [33];
  assign shiftLeftOnePos[33] = \input[32] ;
  assign \input[32]  = \input  [32];
  assign shiftLeftOnePos[32] = \input[31] ;
  assign \input[31]  = \input  [31];
  assign shiftLeftOnePos[31] = \input[30] ;
  assign \input[30]  = \input  [30];
  assign shiftLeftOnePos[30] = \input[29] ;
  assign \input[29]  = \input  [29];
  assign shiftLeftOnePos[29] = \input[28] ;
  assign \input[28]  = \input  [28];
  assign shiftLeftOnePos[28] = \input[27] ;
  assign \input[27]  = \input  [27];
  assign shiftLeftOnePos[27] = \input[26] ;
  assign \input[26]  = \input  [26];
  assign shiftLeftOnePos[26] = \input[25] ;
  assign \input[25]  = \input  [25];
  assign shiftLeftOnePos[25] = \input[24] ;
  assign \input[24]  = \input  [24];
  assign shiftLeftOnePos[24] = \input[23] ;
  assign \input[23]  = \input  [23];
  assign shiftLeftOnePos[23] = \input[22] ;
  assign \input[22]  = \input  [22];
  assign shiftLeftOnePos[22] = \input[21] ;
  assign \input[21]  = \input  [21];
  assign shiftLeftOnePos[21] = \input[20] ;
  assign \input[20]  = \input  [20];
  assign shiftLeftOnePos[20] = \input[19] ;
  assign \input[19]  = \input  [19];
  assign shiftLeftOnePos[19] = \input[18] ;
  assign \input[18]  = \input  [18];
  assign shiftLeftOnePos[18] = \input[17] ;
  assign \input[17]  = \input  [17];
  assign shiftLeftOnePos[17] = \input[16] ;
  assign \input[16]  = \input  [16];
  assign shiftLeftOnePos[16] = \input[15] ;
  assign \input[15]  = \input  [15];
  assign shiftLeftOnePos[15] = \input[14] ;
  assign \input[14]  = \input  [14];
  assign shiftLeftOnePos[14] = \input[13] ;
  assign \input[13]  = \input  [13];
  assign shiftLeftOnePos[13] = \input[12] ;
  assign \input[12]  = \input  [12];
  assign shiftLeftOnePos[12] = \input[11] ;
  assign \input[11]  = \input  [11];
  assign shiftLeftOnePos[11] = \input[10] ;
  assign \input[10]  = \input  [10];
  assign shiftLeftOnePos[10] = \input[9] ;
  assign \input[9]  = \input  [9];
  assign shiftLeftOnePos[9] = \input[8] ;
  assign \input[8]  = \input  [8];
  assign shiftLeftOnePos[8] = \input[7] ;
  assign \input[7]  = \input  [7];
  assign shiftLeftOnePos[7] = \input[6] ;
  assign \input[6]  = \input  [6];
  assign shiftLeftOnePos[6] = \input[5] ;
  assign \input[5]  = \input  [5];
  assign shiftLeftOnePos[5] = \input[4] ;
  assign \input[4]  = \input  [4];
  assign shiftLeftOnePos[4] = \input[3] ;
  assign \input[3]  = \input  [3];
  assign shiftLeftOnePos[3] = \input[2] ;
  assign \input[2]  = \input  [2];
  assign shiftLeftOnePos[2] = \input[1] ;
  assign \input[1]  = \input  [1];
  assign shiftLeftOnePos[1] = \input[0] ;
  assign \input[0]  = \input  [0];

endmodule


module shifter_N64_17 ( \input , shiftLeftOnePos );
  input [63:0] \input ;
  output [63:0] shiftLeftOnePos;
  wire   \input[62] , \input[61] , \input[60] , \input[59] , \input[58] ,
         \input[57] , \input[56] , \input[55] , \input[54] , \input[53] ,
         \input[52] , \input[51] , \input[50] , \input[49] , \input[48] ,
         \input[47] , \input[46] , \input[45] , \input[44] , \input[43] ,
         \input[42] , \input[41] , \input[40] , \input[39] , \input[38] ,
         \input[37] , \input[36] , \input[35] , \input[34] , \input[33] ,
         \input[32] , \input[31] , \input[30] , \input[29] , \input[28] ,
         \input[27] , \input[26] , \input[25] , \input[24] , \input[23] ,
         \input[22] , \input[21] , \input[20] , \input[19] , \input[18] ,
         \input[17] , \input[16] , \input[15] , \input[14] , \input[13] ,
         \input[12] , \input[11] , \input[10] , \input[9] , \input[8] ,
         \input[7] , \input[6] , \input[5] , \input[4] , \input[3] ,
         \input[2] , \input[1] , \input[0] ;
  assign shiftLeftOnePos[0] = 1'b0;
  assign shiftLeftOnePos[63] = \input[62] ;
  assign \input[62]  = \input  [62];
  assign shiftLeftOnePos[62] = \input[61] ;
  assign \input[61]  = \input  [61];
  assign shiftLeftOnePos[61] = \input[60] ;
  assign \input[60]  = \input  [60];
  assign shiftLeftOnePos[60] = \input[59] ;
  assign \input[59]  = \input  [59];
  assign shiftLeftOnePos[59] = \input[58] ;
  assign \input[58]  = \input  [58];
  assign shiftLeftOnePos[58] = \input[57] ;
  assign \input[57]  = \input  [57];
  assign shiftLeftOnePos[57] = \input[56] ;
  assign \input[56]  = \input  [56];
  assign shiftLeftOnePos[56] = \input[55] ;
  assign \input[55]  = \input  [55];
  assign shiftLeftOnePos[55] = \input[54] ;
  assign \input[54]  = \input  [54];
  assign shiftLeftOnePos[54] = \input[53] ;
  assign \input[53]  = \input  [53];
  assign shiftLeftOnePos[53] = \input[52] ;
  assign \input[52]  = \input  [52];
  assign shiftLeftOnePos[52] = \input[51] ;
  assign \input[51]  = \input  [51];
  assign shiftLeftOnePos[51] = \input[50] ;
  assign \input[50]  = \input  [50];
  assign shiftLeftOnePos[50] = \input[49] ;
  assign \input[49]  = \input  [49];
  assign shiftLeftOnePos[49] = \input[48] ;
  assign \input[48]  = \input  [48];
  assign shiftLeftOnePos[48] = \input[47] ;
  assign \input[47]  = \input  [47];
  assign shiftLeftOnePos[47] = \input[46] ;
  assign \input[46]  = \input  [46];
  assign shiftLeftOnePos[46] = \input[45] ;
  assign \input[45]  = \input  [45];
  assign shiftLeftOnePos[45] = \input[44] ;
  assign \input[44]  = \input  [44];
  assign shiftLeftOnePos[44] = \input[43] ;
  assign \input[43]  = \input  [43];
  assign shiftLeftOnePos[43] = \input[42] ;
  assign \input[42]  = \input  [42];
  assign shiftLeftOnePos[42] = \input[41] ;
  assign \input[41]  = \input  [41];
  assign shiftLeftOnePos[41] = \input[40] ;
  assign \input[40]  = \input  [40];
  assign shiftLeftOnePos[40] = \input[39] ;
  assign \input[39]  = \input  [39];
  assign shiftLeftOnePos[39] = \input[38] ;
  assign \input[38]  = \input  [38];
  assign shiftLeftOnePos[38] = \input[37] ;
  assign \input[37]  = \input  [37];
  assign shiftLeftOnePos[37] = \input[36] ;
  assign \input[36]  = \input  [36];
  assign shiftLeftOnePos[36] = \input[35] ;
  assign \input[35]  = \input  [35];
  assign shiftLeftOnePos[35] = \input[34] ;
  assign \input[34]  = \input  [34];
  assign shiftLeftOnePos[34] = \input[33] ;
  assign \input[33]  = \input  [33];
  assign shiftLeftOnePos[33] = \input[32] ;
  assign \input[32]  = \input  [32];
  assign shiftLeftOnePos[32] = \input[31] ;
  assign \input[31]  = \input  [31];
  assign shiftLeftOnePos[31] = \input[30] ;
  assign \input[30]  = \input  [30];
  assign shiftLeftOnePos[30] = \input[29] ;
  assign \input[29]  = \input  [29];
  assign shiftLeftOnePos[29] = \input[28] ;
  assign \input[28]  = \input  [28];
  assign shiftLeftOnePos[28] = \input[27] ;
  assign \input[27]  = \input  [27];
  assign shiftLeftOnePos[27] = \input[26] ;
  assign \input[26]  = \input  [26];
  assign shiftLeftOnePos[26] = \input[25] ;
  assign \input[25]  = \input  [25];
  assign shiftLeftOnePos[25] = \input[24] ;
  assign \input[24]  = \input  [24];
  assign shiftLeftOnePos[24] = \input[23] ;
  assign \input[23]  = \input  [23];
  assign shiftLeftOnePos[23] = \input[22] ;
  assign \input[22]  = \input  [22];
  assign shiftLeftOnePos[22] = \input[21] ;
  assign \input[21]  = \input  [21];
  assign shiftLeftOnePos[21] = \input[20] ;
  assign \input[20]  = \input  [20];
  assign shiftLeftOnePos[20] = \input[19] ;
  assign \input[19]  = \input  [19];
  assign shiftLeftOnePos[19] = \input[18] ;
  assign \input[18]  = \input  [18];
  assign shiftLeftOnePos[18] = \input[17] ;
  assign \input[17]  = \input  [17];
  assign shiftLeftOnePos[17] = \input[16] ;
  assign \input[16]  = \input  [16];
  assign shiftLeftOnePos[16] = \input[15] ;
  assign \input[15]  = \input  [15];
  assign shiftLeftOnePos[15] = \input[14] ;
  assign \input[14]  = \input  [14];
  assign shiftLeftOnePos[14] = \input[13] ;
  assign \input[13]  = \input  [13];
  assign shiftLeftOnePos[13] = \input[12] ;
  assign \input[12]  = \input  [12];
  assign shiftLeftOnePos[12] = \input[11] ;
  assign \input[11]  = \input  [11];
  assign shiftLeftOnePos[11] = \input[10] ;
  assign \input[10]  = \input  [10];
  assign shiftLeftOnePos[10] = \input[9] ;
  assign \input[9]  = \input  [9];
  assign shiftLeftOnePos[9] = \input[8] ;
  assign \input[8]  = \input  [8];
  assign shiftLeftOnePos[8] = \input[7] ;
  assign \input[7]  = \input  [7];
  assign shiftLeftOnePos[7] = \input[6] ;
  assign \input[6]  = \input  [6];
  assign shiftLeftOnePos[6] = \input[5] ;
  assign \input[5]  = \input  [5];
  assign shiftLeftOnePos[5] = \input[4] ;
  assign \input[4]  = \input  [4];
  assign shiftLeftOnePos[4] = \input[3] ;
  assign \input[3]  = \input  [3];
  assign shiftLeftOnePos[3] = \input[2] ;
  assign \input[2]  = \input  [2];
  assign shiftLeftOnePos[2] = \input[1] ;
  assign \input[1]  = \input  [1];
  assign shiftLeftOnePos[1] = \input[0] ;
  assign \input[0]  = \input  [0];

endmodule


module complementer_N64_18_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n190, n191, n192, n193, n194, n196, n197, n198, n199, n200,
         n202, n203, n204, n206, n207, n208, n210, n211, n212, n213, n214,
         n216, n217, n218, n220, n221, n222, n224, n225, n226, n228, n229,
         n230, n232, n233, n234, n235, n237, n238, n239, n241, n242, n243,
         n245, n246, n247, n249, n250, n251, n189, n195, n201, n205, n209,
         n215, n219, n223, n227, n231, n236, n240, n244, n248;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U81 ( .A(n190), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U82 ( .A(n192), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U83 ( .A(n193), .B(B[6]), .Z(DIFF[6]) );
  XOR2_X1 U85 ( .A(n196), .B(B[62]), .Z(DIFF[62]) );
  XOR2_X1 U86 ( .A(n194), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U87 ( .A(n198), .B(B[59]), .Z(DIFF[59]) );
  XOR2_X1 U89 ( .A(n200), .B(B[57]), .Z(DIFF[57]) );
  XOR2_X1 U90 ( .A(n202), .B(B[55]), .Z(DIFF[55]) );
  XOR2_X1 U92 ( .A(n204), .B(B[53]), .Z(DIFF[53]) );
  XOR2_X1 U93 ( .A(n206), .B(B[51]), .Z(DIFF[51]) );
  XOR2_X1 U95 ( .A(n208), .B(B[49]), .Z(DIFF[49]) );
  XOR2_X1 U96 ( .A(n212), .B(B[47]), .Z(DIFF[47]) );
  XOR2_X1 U98 ( .A(n214), .B(B[45]), .Z(DIFF[45]) );
  XOR2_X1 U99 ( .A(n216), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U101 ( .A(n218), .B(B[41]), .Z(DIFF[41]) );
  XOR2_X1 U102 ( .A(n211), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U103 ( .A(n220), .B(B[39]), .Z(DIFF[39]) );
  XOR2_X1 U105 ( .A(n222), .B(B[37]), .Z(DIFF[37]) );
  XOR2_X1 U106 ( .A(n224), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U108 ( .A(n226), .B(B[33]), .Z(DIFF[33]) );
  XOR2_X1 U109 ( .A(n228), .B(B[31]), .Z(DIFF[31]) );
  XOR2_X1 U111 ( .A(n230), .B(B[29]), .Z(DIFF[29]) );
  XOR2_X1 U112 ( .A(n233), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U114 ( .A(n235), .B(B[25]), .Z(DIFF[25]) );
  XOR2_X1 U115 ( .A(n237), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U117 ( .A(n239), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U118 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U119 ( .A(n241), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U121 ( .A(n243), .B(B[17]), .Z(DIFF[17]) );
  XOR2_X1 U122 ( .A(n245), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U124 ( .A(n247), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U125 ( .A(n249), .B(B[11]), .Z(DIFF[11]) );
  XOR2_X1 U126 ( .A(n251), .B(B[10]), .Z(DIFF[10]) );
  XOR2_X1 U1 ( .A(n197), .B(n248), .Z(DIFF[61]) );
  NAND2_X1 U2 ( .A1(n197), .A2(n248), .ZN(n196) );
  NOR3_X1 U3 ( .A1(B[59]), .A2(B[60]), .A3(n198), .ZN(n197) );
  XNOR2_X1 U4 ( .A(B[56]), .B(n203), .ZN(DIFF[56]) );
  NOR2_X1 U5 ( .A1(B[55]), .A2(n202), .ZN(n203) );
  XNOR2_X1 U6 ( .A(B[52]), .B(n207), .ZN(DIFF[52]) );
  NOR2_X1 U7 ( .A1(B[51]), .A2(n206), .ZN(n207) );
  XNOR2_X1 U8 ( .A(B[48]), .B(n213), .ZN(DIFF[48]) );
  NOR2_X1 U9 ( .A1(B[47]), .A2(n212), .ZN(n213) );
  XNOR2_X1 U10 ( .A(B[60]), .B(n199), .ZN(DIFF[60]) );
  NOR2_X1 U11 ( .A1(B[59]), .A2(n198), .ZN(n199) );
  OR3_X1 U12 ( .A1(B[57]), .A2(B[58]), .A3(n200), .ZN(n198) );
  OR3_X1 U13 ( .A1(B[53]), .A2(B[54]), .A3(n204), .ZN(n202) );
  OR3_X1 U14 ( .A1(B[49]), .A2(B[50]), .A3(n208), .ZN(n206) );
  OR3_X1 U15 ( .A1(B[47]), .A2(B[48]), .A3(n212), .ZN(n208) );
  OR3_X1 U16 ( .A1(B[55]), .A2(B[56]), .A3(n202), .ZN(n200) );
  OR3_X1 U17 ( .A1(B[51]), .A2(B[52]), .A3(n206), .ZN(n204) );
  XNOR2_X1 U18 ( .A(n189), .B(B[58]), .ZN(DIFF[58]) );
  NOR2_X1 U19 ( .A1(n200), .A2(B[57]), .ZN(n189) );
  XNOR2_X1 U20 ( .A(n195), .B(B[54]), .ZN(DIFF[54]) );
  NOR2_X1 U21 ( .A1(n204), .A2(B[53]), .ZN(n195) );
  XNOR2_X1 U22 ( .A(n201), .B(B[50]), .ZN(DIFF[50]) );
  NOR2_X1 U23 ( .A1(n208), .A2(B[49]), .ZN(n201) );
  XNOR2_X1 U24 ( .A(n205), .B(B[63]), .ZN(DIFF[63]) );
  NOR2_X1 U25 ( .A1(n196), .A2(B[62]), .ZN(n205) );
  OR3_X1 U26 ( .A1(B[45]), .A2(B[46]), .A3(n214), .ZN(n212) );
  XNOR2_X1 U27 ( .A(n209), .B(B[46]), .ZN(DIFF[46]) );
  NOR2_X1 U28 ( .A1(n214), .A2(B[45]), .ZN(n209) );
  XNOR2_X1 U29 ( .A(B[36]), .B(n225), .ZN(DIFF[36]) );
  NOR2_X1 U30 ( .A1(B[35]), .A2(n224), .ZN(n225) );
  XNOR2_X1 U31 ( .A(B[32]), .B(n229), .ZN(DIFF[32]) );
  NOR2_X1 U32 ( .A1(B[31]), .A2(n228), .ZN(n229) );
  XNOR2_X1 U33 ( .A(B[28]), .B(n234), .ZN(DIFF[28]) );
  NOR2_X1 U34 ( .A1(B[27]), .A2(n233), .ZN(n234) );
  XNOR2_X1 U35 ( .A(B[24]), .B(n238), .ZN(DIFF[24]) );
  NOR2_X1 U36 ( .A1(B[23]), .A2(n237), .ZN(n238) );
  XNOR2_X1 U37 ( .A(B[20]), .B(n242), .ZN(DIFF[20]) );
  NOR2_X1 U38 ( .A1(B[19]), .A2(n241), .ZN(n242) );
  OR3_X1 U39 ( .A1(B[21]), .A2(B[22]), .A3(n239), .ZN(n237) );
  OR3_X1 U40 ( .A1(B[25]), .A2(B[26]), .A3(n235), .ZN(n233) );
  OR3_X1 U41 ( .A1(B[29]), .A2(B[30]), .A3(n230), .ZN(n228) );
  OR3_X1 U42 ( .A1(B[33]), .A2(B[34]), .A3(n226), .ZN(n224) );
  OR3_X1 U43 ( .A1(B[19]), .A2(B[20]), .A3(n241), .ZN(n239) );
  OR3_X1 U44 ( .A1(B[23]), .A2(B[24]), .A3(n237), .ZN(n235) );
  OR3_X1 U45 ( .A1(B[27]), .A2(B[28]), .A3(n233), .ZN(n230) );
  OR3_X1 U46 ( .A1(B[31]), .A2(B[32]), .A3(n228), .ZN(n226) );
  OR3_X1 U47 ( .A1(B[35]), .A2(B[36]), .A3(n224), .ZN(n222) );
  XNOR2_X1 U48 ( .A(n215), .B(B[34]), .ZN(DIFF[34]) );
  NOR2_X1 U49 ( .A1(n226), .A2(B[33]), .ZN(n215) );
  XNOR2_X1 U50 ( .A(n219), .B(B[30]), .ZN(DIFF[30]) );
  NOR2_X1 U51 ( .A1(n230), .A2(B[29]), .ZN(n219) );
  XNOR2_X1 U52 ( .A(n223), .B(B[26]), .ZN(DIFF[26]) );
  NOR2_X1 U53 ( .A1(n235), .A2(B[25]), .ZN(n223) );
  XNOR2_X1 U54 ( .A(n227), .B(B[22]), .ZN(DIFF[22]) );
  NOR2_X1 U55 ( .A1(n239), .A2(B[21]), .ZN(n227) );
  XNOR2_X1 U56 ( .A(B[44]), .B(n217), .ZN(DIFF[44]) );
  NOR2_X1 U57 ( .A1(B[43]), .A2(n216), .ZN(n217) );
  XNOR2_X1 U58 ( .A(B[40]), .B(n221), .ZN(DIFF[40]) );
  NOR2_X1 U59 ( .A1(B[39]), .A2(n220), .ZN(n221) );
  OR3_X1 U60 ( .A1(B[37]), .A2(B[38]), .A3(n222), .ZN(n220) );
  OR3_X1 U61 ( .A1(B[41]), .A2(B[42]), .A3(n218), .ZN(n216) );
  OR3_X1 U62 ( .A1(B[39]), .A2(B[40]), .A3(n220), .ZN(n218) );
  OR3_X1 U63 ( .A1(B[43]), .A2(B[44]), .A3(n216), .ZN(n214) );
  XNOR2_X1 U64 ( .A(n231), .B(B[42]), .ZN(DIFF[42]) );
  NOR2_X1 U65 ( .A1(n218), .A2(B[41]), .ZN(n231) );
  XNOR2_X1 U66 ( .A(n236), .B(B[38]), .ZN(DIFF[38]) );
  NOR2_X1 U67 ( .A1(n222), .A2(B[37]), .ZN(n236) );
  OR3_X1 U68 ( .A1(B[17]), .A2(B[18]), .A3(n243), .ZN(n241) );
  XNOR2_X1 U69 ( .A(n240), .B(B[18]), .ZN(DIFF[18]) );
  NOR2_X1 U70 ( .A1(n243), .A2(B[17]), .ZN(n240) );
  OR3_X1 U71 ( .A1(B[15]), .A2(B[16]), .A3(n245), .ZN(n243) );
  XNOR2_X1 U72 ( .A(B[16]), .B(n246), .ZN(DIFF[16]) );
  NOR2_X1 U73 ( .A1(B[15]), .A2(n245), .ZN(n246) );
  OR3_X1 U74 ( .A1(B[13]), .A2(B[14]), .A3(n247), .ZN(n245) );
  XNOR2_X1 U75 ( .A(n244), .B(B[14]), .ZN(DIFF[14]) );
  NOR2_X1 U76 ( .A1(n247), .A2(B[13]), .ZN(n244) );
  NOR2_X1 U77 ( .A1(B[11]), .A2(n249), .ZN(n250) );
  NOR2_X1 U78 ( .A1(B[7]), .A2(n192), .ZN(n191) );
  NOR2_X1 U79 ( .A1(B[3]), .A2(n211), .ZN(n210) );
  OR3_X1 U80 ( .A1(B[10]), .A2(B[9]), .A3(n190), .ZN(n249) );
  OR3_X1 U84 ( .A1(B[5]), .A2(B[6]), .A3(n194), .ZN(n192) );
  OR3_X1 U88 ( .A1(B[11]), .A2(B[12]), .A3(n249), .ZN(n247) );
  OR3_X1 U91 ( .A1(B[7]), .A2(B[8]), .A3(n192), .ZN(n190) );
  OR3_X1 U94 ( .A1(B[3]), .A2(B[4]), .A3(n211), .ZN(n194) );
  XNOR2_X1 U97 ( .A(B[12]), .B(n250), .ZN(DIFF[12]) );
  XNOR2_X1 U100 ( .A(B[8]), .B(n191), .ZN(DIFF[8]) );
  XNOR2_X1 U104 ( .A(B[4]), .B(n210), .ZN(DIFF[4]) );
  XNOR2_X1 U107 ( .A(B[2]), .B(n232), .ZN(DIFF[2]) );
  OR2_X1 U110 ( .A1(n190), .A2(B[9]), .ZN(n251) );
  OR2_X1 U113 ( .A1(n194), .A2(B[5]), .ZN(n193) );
  OR3_X1 U116 ( .A1(B[1]), .A2(B[2]), .A3(\B[0] ), .ZN(n211) );
  NOR2_X1 U120 ( .A1(\B[0] ), .A2(B[1]), .ZN(n232) );
  INV_X1 U123 ( .A(B[61]), .ZN(n248) );
endmodule


module complementer_N64_18 ( \input , complement2 );
  input [63:0] \input ;
  output [63:0] complement2;


  complementer_N64_18_DW01_sub_0 sub_add_31_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(\input ), .CI(1'b0), .DIFF(complement2) );
endmodule


module complementer_N64_17_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n190, n191, n192, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n189, n193, n251;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U81 ( .A(n190), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U82 ( .A(n192), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U84 ( .A(n195), .B(B[63]), .Z(DIFF[63]) );
  XOR2_X1 U85 ( .A(n196), .B(B[62]), .Z(DIFF[62]) );
  XOR2_X1 U86 ( .A(n194), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U87 ( .A(n198), .B(B[59]), .Z(DIFF[59]) );
  XOR2_X1 U88 ( .A(n201), .B(B[58]), .Z(DIFF[58]) );
  XOR2_X1 U89 ( .A(n200), .B(B[57]), .Z(DIFF[57]) );
  XOR2_X1 U90 ( .A(n202), .B(B[55]), .Z(DIFF[55]) );
  XOR2_X1 U91 ( .A(n205), .B(B[54]), .Z(DIFF[54]) );
  XOR2_X1 U92 ( .A(n204), .B(B[53]), .Z(DIFF[53]) );
  XOR2_X1 U93 ( .A(n206), .B(B[51]), .Z(DIFF[51]) );
  XOR2_X1 U94 ( .A(n209), .B(B[50]), .Z(DIFF[50]) );
  XOR2_X1 U95 ( .A(n208), .B(B[49]), .Z(DIFF[49]) );
  XOR2_X1 U96 ( .A(n212), .B(B[47]), .Z(DIFF[47]) );
  XOR2_X1 U97 ( .A(n215), .B(B[46]), .Z(DIFF[46]) );
  XOR2_X1 U98 ( .A(n214), .B(B[45]), .Z(DIFF[45]) );
  XOR2_X1 U99 ( .A(n216), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U100 ( .A(n219), .B(B[42]), .Z(DIFF[42]) );
  XOR2_X1 U101 ( .A(n218), .B(B[41]), .Z(DIFF[41]) );
  XOR2_X1 U102 ( .A(n211), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U103 ( .A(n220), .B(B[39]), .Z(DIFF[39]) );
  XOR2_X1 U104 ( .A(n223), .B(B[38]), .Z(DIFF[38]) );
  XOR2_X1 U105 ( .A(n222), .B(B[37]), .Z(DIFF[37]) );
  XOR2_X1 U106 ( .A(n224), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U107 ( .A(n227), .B(B[34]), .Z(DIFF[34]) );
  XOR2_X1 U108 ( .A(n226), .B(B[33]), .Z(DIFF[33]) );
  XOR2_X1 U109 ( .A(n228), .B(B[31]), .Z(DIFF[31]) );
  XOR2_X1 U110 ( .A(n231), .B(B[30]), .Z(DIFF[30]) );
  XOR2_X1 U111 ( .A(n230), .B(B[29]), .Z(DIFF[29]) );
  XOR2_X1 U112 ( .A(n233), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U113 ( .A(n236), .B(B[26]), .Z(DIFF[26]) );
  XOR2_X1 U114 ( .A(n235), .B(B[25]), .Z(DIFF[25]) );
  XOR2_X1 U115 ( .A(n237), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U116 ( .A(n240), .B(B[22]), .Z(DIFF[22]) );
  XOR2_X1 U117 ( .A(n239), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U118 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U119 ( .A(n241), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U120 ( .A(n244), .B(B[18]), .Z(DIFF[18]) );
  XOR2_X1 U121 ( .A(n243), .B(B[17]), .Z(DIFF[17]) );
  XOR2_X1 U122 ( .A(n245), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U123 ( .A(n248), .B(B[14]), .Z(DIFF[14]) );
  XOR2_X1 U124 ( .A(n247), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U125 ( .A(n249), .B(B[11]), .Z(DIFF[11]) );
  OR2_X1 U1 ( .A1(n204), .A2(B[53]), .ZN(n205) );
  NAND2_X1 U2 ( .A1(n197), .A2(n251), .ZN(n196) );
  NOR2_X1 U3 ( .A1(B[55]), .A2(n202), .ZN(n203) );
  NOR2_X1 U4 ( .A1(B[51]), .A2(n206), .ZN(n207) );
  OR3_X1 U5 ( .A1(B[57]), .A2(B[58]), .A3(n200), .ZN(n198) );
  OR3_X1 U6 ( .A1(B[53]), .A2(B[54]), .A3(n204), .ZN(n202) );
  OR3_X1 U7 ( .A1(B[49]), .A2(B[50]), .A3(n208), .ZN(n206) );
  OR3_X1 U8 ( .A1(B[55]), .A2(B[56]), .A3(n202), .ZN(n200) );
  OR3_X1 U9 ( .A1(B[51]), .A2(B[52]), .A3(n206), .ZN(n204) );
  OR2_X1 U10 ( .A1(n200), .A2(B[57]), .ZN(n201) );
  OR2_X1 U11 ( .A1(n208), .A2(B[49]), .ZN(n209) );
  NOR3_X1 U12 ( .A1(B[59]), .A2(B[60]), .A3(n198), .ZN(n197) );
  NOR2_X1 U13 ( .A1(B[59]), .A2(n198), .ZN(n199) );
  OR2_X1 U14 ( .A1(n196), .A2(B[62]), .ZN(n195) );
  NOR2_X1 U15 ( .A1(B[47]), .A2(n212), .ZN(n213) );
  OR3_X1 U16 ( .A1(B[47]), .A2(B[48]), .A3(n212), .ZN(n208) );
  XNOR2_X1 U17 ( .A(B[24]), .B(n238), .ZN(DIFF[24]) );
  XNOR2_X1 U18 ( .A(B[20]), .B(n242), .ZN(DIFF[20]) );
  NOR2_X1 U19 ( .A1(B[31]), .A2(n228), .ZN(n229) );
  NOR2_X1 U20 ( .A1(B[27]), .A2(n233), .ZN(n234) );
  NOR2_X1 U21 ( .A1(B[23]), .A2(n237), .ZN(n238) );
  NOR2_X1 U22 ( .A1(B[19]), .A2(n241), .ZN(n242) );
  OR3_X1 U23 ( .A1(B[29]), .A2(B[30]), .A3(n230), .ZN(n228) );
  OR3_X1 U24 ( .A1(B[25]), .A2(B[26]), .A3(n235), .ZN(n233) );
  OR3_X1 U25 ( .A1(B[21]), .A2(B[22]), .A3(n239), .ZN(n237) );
  OR3_X1 U26 ( .A1(B[31]), .A2(B[32]), .A3(n228), .ZN(n226) );
  OR3_X1 U27 ( .A1(B[27]), .A2(B[28]), .A3(n233), .ZN(n230) );
  OR3_X1 U28 ( .A1(B[23]), .A2(B[24]), .A3(n237), .ZN(n235) );
  OR3_X1 U29 ( .A1(B[19]), .A2(B[20]), .A3(n241), .ZN(n239) );
  XNOR2_X1 U30 ( .A(B[36]), .B(n225), .ZN(DIFF[36]) );
  XNOR2_X1 U31 ( .A(B[32]), .B(n229), .ZN(DIFF[32]) );
  XNOR2_X1 U32 ( .A(B[28]), .B(n234), .ZN(DIFF[28]) );
  OR2_X1 U33 ( .A1(n226), .A2(B[33]), .ZN(n227) );
  OR2_X1 U34 ( .A1(n230), .A2(B[29]), .ZN(n231) );
  OR2_X1 U35 ( .A1(n235), .A2(B[25]), .ZN(n236) );
  OR2_X1 U36 ( .A1(n239), .A2(B[21]), .ZN(n240) );
  NOR2_X1 U37 ( .A1(B[43]), .A2(n216), .ZN(n217) );
  NOR2_X1 U38 ( .A1(B[39]), .A2(n220), .ZN(n221) );
  NOR2_X1 U39 ( .A1(B[35]), .A2(n224), .ZN(n225) );
  OR3_X1 U40 ( .A1(B[41]), .A2(B[42]), .A3(n218), .ZN(n216) );
  OR3_X1 U41 ( .A1(B[37]), .A2(B[38]), .A3(n222), .ZN(n220) );
  OR3_X1 U42 ( .A1(B[33]), .A2(B[34]), .A3(n226), .ZN(n224) );
  OR3_X1 U43 ( .A1(B[45]), .A2(B[46]), .A3(n214), .ZN(n212) );
  OR3_X1 U44 ( .A1(B[43]), .A2(B[44]), .A3(n216), .ZN(n214) );
  OR3_X1 U45 ( .A1(B[39]), .A2(B[40]), .A3(n220), .ZN(n218) );
  OR3_X1 U46 ( .A1(B[35]), .A2(B[36]), .A3(n224), .ZN(n222) );
  XNOR2_X1 U47 ( .A(B[56]), .B(n203), .ZN(DIFF[56]) );
  XNOR2_X1 U48 ( .A(B[44]), .B(n217), .ZN(DIFF[44]) );
  XNOR2_X1 U49 ( .A(B[40]), .B(n221), .ZN(DIFF[40]) );
  XNOR2_X1 U50 ( .A(B[52]), .B(n207), .ZN(DIFF[52]) );
  XNOR2_X1 U51 ( .A(B[48]), .B(n213), .ZN(DIFF[48]) );
  XNOR2_X1 U52 ( .A(n197), .B(B[61]), .ZN(DIFF[61]) );
  XNOR2_X1 U53 ( .A(B[60]), .B(n199), .ZN(DIFF[60]) );
  OR2_X1 U54 ( .A1(n214), .A2(B[45]), .ZN(n215) );
  OR2_X1 U55 ( .A1(n218), .A2(B[41]), .ZN(n219) );
  OR2_X1 U56 ( .A1(n222), .A2(B[37]), .ZN(n223) );
  XNOR2_X1 U57 ( .A(B[16]), .B(n246), .ZN(DIFF[16]) );
  OR3_X1 U58 ( .A1(B[17]), .A2(B[18]), .A3(n243), .ZN(n241) );
  OR2_X1 U59 ( .A1(n243), .A2(B[17]), .ZN(n244) );
  OR3_X1 U60 ( .A1(B[15]), .A2(B[16]), .A3(n245), .ZN(n243) );
  NOR2_X1 U61 ( .A1(B[15]), .A2(n245), .ZN(n246) );
  XNOR2_X1 U62 ( .A(n189), .B(B[10]), .ZN(DIFF[10]) );
  NOR2_X1 U63 ( .A1(n190), .A2(B[9]), .ZN(n189) );
  XNOR2_X1 U64 ( .A(n193), .B(B[6]), .ZN(DIFF[6]) );
  NOR2_X1 U65 ( .A1(n194), .A2(B[5]), .ZN(n193) );
  XNOR2_X1 U66 ( .A(B[12]), .B(n250), .ZN(DIFF[12]) );
  NOR2_X1 U67 ( .A1(B[11]), .A2(n249), .ZN(n250) );
  XNOR2_X1 U68 ( .A(B[8]), .B(n191), .ZN(DIFF[8]) );
  NOR2_X1 U69 ( .A1(B[7]), .A2(n192), .ZN(n191) );
  XNOR2_X1 U70 ( .A(B[2]), .B(n232), .ZN(DIFF[2]) );
  NOR2_X1 U71 ( .A1(\B[0] ), .A2(B[1]), .ZN(n232) );
  XNOR2_X1 U72 ( .A(B[4]), .B(n210), .ZN(DIFF[4]) );
  NOR2_X1 U73 ( .A1(B[3]), .A2(n211), .ZN(n210) );
  OR3_X1 U74 ( .A1(B[5]), .A2(B[6]), .A3(n194), .ZN(n192) );
  OR3_X1 U75 ( .A1(B[10]), .A2(B[9]), .A3(n190), .ZN(n249) );
  OR3_X1 U76 ( .A1(B[13]), .A2(B[14]), .A3(n247), .ZN(n245) );
  OR3_X1 U77 ( .A1(B[7]), .A2(B[8]), .A3(n192), .ZN(n190) );
  OR3_X1 U78 ( .A1(B[11]), .A2(B[12]), .A3(n249), .ZN(n247) );
  OR3_X1 U79 ( .A1(B[3]), .A2(B[4]), .A3(n211), .ZN(n194) );
  OR2_X1 U80 ( .A1(n247), .A2(B[13]), .ZN(n248) );
  OR3_X1 U83 ( .A1(B[1]), .A2(B[2]), .A3(\B[0] ), .ZN(n211) );
  INV_X1 U126 ( .A(B[61]), .ZN(n251) );
endmodule


module complementer_N64_17 ( \input , complement2 );
  input [63:0] \input ;
  output [63:0] complement2;


  complementer_N64_17_DW01_sub_0 sub_add_31_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(\input ), .CI(1'b0), .DIFF(complement2) );
endmodule


module ShiftnCompl_N64_9 ( plusA, plus2A_out, minus2A_out, plus4A_out, 
        minus4A_out );
  input [63:0] plusA;
  output [63:0] plus2A_out;
  output [63:0] minus2A_out;
  output [63:0] plus4A_out;
  output [63:0] minus4A_out;
  wire   n9, n10, n2, n11, n12, n13, n14;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign plus2A_out[0] = 1'b0;
  assign plus2A_out[51] = n2;
  assign plus4A_out[0] = 1'b0;

  shifter_N64_18 shifter_1 ( .\input (plusA), .shiftLeftOnePos({
        plus2A_out[63:59], n9, plus2A_out[57:54], n10, plus2A_out[52], n2, 
        plus2A_out[50:49], n11, plus2A_out[47:1], SYNOPSYS_UNCONNECTED__0}) );
  shifter_N64_17 shifter_2 ( .\input ({plus2A_out[63:52], n2, plus2A_out[50:1], 
        1'b0}), .shiftLeftOnePos({plus4A_out[63:59], n12, plus4A_out[57:54], 
        n13, plus4A_out[52:49], n14, plus4A_out[47:1], SYNOPSYS_UNCONNECTED__1}) );
  complementer_N64_18 complementer_1 ( .\input ({plus2A_out[63:52], n2, 
        plus2A_out[50:1], 1'b0}), .complement2(minus2A_out) );
  complementer_N64_17 complementer_2 ( .\input ({plus4A_out[63:1], 1'b0}), 
        .complement2(minus4A_out) );
  BUF_X1 U1 ( .A(n13), .Z(plus4A_out[53]) );
  BUF_X1 U4 ( .A(n10), .Z(plus2A_out[53]) );
  BUF_X1 U5 ( .A(n14), .Z(plus4A_out[48]) );
  BUF_X1 U6 ( .A(n12), .Z(plus4A_out[58]) );
  BUF_X1 U7 ( .A(n11), .Z(plus2A_out[48]) );
  BUF_X1 U8 ( .A(n9), .Z(plus2A_out[58]) );
endmodule


module MUX_GENERIC_N64_RADIX3_9 ( plusA, minusA, plus2A, minus2A, SEL, Y );
  input [63:0] plusA;
  input [63:0] minusA;
  input [63:0] plus2A;
  input [63:0] minus2A;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502;
  tri   [63:0] Y;

  TBUF_X1 \Y_tri[55]  ( .A(n446), .EN(n301), .Z(Y[55]) );
  TBUF_X1 \Y_tri[56]  ( .A(n445), .EN(n301), .Z(Y[56]) );
  TBUF_X1 \Y_tri[57]  ( .A(n444), .EN(n301), .Z(Y[57]) );
  TBUF_X1 \Y_tri[58]  ( .A(n443), .EN(n301), .Z(Y[58]) );
  TBUF_X1 \Y_tri[59]  ( .A(n442), .EN(n301), .Z(Y[59]) );
  TBUF_X1 \Y_tri[60]  ( .A(n441), .EN(n301), .Z(Y[60]) );
  TBUF_X1 \Y_tri[61]  ( .A(n440), .EN(n301), .Z(Y[61]) );
  TBUF_X1 \Y_tri[62]  ( .A(n439), .EN(n301), .Z(Y[62]) );
  TBUF_X1 \Y_tri[63]  ( .A(n438), .EN(n301), .Z(Y[63]) );
  TBUF_X1 \Y_tri[38]  ( .A(n463), .EN(n299), .Z(Y[38]) );
  TBUF_X1 \Y_tri[39]  ( .A(n462), .EN(n299), .Z(Y[39]) );
  TBUF_X1 \Y_tri[40]  ( .A(n461), .EN(n299), .Z(Y[40]) );
  TBUF_X1 \Y_tri[41]  ( .A(n460), .EN(n299), .Z(Y[41]) );
  TBUF_X1 \Y_tri[42]  ( .A(n459), .EN(n299), .Z(Y[42]) );
  TBUF_X1 \Y_tri[43]  ( .A(n458), .EN(n299), .Z(Y[43]) );
  TBUF_X1 \Y_tri[44]  ( .A(n457), .EN(n300), .Z(Y[44]) );
  TBUF_X1 \Y_tri[45]  ( .A(n456), .EN(n300), .Z(Y[45]) );
  TBUF_X1 \Y_tri[46]  ( .A(n455), .EN(n300), .Z(Y[46]) );
  TBUF_X1 \Y_tri[47]  ( .A(n454), .EN(n300), .Z(Y[47]) );
  TBUF_X1 \Y_tri[48]  ( .A(n453), .EN(n300), .Z(Y[48]) );
  TBUF_X1 \Y_tri[49]  ( .A(n452), .EN(n300), .Z(Y[49]) );
  TBUF_X1 \Y_tri[50]  ( .A(n451), .EN(n300), .Z(Y[50]) );
  TBUF_X1 \Y_tri[51]  ( .A(n450), .EN(n300), .Z(Y[51]) );
  TBUF_X1 \Y_tri[52]  ( .A(n449), .EN(n300), .Z(Y[52]) );
  TBUF_X1 \Y_tri[53]  ( .A(n448), .EN(n300), .Z(Y[53]) );
  TBUF_X1 \Y_tri[54]  ( .A(n447), .EN(n300), .Z(Y[54]) );
  TBUF_X1 \Y_tri[12]  ( .A(n489), .EN(n297), .Z(Y[12]) );
  TBUF_X1 \Y_tri[13]  ( .A(n488), .EN(n297), .Z(Y[13]) );
  TBUF_X1 \Y_tri[14]  ( .A(n487), .EN(n297), .Z(Y[14]) );
  TBUF_X1 \Y_tri[15]  ( .A(n486), .EN(n297), .Z(Y[15]) );
  TBUF_X1 \Y_tri[16]  ( .A(n485), .EN(n297), .Z(Y[16]) );
  TBUF_X1 \Y_tri[18]  ( .A(n483), .EN(n297), .Z(Y[18]) );
  TBUF_X1 \Y_tri[19]  ( .A(n482), .EN(n297), .Z(Y[19]) );
  TBUF_X1 \Y_tri[20]  ( .A(n481), .EN(n297), .Z(Y[20]) );
  TBUF_X1 \Y_tri[21]  ( .A(n480), .EN(n297), .Z(Y[21]) );
  TBUF_X1 \Y_tri[22]  ( .A(n479), .EN(n298), .Z(Y[22]) );
  TBUF_X1 \Y_tri[23]  ( .A(n478), .EN(n298), .Z(Y[23]) );
  TBUF_X1 \Y_tri[24]  ( .A(n477), .EN(n298), .Z(Y[24]) );
  TBUF_X1 \Y_tri[25]  ( .A(n476), .EN(n298), .Z(Y[25]) );
  TBUF_X1 \Y_tri[26]  ( .A(n475), .EN(n298), .Z(Y[26]) );
  TBUF_X1 \Y_tri[27]  ( .A(n474), .EN(n298), .Z(Y[27]) );
  TBUF_X1 \Y_tri[28]  ( .A(n473), .EN(n298), .Z(Y[28]) );
  TBUF_X1 \Y_tri[29]  ( .A(n472), .EN(n298), .Z(Y[29]) );
  TBUF_X1 \Y_tri[30]  ( .A(n471), .EN(n298), .Z(Y[30]) );
  TBUF_X1 \Y_tri[31]  ( .A(n470), .EN(n298), .Z(Y[31]) );
  TBUF_X1 \Y_tri[32]  ( .A(n469), .EN(n298), .Z(Y[32]) );
  TBUF_X1 \Y_tri[33]  ( .A(n468), .EN(n299), .Z(Y[33]) );
  TBUF_X1 \Y_tri[34]  ( .A(n467), .EN(n299), .Z(Y[34]) );
  TBUF_X1 \Y_tri[35]  ( .A(n466), .EN(n299), .Z(Y[35]) );
  TBUF_X1 \Y_tri[36]  ( .A(n465), .EN(n299), .Z(Y[36]) );
  TBUF_X1 \Y_tri[37]  ( .A(n464), .EN(n299), .Z(Y[37]) );
  TBUF_X1 \Y_tri[2]  ( .A(n500), .EN(n296), .Z(Y[2]) );
  TBUF_X1 \Y_tri[3]  ( .A(n499), .EN(n296), .Z(Y[3]) );
  TBUF_X1 \Y_tri[4]  ( .A(n498), .EN(n296), .Z(Y[4]) );
  TBUF_X1 \Y_tri[5]  ( .A(n497), .EN(n296), .Z(Y[5]) );
  TBUF_X1 \Y_tri[6]  ( .A(n496), .EN(n296), .Z(Y[6]) );
  TBUF_X1 \Y_tri[7]  ( .A(n495), .EN(n296), .Z(Y[7]) );
  TBUF_X1 \Y_tri[8]  ( .A(n494), .EN(n296), .Z(Y[8]) );
  TBUF_X1 \Y_tri[9]  ( .A(n492), .EN(n296), .Z(Y[9]) );
  TBUF_X1 \Y_tri[10]  ( .A(n491), .EN(n296), .Z(Y[10]) );
  TBUF_X1 \Y_tri[11]  ( .A(n490), .EN(n297), .Z(Y[11]) );
  TBUF_X1 \Y_tri[0]  ( .A(n502), .EN(n296), .Z(Y[0]) );
  TBUF_X1 \Y_tri[1]  ( .A(n501), .EN(n296), .Z(Y[1]) );
  TBUF_X1 \Y_tri[17]  ( .A(n484), .EN(n297), .Z(Y[17]) );
  NAND2_X1 U2 ( .A1(n359), .A2(n358), .ZN(n475) );
  AOI22_X1 U3 ( .A1(plusA[26]), .A2(n280), .B1(plus2A[26]), .B2(n274), .ZN(
        n359) );
  AOI22_X1 U4 ( .A1(minus2A[26]), .A2(n292), .B1(minusA[26]), .B2(n286), .ZN(
        n358) );
  NAND2_X1 U5 ( .A1(n355), .A2(n354), .ZN(n477) );
  AOI22_X1 U6 ( .A1(plusA[24]), .A2(n280), .B1(plus2A[24]), .B2(n274), .ZN(
        n355) );
  AOI22_X1 U7 ( .A1(minus2A[24]), .A2(n292), .B1(minusA[24]), .B2(n286), .ZN(
        n354) );
  NAND2_X1 U8 ( .A1(n353), .A2(n352), .ZN(n478) );
  AOI22_X1 U9 ( .A1(plusA[23]), .A2(n279), .B1(plus2A[23]), .B2(n273), .ZN(
        n353) );
  AOI22_X1 U10 ( .A1(minus2A[23]), .A2(n291), .B1(minusA[23]), .B2(n285), .ZN(
        n352) );
  NAND2_X1 U11 ( .A1(n351), .A2(n350), .ZN(n479) );
  AOI22_X1 U12 ( .A1(plusA[22]), .A2(n279), .B1(plus2A[22]), .B2(n273), .ZN(
        n351) );
  AOI22_X1 U13 ( .A1(minus2A[22]), .A2(n291), .B1(minusA[22]), .B2(n285), .ZN(
        n350) );
  NAND2_X1 U14 ( .A1(n347), .A2(n346), .ZN(n481) );
  AOI22_X1 U15 ( .A1(plusA[20]), .A2(n279), .B1(plus2A[20]), .B2(n273), .ZN(
        n347) );
  AOI22_X1 U16 ( .A1(minus2A[20]), .A2(n291), .B1(minusA[20]), .B2(n285), .ZN(
        n346) );
  NAND2_X1 U17 ( .A1(n345), .A2(n344), .ZN(n482) );
  AOI22_X1 U18 ( .A1(plusA[19]), .A2(n279), .B1(plus2A[19]), .B2(n273), .ZN(
        n345) );
  AOI22_X1 U19 ( .A1(minus2A[19]), .A2(n291), .B1(minusA[19]), .B2(n285), .ZN(
        n344) );
  NAND2_X1 U20 ( .A1(n343), .A2(n342), .ZN(n483) );
  AOI22_X1 U21 ( .A1(plusA[18]), .A2(n279), .B1(plus2A[18]), .B2(n273), .ZN(
        n343) );
  AOI22_X1 U22 ( .A1(minus2A[18]), .A2(n291), .B1(minusA[18]), .B2(n285), .ZN(
        n342) );
  NAND2_X1 U23 ( .A1(n375), .A2(n374), .ZN(n467) );
  AOI22_X1 U24 ( .A1(plusA[34]), .A2(n280), .B1(plus2A[34]), .B2(n274), .ZN(
        n375) );
  AOI22_X1 U25 ( .A1(minus2A[34]), .A2(n292), .B1(minusA[34]), .B2(n286), .ZN(
        n374) );
  NAND2_X1 U26 ( .A1(n367), .A2(n366), .ZN(n471) );
  AOI22_X1 U27 ( .A1(plusA[30]), .A2(n280), .B1(plus2A[30]), .B2(n274), .ZN(
        n367) );
  AOI22_X1 U28 ( .A1(minus2A[30]), .A2(n292), .B1(minusA[30]), .B2(n286), .ZN(
        n366) );
  NAND2_X1 U29 ( .A1(n379), .A2(n378), .ZN(n465) );
  AOI22_X1 U30 ( .A1(plusA[36]), .A2(n281), .B1(plus2A[36]), .B2(n275), .ZN(
        n379) );
  AOI22_X1 U31 ( .A1(minus2A[36]), .A2(n293), .B1(minusA[36]), .B2(n287), .ZN(
        n378) );
  NAND2_X1 U32 ( .A1(n371), .A2(n370), .ZN(n469) );
  AOI22_X1 U33 ( .A1(plusA[32]), .A2(n280), .B1(plus2A[32]), .B2(n274), .ZN(
        n371) );
  AOI22_X1 U34 ( .A1(minus2A[32]), .A2(n292), .B1(minusA[32]), .B2(n286), .ZN(
        n370) );
  NAND2_X1 U35 ( .A1(n363), .A2(n362), .ZN(n473) );
  AOI22_X1 U36 ( .A1(plusA[28]), .A2(n280), .B1(plus2A[28]), .B2(n274), .ZN(
        n363) );
  AOI22_X1 U37 ( .A1(minus2A[28]), .A2(n292), .B1(minusA[28]), .B2(n286), .ZN(
        n362) );
  NAND2_X1 U38 ( .A1(n377), .A2(n376), .ZN(n466) );
  AOI22_X1 U39 ( .A1(plusA[35]), .A2(n280), .B1(plus2A[35]), .B2(n274), .ZN(
        n377) );
  AOI22_X1 U40 ( .A1(minus2A[35]), .A2(n292), .B1(minusA[35]), .B2(n286), .ZN(
        n376) );
  NAND2_X1 U41 ( .A1(n369), .A2(n368), .ZN(n470) );
  AOI22_X1 U42 ( .A1(plusA[31]), .A2(n280), .B1(plus2A[31]), .B2(n274), .ZN(
        n369) );
  AOI22_X1 U43 ( .A1(minus2A[31]), .A2(n292), .B1(minusA[31]), .B2(n286), .ZN(
        n368) );
  NAND2_X1 U44 ( .A1(n361), .A2(n360), .ZN(n474) );
  AOI22_X1 U45 ( .A1(plusA[27]), .A2(n280), .B1(plus2A[27]), .B2(n274), .ZN(
        n361) );
  AOI22_X1 U46 ( .A1(minus2A[27]), .A2(n292), .B1(minusA[27]), .B2(n286), .ZN(
        n360) );
  NAND2_X1 U47 ( .A1(n381), .A2(n380), .ZN(n464) );
  AOI22_X1 U48 ( .A1(plusA[37]), .A2(n281), .B1(plus2A[37]), .B2(n275), .ZN(
        n381) );
  AOI22_X1 U49 ( .A1(minus2A[37]), .A2(n293), .B1(minusA[37]), .B2(n287), .ZN(
        n380) );
  NAND2_X1 U50 ( .A1(n373), .A2(n372), .ZN(n468) );
  AOI22_X1 U51 ( .A1(plusA[33]), .A2(n280), .B1(plus2A[33]), .B2(n274), .ZN(
        n373) );
  AOI22_X1 U52 ( .A1(minus2A[33]), .A2(n292), .B1(minusA[33]), .B2(n286), .ZN(
        n372) );
  NAND2_X1 U53 ( .A1(n365), .A2(n364), .ZN(n472) );
  AOI22_X1 U54 ( .A1(plusA[29]), .A2(n280), .B1(plus2A[29]), .B2(n274), .ZN(
        n365) );
  AOI22_X1 U55 ( .A1(minus2A[29]), .A2(n292), .B1(minusA[29]), .B2(n286), .ZN(
        n364) );
  NAND2_X1 U56 ( .A1(n357), .A2(n356), .ZN(n476) );
  AOI22_X1 U57 ( .A1(plusA[25]), .A2(n280), .B1(plus2A[25]), .B2(n274), .ZN(
        n357) );
  AOI22_X1 U58 ( .A1(minus2A[25]), .A2(n292), .B1(minusA[25]), .B2(n286), .ZN(
        n356) );
  NAND2_X1 U59 ( .A1(n349), .A2(n348), .ZN(n480) );
  AOI22_X1 U60 ( .A1(plusA[21]), .A2(n279), .B1(plus2A[21]), .B2(n273), .ZN(
        n349) );
  AOI22_X1 U61 ( .A1(minus2A[21]), .A2(n291), .B1(minusA[21]), .B2(n285), .ZN(
        n348) );
  NAND2_X1 U62 ( .A1(n391), .A2(n390), .ZN(n459) );
  AOI22_X1 U63 ( .A1(plusA[42]), .A2(n281), .B1(plus2A[42]), .B2(n275), .ZN(
        n391) );
  AOI22_X1 U64 ( .A1(minus2A[42]), .A2(n293), .B1(minusA[42]), .B2(n287), .ZN(
        n390) );
  NAND2_X1 U65 ( .A1(n383), .A2(n382), .ZN(n463) );
  AOI22_X1 U66 ( .A1(plusA[38]), .A2(n281), .B1(plus2A[38]), .B2(n275), .ZN(
        n383) );
  AOI22_X1 U67 ( .A1(minus2A[38]), .A2(n293), .B1(minusA[38]), .B2(n287), .ZN(
        n382) );
  NAND2_X1 U68 ( .A1(n401), .A2(n400), .ZN(n454) );
  AOI22_X1 U69 ( .A1(plusA[47]), .A2(n281), .B1(plus2A[47]), .B2(n275), .ZN(
        n401) );
  AOI22_X1 U70 ( .A1(minus2A[47]), .A2(n293), .B1(minusA[47]), .B2(n287), .ZN(
        n400) );
  NAND2_X1 U71 ( .A1(n419), .A2(n418), .ZN(n445) );
  AOI22_X1 U72 ( .A1(plusA[56]), .A2(n282), .B1(plus2A[56]), .B2(n276), .ZN(
        n419) );
  AOI22_X1 U73 ( .A1(minus2A[56]), .A2(n294), .B1(minusA[56]), .B2(n288), .ZN(
        n418) );
  NAND2_X1 U74 ( .A1(n415), .A2(n414), .ZN(n447) );
  AOI22_X1 U75 ( .A1(plusA[54]), .A2(n282), .B1(plus2A[54]), .B2(n276), .ZN(
        n415) );
  AOI22_X1 U76 ( .A1(minus2A[54]), .A2(n294), .B1(minusA[54]), .B2(n288), .ZN(
        n414) );
  NAND2_X1 U77 ( .A1(n395), .A2(n394), .ZN(n457) );
  AOI22_X1 U78 ( .A1(plusA[44]), .A2(n281), .B1(plus2A[44]), .B2(n275), .ZN(
        n395) );
  AOI22_X1 U79 ( .A1(minus2A[44]), .A2(n293), .B1(minusA[44]), .B2(n287), .ZN(
        n394) );
  NAND2_X1 U80 ( .A1(n387), .A2(n386), .ZN(n461) );
  AOI22_X1 U81 ( .A1(plusA[40]), .A2(n281), .B1(plus2A[40]), .B2(n275), .ZN(
        n387) );
  AOI22_X1 U82 ( .A1(minus2A[40]), .A2(n293), .B1(minusA[40]), .B2(n287), .ZN(
        n386) );
  NAND2_X1 U83 ( .A1(n421), .A2(n420), .ZN(n444) );
  AOI22_X1 U84 ( .A1(plusA[57]), .A2(n282), .B1(plus2A[57]), .B2(n276), .ZN(
        n421) );
  AOI22_X1 U85 ( .A1(minus2A[57]), .A2(n294), .B1(minusA[57]), .B2(n288), .ZN(
        n420) );
  NAND2_X1 U86 ( .A1(n417), .A2(n416), .ZN(n446) );
  AOI22_X1 U87 ( .A1(plusA[55]), .A2(n282), .B1(plus2A[55]), .B2(n276), .ZN(
        n417) );
  AOI22_X1 U88 ( .A1(minus2A[55]), .A2(n294), .B1(minusA[55]), .B2(n288), .ZN(
        n416) );
  NAND2_X1 U89 ( .A1(n413), .A2(n412), .ZN(n448) );
  AOI22_X1 U90 ( .A1(plusA[53]), .A2(n282), .B1(plus2A[53]), .B2(n276), .ZN(
        n413) );
  AOI22_X1 U91 ( .A1(minus2A[53]), .A2(n294), .B1(minusA[53]), .B2(n288), .ZN(
        n412) );
  NAND2_X1 U92 ( .A1(n397), .A2(n396), .ZN(n456) );
  AOI22_X1 U93 ( .A1(plusA[45]), .A2(n281), .B1(plus2A[45]), .B2(n275), .ZN(
        n397) );
  AOI22_X1 U94 ( .A1(minus2A[45]), .A2(n293), .B1(minusA[45]), .B2(n287), .ZN(
        n396) );
  NAND2_X1 U95 ( .A1(n409), .A2(n408), .ZN(n450) );
  AOI22_X1 U96 ( .A1(plusA[51]), .A2(n282), .B1(plus2A[51]), .B2(n276), .ZN(
        n409) );
  AOI22_X1 U97 ( .A1(minus2A[51]), .A2(n294), .B1(minusA[51]), .B2(n288), .ZN(
        n408) );
  NAND2_X1 U98 ( .A1(n405), .A2(n404), .ZN(n452) );
  AOI22_X1 U99 ( .A1(plusA[49]), .A2(n282), .B1(plus2A[49]), .B2(n276), .ZN(
        n405) );
  AOI22_X1 U100 ( .A1(minus2A[49]), .A2(n294), .B1(minusA[49]), .B2(n288), 
        .ZN(n404) );
  NAND2_X1 U101 ( .A1(n393), .A2(n392), .ZN(n458) );
  AOI22_X1 U102 ( .A1(plusA[43]), .A2(n281), .B1(plus2A[43]), .B2(n275), .ZN(
        n393) );
  AOI22_X1 U103 ( .A1(minus2A[43]), .A2(n293), .B1(minusA[43]), .B2(n287), 
        .ZN(n392) );
  NAND2_X1 U104 ( .A1(n385), .A2(n384), .ZN(n462) );
  AOI22_X1 U105 ( .A1(plusA[39]), .A2(n281), .B1(plus2A[39]), .B2(n275), .ZN(
        n385) );
  AOI22_X1 U106 ( .A1(minus2A[39]), .A2(n293), .B1(minusA[39]), .B2(n287), 
        .ZN(n384) );
  NAND2_X1 U107 ( .A1(n411), .A2(n410), .ZN(n449) );
  AOI22_X1 U108 ( .A1(plusA[52]), .A2(n282), .B1(plus2A[52]), .B2(n276), .ZN(
        n411) );
  AOI22_X1 U109 ( .A1(minus2A[52]), .A2(n294), .B1(minusA[52]), .B2(n288), 
        .ZN(n410) );
  NAND2_X1 U110 ( .A1(n407), .A2(n406), .ZN(n451) );
  AOI22_X1 U111 ( .A1(plusA[50]), .A2(n282), .B1(plus2A[50]), .B2(n276), .ZN(
        n407) );
  AOI22_X1 U112 ( .A1(minus2A[50]), .A2(n294), .B1(minusA[50]), .B2(n288), 
        .ZN(n406) );
  NAND2_X1 U113 ( .A1(n403), .A2(n402), .ZN(n453) );
  AOI22_X1 U114 ( .A1(plusA[48]), .A2(n282), .B1(plus2A[48]), .B2(n276), .ZN(
        n403) );
  AOI22_X1 U115 ( .A1(minus2A[48]), .A2(n294), .B1(minusA[48]), .B2(n288), 
        .ZN(n402) );
  NAND2_X1 U116 ( .A1(n389), .A2(n388), .ZN(n460) );
  AOI22_X1 U117 ( .A1(plusA[41]), .A2(n281), .B1(plus2A[41]), .B2(n275), .ZN(
        n389) );
  AOI22_X1 U118 ( .A1(minus2A[41]), .A2(n293), .B1(minusA[41]), .B2(n287), 
        .ZN(n388) );
  NAND2_X1 U119 ( .A1(n399), .A2(n398), .ZN(n455) );
  AOI22_X1 U120 ( .A1(plusA[46]), .A2(n281), .B1(plus2A[46]), .B2(n275), .ZN(
        n399) );
  AOI22_X1 U121 ( .A1(minus2A[46]), .A2(n293), .B1(minusA[46]), .B2(n287), 
        .ZN(n398) );
  NAND2_X1 U122 ( .A1(n437), .A2(n436), .ZN(n438) );
  AOI22_X1 U123 ( .A1(plusA[63]), .A2(n283), .B1(plus2A[63]), .B2(n277), .ZN(
        n437) );
  AOI22_X1 U124 ( .A1(minus2A[63]), .A2(n295), .B1(minusA[63]), .B2(n289), 
        .ZN(n436) );
  NAND2_X1 U125 ( .A1(n431), .A2(n430), .ZN(n439) );
  AOI22_X1 U126 ( .A1(plusA[62]), .A2(n283), .B1(plus2A[62]), .B2(n277), .ZN(
        n431) );
  AOI22_X1 U127 ( .A1(minus2A[62]), .A2(n295), .B1(minusA[62]), .B2(n289), 
        .ZN(n430) );
  NAND2_X1 U128 ( .A1(n429), .A2(n428), .ZN(n440) );
  AOI22_X1 U129 ( .A1(plusA[61]), .A2(n283), .B1(plus2A[61]), .B2(n277), .ZN(
        n429) );
  AOI22_X1 U130 ( .A1(minus2A[61]), .A2(n295), .B1(minusA[61]), .B2(n289), 
        .ZN(n428) );
  NAND2_X1 U131 ( .A1(n427), .A2(n426), .ZN(n441) );
  AOI22_X1 U132 ( .A1(plusA[60]), .A2(n283), .B1(plus2A[60]), .B2(n277), .ZN(
        n427) );
  AOI22_X1 U133 ( .A1(minus2A[60]), .A2(n295), .B1(minusA[60]), .B2(n289), 
        .ZN(n426) );
  NAND2_X1 U134 ( .A1(n425), .A2(n424), .ZN(n442) );
  AOI22_X1 U135 ( .A1(plusA[59]), .A2(n282), .B1(plus2A[59]), .B2(n276), .ZN(
        n425) );
  AOI22_X1 U136 ( .A1(minus2A[59]), .A2(n294), .B1(minusA[59]), .B2(n288), 
        .ZN(n424) );
  NAND2_X1 U137 ( .A1(n423), .A2(n422), .ZN(n443) );
  AOI22_X1 U138 ( .A1(plusA[58]), .A2(n282), .B1(plus2A[58]), .B2(n276), .ZN(
        n423) );
  AOI22_X1 U139 ( .A1(minus2A[58]), .A2(n294), .B1(minusA[58]), .B2(n288), 
        .ZN(n422) );
  BUF_X1 U140 ( .A(n493), .Z(n296) );
  BUF_X1 U141 ( .A(n434), .Z(n285) );
  BUF_X1 U142 ( .A(n432), .Z(n273) );
  BUF_X1 U143 ( .A(n493), .Z(n297) );
  NAND2_X1 U144 ( .A1(n341), .A2(n340), .ZN(n484) );
  AOI22_X1 U145 ( .A1(plusA[17]), .A2(n279), .B1(plus2A[17]), .B2(n273), .ZN(
        n341) );
  AOI22_X1 U146 ( .A1(minus2A[17]), .A2(n291), .B1(minusA[17]), .B2(n285), 
        .ZN(n340) );
  BUF_X1 U147 ( .A(n433), .Z(n279) );
  BUF_X1 U148 ( .A(n435), .Z(n291) );
  BUF_X1 U149 ( .A(n493), .Z(n298) );
  NAND2_X1 U150 ( .A1(n339), .A2(n338), .ZN(n485) );
  AOI22_X1 U151 ( .A1(plusA[16]), .A2(n279), .B1(plus2A[16]), .B2(n273), .ZN(
        n339) );
  AOI22_X1 U152 ( .A1(minus2A[16]), .A2(n291), .B1(minusA[16]), .B2(n285), 
        .ZN(n338) );
  BUF_X1 U153 ( .A(n433), .Z(n280) );
  BUF_X1 U154 ( .A(n435), .Z(n292) );
  BUF_X1 U155 ( .A(n434), .Z(n286) );
  BUF_X1 U156 ( .A(n432), .Z(n274) );
  BUF_X1 U157 ( .A(n433), .Z(n281) );
  BUF_X1 U158 ( .A(n435), .Z(n293) );
  BUF_X1 U159 ( .A(n434), .Z(n287) );
  BUF_X1 U160 ( .A(n432), .Z(n275) );
  BUF_X1 U161 ( .A(n493), .Z(n299) );
  BUF_X1 U162 ( .A(n433), .Z(n282) );
  BUF_X1 U163 ( .A(n435), .Z(n294) );
  BUF_X1 U164 ( .A(n434), .Z(n288) );
  BUF_X1 U165 ( .A(n432), .Z(n276) );
  BUF_X1 U166 ( .A(n493), .Z(n300) );
  BUF_X1 U167 ( .A(n493), .Z(n301) );
  BUF_X1 U168 ( .A(n433), .Z(n278) );
  BUF_X1 U169 ( .A(n435), .Z(n290) );
  BUF_X1 U170 ( .A(n434), .Z(n284) );
  BUF_X1 U171 ( .A(n432), .Z(n272) );
  NOR2_X1 U172 ( .A1(n323), .A2(n304), .ZN(n493) );
  INV_X1 U173 ( .A(SEL[2]), .ZN(n304) );
  NOR2_X1 U174 ( .A1(SEL[1]), .A2(SEL[0]), .ZN(n323) );
  NOR3_X1 U175 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n302), .ZN(n434) );
  NOR3_X1 U176 ( .A1(n302), .A2(SEL[2]), .A3(n303), .ZN(n432) );
  INV_X1 U177 ( .A(SEL[1]), .ZN(n302) );
  INV_X1 U178 ( .A(SEL[0]), .ZN(n303) );
  NOR3_X1 U179 ( .A1(SEL[1]), .A2(SEL[2]), .A3(n303), .ZN(n433) );
  NAND2_X1 U180 ( .A1(n337), .A2(n336), .ZN(n486) );
  AOI22_X1 U181 ( .A1(plusA[15]), .A2(n279), .B1(plus2A[15]), .B2(n273), .ZN(
        n337) );
  AOI22_X1 U182 ( .A1(minus2A[15]), .A2(n291), .B1(minusA[15]), .B2(n285), 
        .ZN(n336) );
  AND2_X1 U183 ( .A1(SEL[2]), .A2(n323), .ZN(n435) );
  NAND2_X1 U184 ( .A1(n335), .A2(n334), .ZN(n487) );
  AOI22_X1 U185 ( .A1(plusA[14]), .A2(n279), .B1(plus2A[14]), .B2(n273), .ZN(
        n335) );
  AOI22_X1 U186 ( .A1(minus2A[14]), .A2(n291), .B1(minusA[14]), .B2(n285), 
        .ZN(n334) );
  NAND2_X1 U187 ( .A1(n333), .A2(n332), .ZN(n488) );
  AOI22_X1 U188 ( .A1(plusA[13]), .A2(n279), .B1(plus2A[13]), .B2(n273), .ZN(
        n333) );
  AOI22_X1 U189 ( .A1(minus2A[13]), .A2(n291), .B1(minusA[13]), .B2(n285), 
        .ZN(n332) );
  NAND2_X1 U190 ( .A1(n329), .A2(n328), .ZN(n490) );
  AOI22_X1 U191 ( .A1(plusA[11]), .A2(n278), .B1(plus2A[11]), .B2(n272), .ZN(
        n329) );
  AOI22_X1 U192 ( .A1(minus2A[11]), .A2(n290), .B1(minusA[11]), .B2(n284), 
        .ZN(n328) );
  NAND2_X1 U193 ( .A1(n327), .A2(n326), .ZN(n491) );
  AOI22_X1 U194 ( .A1(plusA[10]), .A2(n278), .B1(plus2A[10]), .B2(n272), .ZN(
        n327) );
  AOI22_X1 U195 ( .A1(minus2A[10]), .A2(n290), .B1(minusA[10]), .B2(n284), 
        .ZN(n326) );
  NAND2_X1 U196 ( .A1(n325), .A2(n324), .ZN(n492) );
  AOI22_X1 U197 ( .A1(plusA[9]), .A2(n278), .B1(plus2A[9]), .B2(n272), .ZN(
        n325) );
  AOI22_X1 U198 ( .A1(minus2A[9]), .A2(n290), .B1(minusA[9]), .B2(n284), .ZN(
        n324) );
  NAND2_X1 U199 ( .A1(n320), .A2(n319), .ZN(n495) );
  AOI22_X1 U200 ( .A1(plusA[7]), .A2(n278), .B1(plus2A[7]), .B2(n272), .ZN(
        n320) );
  AOI22_X1 U201 ( .A1(minus2A[7]), .A2(n290), .B1(minusA[7]), .B2(n284), .ZN(
        n319) );
  NAND2_X1 U202 ( .A1(n318), .A2(n317), .ZN(n496) );
  AOI22_X1 U203 ( .A1(plusA[6]), .A2(n278), .B1(plus2A[6]), .B2(n272), .ZN(
        n318) );
  AOI22_X1 U204 ( .A1(minus2A[6]), .A2(n290), .B1(minusA[6]), .B2(n284), .ZN(
        n317) );
  NAND2_X1 U205 ( .A1(n316), .A2(n315), .ZN(n497) );
  AOI22_X1 U206 ( .A1(plusA[5]), .A2(n278), .B1(plus2A[5]), .B2(n272), .ZN(
        n316) );
  AOI22_X1 U207 ( .A1(minus2A[5]), .A2(n290), .B1(minusA[5]), .B2(n284), .ZN(
        n315) );
  NAND2_X1 U208 ( .A1(n312), .A2(n311), .ZN(n499) );
  AOI22_X1 U209 ( .A1(plusA[3]), .A2(n278), .B1(plus2A[3]), .B2(n272), .ZN(
        n312) );
  AOI22_X1 U210 ( .A1(minus2A[3]), .A2(n290), .B1(minusA[3]), .B2(n284), .ZN(
        n311) );
  NAND2_X1 U211 ( .A1(n331), .A2(n330), .ZN(n489) );
  AOI22_X1 U212 ( .A1(plusA[12]), .A2(n279), .B1(plus2A[12]), .B2(n273), .ZN(
        n331) );
  AOI22_X1 U213 ( .A1(minus2A[12]), .A2(n291), .B1(minusA[12]), .B2(n285), 
        .ZN(n330) );
  NAND2_X1 U214 ( .A1(n322), .A2(n321), .ZN(n494) );
  AOI22_X1 U215 ( .A1(plusA[8]), .A2(n278), .B1(plus2A[8]), .B2(n272), .ZN(
        n322) );
  AOI22_X1 U216 ( .A1(minus2A[8]), .A2(n290), .B1(minusA[8]), .B2(n284), .ZN(
        n321) );
  NAND2_X1 U217 ( .A1(n314), .A2(n313), .ZN(n498) );
  AOI22_X1 U218 ( .A1(plusA[4]), .A2(n278), .B1(plus2A[4]), .B2(n272), .ZN(
        n314) );
  AOI22_X1 U219 ( .A1(minus2A[4]), .A2(n290), .B1(minusA[4]), .B2(n284), .ZN(
        n313) );
  NAND2_X1 U220 ( .A1(n310), .A2(n309), .ZN(n500) );
  AOI22_X1 U221 ( .A1(plusA[2]), .A2(n278), .B1(plus2A[2]), .B2(n272), .ZN(
        n310) );
  AOI22_X1 U222 ( .A1(minus2A[2]), .A2(n290), .B1(minusA[2]), .B2(n284), .ZN(
        n309) );
  NAND2_X1 U223 ( .A1(n308), .A2(n307), .ZN(n501) );
  AOI22_X1 U224 ( .A1(plusA[1]), .A2(n278), .B1(plus2A[1]), .B2(n272), .ZN(
        n308) );
  AOI22_X1 U225 ( .A1(minus2A[1]), .A2(n290), .B1(minusA[1]), .B2(n284), .ZN(
        n307) );
  NAND2_X1 U226 ( .A1(n306), .A2(n305), .ZN(n502) );
  AOI22_X1 U227 ( .A1(plusA[0]), .A2(n278), .B1(plus2A[0]), .B2(n272), .ZN(
        n306) );
  AOI22_X1 U228 ( .A1(minus2A[0]), .A2(n290), .B1(minusA[0]), .B2(n284), .ZN(
        n305) );
  CLKBUF_X1 U229 ( .A(n432), .Z(n277) );
  CLKBUF_X1 U230 ( .A(n433), .Z(n283) );
  CLKBUF_X1 U231 ( .A(n434), .Z(n289) );
  CLKBUF_X1 U232 ( .A(n435), .Z(n295) );
endmodule


module FA_576 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_575 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_574 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_573 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_572 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_571 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_570 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_569 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_568 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_567 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_566 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_565 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_564 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_563 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_562 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_561 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_560 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_559 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_558 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_557 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_556 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_555 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_554 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_553 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_552 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_551 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_550 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_549 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_548 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_547 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_546 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_545 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_544 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_543 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_542 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_541 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_540 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_539 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_538 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_537 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_536 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_535 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_534 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_533 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_532 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_531 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_530 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_529 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_528 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_527 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_526 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_525 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_524 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_523 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_522 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_521 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_520 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_519 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_518 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_517 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_516 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_515 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_514 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_513 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N64_9 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Ci;
  output Co;

  wire   [63:1] CTMP;
  tri   [63:0] A;

  FA_576 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_575 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_574 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_573 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(CTMP[4]) );
  FA_572 FAI_5 ( .A(A[4]), .B(B[4]), .Ci(CTMP[4]), .S(S[4]), .Co(CTMP[5]) );
  FA_571 FAI_6 ( .A(A[5]), .B(B[5]), .Ci(CTMP[5]), .S(S[5]), .Co(CTMP[6]) );
  FA_570 FAI_7 ( .A(A[6]), .B(B[6]), .Ci(CTMP[6]), .S(S[6]), .Co(CTMP[7]) );
  FA_569 FAI_8 ( .A(A[7]), .B(B[7]), .Ci(CTMP[7]), .S(S[7]), .Co(CTMP[8]) );
  FA_568 FAI_9 ( .A(A[8]), .B(B[8]), .Ci(CTMP[8]), .S(S[8]), .Co(CTMP[9]) );
  FA_567 FAI_10 ( .A(A[9]), .B(B[9]), .Ci(CTMP[9]), .S(S[9]), .Co(CTMP[10]) );
  FA_566 FAI_11 ( .A(A[10]), .B(B[10]), .Ci(CTMP[10]), .S(S[10]), .Co(CTMP[11]) );
  FA_565 FAI_12 ( .A(A[11]), .B(B[11]), .Ci(CTMP[11]), .S(S[11]), .Co(CTMP[12]) );
  FA_564 FAI_13 ( .A(A[12]), .B(B[12]), .Ci(CTMP[12]), .S(S[12]), .Co(CTMP[13]) );
  FA_563 FAI_14 ( .A(A[13]), .B(B[13]), .Ci(CTMP[13]), .S(S[13]), .Co(CTMP[14]) );
  FA_562 FAI_15 ( .A(A[14]), .B(B[14]), .Ci(CTMP[14]), .S(S[14]), .Co(CTMP[15]) );
  FA_561 FAI_16 ( .A(A[15]), .B(B[15]), .Ci(CTMP[15]), .S(S[15]), .Co(CTMP[16]) );
  FA_560 FAI_17 ( .A(A[16]), .B(B[16]), .Ci(CTMP[16]), .S(S[16]), .Co(CTMP[17]) );
  FA_559 FAI_18 ( .A(A[17]), .B(B[17]), .Ci(CTMP[17]), .S(S[17]), .Co(CTMP[18]) );
  FA_558 FAI_19 ( .A(A[18]), .B(B[18]), .Ci(CTMP[18]), .S(S[18]), .Co(CTMP[19]) );
  FA_557 FAI_20 ( .A(A[19]), .B(B[19]), .Ci(CTMP[19]), .S(S[19]), .Co(CTMP[20]) );
  FA_556 FAI_21 ( .A(A[20]), .B(B[20]), .Ci(CTMP[20]), .S(S[20]), .Co(CTMP[21]) );
  FA_555 FAI_22 ( .A(A[21]), .B(B[21]), .Ci(CTMP[21]), .S(S[21]), .Co(CTMP[22]) );
  FA_554 FAI_23 ( .A(A[22]), .B(B[22]), .Ci(CTMP[22]), .S(S[22]), .Co(CTMP[23]) );
  FA_553 FAI_24 ( .A(A[23]), .B(B[23]), .Ci(CTMP[23]), .S(S[23]), .Co(CTMP[24]) );
  FA_552 FAI_25 ( .A(A[24]), .B(B[24]), .Ci(CTMP[24]), .S(S[24]), .Co(CTMP[25]) );
  FA_551 FAI_26 ( .A(A[25]), .B(B[25]), .Ci(CTMP[25]), .S(S[25]), .Co(CTMP[26]) );
  FA_550 FAI_27 ( .A(A[26]), .B(B[26]), .Ci(CTMP[26]), .S(S[26]), .Co(CTMP[27]) );
  FA_549 FAI_28 ( .A(A[27]), .B(B[27]), .Ci(CTMP[27]), .S(S[27]), .Co(CTMP[28]) );
  FA_548 FAI_29 ( .A(A[28]), .B(B[28]), .Ci(CTMP[28]), .S(S[28]), .Co(CTMP[29]) );
  FA_547 FAI_30 ( .A(A[29]), .B(B[29]), .Ci(CTMP[29]), .S(S[29]), .Co(CTMP[30]) );
  FA_546 FAI_31 ( .A(A[30]), .B(B[30]), .Ci(CTMP[30]), .S(S[30]), .Co(CTMP[31]) );
  FA_545 FAI_32 ( .A(A[31]), .B(B[31]), .Ci(CTMP[31]), .S(S[31]), .Co(CTMP[32]) );
  FA_544 FAI_33 ( .A(A[32]), .B(B[32]), .Ci(CTMP[32]), .S(S[32]), .Co(CTMP[33]) );
  FA_543 FAI_34 ( .A(A[33]), .B(B[33]), .Ci(CTMP[33]), .S(S[33]), .Co(CTMP[34]) );
  FA_542 FAI_35 ( .A(A[34]), .B(B[34]), .Ci(CTMP[34]), .S(S[34]), .Co(CTMP[35]) );
  FA_541 FAI_36 ( .A(A[35]), .B(B[35]), .Ci(CTMP[35]), .S(S[35]), .Co(CTMP[36]) );
  FA_540 FAI_37 ( .A(A[36]), .B(B[36]), .Ci(CTMP[36]), .S(S[36]), .Co(CTMP[37]) );
  FA_539 FAI_38 ( .A(A[37]), .B(B[37]), .Ci(CTMP[37]), .S(S[37]), .Co(CTMP[38]) );
  FA_538 FAI_39 ( .A(A[38]), .B(B[38]), .Ci(CTMP[38]), .S(S[38]), .Co(CTMP[39]) );
  FA_537 FAI_40 ( .A(A[39]), .B(B[39]), .Ci(CTMP[39]), .S(S[39]), .Co(CTMP[40]) );
  FA_536 FAI_41 ( .A(A[40]), .B(B[40]), .Ci(CTMP[40]), .S(S[40]), .Co(CTMP[41]) );
  FA_535 FAI_42 ( .A(A[41]), .B(B[41]), .Ci(CTMP[41]), .S(S[41]), .Co(CTMP[42]) );
  FA_534 FAI_43 ( .A(A[42]), .B(B[42]), .Ci(CTMP[42]), .S(S[42]), .Co(CTMP[43]) );
  FA_533 FAI_44 ( .A(A[43]), .B(B[43]), .Ci(CTMP[43]), .S(S[43]), .Co(CTMP[44]) );
  FA_532 FAI_45 ( .A(A[44]), .B(B[44]), .Ci(CTMP[44]), .S(S[44]), .Co(CTMP[45]) );
  FA_531 FAI_46 ( .A(A[45]), .B(B[45]), .Ci(CTMP[45]), .S(S[45]), .Co(CTMP[46]) );
  FA_530 FAI_47 ( .A(A[46]), .B(B[46]), .Ci(CTMP[46]), .S(S[46]), .Co(CTMP[47]) );
  FA_529 FAI_48 ( .A(A[47]), .B(B[47]), .Ci(CTMP[47]), .S(S[47]), .Co(CTMP[48]) );
  FA_528 FAI_49 ( .A(A[48]), .B(B[48]), .Ci(CTMP[48]), .S(S[48]), .Co(CTMP[49]) );
  FA_527 FAI_50 ( .A(A[49]), .B(B[49]), .Ci(CTMP[49]), .S(S[49]), .Co(CTMP[50]) );
  FA_526 FAI_51 ( .A(A[50]), .B(B[50]), .Ci(CTMP[50]), .S(S[50]), .Co(CTMP[51]) );
  FA_525 FAI_52 ( .A(A[51]), .B(B[51]), .Ci(CTMP[51]), .S(S[51]), .Co(CTMP[52]) );
  FA_524 FAI_53 ( .A(A[52]), .B(B[52]), .Ci(CTMP[52]), .S(S[52]), .Co(CTMP[53]) );
  FA_523 FAI_54 ( .A(A[53]), .B(B[53]), .Ci(CTMP[53]), .S(S[53]), .Co(CTMP[54]) );
  FA_522 FAI_55 ( .A(A[54]), .B(B[54]), .Ci(CTMP[54]), .S(S[54]), .Co(CTMP[55]) );
  FA_521 FAI_56 ( .A(A[55]), .B(B[55]), .Ci(CTMP[55]), .S(S[55]), .Co(CTMP[56]) );
  FA_520 FAI_57 ( .A(A[56]), .B(B[56]), .Ci(CTMP[56]), .S(S[56]), .Co(CTMP[57]) );
  FA_519 FAI_58 ( .A(A[57]), .B(B[57]), .Ci(CTMP[57]), .S(S[57]), .Co(CTMP[58]) );
  FA_518 FAI_59 ( .A(A[58]), .B(B[58]), .Ci(CTMP[58]), .S(S[58]), .Co(CTMP[59]) );
  FA_517 FAI_60 ( .A(A[59]), .B(B[59]), .Ci(CTMP[59]), .S(S[59]), .Co(CTMP[60]) );
  FA_516 FAI_61 ( .A(A[60]), .B(B[60]), .Ci(CTMP[60]), .S(S[60]), .Co(CTMP[61]) );
  FA_515 FAI_62 ( .A(A[61]), .B(B[61]), .Ci(CTMP[61]), .S(S[61]), .Co(CTMP[62]) );
  FA_514 FAI_63 ( .A(A[62]), .B(B[62]), .Ci(CTMP[62]), .S(S[62]), .Co(CTMP[63]) );
  FA_513 FAI_64 ( .A(A[63]), .B(B[63]), .Ci(CTMP[63]), .S(S[63]), .Co(Co) );
endmodule


module booth_mul_row_N64_RADIX3_9 ( prevA, prevSum, encoderIn, nextA, nextSum
 );
  input [63:0] prevA;
  input [63:0] prevSum;
  input [2:0] encoderIn;
  output [63:0] nextA;
  output [63:0] nextSum;
  wire   n3;
  wire   [2:0] encoder_to_mux;
  wire   [63:0] plus2A_s;
  wire   [63:0] minus2A_s;
  wire   [63:0] minus4A_s;
  tri   [63:0] mux_to_adder;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign nextA[51] = n3;
  assign nextA[0] = 1'b0;

  encoder_N64_RADIX3_9 encoder_1 ( .X(encoderIn), .Z(encoder_to_mux) );
  ShiftnCompl_N64_9 ShiftnCompl_1 ( .plusA(prevA), .plus2A_out({plus2A_s[63:1], 
        SYNOPSYS_UNCONNECTED__0}), .minus2A_out(minus2A_s), .plus4A_out({
        nextA[63:52], n3, nextA[50:1], SYNOPSYS_UNCONNECTED__1}), 
        .minus4A_out(minus4A_s) );
  MUX_GENERIC_N64_RADIX3_9 mux_1 ( .plusA({plus2A_s[63:1], 1'b0}), .minusA(
        minus2A_s), .plus2A({nextA[63:52], n3, nextA[50:1], 1'b0}), .minus2A(
        minus4A_s), .SEL(encoder_to_mux), .Y(mux_to_adder) );
  RCA_N64_9 rca_1 ( .A(mux_to_adder), .B(prevSum), .Ci(1'b0), .S(nextSum) );
endmodule


module encoder_N64_RADIX3_8 ( X, Z );
  input [2:0] X;
  output [2:0] Z;
  wire   n5, n7, n8;

  OAI22_X1 U1 ( .A1(n8), .A2(n5), .B1(X[2]), .B2(n7), .ZN(Z[1]) );
  INV_X1 U2 ( .A(X[2]), .ZN(n5) );
  AOI21_X1 U3 ( .B1(n8), .B2(n7), .A(X[2]), .ZN(Z[0]) );
  OAI21_X1 U4 ( .B1(X[1]), .B2(X[0]), .A(n7), .ZN(n8) );
  AND3_X1 U5 ( .A1(X[2]), .A2(n7), .A3(n8), .ZN(Z[2]) );
  NAND2_X1 U6 ( .A1(X[1]), .A2(X[0]), .ZN(n7) );
endmodule


module shifter_N64_16 ( \input , shiftLeftOnePos );
  input [63:0] \input ;
  output [63:0] shiftLeftOnePos;
  wire   \input[62] , \input[61] , \input[60] , \input[59] , \input[58] ,
         \input[57] , \input[56] , \input[55] , \input[54] , \input[53] ,
         \input[52] , \input[51] , \input[50] , \input[49] , \input[48] ,
         \input[47] , \input[46] , \input[45] , \input[44] , \input[43] ,
         \input[42] , \input[41] , \input[40] , \input[39] , \input[38] ,
         \input[37] , \input[36] , \input[35] , \input[34] , \input[33] ,
         \input[32] , \input[31] , \input[30] , \input[29] , \input[28] ,
         \input[27] , \input[26] , \input[25] , \input[24] , \input[23] ,
         \input[22] , \input[21] , \input[20] , \input[19] , \input[18] ,
         \input[17] , \input[16] , \input[15] , \input[14] , \input[13] ,
         \input[12] , \input[11] , \input[10] , \input[9] , \input[8] ,
         \input[7] , \input[6] , \input[5] , \input[4] , \input[3] ,
         \input[2] , \input[1] , \input[0] ;
  assign shiftLeftOnePos[0] = 1'b0;
  assign shiftLeftOnePos[63] = \input[62] ;
  assign \input[62]  = \input  [62];
  assign shiftLeftOnePos[62] = \input[61] ;
  assign \input[61]  = \input  [61];
  assign shiftLeftOnePos[61] = \input[60] ;
  assign \input[60]  = \input  [60];
  assign shiftLeftOnePos[60] = \input[59] ;
  assign \input[59]  = \input  [59];
  assign shiftLeftOnePos[59] = \input[58] ;
  assign \input[58]  = \input  [58];
  assign shiftLeftOnePos[58] = \input[57] ;
  assign \input[57]  = \input  [57];
  assign shiftLeftOnePos[57] = \input[56] ;
  assign \input[56]  = \input  [56];
  assign shiftLeftOnePos[56] = \input[55] ;
  assign \input[55]  = \input  [55];
  assign shiftLeftOnePos[55] = \input[54] ;
  assign \input[54]  = \input  [54];
  assign shiftLeftOnePos[54] = \input[53] ;
  assign \input[53]  = \input  [53];
  assign shiftLeftOnePos[53] = \input[52] ;
  assign \input[52]  = \input  [52];
  assign shiftLeftOnePos[52] = \input[51] ;
  assign \input[51]  = \input  [51];
  assign shiftLeftOnePos[51] = \input[50] ;
  assign \input[50]  = \input  [50];
  assign shiftLeftOnePos[50] = \input[49] ;
  assign \input[49]  = \input  [49];
  assign shiftLeftOnePos[49] = \input[48] ;
  assign \input[48]  = \input  [48];
  assign shiftLeftOnePos[48] = \input[47] ;
  assign \input[47]  = \input  [47];
  assign shiftLeftOnePos[47] = \input[46] ;
  assign \input[46]  = \input  [46];
  assign shiftLeftOnePos[46] = \input[45] ;
  assign \input[45]  = \input  [45];
  assign shiftLeftOnePos[45] = \input[44] ;
  assign \input[44]  = \input  [44];
  assign shiftLeftOnePos[44] = \input[43] ;
  assign \input[43]  = \input  [43];
  assign shiftLeftOnePos[43] = \input[42] ;
  assign \input[42]  = \input  [42];
  assign shiftLeftOnePos[42] = \input[41] ;
  assign \input[41]  = \input  [41];
  assign shiftLeftOnePos[41] = \input[40] ;
  assign \input[40]  = \input  [40];
  assign shiftLeftOnePos[40] = \input[39] ;
  assign \input[39]  = \input  [39];
  assign shiftLeftOnePos[39] = \input[38] ;
  assign \input[38]  = \input  [38];
  assign shiftLeftOnePos[38] = \input[37] ;
  assign \input[37]  = \input  [37];
  assign shiftLeftOnePos[37] = \input[36] ;
  assign \input[36]  = \input  [36];
  assign shiftLeftOnePos[36] = \input[35] ;
  assign \input[35]  = \input  [35];
  assign shiftLeftOnePos[35] = \input[34] ;
  assign \input[34]  = \input  [34];
  assign shiftLeftOnePos[34] = \input[33] ;
  assign \input[33]  = \input  [33];
  assign shiftLeftOnePos[33] = \input[32] ;
  assign \input[32]  = \input  [32];
  assign shiftLeftOnePos[32] = \input[31] ;
  assign \input[31]  = \input  [31];
  assign shiftLeftOnePos[31] = \input[30] ;
  assign \input[30]  = \input  [30];
  assign shiftLeftOnePos[30] = \input[29] ;
  assign \input[29]  = \input  [29];
  assign shiftLeftOnePos[29] = \input[28] ;
  assign \input[28]  = \input  [28];
  assign shiftLeftOnePos[28] = \input[27] ;
  assign \input[27]  = \input  [27];
  assign shiftLeftOnePos[27] = \input[26] ;
  assign \input[26]  = \input  [26];
  assign shiftLeftOnePos[26] = \input[25] ;
  assign \input[25]  = \input  [25];
  assign shiftLeftOnePos[25] = \input[24] ;
  assign \input[24]  = \input  [24];
  assign shiftLeftOnePos[24] = \input[23] ;
  assign \input[23]  = \input  [23];
  assign shiftLeftOnePos[23] = \input[22] ;
  assign \input[22]  = \input  [22];
  assign shiftLeftOnePos[22] = \input[21] ;
  assign \input[21]  = \input  [21];
  assign shiftLeftOnePos[21] = \input[20] ;
  assign \input[20]  = \input  [20];
  assign shiftLeftOnePos[20] = \input[19] ;
  assign \input[19]  = \input  [19];
  assign shiftLeftOnePos[19] = \input[18] ;
  assign \input[18]  = \input  [18];
  assign shiftLeftOnePos[18] = \input[17] ;
  assign \input[17]  = \input  [17];
  assign shiftLeftOnePos[17] = \input[16] ;
  assign \input[16]  = \input  [16];
  assign shiftLeftOnePos[16] = \input[15] ;
  assign \input[15]  = \input  [15];
  assign shiftLeftOnePos[15] = \input[14] ;
  assign \input[14]  = \input  [14];
  assign shiftLeftOnePos[14] = \input[13] ;
  assign \input[13]  = \input  [13];
  assign shiftLeftOnePos[13] = \input[12] ;
  assign \input[12]  = \input  [12];
  assign shiftLeftOnePos[12] = \input[11] ;
  assign \input[11]  = \input  [11];
  assign shiftLeftOnePos[11] = \input[10] ;
  assign \input[10]  = \input  [10];
  assign shiftLeftOnePos[10] = \input[9] ;
  assign \input[9]  = \input  [9];
  assign shiftLeftOnePos[9] = \input[8] ;
  assign \input[8]  = \input  [8];
  assign shiftLeftOnePos[8] = \input[7] ;
  assign \input[7]  = \input  [7];
  assign shiftLeftOnePos[7] = \input[6] ;
  assign \input[6]  = \input  [6];
  assign shiftLeftOnePos[6] = \input[5] ;
  assign \input[5]  = \input  [5];
  assign shiftLeftOnePos[5] = \input[4] ;
  assign \input[4]  = \input  [4];
  assign shiftLeftOnePos[4] = \input[3] ;
  assign \input[3]  = \input  [3];
  assign shiftLeftOnePos[3] = \input[2] ;
  assign \input[2]  = \input  [2];
  assign shiftLeftOnePos[2] = \input[1] ;
  assign \input[1]  = \input  [1];
  assign shiftLeftOnePos[1] = \input[0] ;
  assign \input[0]  = \input  [0];

endmodule


module shifter_N64_15 ( \input , shiftLeftOnePos );
  input [63:0] \input ;
  output [63:0] shiftLeftOnePos;
  wire   \input[62] , \input[61] , \input[60] , \input[59] , \input[58] ,
         \input[57] , \input[56] , \input[55] , \input[54] , \input[53] ,
         \input[52] , \input[51] , \input[50] , \input[49] , \input[48] ,
         \input[47] , \input[46] , \input[45] , \input[44] , \input[43] ,
         \input[42] , \input[41] , \input[40] , \input[39] , \input[38] ,
         \input[37] , \input[36] , \input[35] , \input[34] , \input[33] ,
         \input[32] , \input[31] , \input[30] , \input[29] , \input[28] ,
         \input[27] , \input[26] , \input[25] , \input[24] , \input[23] ,
         \input[22] , \input[21] , \input[20] , \input[19] , \input[18] ,
         \input[17] , \input[16] , \input[15] , \input[14] , \input[13] ,
         \input[12] , \input[11] , \input[10] , \input[9] , \input[8] ,
         \input[7] , \input[6] , \input[5] , \input[4] , \input[3] ,
         \input[2] , \input[1] , \input[0] ;
  assign shiftLeftOnePos[0] = 1'b0;
  assign shiftLeftOnePos[63] = \input[62] ;
  assign \input[62]  = \input  [62];
  assign shiftLeftOnePos[62] = \input[61] ;
  assign \input[61]  = \input  [61];
  assign shiftLeftOnePos[61] = \input[60] ;
  assign \input[60]  = \input  [60];
  assign shiftLeftOnePos[60] = \input[59] ;
  assign \input[59]  = \input  [59];
  assign shiftLeftOnePos[59] = \input[58] ;
  assign \input[58]  = \input  [58];
  assign shiftLeftOnePos[58] = \input[57] ;
  assign \input[57]  = \input  [57];
  assign shiftLeftOnePos[57] = \input[56] ;
  assign \input[56]  = \input  [56];
  assign shiftLeftOnePos[56] = \input[55] ;
  assign \input[55]  = \input  [55];
  assign shiftLeftOnePos[55] = \input[54] ;
  assign \input[54]  = \input  [54];
  assign shiftLeftOnePos[54] = \input[53] ;
  assign \input[53]  = \input  [53];
  assign shiftLeftOnePos[53] = \input[52] ;
  assign \input[52]  = \input  [52];
  assign shiftLeftOnePos[52] = \input[51] ;
  assign \input[51]  = \input  [51];
  assign shiftLeftOnePos[51] = \input[50] ;
  assign \input[50]  = \input  [50];
  assign shiftLeftOnePos[50] = \input[49] ;
  assign \input[49]  = \input  [49];
  assign shiftLeftOnePos[49] = \input[48] ;
  assign \input[48]  = \input  [48];
  assign shiftLeftOnePos[48] = \input[47] ;
  assign \input[47]  = \input  [47];
  assign shiftLeftOnePos[47] = \input[46] ;
  assign \input[46]  = \input  [46];
  assign shiftLeftOnePos[46] = \input[45] ;
  assign \input[45]  = \input  [45];
  assign shiftLeftOnePos[45] = \input[44] ;
  assign \input[44]  = \input  [44];
  assign shiftLeftOnePos[44] = \input[43] ;
  assign \input[43]  = \input  [43];
  assign shiftLeftOnePos[43] = \input[42] ;
  assign \input[42]  = \input  [42];
  assign shiftLeftOnePos[42] = \input[41] ;
  assign \input[41]  = \input  [41];
  assign shiftLeftOnePos[41] = \input[40] ;
  assign \input[40]  = \input  [40];
  assign shiftLeftOnePos[40] = \input[39] ;
  assign \input[39]  = \input  [39];
  assign shiftLeftOnePos[39] = \input[38] ;
  assign \input[38]  = \input  [38];
  assign shiftLeftOnePos[38] = \input[37] ;
  assign \input[37]  = \input  [37];
  assign shiftLeftOnePos[37] = \input[36] ;
  assign \input[36]  = \input  [36];
  assign shiftLeftOnePos[36] = \input[35] ;
  assign \input[35]  = \input  [35];
  assign shiftLeftOnePos[35] = \input[34] ;
  assign \input[34]  = \input  [34];
  assign shiftLeftOnePos[34] = \input[33] ;
  assign \input[33]  = \input  [33];
  assign shiftLeftOnePos[33] = \input[32] ;
  assign \input[32]  = \input  [32];
  assign shiftLeftOnePos[32] = \input[31] ;
  assign \input[31]  = \input  [31];
  assign shiftLeftOnePos[31] = \input[30] ;
  assign \input[30]  = \input  [30];
  assign shiftLeftOnePos[30] = \input[29] ;
  assign \input[29]  = \input  [29];
  assign shiftLeftOnePos[29] = \input[28] ;
  assign \input[28]  = \input  [28];
  assign shiftLeftOnePos[28] = \input[27] ;
  assign \input[27]  = \input  [27];
  assign shiftLeftOnePos[27] = \input[26] ;
  assign \input[26]  = \input  [26];
  assign shiftLeftOnePos[26] = \input[25] ;
  assign \input[25]  = \input  [25];
  assign shiftLeftOnePos[25] = \input[24] ;
  assign \input[24]  = \input  [24];
  assign shiftLeftOnePos[24] = \input[23] ;
  assign \input[23]  = \input  [23];
  assign shiftLeftOnePos[23] = \input[22] ;
  assign \input[22]  = \input  [22];
  assign shiftLeftOnePos[22] = \input[21] ;
  assign \input[21]  = \input  [21];
  assign shiftLeftOnePos[21] = \input[20] ;
  assign \input[20]  = \input  [20];
  assign shiftLeftOnePos[20] = \input[19] ;
  assign \input[19]  = \input  [19];
  assign shiftLeftOnePos[19] = \input[18] ;
  assign \input[18]  = \input  [18];
  assign shiftLeftOnePos[18] = \input[17] ;
  assign \input[17]  = \input  [17];
  assign shiftLeftOnePos[17] = \input[16] ;
  assign \input[16]  = \input  [16];
  assign shiftLeftOnePos[16] = \input[15] ;
  assign \input[15]  = \input  [15];
  assign shiftLeftOnePos[15] = \input[14] ;
  assign \input[14]  = \input  [14];
  assign shiftLeftOnePos[14] = \input[13] ;
  assign \input[13]  = \input  [13];
  assign shiftLeftOnePos[13] = \input[12] ;
  assign \input[12]  = \input  [12];
  assign shiftLeftOnePos[12] = \input[11] ;
  assign \input[11]  = \input  [11];
  assign shiftLeftOnePos[11] = \input[10] ;
  assign \input[10]  = \input  [10];
  assign shiftLeftOnePos[10] = \input[9] ;
  assign \input[9]  = \input  [9];
  assign shiftLeftOnePos[9] = \input[8] ;
  assign \input[8]  = \input  [8];
  assign shiftLeftOnePos[8] = \input[7] ;
  assign \input[7]  = \input  [7];
  assign shiftLeftOnePos[7] = \input[6] ;
  assign \input[6]  = \input  [6];
  assign shiftLeftOnePos[6] = \input[5] ;
  assign \input[5]  = \input  [5];
  assign shiftLeftOnePos[5] = \input[4] ;
  assign \input[4]  = \input  [4];
  assign shiftLeftOnePos[4] = \input[3] ;
  assign \input[3]  = \input  [3];
  assign shiftLeftOnePos[3] = \input[2] ;
  assign \input[2]  = \input  [2];
  assign shiftLeftOnePos[2] = \input[1] ;
  assign \input[1]  = \input  [1];
  assign shiftLeftOnePos[1] = \input[0] ;
  assign \input[0]  = \input  [0];

endmodule


module complementer_N64_16_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n189;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U81 ( .A(n190), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U82 ( .A(n192), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U83 ( .A(n193), .B(B[6]), .Z(DIFF[6]) );
  XOR2_X1 U84 ( .A(n195), .B(B[63]), .Z(DIFF[63]) );
  XOR2_X1 U85 ( .A(n196), .B(B[62]), .Z(DIFF[62]) );
  XOR2_X1 U86 ( .A(n194), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U87 ( .A(n198), .B(B[59]), .Z(DIFF[59]) );
  XOR2_X1 U88 ( .A(n201), .B(B[58]), .Z(DIFF[58]) );
  XOR2_X1 U89 ( .A(n200), .B(B[57]), .Z(DIFF[57]) );
  XOR2_X1 U90 ( .A(n202), .B(B[55]), .Z(DIFF[55]) );
  XOR2_X1 U91 ( .A(n205), .B(B[54]), .Z(DIFF[54]) );
  XOR2_X1 U92 ( .A(n204), .B(B[53]), .Z(DIFF[53]) );
  XOR2_X1 U93 ( .A(n206), .B(B[51]), .Z(DIFF[51]) );
  XOR2_X1 U94 ( .A(n209), .B(B[50]), .Z(DIFF[50]) );
  XOR2_X1 U95 ( .A(n208), .B(B[49]), .Z(DIFF[49]) );
  XOR2_X1 U96 ( .A(n212), .B(B[47]), .Z(DIFF[47]) );
  XOR2_X1 U97 ( .A(n215), .B(B[46]), .Z(DIFF[46]) );
  XOR2_X1 U98 ( .A(n214), .B(B[45]), .Z(DIFF[45]) );
  XOR2_X1 U99 ( .A(n216), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U100 ( .A(n219), .B(B[42]), .Z(DIFF[42]) );
  XOR2_X1 U101 ( .A(n218), .B(B[41]), .Z(DIFF[41]) );
  XOR2_X1 U102 ( .A(n211), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U103 ( .A(n220), .B(B[39]), .Z(DIFF[39]) );
  XOR2_X1 U104 ( .A(n223), .B(B[38]), .Z(DIFF[38]) );
  XOR2_X1 U105 ( .A(n222), .B(B[37]), .Z(DIFF[37]) );
  XOR2_X1 U106 ( .A(n224), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U107 ( .A(n227), .B(B[34]), .Z(DIFF[34]) );
  XOR2_X1 U108 ( .A(n226), .B(B[33]), .Z(DIFF[33]) );
  XOR2_X1 U109 ( .A(n228), .B(B[31]), .Z(DIFF[31]) );
  XOR2_X1 U110 ( .A(n231), .B(B[30]), .Z(DIFF[30]) );
  XOR2_X1 U111 ( .A(n230), .B(B[29]), .Z(DIFF[29]) );
  XOR2_X1 U112 ( .A(n233), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U113 ( .A(n236), .B(B[26]), .Z(DIFF[26]) );
  XOR2_X1 U114 ( .A(n235), .B(B[25]), .Z(DIFF[25]) );
  XOR2_X1 U115 ( .A(n237), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U116 ( .A(n240), .B(B[22]), .Z(DIFF[22]) );
  XOR2_X1 U117 ( .A(n239), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U118 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U119 ( .A(n241), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U120 ( .A(n244), .B(B[18]), .Z(DIFF[18]) );
  XOR2_X1 U121 ( .A(n243), .B(B[17]), .Z(DIFF[17]) );
  XOR2_X1 U122 ( .A(n245), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U123 ( .A(n248), .B(B[14]), .Z(DIFF[14]) );
  XOR2_X1 U124 ( .A(n247), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U125 ( .A(n249), .B(B[11]), .Z(DIFF[11]) );
  XOR2_X1 U126 ( .A(n251), .B(B[10]), .Z(DIFF[10]) );
  OR3_X1 U1 ( .A1(B[53]), .A2(B[54]), .A3(n204), .ZN(n202) );
  OR2_X1 U2 ( .A1(n204), .A2(B[53]), .ZN(n205) );
  NOR2_X1 U3 ( .A1(B[59]), .A2(n198), .ZN(n199) );
  NAND2_X1 U4 ( .A1(n197), .A2(n189), .ZN(n196) );
  NOR2_X1 U5 ( .A1(B[51]), .A2(n206), .ZN(n207) );
  OR3_X1 U6 ( .A1(B[49]), .A2(B[50]), .A3(n208), .ZN(n206) );
  OR3_X1 U7 ( .A1(B[51]), .A2(B[52]), .A3(n206), .ZN(n204) );
  OR2_X1 U8 ( .A1(n208), .A2(B[49]), .ZN(n209) );
  NOR3_X1 U9 ( .A1(B[59]), .A2(B[60]), .A3(n198), .ZN(n197) );
  NOR2_X1 U10 ( .A1(B[55]), .A2(n202), .ZN(n203) );
  OR3_X1 U11 ( .A1(B[57]), .A2(B[58]), .A3(n200), .ZN(n198) );
  OR3_X1 U12 ( .A1(B[55]), .A2(B[56]), .A3(n202), .ZN(n200) );
  OR2_X1 U13 ( .A1(n200), .A2(B[57]), .ZN(n201) );
  OR2_X1 U14 ( .A1(n196), .A2(B[62]), .ZN(n195) );
  NOR2_X1 U15 ( .A1(B[47]), .A2(n212), .ZN(n213) );
  OR3_X1 U16 ( .A1(B[47]), .A2(B[48]), .A3(n212), .ZN(n208) );
  XNOR2_X1 U17 ( .A(B[24]), .B(n238), .ZN(DIFF[24]) );
  XNOR2_X1 U18 ( .A(B[20]), .B(n242), .ZN(DIFF[20]) );
  NOR2_X1 U19 ( .A1(B[27]), .A2(n233), .ZN(n234) );
  NOR2_X1 U20 ( .A1(B[23]), .A2(n237), .ZN(n238) );
  OR3_X1 U21 ( .A1(B[25]), .A2(B[26]), .A3(n235), .ZN(n233) );
  OR3_X1 U22 ( .A1(B[21]), .A2(B[22]), .A3(n239), .ZN(n237) );
  OR3_X1 U23 ( .A1(B[27]), .A2(B[28]), .A3(n233), .ZN(n230) );
  OR3_X1 U24 ( .A1(B[23]), .A2(B[24]), .A3(n237), .ZN(n235) );
  XNOR2_X1 U25 ( .A(B[28]), .B(n234), .ZN(DIFF[28]) );
  OR2_X1 U26 ( .A1(n230), .A2(B[29]), .ZN(n231) );
  OR2_X1 U27 ( .A1(n235), .A2(B[25]), .ZN(n236) );
  OR2_X1 U28 ( .A1(n239), .A2(B[21]), .ZN(n240) );
  NOR2_X1 U29 ( .A1(B[43]), .A2(n216), .ZN(n217) );
  NOR2_X1 U30 ( .A1(B[39]), .A2(n220), .ZN(n221) );
  NOR2_X1 U31 ( .A1(B[35]), .A2(n224), .ZN(n225) );
  NOR2_X1 U32 ( .A1(B[31]), .A2(n228), .ZN(n229) );
  OR3_X1 U33 ( .A1(B[45]), .A2(B[46]), .A3(n214), .ZN(n212) );
  OR3_X1 U34 ( .A1(B[41]), .A2(B[42]), .A3(n218), .ZN(n216) );
  OR3_X1 U35 ( .A1(B[37]), .A2(B[38]), .A3(n222), .ZN(n220) );
  OR3_X1 U36 ( .A1(B[33]), .A2(B[34]), .A3(n226), .ZN(n224) );
  OR3_X1 U37 ( .A1(B[29]), .A2(B[30]), .A3(n230), .ZN(n228) );
  OR3_X1 U38 ( .A1(B[43]), .A2(B[44]), .A3(n216), .ZN(n214) );
  OR3_X1 U39 ( .A1(B[39]), .A2(B[40]), .A3(n220), .ZN(n218) );
  OR3_X1 U40 ( .A1(B[35]), .A2(B[36]), .A3(n224), .ZN(n222) );
  OR3_X1 U41 ( .A1(B[31]), .A2(B[32]), .A3(n228), .ZN(n226) );
  XNOR2_X1 U42 ( .A(B[48]), .B(n213), .ZN(DIFF[48]) );
  XNOR2_X1 U43 ( .A(B[56]), .B(n203), .ZN(DIFF[56]) );
  XNOR2_X1 U44 ( .A(B[52]), .B(n207), .ZN(DIFF[52]) );
  XNOR2_X1 U45 ( .A(B[44]), .B(n217), .ZN(DIFF[44]) );
  XNOR2_X1 U46 ( .A(B[40]), .B(n221), .ZN(DIFF[40]) );
  XNOR2_X1 U47 ( .A(B[36]), .B(n225), .ZN(DIFF[36]) );
  XNOR2_X1 U48 ( .A(B[32]), .B(n229), .ZN(DIFF[32]) );
  OR2_X1 U49 ( .A1(n214), .A2(B[45]), .ZN(n215) );
  OR2_X1 U50 ( .A1(n218), .A2(B[41]), .ZN(n219) );
  OR2_X1 U51 ( .A1(n222), .A2(B[37]), .ZN(n223) );
  OR2_X1 U52 ( .A1(n226), .A2(B[33]), .ZN(n227) );
  XNOR2_X1 U53 ( .A(n197), .B(B[61]), .ZN(DIFF[61]) );
  XNOR2_X1 U54 ( .A(B[60]), .B(n199), .ZN(DIFF[60]) );
  NOR2_X1 U55 ( .A1(B[19]), .A2(n241), .ZN(n242) );
  OR3_X1 U56 ( .A1(B[19]), .A2(B[20]), .A3(n241), .ZN(n239) );
  OR3_X1 U57 ( .A1(B[17]), .A2(B[18]), .A3(n243), .ZN(n241) );
  OR2_X1 U58 ( .A1(n243), .A2(B[17]), .ZN(n244) );
  OR3_X1 U59 ( .A1(B[15]), .A2(B[16]), .A3(n245), .ZN(n243) );
  XNOR2_X1 U60 ( .A(B[16]), .B(n246), .ZN(DIFF[16]) );
  NOR2_X1 U61 ( .A1(B[15]), .A2(n245), .ZN(n246) );
  NOR2_X1 U62 ( .A1(B[11]), .A2(n249), .ZN(n250) );
  NOR2_X1 U63 ( .A1(B[7]), .A2(n192), .ZN(n191) );
  NOR2_X1 U64 ( .A1(B[3]), .A2(n211), .ZN(n210) );
  OR3_X1 U65 ( .A1(B[13]), .A2(B[14]), .A3(n247), .ZN(n245) );
  OR3_X1 U66 ( .A1(B[10]), .A2(B[9]), .A3(n190), .ZN(n249) );
  OR3_X1 U67 ( .A1(B[5]), .A2(B[6]), .A3(n194), .ZN(n192) );
  OR3_X1 U68 ( .A1(B[11]), .A2(B[12]), .A3(n249), .ZN(n247) );
  OR3_X1 U69 ( .A1(B[7]), .A2(B[8]), .A3(n192), .ZN(n190) );
  OR3_X1 U70 ( .A1(B[3]), .A2(B[4]), .A3(n211), .ZN(n194) );
  XNOR2_X1 U71 ( .A(B[12]), .B(n250), .ZN(DIFF[12]) );
  XNOR2_X1 U72 ( .A(B[8]), .B(n191), .ZN(DIFF[8]) );
  XNOR2_X1 U73 ( .A(B[4]), .B(n210), .ZN(DIFF[4]) );
  XNOR2_X1 U74 ( .A(B[2]), .B(n232), .ZN(DIFF[2]) );
  OR2_X1 U75 ( .A1(n247), .A2(B[13]), .ZN(n248) );
  OR2_X1 U76 ( .A1(n190), .A2(B[9]), .ZN(n251) );
  OR2_X1 U77 ( .A1(n194), .A2(B[5]), .ZN(n193) );
  OR3_X1 U78 ( .A1(B[1]), .A2(B[2]), .A3(\B[0] ), .ZN(n211) );
  NOR2_X1 U79 ( .A1(\B[0] ), .A2(B[1]), .ZN(n232) );
  INV_X1 U80 ( .A(B[61]), .ZN(n189) );
endmodule


module complementer_N64_16 ( \input , complement2 );
  input [63:0] \input ;
  output [63:0] complement2;


  complementer_N64_16_DW01_sub_0 sub_add_31_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(\input ), .CI(1'b0), .DIFF(complement2) );
endmodule


module complementer_N64_15_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n190, n191, n192, n194, n196, n197, n198, n199, n200, n202,
         n203, n204, n206, n207, n208, n210, n211, n212, n213, n214, n216,
         n217, n218, n220, n221, n222, n224, n225, n226, n228, n229, n230,
         n232, n233, n234, n235, n237, n238, n239, n241, n242, n243, n245,
         n246, n247, n249, n250, n189, n193, n195, n201, n205, n209, n215,
         n219, n223, n227, n231, n236, n240, n244, n248, n251;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U81 ( .A(n190), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U82 ( .A(n192), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U85 ( .A(n196), .B(B[62]), .Z(DIFF[62]) );
  XOR2_X1 U86 ( .A(n194), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U87 ( .A(n198), .B(B[59]), .Z(DIFF[59]) );
  XOR2_X1 U89 ( .A(n200), .B(B[57]), .Z(DIFF[57]) );
  XOR2_X1 U90 ( .A(n202), .B(B[55]), .Z(DIFF[55]) );
  XOR2_X1 U92 ( .A(n204), .B(B[53]), .Z(DIFF[53]) );
  XOR2_X1 U93 ( .A(n206), .B(B[51]), .Z(DIFF[51]) );
  XOR2_X1 U95 ( .A(n208), .B(B[49]), .Z(DIFF[49]) );
  XOR2_X1 U96 ( .A(n212), .B(B[47]), .Z(DIFF[47]) );
  XOR2_X1 U98 ( .A(n214), .B(B[45]), .Z(DIFF[45]) );
  XOR2_X1 U99 ( .A(n216), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U101 ( .A(n218), .B(B[41]), .Z(DIFF[41]) );
  XOR2_X1 U102 ( .A(n211), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U103 ( .A(n220), .B(B[39]), .Z(DIFF[39]) );
  XOR2_X1 U105 ( .A(n222), .B(B[37]), .Z(DIFF[37]) );
  XOR2_X1 U106 ( .A(n224), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U108 ( .A(n226), .B(B[33]), .Z(DIFF[33]) );
  XOR2_X1 U109 ( .A(n228), .B(B[31]), .Z(DIFF[31]) );
  XOR2_X1 U111 ( .A(n230), .B(B[29]), .Z(DIFF[29]) );
  XOR2_X1 U112 ( .A(n233), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U114 ( .A(n235), .B(B[25]), .Z(DIFF[25]) );
  XOR2_X1 U115 ( .A(n237), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U117 ( .A(n239), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U118 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U119 ( .A(n241), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U121 ( .A(n243), .B(B[17]), .Z(DIFF[17]) );
  XOR2_X1 U122 ( .A(n245), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U124 ( .A(n247), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U125 ( .A(n249), .B(B[11]), .Z(DIFF[11]) );
  OR3_X1 U1 ( .A1(B[53]), .A2(B[54]), .A3(n204), .ZN(n202) );
  XNOR2_X1 U2 ( .A(n189), .B(B[54]), .ZN(DIFF[54]) );
  NOR2_X1 U3 ( .A1(n204), .A2(B[53]), .ZN(n189) );
  NOR3_X1 U4 ( .A1(B[59]), .A2(B[60]), .A3(n198), .ZN(n197) );
  XNOR2_X1 U5 ( .A(B[60]), .B(n199), .ZN(DIFF[60]) );
  NOR2_X1 U6 ( .A1(B[59]), .A2(n198), .ZN(n199) );
  XOR2_X1 U7 ( .A(n197), .B(n251), .Z(DIFF[61]) );
  NAND2_X1 U8 ( .A1(n197), .A2(n251), .ZN(n196) );
  XNOR2_X1 U9 ( .A(B[56]), .B(n203), .ZN(DIFF[56]) );
  NOR2_X1 U10 ( .A1(B[55]), .A2(n202), .ZN(n203) );
  XNOR2_X1 U11 ( .A(B[52]), .B(n207), .ZN(DIFF[52]) );
  NOR2_X1 U12 ( .A1(B[51]), .A2(n206), .ZN(n207) );
  OR3_X1 U13 ( .A1(B[49]), .A2(B[50]), .A3(n208), .ZN(n206) );
  OR3_X1 U14 ( .A1(B[51]), .A2(B[52]), .A3(n206), .ZN(n204) );
  XNOR2_X1 U15 ( .A(n193), .B(B[50]), .ZN(DIFF[50]) );
  NOR2_X1 U16 ( .A1(n208), .A2(B[49]), .ZN(n193) );
  OR3_X1 U17 ( .A1(B[57]), .A2(B[58]), .A3(n200), .ZN(n198) );
  OR3_X1 U18 ( .A1(B[55]), .A2(B[56]), .A3(n202), .ZN(n200) );
  XNOR2_X1 U19 ( .A(n195), .B(B[58]), .ZN(DIFF[58]) );
  NOR2_X1 U20 ( .A1(n200), .A2(B[57]), .ZN(n195) );
  XNOR2_X1 U21 ( .A(n201), .B(B[63]), .ZN(DIFF[63]) );
  NOR2_X1 U22 ( .A1(n196), .A2(B[62]), .ZN(n201) );
  XNOR2_X1 U23 ( .A(B[28]), .B(n234), .ZN(DIFF[28]) );
  NOR2_X1 U24 ( .A1(B[27]), .A2(n233), .ZN(n234) );
  XNOR2_X1 U25 ( .A(B[24]), .B(n238), .ZN(DIFF[24]) );
  NOR2_X1 U26 ( .A1(B[23]), .A2(n237), .ZN(n238) );
  OR3_X1 U27 ( .A1(B[25]), .A2(B[26]), .A3(n235), .ZN(n233) );
  OR3_X1 U28 ( .A1(B[29]), .A2(B[30]), .A3(n230), .ZN(n228) );
  OR3_X1 U29 ( .A1(B[23]), .A2(B[24]), .A3(n237), .ZN(n235) );
  OR3_X1 U30 ( .A1(B[27]), .A2(B[28]), .A3(n233), .ZN(n230) );
  XNOR2_X1 U31 ( .A(n205), .B(B[30]), .ZN(DIFF[30]) );
  NOR2_X1 U32 ( .A1(n230), .A2(B[29]), .ZN(n205) );
  XNOR2_X1 U33 ( .A(n209), .B(B[26]), .ZN(DIFF[26]) );
  NOR2_X1 U34 ( .A1(n235), .A2(B[25]), .ZN(n209) );
  XNOR2_X1 U35 ( .A(B[48]), .B(n213), .ZN(DIFF[48]) );
  NOR2_X1 U36 ( .A1(B[47]), .A2(n212), .ZN(n213) );
  XNOR2_X1 U37 ( .A(B[44]), .B(n217), .ZN(DIFF[44]) );
  NOR2_X1 U38 ( .A1(B[43]), .A2(n216), .ZN(n217) );
  XNOR2_X1 U39 ( .A(B[40]), .B(n221), .ZN(DIFF[40]) );
  NOR2_X1 U40 ( .A1(B[39]), .A2(n220), .ZN(n221) );
  XNOR2_X1 U41 ( .A(B[36]), .B(n225), .ZN(DIFF[36]) );
  NOR2_X1 U42 ( .A1(B[35]), .A2(n224), .ZN(n225) );
  XNOR2_X1 U43 ( .A(B[32]), .B(n229), .ZN(DIFF[32]) );
  NOR2_X1 U44 ( .A1(B[31]), .A2(n228), .ZN(n229) );
  OR3_X1 U45 ( .A1(B[33]), .A2(B[34]), .A3(n226), .ZN(n224) );
  OR3_X1 U46 ( .A1(B[37]), .A2(B[38]), .A3(n222), .ZN(n220) );
  OR3_X1 U47 ( .A1(B[41]), .A2(B[42]), .A3(n218), .ZN(n216) );
  OR3_X1 U48 ( .A1(B[45]), .A2(B[46]), .A3(n214), .ZN(n212) );
  OR3_X1 U49 ( .A1(B[31]), .A2(B[32]), .A3(n228), .ZN(n226) );
  OR3_X1 U50 ( .A1(B[35]), .A2(B[36]), .A3(n224), .ZN(n222) );
  OR3_X1 U51 ( .A1(B[39]), .A2(B[40]), .A3(n220), .ZN(n218) );
  OR3_X1 U52 ( .A1(B[43]), .A2(B[44]), .A3(n216), .ZN(n214) );
  OR3_X1 U53 ( .A1(B[47]), .A2(B[48]), .A3(n212), .ZN(n208) );
  XNOR2_X1 U54 ( .A(n215), .B(B[46]), .ZN(DIFF[46]) );
  NOR2_X1 U55 ( .A1(n214), .A2(B[45]), .ZN(n215) );
  XNOR2_X1 U56 ( .A(n219), .B(B[42]), .ZN(DIFF[42]) );
  NOR2_X1 U57 ( .A1(n218), .A2(B[41]), .ZN(n219) );
  XNOR2_X1 U58 ( .A(n223), .B(B[38]), .ZN(DIFF[38]) );
  NOR2_X1 U59 ( .A1(n222), .A2(B[37]), .ZN(n223) );
  XNOR2_X1 U60 ( .A(n227), .B(B[34]), .ZN(DIFF[34]) );
  NOR2_X1 U61 ( .A1(n226), .A2(B[33]), .ZN(n227) );
  XNOR2_X1 U62 ( .A(n231), .B(B[22]), .ZN(DIFF[22]) );
  NOR2_X1 U63 ( .A1(n239), .A2(B[21]), .ZN(n231) );
  OR3_X1 U64 ( .A1(B[21]), .A2(B[22]), .A3(n239), .ZN(n237) );
  XNOR2_X1 U65 ( .A(B[20]), .B(n242), .ZN(DIFF[20]) );
  NOR2_X1 U66 ( .A1(B[19]), .A2(n241), .ZN(n242) );
  OR3_X1 U67 ( .A1(B[19]), .A2(B[20]), .A3(n241), .ZN(n239) );
  XNOR2_X1 U68 ( .A(n236), .B(B[18]), .ZN(DIFF[18]) );
  NOR2_X1 U69 ( .A1(n243), .A2(B[17]), .ZN(n236) );
  OR3_X1 U70 ( .A1(B[17]), .A2(B[18]), .A3(n243), .ZN(n241) );
  XNOR2_X1 U71 ( .A(B[16]), .B(n246), .ZN(DIFF[16]) );
  XNOR2_X1 U72 ( .A(n240), .B(B[14]), .ZN(DIFF[14]) );
  NOR2_X1 U73 ( .A1(n247), .A2(B[13]), .ZN(n240) );
  XNOR2_X1 U74 ( .A(n244), .B(B[10]), .ZN(DIFF[10]) );
  NOR2_X1 U75 ( .A1(n190), .A2(B[9]), .ZN(n244) );
  XNOR2_X1 U76 ( .A(n248), .B(B[6]), .ZN(DIFF[6]) );
  NOR2_X1 U77 ( .A1(n194), .A2(B[5]), .ZN(n248) );
  NOR2_X1 U78 ( .A1(B[15]), .A2(n245), .ZN(n246) );
  XNOR2_X1 U79 ( .A(B[12]), .B(n250), .ZN(DIFF[12]) );
  NOR2_X1 U80 ( .A1(B[11]), .A2(n249), .ZN(n250) );
  XNOR2_X1 U83 ( .A(B[8]), .B(n191), .ZN(DIFF[8]) );
  NOR2_X1 U84 ( .A1(B[7]), .A2(n192), .ZN(n191) );
  XNOR2_X1 U88 ( .A(B[2]), .B(n232), .ZN(DIFF[2]) );
  NOR2_X1 U91 ( .A1(\B[0] ), .A2(B[1]), .ZN(n232) );
  XNOR2_X1 U94 ( .A(B[4]), .B(n210), .ZN(DIFF[4]) );
  NOR2_X1 U97 ( .A1(B[3]), .A2(n211), .ZN(n210) );
  OR3_X1 U100 ( .A1(B[5]), .A2(B[6]), .A3(n194), .ZN(n192) );
  OR3_X1 U104 ( .A1(B[10]), .A2(B[9]), .A3(n190), .ZN(n249) );
  OR3_X1 U107 ( .A1(B[13]), .A2(B[14]), .A3(n247), .ZN(n245) );
  OR3_X1 U110 ( .A1(B[7]), .A2(B[8]), .A3(n192), .ZN(n190) );
  OR3_X1 U113 ( .A1(B[11]), .A2(B[12]), .A3(n249), .ZN(n247) );
  OR3_X1 U116 ( .A1(B[15]), .A2(B[16]), .A3(n245), .ZN(n243) );
  OR3_X1 U120 ( .A1(B[3]), .A2(B[4]), .A3(n211), .ZN(n194) );
  OR3_X1 U123 ( .A1(B[1]), .A2(B[2]), .A3(\B[0] ), .ZN(n211) );
  INV_X1 U126 ( .A(B[61]), .ZN(n251) );
endmodule


module complementer_N64_15 ( \input , complement2 );
  input [63:0] \input ;
  output [63:0] complement2;


  complementer_N64_15_DW01_sub_0 sub_add_31_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(\input ), .CI(1'b0), .DIFF(complement2) );
endmodule


module ShiftnCompl_N64_8 ( plusA, plus2A_out, minus2A_out, plus4A_out, 
        minus4A_out );
  input [63:0] plusA;
  output [63:0] plus2A_out;
  output [63:0] minus2A_out;
  output [63:0] plus4A_out;
  output [63:0] minus4A_out;
  wire   n40, n41, n2, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign plus2A_out[0] = 1'b0;
  assign plus2A_out[51] = n2;
  assign plus4A_out[0] = 1'b0;

  shifter_N64_16 shifter_1 ( .\input (plusA), .shiftLeftOnePos({
        plus2A_out[63:59], n40, plus2A_out[57:54], n41, plus2A_out[52], n2, 
        plus2A_out[50:49], n42, n43, n44, plus2A_out[45:1], 
        SYNOPSYS_UNCONNECTED__0}) );
  shifter_N64_15 shifter_2 ( .\input ({plus2A_out[63:52], n2, plus2A_out[50:1], 
        1'b0}), .shiftLeftOnePos({plus4A_out[63:59], n45, plus4A_out[57:54], 
        n46, plus4A_out[52:47], n47, n48, n49, n50, n51, n52, n53, n54, n55, 
        n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, 
        n70, n71, n72, n73, n74, n75, n76, plus4A_out[16:1], 
        SYNOPSYS_UNCONNECTED__1}) );
  complementer_N64_16 complementer_1 ( .\input ({plus2A_out[63:52], n2, 
        plus2A_out[50:1], 1'b0}), .complement2(minus2A_out) );
  complementer_N64_15 complementer_2 ( .\input ({plus4A_out[63:1], 1'b0}), 
        .complement2(minus4A_out) );
  BUF_X1 U1 ( .A(n46), .Z(plus4A_out[53]) );
  BUF_X1 U4 ( .A(n62), .Z(plus4A_out[31]) );
  BUF_X1 U5 ( .A(n66), .Z(plus4A_out[27]) );
  BUF_X1 U6 ( .A(n64), .Z(plus4A_out[29]) );
  BUF_X1 U7 ( .A(n68), .Z(plus4A_out[25]) );
  BUF_X1 U8 ( .A(n69), .Z(plus4A_out[24]) );
  BUF_X1 U9 ( .A(n54), .Z(plus4A_out[39]) );
  BUF_X1 U10 ( .A(n58), .Z(plus4A_out[35]) );
  BUF_X1 U11 ( .A(n52), .Z(plus4A_out[41]) );
  BUF_X1 U12 ( .A(n56), .Z(plus4A_out[37]) );
  BUF_X1 U13 ( .A(n60), .Z(plus4A_out[33]) );
  BUF_X1 U14 ( .A(n51), .Z(plus4A_out[42]) );
  BUF_X1 U15 ( .A(n55), .Z(plus4A_out[38]) );
  BUF_X1 U16 ( .A(n59), .Z(plus4A_out[34]) );
  BUF_X1 U17 ( .A(n53), .Z(plus4A_out[40]) );
  BUF_X1 U18 ( .A(n57), .Z(plus4A_out[36]) );
  BUF_X1 U19 ( .A(n50), .Z(plus4A_out[43]) );
  BUF_X1 U20 ( .A(n48), .Z(plus4A_out[45]) );
  BUF_X1 U21 ( .A(n47), .Z(plus4A_out[46]) );
  BUF_X1 U22 ( .A(n44), .Z(plus2A_out[46]) );
  BUF_X1 U23 ( .A(n49), .Z(plus4A_out[44]) );
  BUF_X1 U24 ( .A(n43), .Z(plus2A_out[47]) );
  BUF_X1 U25 ( .A(n41), .Z(plus2A_out[53]) );
  BUF_X1 U26 ( .A(n42), .Z(plus2A_out[48]) );
  BUF_X1 U27 ( .A(n45), .Z(plus4A_out[58]) );
  BUF_X1 U28 ( .A(n40), .Z(plus2A_out[58]) );
  BUF_X1 U29 ( .A(n70), .Z(plus4A_out[23]) );
  BUF_X1 U30 ( .A(n74), .Z(plus4A_out[19]) );
  BUF_X1 U31 ( .A(n72), .Z(plus4A_out[21]) );
  BUF_X1 U32 ( .A(n76), .Z(plus4A_out[17]) );
  BUF_X1 U33 ( .A(n73), .Z(plus4A_out[20]) );
  BUF_X1 U34 ( .A(n71), .Z(plus4A_out[22]) );
  BUF_X1 U35 ( .A(n75), .Z(plus4A_out[18]) );
  BUF_X1 U36 ( .A(n61), .Z(plus4A_out[32]) );
  BUF_X1 U37 ( .A(n65), .Z(plus4A_out[28]) );
  BUF_X1 U38 ( .A(n63), .Z(plus4A_out[30]) );
  BUF_X1 U39 ( .A(n67), .Z(plus4A_out[26]) );
endmodule


module MUX_GENERIC_N64_RADIX3_8 ( plusA, minusA, plus2A, minus2A, SEL, Y );
  input [63:0] plusA;
  input [63:0] minusA;
  input [63:0] plus2A;
  input [63:0] minus2A;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502;
  tri   [63:0] Y;

  TBUF_X1 \Y_tri[57]  ( .A(n444), .EN(n301), .Z(Y[57]) );
  TBUF_X1 \Y_tri[58]  ( .A(n443), .EN(n301), .Z(Y[58]) );
  TBUF_X1 \Y_tri[59]  ( .A(n442), .EN(n301), .Z(Y[59]) );
  TBUF_X1 \Y_tri[60]  ( .A(n441), .EN(n301), .Z(Y[60]) );
  TBUF_X1 \Y_tri[61]  ( .A(n440), .EN(n301), .Z(Y[61]) );
  TBUF_X1 \Y_tri[62]  ( .A(n439), .EN(n301), .Z(Y[62]) );
  TBUF_X1 \Y_tri[63]  ( .A(n438), .EN(n301), .Z(Y[63]) );
  TBUF_X1 \Y_tri[55]  ( .A(n446), .EN(n301), .Z(Y[55]) );
  TBUF_X1 \Y_tri[56]  ( .A(n445), .EN(n301), .Z(Y[56]) );
  TBUF_X1 \Y_tri[32]  ( .A(n469), .EN(n298), .Z(Y[32]) );
  TBUF_X1 \Y_tri[33]  ( .A(n468), .EN(n299), .Z(Y[33]) );
  TBUF_X1 \Y_tri[34]  ( .A(n467), .EN(n299), .Z(Y[34]) );
  TBUF_X1 \Y_tri[35]  ( .A(n466), .EN(n299), .Z(Y[35]) );
  TBUF_X1 \Y_tri[36]  ( .A(n465), .EN(n299), .Z(Y[36]) );
  TBUF_X1 \Y_tri[37]  ( .A(n464), .EN(n299), .Z(Y[37]) );
  TBUF_X1 \Y_tri[38]  ( .A(n463), .EN(n299), .Z(Y[38]) );
  TBUF_X1 \Y_tri[39]  ( .A(n462), .EN(n299), .Z(Y[39]) );
  TBUF_X1 \Y_tri[40]  ( .A(n461), .EN(n299), .Z(Y[40]) );
  TBUF_X1 \Y_tri[41]  ( .A(n460), .EN(n299), .Z(Y[41]) );
  TBUF_X1 \Y_tri[42]  ( .A(n459), .EN(n299), .Z(Y[42]) );
  TBUF_X1 \Y_tri[43]  ( .A(n458), .EN(n299), .Z(Y[43]) );
  TBUF_X1 \Y_tri[44]  ( .A(n457), .EN(n300), .Z(Y[44]) );
  TBUF_X1 \Y_tri[45]  ( .A(n456), .EN(n300), .Z(Y[45]) );
  TBUF_X1 \Y_tri[46]  ( .A(n455), .EN(n300), .Z(Y[46]) );
  TBUF_X1 \Y_tri[47]  ( .A(n454), .EN(n300), .Z(Y[47]) );
  TBUF_X1 \Y_tri[48]  ( .A(n453), .EN(n300), .Z(Y[48]) );
  TBUF_X1 \Y_tri[49]  ( .A(n452), .EN(n300), .Z(Y[49]) );
  TBUF_X1 \Y_tri[50]  ( .A(n451), .EN(n300), .Z(Y[50]) );
  TBUF_X1 \Y_tri[51]  ( .A(n450), .EN(n300), .Z(Y[51]) );
  TBUF_X1 \Y_tri[52]  ( .A(n449), .EN(n300), .Z(Y[52]) );
  TBUF_X1 \Y_tri[53]  ( .A(n448), .EN(n300), .Z(Y[53]) );
  TBUF_X1 \Y_tri[54]  ( .A(n447), .EN(n300), .Z(Y[54]) );
  TBUF_X1 \Y_tri[11]  ( .A(n490), .EN(n297), .Z(Y[11]) );
  TBUF_X1 \Y_tri[12]  ( .A(n489), .EN(n297), .Z(Y[12]) );
  TBUF_X1 \Y_tri[13]  ( .A(n488), .EN(n297), .Z(Y[13]) );
  TBUF_X1 \Y_tri[14]  ( .A(n487), .EN(n297), .Z(Y[14]) );
  TBUF_X1 \Y_tri[15]  ( .A(n486), .EN(n297), .Z(Y[15]) );
  TBUF_X1 \Y_tri[16]  ( .A(n485), .EN(n297), .Z(Y[16]) );
  TBUF_X1 \Y_tri[17]  ( .A(n484), .EN(n297), .Z(Y[17]) );
  TBUF_X1 \Y_tri[18]  ( .A(n483), .EN(n297), .Z(Y[18]) );
  TBUF_X1 \Y_tri[19]  ( .A(n482), .EN(n297), .Z(Y[19]) );
  TBUF_X1 \Y_tri[20]  ( .A(n481), .EN(n297), .Z(Y[20]) );
  TBUF_X1 \Y_tri[21]  ( .A(n480), .EN(n297), .Z(Y[21]) );
  TBUF_X1 \Y_tri[22]  ( .A(n479), .EN(n298), .Z(Y[22]) );
  TBUF_X1 \Y_tri[23]  ( .A(n478), .EN(n298), .Z(Y[23]) );
  TBUF_X1 \Y_tri[24]  ( .A(n477), .EN(n298), .Z(Y[24]) );
  TBUF_X1 \Y_tri[25]  ( .A(n476), .EN(n298), .Z(Y[25]) );
  TBUF_X1 \Y_tri[26]  ( .A(n475), .EN(n298), .Z(Y[26]) );
  TBUF_X1 \Y_tri[27]  ( .A(n474), .EN(n298), .Z(Y[27]) );
  TBUF_X1 \Y_tri[28]  ( .A(n473), .EN(n298), .Z(Y[28]) );
  TBUF_X1 \Y_tri[29]  ( .A(n472), .EN(n298), .Z(Y[29]) );
  TBUF_X1 \Y_tri[30]  ( .A(n471), .EN(n298), .Z(Y[30]) );
  TBUF_X1 \Y_tri[31]  ( .A(n470), .EN(n298), .Z(Y[31]) );
  TBUF_X1 \Y_tri[0]  ( .A(n502), .EN(n296), .Z(Y[0]) );
  TBUF_X1 \Y_tri[1]  ( .A(n501), .EN(n296), .Z(Y[1]) );
  TBUF_X1 \Y_tri[3]  ( .A(n499), .EN(n296), .Z(Y[3]) );
  TBUF_X1 \Y_tri[4]  ( .A(n498), .EN(n296), .Z(Y[4]) );
  TBUF_X1 \Y_tri[5]  ( .A(n497), .EN(n296), .Z(Y[5]) );
  TBUF_X1 \Y_tri[6]  ( .A(n496), .EN(n296), .Z(Y[6]) );
  TBUF_X1 \Y_tri[7]  ( .A(n495), .EN(n296), .Z(Y[7]) );
  TBUF_X1 \Y_tri[8]  ( .A(n494), .EN(n296), .Z(Y[8]) );
  TBUF_X1 \Y_tri[9]  ( .A(n492), .EN(n296), .Z(Y[9]) );
  TBUF_X1 \Y_tri[10]  ( .A(n491), .EN(n296), .Z(Y[10]) );
  TBUF_X1 \Y_tri[2]  ( .A(n500), .EN(n296), .Z(Y[2]) );
  NAND2_X1 U2 ( .A1(n355), .A2(n354), .ZN(n477) );
  AOI22_X1 U3 ( .A1(plusA[24]), .A2(n280), .B1(plus2A[24]), .B2(n274), .ZN(
        n355) );
  AOI22_X1 U4 ( .A1(minus2A[24]), .A2(n292), .B1(minusA[24]), .B2(n286), .ZN(
        n354) );
  NAND2_X1 U5 ( .A1(n347), .A2(n346), .ZN(n481) );
  AOI22_X1 U6 ( .A1(plusA[20]), .A2(n279), .B1(plus2A[20]), .B2(n273), .ZN(
        n347) );
  AOI22_X1 U7 ( .A1(minus2A[20]), .A2(n291), .B1(minusA[20]), .B2(n285), .ZN(
        n346) );
  NAND2_X1 U8 ( .A1(n369), .A2(n368), .ZN(n470) );
  AOI22_X1 U9 ( .A1(plusA[31]), .A2(n280), .B1(plus2A[31]), .B2(n274), .ZN(
        n369) );
  AOI22_X1 U10 ( .A1(minus2A[31]), .A2(n292), .B1(minusA[31]), .B2(n286), .ZN(
        n368) );
  NAND2_X1 U11 ( .A1(n361), .A2(n360), .ZN(n474) );
  AOI22_X1 U12 ( .A1(plusA[27]), .A2(n280), .B1(plus2A[27]), .B2(n274), .ZN(
        n361) );
  AOI22_X1 U13 ( .A1(minus2A[27]), .A2(n292), .B1(minusA[27]), .B2(n286), .ZN(
        n360) );
  NAND2_X1 U14 ( .A1(n353), .A2(n352), .ZN(n478) );
  AOI22_X1 U15 ( .A1(plusA[23]), .A2(n279), .B1(plus2A[23]), .B2(n273), .ZN(
        n353) );
  AOI22_X1 U16 ( .A1(minus2A[23]), .A2(n291), .B1(minusA[23]), .B2(n285), .ZN(
        n352) );
  NAND2_X1 U17 ( .A1(n365), .A2(n364), .ZN(n472) );
  AOI22_X1 U18 ( .A1(plusA[29]), .A2(n280), .B1(plus2A[29]), .B2(n274), .ZN(
        n365) );
  AOI22_X1 U19 ( .A1(minus2A[29]), .A2(n292), .B1(minusA[29]), .B2(n286), .ZN(
        n364) );
  NAND2_X1 U20 ( .A1(n357), .A2(n356), .ZN(n476) );
  AOI22_X1 U21 ( .A1(plusA[25]), .A2(n280), .B1(plus2A[25]), .B2(n274), .ZN(
        n357) );
  AOI22_X1 U22 ( .A1(minus2A[25]), .A2(n292), .B1(minusA[25]), .B2(n286), .ZN(
        n356) );
  NAND2_X1 U23 ( .A1(n349), .A2(n348), .ZN(n480) );
  AOI22_X1 U24 ( .A1(plusA[21]), .A2(n279), .B1(plus2A[21]), .B2(n273), .ZN(
        n349) );
  AOI22_X1 U25 ( .A1(minus2A[21]), .A2(n291), .B1(minusA[21]), .B2(n285), .ZN(
        n348) );
  NAND2_X1 U26 ( .A1(n363), .A2(n362), .ZN(n473) );
  AOI22_X1 U27 ( .A1(plusA[28]), .A2(n280), .B1(plus2A[28]), .B2(n274), .ZN(
        n363) );
  AOI22_X1 U28 ( .A1(minus2A[28]), .A2(n292), .B1(minusA[28]), .B2(n286), .ZN(
        n362) );
  NAND2_X1 U29 ( .A1(n367), .A2(n366), .ZN(n471) );
  AOI22_X1 U30 ( .A1(plusA[30]), .A2(n280), .B1(plus2A[30]), .B2(n274), .ZN(
        n367) );
  AOI22_X1 U31 ( .A1(minus2A[30]), .A2(n292), .B1(minusA[30]), .B2(n286), .ZN(
        n366) );
  NAND2_X1 U32 ( .A1(n359), .A2(n358), .ZN(n475) );
  AOI22_X1 U33 ( .A1(plusA[26]), .A2(n280), .B1(plus2A[26]), .B2(n274), .ZN(
        n359) );
  AOI22_X1 U34 ( .A1(minus2A[26]), .A2(n292), .B1(minusA[26]), .B2(n286), .ZN(
        n358) );
  NAND2_X1 U35 ( .A1(n351), .A2(n350), .ZN(n479) );
  AOI22_X1 U36 ( .A1(plusA[22]), .A2(n279), .B1(plus2A[22]), .B2(n273), .ZN(
        n351) );
  AOI22_X1 U37 ( .A1(minus2A[22]), .A2(n291), .B1(minusA[22]), .B2(n285), .ZN(
        n350) );
  NAND2_X1 U38 ( .A1(n403), .A2(n402), .ZN(n453) );
  AOI22_X1 U39 ( .A1(plusA[48]), .A2(n282), .B1(plus2A[48]), .B2(n276), .ZN(
        n403) );
  AOI22_X1 U40 ( .A1(minus2A[48]), .A2(n294), .B1(minusA[48]), .B2(n288), .ZN(
        n402) );
  NAND2_X1 U41 ( .A1(n393), .A2(n392), .ZN(n458) );
  AOI22_X1 U42 ( .A1(plusA[43]), .A2(n281), .B1(plus2A[43]), .B2(n275), .ZN(
        n393) );
  AOI22_X1 U43 ( .A1(minus2A[43]), .A2(n293), .B1(minusA[43]), .B2(n287), .ZN(
        n392) );
  NAND2_X1 U44 ( .A1(n385), .A2(n384), .ZN(n462) );
  AOI22_X1 U45 ( .A1(plusA[39]), .A2(n281), .B1(plus2A[39]), .B2(n275), .ZN(
        n385) );
  AOI22_X1 U46 ( .A1(minus2A[39]), .A2(n293), .B1(minusA[39]), .B2(n287), .ZN(
        n384) );
  NAND2_X1 U47 ( .A1(n377), .A2(n376), .ZN(n466) );
  AOI22_X1 U48 ( .A1(plusA[35]), .A2(n280), .B1(plus2A[35]), .B2(n274), .ZN(
        n377) );
  AOI22_X1 U49 ( .A1(minus2A[35]), .A2(n292), .B1(minusA[35]), .B2(n286), .ZN(
        n376) );
  NAND2_X1 U50 ( .A1(n419), .A2(n418), .ZN(n445) );
  AOI22_X1 U51 ( .A1(plusA[56]), .A2(n282), .B1(plus2A[56]), .B2(n276), .ZN(
        n419) );
  AOI22_X1 U52 ( .A1(minus2A[56]), .A2(n294), .B1(minusA[56]), .B2(n288), .ZN(
        n418) );
  NAND2_X1 U53 ( .A1(n415), .A2(n414), .ZN(n447) );
  AOI22_X1 U54 ( .A1(plusA[54]), .A2(n282), .B1(plus2A[54]), .B2(n276), .ZN(
        n415) );
  AOI22_X1 U55 ( .A1(minus2A[54]), .A2(n294), .B1(minusA[54]), .B2(n288), .ZN(
        n414) );
  NAND2_X1 U56 ( .A1(n417), .A2(n416), .ZN(n446) );
  AOI22_X1 U57 ( .A1(plusA[55]), .A2(n282), .B1(plus2A[55]), .B2(n276), .ZN(
        n417) );
  AOI22_X1 U58 ( .A1(minus2A[55]), .A2(n294), .B1(minusA[55]), .B2(n288), .ZN(
        n416) );
  NAND2_X1 U59 ( .A1(n413), .A2(n412), .ZN(n448) );
  AOI22_X1 U60 ( .A1(plusA[53]), .A2(n282), .B1(plus2A[53]), .B2(n276), .ZN(
        n413) );
  AOI22_X1 U61 ( .A1(minus2A[53]), .A2(n294), .B1(minusA[53]), .B2(n288), .ZN(
        n412) );
  NAND2_X1 U62 ( .A1(n397), .A2(n396), .ZN(n456) );
  AOI22_X1 U63 ( .A1(plusA[45]), .A2(n281), .B1(plus2A[45]), .B2(n275), .ZN(
        n397) );
  AOI22_X1 U64 ( .A1(minus2A[45]), .A2(n293), .B1(minusA[45]), .B2(n287), .ZN(
        n396) );
  NAND2_X1 U65 ( .A1(n389), .A2(n388), .ZN(n460) );
  AOI22_X1 U66 ( .A1(plusA[41]), .A2(n281), .B1(plus2A[41]), .B2(n275), .ZN(
        n389) );
  AOI22_X1 U67 ( .A1(minus2A[41]), .A2(n293), .B1(minusA[41]), .B2(n287), .ZN(
        n388) );
  NAND2_X1 U68 ( .A1(n381), .A2(n380), .ZN(n464) );
  AOI22_X1 U69 ( .A1(plusA[37]), .A2(n281), .B1(plus2A[37]), .B2(n275), .ZN(
        n381) );
  AOI22_X1 U70 ( .A1(minus2A[37]), .A2(n293), .B1(minusA[37]), .B2(n287), .ZN(
        n380) );
  NAND2_X1 U71 ( .A1(n373), .A2(n372), .ZN(n468) );
  AOI22_X1 U72 ( .A1(plusA[33]), .A2(n280), .B1(plus2A[33]), .B2(n274), .ZN(
        n373) );
  AOI22_X1 U73 ( .A1(minus2A[33]), .A2(n292), .B1(minusA[33]), .B2(n286), .ZN(
        n372) );
  NAND2_X1 U74 ( .A1(n409), .A2(n408), .ZN(n450) );
  AOI22_X1 U75 ( .A1(plusA[51]), .A2(n282), .B1(plus2A[51]), .B2(n276), .ZN(
        n409) );
  AOI22_X1 U76 ( .A1(minus2A[51]), .A2(n294), .B1(minusA[51]), .B2(n288), .ZN(
        n408) );
  NAND2_X1 U77 ( .A1(n405), .A2(n404), .ZN(n452) );
  AOI22_X1 U78 ( .A1(plusA[49]), .A2(n282), .B1(plus2A[49]), .B2(n276), .ZN(
        n405) );
  AOI22_X1 U79 ( .A1(minus2A[49]), .A2(n294), .B1(minusA[49]), .B2(n288), .ZN(
        n404) );
  NAND2_X1 U80 ( .A1(n411), .A2(n410), .ZN(n449) );
  AOI22_X1 U81 ( .A1(plusA[52]), .A2(n282), .B1(plus2A[52]), .B2(n276), .ZN(
        n411) );
  AOI22_X1 U82 ( .A1(minus2A[52]), .A2(n294), .B1(minusA[52]), .B2(n288), .ZN(
        n410) );
  NAND2_X1 U83 ( .A1(n407), .A2(n406), .ZN(n451) );
  AOI22_X1 U84 ( .A1(plusA[50]), .A2(n282), .B1(plus2A[50]), .B2(n276), .ZN(
        n407) );
  AOI22_X1 U85 ( .A1(minus2A[50]), .A2(n294), .B1(minusA[50]), .B2(n288), .ZN(
        n406) );
  NAND2_X1 U86 ( .A1(n395), .A2(n394), .ZN(n457) );
  AOI22_X1 U87 ( .A1(plusA[44]), .A2(n281), .B1(plus2A[44]), .B2(n275), .ZN(
        n395) );
  AOI22_X1 U88 ( .A1(minus2A[44]), .A2(n293), .B1(minusA[44]), .B2(n287), .ZN(
        n394) );
  NAND2_X1 U89 ( .A1(n387), .A2(n386), .ZN(n461) );
  AOI22_X1 U90 ( .A1(plusA[40]), .A2(n281), .B1(plus2A[40]), .B2(n275), .ZN(
        n387) );
  AOI22_X1 U91 ( .A1(minus2A[40]), .A2(n293), .B1(minusA[40]), .B2(n287), .ZN(
        n386) );
  NAND2_X1 U92 ( .A1(n379), .A2(n378), .ZN(n465) );
  AOI22_X1 U93 ( .A1(plusA[36]), .A2(n281), .B1(plus2A[36]), .B2(n275), .ZN(
        n379) );
  AOI22_X1 U94 ( .A1(minus2A[36]), .A2(n293), .B1(minusA[36]), .B2(n287), .ZN(
        n378) );
  NAND2_X1 U95 ( .A1(n371), .A2(n370), .ZN(n469) );
  AOI22_X1 U96 ( .A1(plusA[32]), .A2(n280), .B1(plus2A[32]), .B2(n274), .ZN(
        n371) );
  AOI22_X1 U97 ( .A1(minus2A[32]), .A2(n292), .B1(minusA[32]), .B2(n286), .ZN(
        n370) );
  NAND2_X1 U98 ( .A1(n401), .A2(n400), .ZN(n454) );
  AOI22_X1 U99 ( .A1(plusA[47]), .A2(n281), .B1(plus2A[47]), .B2(n275), .ZN(
        n401) );
  AOI22_X1 U100 ( .A1(minus2A[47]), .A2(n293), .B1(minusA[47]), .B2(n287), 
        .ZN(n400) );
  NAND2_X1 U101 ( .A1(n399), .A2(n398), .ZN(n455) );
  AOI22_X1 U102 ( .A1(plusA[46]), .A2(n281), .B1(plus2A[46]), .B2(n275), .ZN(
        n399) );
  AOI22_X1 U103 ( .A1(minus2A[46]), .A2(n293), .B1(minusA[46]), .B2(n287), 
        .ZN(n398) );
  NAND2_X1 U104 ( .A1(n391), .A2(n390), .ZN(n459) );
  AOI22_X1 U105 ( .A1(plusA[42]), .A2(n281), .B1(plus2A[42]), .B2(n275), .ZN(
        n391) );
  AOI22_X1 U106 ( .A1(minus2A[42]), .A2(n293), .B1(minusA[42]), .B2(n287), 
        .ZN(n390) );
  NAND2_X1 U107 ( .A1(n383), .A2(n382), .ZN(n463) );
  AOI22_X1 U108 ( .A1(plusA[38]), .A2(n281), .B1(plus2A[38]), .B2(n275), .ZN(
        n383) );
  AOI22_X1 U109 ( .A1(minus2A[38]), .A2(n293), .B1(minusA[38]), .B2(n287), 
        .ZN(n382) );
  NAND2_X1 U110 ( .A1(n375), .A2(n374), .ZN(n467) );
  AOI22_X1 U111 ( .A1(plusA[34]), .A2(n280), .B1(plus2A[34]), .B2(n274), .ZN(
        n375) );
  AOI22_X1 U112 ( .A1(minus2A[34]), .A2(n292), .B1(minusA[34]), .B2(n286), 
        .ZN(n374) );
  NAND2_X1 U113 ( .A1(n421), .A2(n420), .ZN(n444) );
  AOI22_X1 U114 ( .A1(plusA[57]), .A2(n282), .B1(plus2A[57]), .B2(n276), .ZN(
        n421) );
  AOI22_X1 U115 ( .A1(minus2A[57]), .A2(n294), .B1(minusA[57]), .B2(n288), 
        .ZN(n420) );
  NAND2_X1 U116 ( .A1(n437), .A2(n436), .ZN(n438) );
  AOI22_X1 U117 ( .A1(plusA[63]), .A2(n283), .B1(plus2A[63]), .B2(n277), .ZN(
        n437) );
  AOI22_X1 U118 ( .A1(minus2A[63]), .A2(n295), .B1(minusA[63]), .B2(n289), 
        .ZN(n436) );
  NAND2_X1 U119 ( .A1(n431), .A2(n430), .ZN(n439) );
  AOI22_X1 U120 ( .A1(plusA[62]), .A2(n283), .B1(plus2A[62]), .B2(n277), .ZN(
        n431) );
  AOI22_X1 U121 ( .A1(minus2A[62]), .A2(n295), .B1(minusA[62]), .B2(n289), 
        .ZN(n430) );
  NAND2_X1 U122 ( .A1(n429), .A2(n428), .ZN(n440) );
  AOI22_X1 U123 ( .A1(plusA[61]), .A2(n283), .B1(plus2A[61]), .B2(n277), .ZN(
        n429) );
  AOI22_X1 U124 ( .A1(minus2A[61]), .A2(n295), .B1(minusA[61]), .B2(n289), 
        .ZN(n428) );
  NAND2_X1 U125 ( .A1(n427), .A2(n426), .ZN(n441) );
  AOI22_X1 U126 ( .A1(plusA[60]), .A2(n283), .B1(plus2A[60]), .B2(n277), .ZN(
        n427) );
  AOI22_X1 U127 ( .A1(minus2A[60]), .A2(n295), .B1(minusA[60]), .B2(n289), 
        .ZN(n426) );
  NAND2_X1 U128 ( .A1(n425), .A2(n424), .ZN(n442) );
  AOI22_X1 U129 ( .A1(plusA[59]), .A2(n282), .B1(plus2A[59]), .B2(n276), .ZN(
        n425) );
  AOI22_X1 U130 ( .A1(minus2A[59]), .A2(n294), .B1(minusA[59]), .B2(n288), 
        .ZN(n424) );
  NAND2_X1 U131 ( .A1(n423), .A2(n422), .ZN(n443) );
  AOI22_X1 U132 ( .A1(plusA[58]), .A2(n282), .B1(plus2A[58]), .B2(n276), .ZN(
        n423) );
  AOI22_X1 U133 ( .A1(minus2A[58]), .A2(n294), .B1(minusA[58]), .B2(n288), 
        .ZN(n422) );
  BUF_X1 U134 ( .A(n493), .Z(n296) );
  BUF_X1 U135 ( .A(n433), .Z(n279) );
  BUF_X1 U136 ( .A(n435), .Z(n291) );
  BUF_X1 U137 ( .A(n434), .Z(n285) );
  BUF_X1 U138 ( .A(n432), .Z(n273) );
  BUF_X1 U139 ( .A(n493), .Z(n297) );
  NAND2_X1 U140 ( .A1(n345), .A2(n344), .ZN(n482) );
  AOI22_X1 U141 ( .A1(plusA[19]), .A2(n279), .B1(plus2A[19]), .B2(n273), .ZN(
        n345) );
  AOI22_X1 U142 ( .A1(minus2A[19]), .A2(n291), .B1(minusA[19]), .B2(n285), 
        .ZN(n344) );
  NAND2_X1 U143 ( .A1(n343), .A2(n342), .ZN(n483) );
  AOI22_X1 U144 ( .A1(plusA[18]), .A2(n279), .B1(plus2A[18]), .B2(n273), .ZN(
        n343) );
  AOI22_X1 U145 ( .A1(minus2A[18]), .A2(n291), .B1(minusA[18]), .B2(n285), 
        .ZN(n342) );
  BUF_X1 U146 ( .A(n433), .Z(n280) );
  BUF_X1 U147 ( .A(n435), .Z(n292) );
  BUF_X1 U148 ( .A(n434), .Z(n286) );
  BUF_X1 U149 ( .A(n432), .Z(n274) );
  BUF_X1 U150 ( .A(n493), .Z(n298) );
  BUF_X1 U151 ( .A(n433), .Z(n281) );
  BUF_X1 U152 ( .A(n435), .Z(n293) );
  BUF_X1 U153 ( .A(n434), .Z(n287) );
  BUF_X1 U154 ( .A(n432), .Z(n275) );
  BUF_X1 U155 ( .A(n493), .Z(n299) );
  BUF_X1 U156 ( .A(n433), .Z(n282) );
  BUF_X1 U157 ( .A(n435), .Z(n294) );
  BUF_X1 U158 ( .A(n434), .Z(n288) );
  BUF_X1 U159 ( .A(n432), .Z(n276) );
  BUF_X1 U160 ( .A(n493), .Z(n300) );
  BUF_X1 U161 ( .A(n493), .Z(n301) );
  BUF_X1 U162 ( .A(n433), .Z(n278) );
  BUF_X1 U163 ( .A(n435), .Z(n290) );
  BUF_X1 U164 ( .A(n434), .Z(n284) );
  BUF_X1 U165 ( .A(n432), .Z(n272) );
  NOR2_X1 U166 ( .A1(n323), .A2(n304), .ZN(n493) );
  INV_X1 U167 ( .A(SEL[2]), .ZN(n304) );
  NOR2_X1 U168 ( .A1(SEL[1]), .A2(SEL[0]), .ZN(n323) );
  NOR3_X1 U169 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n302), .ZN(n434) );
  NOR3_X1 U170 ( .A1(SEL[1]), .A2(SEL[2]), .A3(n303), .ZN(n433) );
  NOR3_X1 U171 ( .A1(n302), .A2(SEL[2]), .A3(n303), .ZN(n432) );
  NAND2_X1 U172 ( .A1(n341), .A2(n340), .ZN(n484) );
  AOI22_X1 U173 ( .A1(plusA[17]), .A2(n279), .B1(plus2A[17]), .B2(n273), .ZN(
        n341) );
  AOI22_X1 U174 ( .A1(minus2A[17]), .A2(n291), .B1(minusA[17]), .B2(n285), 
        .ZN(n340) );
  AND2_X1 U175 ( .A1(SEL[2]), .A2(n323), .ZN(n435) );
  INV_X1 U176 ( .A(SEL[1]), .ZN(n302) );
  INV_X1 U177 ( .A(SEL[0]), .ZN(n303) );
  NAND2_X1 U178 ( .A1(n339), .A2(n338), .ZN(n485) );
  AOI22_X1 U179 ( .A1(plusA[16]), .A2(n279), .B1(plus2A[16]), .B2(n273), .ZN(
        n339) );
  AOI22_X1 U180 ( .A1(minus2A[16]), .A2(n291), .B1(minusA[16]), .B2(n285), 
        .ZN(n338) );
  NAND2_X1 U181 ( .A1(n337), .A2(n336), .ZN(n486) );
  AOI22_X1 U182 ( .A1(plusA[15]), .A2(n279), .B1(plus2A[15]), .B2(n273), .ZN(
        n337) );
  AOI22_X1 U183 ( .A1(minus2A[15]), .A2(n291), .B1(minusA[15]), .B2(n285), 
        .ZN(n336) );
  NAND2_X1 U184 ( .A1(n335), .A2(n334), .ZN(n487) );
  AOI22_X1 U185 ( .A1(plusA[14]), .A2(n279), .B1(plus2A[14]), .B2(n273), .ZN(
        n335) );
  AOI22_X1 U186 ( .A1(minus2A[14]), .A2(n291), .B1(minusA[14]), .B2(n285), 
        .ZN(n334) );
  NAND2_X1 U187 ( .A1(n333), .A2(n332), .ZN(n488) );
  AOI22_X1 U188 ( .A1(plusA[13]), .A2(n279), .B1(plus2A[13]), .B2(n273), .ZN(
        n333) );
  AOI22_X1 U189 ( .A1(minus2A[13]), .A2(n291), .B1(minusA[13]), .B2(n285), 
        .ZN(n332) );
  NAND2_X1 U190 ( .A1(n329), .A2(n328), .ZN(n490) );
  AOI22_X1 U191 ( .A1(plusA[11]), .A2(n278), .B1(plus2A[11]), .B2(n272), .ZN(
        n329) );
  AOI22_X1 U192 ( .A1(minus2A[11]), .A2(n290), .B1(minusA[11]), .B2(n284), 
        .ZN(n328) );
  NAND2_X1 U193 ( .A1(n327), .A2(n326), .ZN(n491) );
  AOI22_X1 U194 ( .A1(plusA[10]), .A2(n278), .B1(plus2A[10]), .B2(n272), .ZN(
        n327) );
  AOI22_X1 U195 ( .A1(minus2A[10]), .A2(n290), .B1(minusA[10]), .B2(n284), 
        .ZN(n326) );
  NAND2_X1 U196 ( .A1(n325), .A2(n324), .ZN(n492) );
  AOI22_X1 U197 ( .A1(plusA[9]), .A2(n278), .B1(plus2A[9]), .B2(n272), .ZN(
        n325) );
  AOI22_X1 U198 ( .A1(minus2A[9]), .A2(n290), .B1(minusA[9]), .B2(n284), .ZN(
        n324) );
  NAND2_X1 U199 ( .A1(n320), .A2(n319), .ZN(n495) );
  AOI22_X1 U200 ( .A1(plusA[7]), .A2(n278), .B1(plus2A[7]), .B2(n272), .ZN(
        n320) );
  AOI22_X1 U201 ( .A1(minus2A[7]), .A2(n290), .B1(minusA[7]), .B2(n284), .ZN(
        n319) );
  NAND2_X1 U202 ( .A1(n318), .A2(n317), .ZN(n496) );
  AOI22_X1 U203 ( .A1(plusA[6]), .A2(n278), .B1(plus2A[6]), .B2(n272), .ZN(
        n318) );
  AOI22_X1 U204 ( .A1(minus2A[6]), .A2(n290), .B1(minusA[6]), .B2(n284), .ZN(
        n317) );
  NAND2_X1 U205 ( .A1(n316), .A2(n315), .ZN(n497) );
  AOI22_X1 U206 ( .A1(plusA[5]), .A2(n278), .B1(plus2A[5]), .B2(n272), .ZN(
        n316) );
  AOI22_X1 U207 ( .A1(minus2A[5]), .A2(n290), .B1(minusA[5]), .B2(n284), .ZN(
        n315) );
  NAND2_X1 U208 ( .A1(n312), .A2(n311), .ZN(n499) );
  AOI22_X1 U209 ( .A1(plusA[3]), .A2(n278), .B1(plus2A[3]), .B2(n272), .ZN(
        n312) );
  AOI22_X1 U210 ( .A1(minus2A[3]), .A2(n290), .B1(minusA[3]), .B2(n284), .ZN(
        n311) );
  NAND2_X1 U211 ( .A1(n331), .A2(n330), .ZN(n489) );
  AOI22_X1 U212 ( .A1(plusA[12]), .A2(n279), .B1(plus2A[12]), .B2(n273), .ZN(
        n331) );
  AOI22_X1 U213 ( .A1(minus2A[12]), .A2(n291), .B1(minusA[12]), .B2(n285), 
        .ZN(n330) );
  NAND2_X1 U214 ( .A1(n322), .A2(n321), .ZN(n494) );
  AOI22_X1 U215 ( .A1(plusA[8]), .A2(n278), .B1(plus2A[8]), .B2(n272), .ZN(
        n322) );
  AOI22_X1 U216 ( .A1(minus2A[8]), .A2(n290), .B1(minusA[8]), .B2(n284), .ZN(
        n321) );
  NAND2_X1 U217 ( .A1(n314), .A2(n313), .ZN(n498) );
  AOI22_X1 U218 ( .A1(plusA[4]), .A2(n278), .B1(plus2A[4]), .B2(n272), .ZN(
        n314) );
  AOI22_X1 U219 ( .A1(minus2A[4]), .A2(n290), .B1(minusA[4]), .B2(n284), .ZN(
        n313) );
  NAND2_X1 U220 ( .A1(n310), .A2(n309), .ZN(n500) );
  AOI22_X1 U221 ( .A1(plusA[2]), .A2(n278), .B1(plus2A[2]), .B2(n272), .ZN(
        n310) );
  AOI22_X1 U222 ( .A1(minus2A[2]), .A2(n290), .B1(minusA[2]), .B2(n284), .ZN(
        n309) );
  NAND2_X1 U223 ( .A1(n308), .A2(n307), .ZN(n501) );
  AOI22_X1 U224 ( .A1(plusA[1]), .A2(n278), .B1(plus2A[1]), .B2(n272), .ZN(
        n308) );
  AOI22_X1 U225 ( .A1(minus2A[1]), .A2(n290), .B1(minusA[1]), .B2(n284), .ZN(
        n307) );
  NAND2_X1 U226 ( .A1(n306), .A2(n305), .ZN(n502) );
  AOI22_X1 U227 ( .A1(plusA[0]), .A2(n278), .B1(plus2A[0]), .B2(n272), .ZN(
        n306) );
  AOI22_X1 U228 ( .A1(minus2A[0]), .A2(n290), .B1(minusA[0]), .B2(n284), .ZN(
        n305) );
  CLKBUF_X1 U229 ( .A(n432), .Z(n277) );
  CLKBUF_X1 U230 ( .A(n433), .Z(n283) );
  CLKBUF_X1 U231 ( .A(n434), .Z(n289) );
  CLKBUF_X1 U232 ( .A(n435), .Z(n295) );
endmodule


module FA_512 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_511 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_510 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_509 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_508 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_507 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_506 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_505 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_504 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_503 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_502 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_501 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_500 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_499 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_498 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_497 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_496 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_495 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_494 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_493 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_492 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_491 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_490 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_489 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_488 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_487 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_486 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_485 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_484 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_483 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_482 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_481 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_480 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_479 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_478 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_477 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_476 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_475 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_474 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_473 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_472 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_471 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_470 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_469 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_468 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_467 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_466 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_465 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_464 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_463 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_462 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_461 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_460 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_459 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_458 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_457 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_456 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_455 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_454 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_453 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_452 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_451 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_450 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_449 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N64_8 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Ci;
  output Co;

  wire   [63:1] CTMP;
  tri   [63:0] A;

  FA_512 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_511 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_510 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_509 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(CTMP[4]) );
  FA_508 FAI_5 ( .A(A[4]), .B(B[4]), .Ci(CTMP[4]), .S(S[4]), .Co(CTMP[5]) );
  FA_507 FAI_6 ( .A(A[5]), .B(B[5]), .Ci(CTMP[5]), .S(S[5]), .Co(CTMP[6]) );
  FA_506 FAI_7 ( .A(A[6]), .B(B[6]), .Ci(CTMP[6]), .S(S[6]), .Co(CTMP[7]) );
  FA_505 FAI_8 ( .A(A[7]), .B(B[7]), .Ci(CTMP[7]), .S(S[7]), .Co(CTMP[8]) );
  FA_504 FAI_9 ( .A(A[8]), .B(B[8]), .Ci(CTMP[8]), .S(S[8]), .Co(CTMP[9]) );
  FA_503 FAI_10 ( .A(A[9]), .B(B[9]), .Ci(CTMP[9]), .S(S[9]), .Co(CTMP[10]) );
  FA_502 FAI_11 ( .A(A[10]), .B(B[10]), .Ci(CTMP[10]), .S(S[10]), .Co(CTMP[11]) );
  FA_501 FAI_12 ( .A(A[11]), .B(B[11]), .Ci(CTMP[11]), .S(S[11]), .Co(CTMP[12]) );
  FA_500 FAI_13 ( .A(A[12]), .B(B[12]), .Ci(CTMP[12]), .S(S[12]), .Co(CTMP[13]) );
  FA_499 FAI_14 ( .A(A[13]), .B(B[13]), .Ci(CTMP[13]), .S(S[13]), .Co(CTMP[14]) );
  FA_498 FAI_15 ( .A(A[14]), .B(B[14]), .Ci(CTMP[14]), .S(S[14]), .Co(CTMP[15]) );
  FA_497 FAI_16 ( .A(A[15]), .B(B[15]), .Ci(CTMP[15]), .S(S[15]), .Co(CTMP[16]) );
  FA_496 FAI_17 ( .A(A[16]), .B(B[16]), .Ci(CTMP[16]), .S(S[16]), .Co(CTMP[17]) );
  FA_495 FAI_18 ( .A(A[17]), .B(B[17]), .Ci(CTMP[17]), .S(S[17]), .Co(CTMP[18]) );
  FA_494 FAI_19 ( .A(A[18]), .B(B[18]), .Ci(CTMP[18]), .S(S[18]), .Co(CTMP[19]) );
  FA_493 FAI_20 ( .A(A[19]), .B(B[19]), .Ci(CTMP[19]), .S(S[19]), .Co(CTMP[20]) );
  FA_492 FAI_21 ( .A(A[20]), .B(B[20]), .Ci(CTMP[20]), .S(S[20]), .Co(CTMP[21]) );
  FA_491 FAI_22 ( .A(A[21]), .B(B[21]), .Ci(CTMP[21]), .S(S[21]), .Co(CTMP[22]) );
  FA_490 FAI_23 ( .A(A[22]), .B(B[22]), .Ci(CTMP[22]), .S(S[22]), .Co(CTMP[23]) );
  FA_489 FAI_24 ( .A(A[23]), .B(B[23]), .Ci(CTMP[23]), .S(S[23]), .Co(CTMP[24]) );
  FA_488 FAI_25 ( .A(A[24]), .B(B[24]), .Ci(CTMP[24]), .S(S[24]), .Co(CTMP[25]) );
  FA_487 FAI_26 ( .A(A[25]), .B(B[25]), .Ci(CTMP[25]), .S(S[25]), .Co(CTMP[26]) );
  FA_486 FAI_27 ( .A(A[26]), .B(B[26]), .Ci(CTMP[26]), .S(S[26]), .Co(CTMP[27]) );
  FA_485 FAI_28 ( .A(A[27]), .B(B[27]), .Ci(CTMP[27]), .S(S[27]), .Co(CTMP[28]) );
  FA_484 FAI_29 ( .A(A[28]), .B(B[28]), .Ci(CTMP[28]), .S(S[28]), .Co(CTMP[29]) );
  FA_483 FAI_30 ( .A(A[29]), .B(B[29]), .Ci(CTMP[29]), .S(S[29]), .Co(CTMP[30]) );
  FA_482 FAI_31 ( .A(A[30]), .B(B[30]), .Ci(CTMP[30]), .S(S[30]), .Co(CTMP[31]) );
  FA_481 FAI_32 ( .A(A[31]), .B(B[31]), .Ci(CTMP[31]), .S(S[31]), .Co(CTMP[32]) );
  FA_480 FAI_33 ( .A(A[32]), .B(B[32]), .Ci(CTMP[32]), .S(S[32]), .Co(CTMP[33]) );
  FA_479 FAI_34 ( .A(A[33]), .B(B[33]), .Ci(CTMP[33]), .S(S[33]), .Co(CTMP[34]) );
  FA_478 FAI_35 ( .A(A[34]), .B(B[34]), .Ci(CTMP[34]), .S(S[34]), .Co(CTMP[35]) );
  FA_477 FAI_36 ( .A(A[35]), .B(B[35]), .Ci(CTMP[35]), .S(S[35]), .Co(CTMP[36]) );
  FA_476 FAI_37 ( .A(A[36]), .B(B[36]), .Ci(CTMP[36]), .S(S[36]), .Co(CTMP[37]) );
  FA_475 FAI_38 ( .A(A[37]), .B(B[37]), .Ci(CTMP[37]), .S(S[37]), .Co(CTMP[38]) );
  FA_474 FAI_39 ( .A(A[38]), .B(B[38]), .Ci(CTMP[38]), .S(S[38]), .Co(CTMP[39]) );
  FA_473 FAI_40 ( .A(A[39]), .B(B[39]), .Ci(CTMP[39]), .S(S[39]), .Co(CTMP[40]) );
  FA_472 FAI_41 ( .A(A[40]), .B(B[40]), .Ci(CTMP[40]), .S(S[40]), .Co(CTMP[41]) );
  FA_471 FAI_42 ( .A(A[41]), .B(B[41]), .Ci(CTMP[41]), .S(S[41]), .Co(CTMP[42]) );
  FA_470 FAI_43 ( .A(A[42]), .B(B[42]), .Ci(CTMP[42]), .S(S[42]), .Co(CTMP[43]) );
  FA_469 FAI_44 ( .A(A[43]), .B(B[43]), .Ci(CTMP[43]), .S(S[43]), .Co(CTMP[44]) );
  FA_468 FAI_45 ( .A(A[44]), .B(B[44]), .Ci(CTMP[44]), .S(S[44]), .Co(CTMP[45]) );
  FA_467 FAI_46 ( .A(A[45]), .B(B[45]), .Ci(CTMP[45]), .S(S[45]), .Co(CTMP[46]) );
  FA_466 FAI_47 ( .A(A[46]), .B(B[46]), .Ci(CTMP[46]), .S(S[46]), .Co(CTMP[47]) );
  FA_465 FAI_48 ( .A(A[47]), .B(B[47]), .Ci(CTMP[47]), .S(S[47]), .Co(CTMP[48]) );
  FA_464 FAI_49 ( .A(A[48]), .B(B[48]), .Ci(CTMP[48]), .S(S[48]), .Co(CTMP[49]) );
  FA_463 FAI_50 ( .A(A[49]), .B(B[49]), .Ci(CTMP[49]), .S(S[49]), .Co(CTMP[50]) );
  FA_462 FAI_51 ( .A(A[50]), .B(B[50]), .Ci(CTMP[50]), .S(S[50]), .Co(CTMP[51]) );
  FA_461 FAI_52 ( .A(A[51]), .B(B[51]), .Ci(CTMP[51]), .S(S[51]), .Co(CTMP[52]) );
  FA_460 FAI_53 ( .A(A[52]), .B(B[52]), .Ci(CTMP[52]), .S(S[52]), .Co(CTMP[53]) );
  FA_459 FAI_54 ( .A(A[53]), .B(B[53]), .Ci(CTMP[53]), .S(S[53]), .Co(CTMP[54]) );
  FA_458 FAI_55 ( .A(A[54]), .B(B[54]), .Ci(CTMP[54]), .S(S[54]), .Co(CTMP[55]) );
  FA_457 FAI_56 ( .A(A[55]), .B(B[55]), .Ci(CTMP[55]), .S(S[55]), .Co(CTMP[56]) );
  FA_456 FAI_57 ( .A(A[56]), .B(B[56]), .Ci(CTMP[56]), .S(S[56]), .Co(CTMP[57]) );
  FA_455 FAI_58 ( .A(A[57]), .B(B[57]), .Ci(CTMP[57]), .S(S[57]), .Co(CTMP[58]) );
  FA_454 FAI_59 ( .A(A[58]), .B(B[58]), .Ci(CTMP[58]), .S(S[58]), .Co(CTMP[59]) );
  FA_453 FAI_60 ( .A(A[59]), .B(B[59]), .Ci(CTMP[59]), .S(S[59]), .Co(CTMP[60]) );
  FA_452 FAI_61 ( .A(A[60]), .B(B[60]), .Ci(CTMP[60]), .S(S[60]), .Co(CTMP[61]) );
  FA_451 FAI_62 ( .A(A[61]), .B(B[61]), .Ci(CTMP[61]), .S(S[61]), .Co(CTMP[62]) );
  FA_450 FAI_63 ( .A(A[62]), .B(B[62]), .Ci(CTMP[62]), .S(S[62]), .Co(CTMP[63]) );
  FA_449 FAI_64 ( .A(A[63]), .B(B[63]), .Ci(CTMP[63]), .S(S[63]), .Co(Co) );
endmodule


module booth_mul_row_N64_RADIX3_8 ( prevA, prevSum, encoderIn, nextA, nextSum
 );
  input [63:0] prevA;
  input [63:0] prevSum;
  input [2:0] encoderIn;
  output [63:0] nextA;
  output [63:0] nextSum;
  wire   n3;
  wire   [2:0] encoder_to_mux;
  wire   [63:0] plus2A_s;
  wire   [63:0] minus2A_s;
  wire   [63:0] minus4A_s;
  tri   [63:0] mux_to_adder;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign nextA[51] = n3;
  assign nextA[0] = 1'b0;

  encoder_N64_RADIX3_8 encoder_1 ( .X(encoderIn), .Z(encoder_to_mux) );
  ShiftnCompl_N64_8 ShiftnCompl_1 ( .plusA(prevA), .plus2A_out({plus2A_s[63:1], 
        SYNOPSYS_UNCONNECTED__0}), .minus2A_out(minus2A_s), .plus4A_out({
        nextA[63:52], n3, nextA[50:1], SYNOPSYS_UNCONNECTED__1}), 
        .minus4A_out(minus4A_s) );
  MUX_GENERIC_N64_RADIX3_8 mux_1 ( .plusA({plus2A_s[63:1], 1'b0}), .minusA(
        minus2A_s), .plus2A({nextA[63:52], n3, nextA[50:1], 1'b0}), .minus2A(
        minus4A_s), .SEL(encoder_to_mux), .Y(mux_to_adder) );
  RCA_N64_8 rca_1 ( .A(mux_to_adder), .B(prevSum), .Ci(1'b0), .S(nextSum) );
endmodule


module encoder_N64_RADIX3_7 ( X, Z );
  input [2:0] X;
  output [2:0] Z;
  wire   n5, n7, n8;

  OAI22_X1 U1 ( .A1(n8), .A2(n5), .B1(X[2]), .B2(n7), .ZN(Z[1]) );
  INV_X1 U2 ( .A(X[2]), .ZN(n5) );
  AOI21_X1 U3 ( .B1(n8), .B2(n7), .A(X[2]), .ZN(Z[0]) );
  OAI21_X1 U4 ( .B1(X[1]), .B2(X[0]), .A(n7), .ZN(n8) );
  AND3_X1 U5 ( .A1(X[2]), .A2(n7), .A3(n8), .ZN(Z[2]) );
  NAND2_X1 U6 ( .A1(X[1]), .A2(X[0]), .ZN(n7) );
endmodule


module shifter_N64_14 ( \input , shiftLeftOnePos );
  input [63:0] \input ;
  output [63:0] shiftLeftOnePos;
  wire   \input[62] , \input[61] , \input[60] , \input[59] , \input[58] ,
         \input[57] , \input[56] , \input[55] , \input[54] , \input[53] ,
         \input[52] , \input[51] , \input[50] , \input[49] , \input[48] ,
         \input[47] , \input[46] , \input[45] , \input[44] , \input[43] ,
         \input[42] , \input[41] , \input[40] , \input[39] , \input[38] ,
         \input[37] , \input[36] , \input[35] , \input[34] , \input[33] ,
         \input[32] , \input[31] , \input[30] , \input[29] , \input[28] ,
         \input[27] , \input[26] , \input[25] , \input[24] , \input[23] ,
         \input[22] , \input[21] , \input[20] , \input[19] , \input[18] ,
         \input[17] , \input[16] , \input[15] , \input[14] , \input[13] ,
         \input[12] , \input[11] , \input[10] , \input[9] , \input[8] ,
         \input[7] , \input[6] , \input[5] , \input[4] , \input[3] ,
         \input[2] , \input[1] , \input[0] ;
  assign shiftLeftOnePos[0] = 1'b0;
  assign shiftLeftOnePos[63] = \input[62] ;
  assign \input[62]  = \input  [62];
  assign shiftLeftOnePos[62] = \input[61] ;
  assign \input[61]  = \input  [61];
  assign shiftLeftOnePos[61] = \input[60] ;
  assign \input[60]  = \input  [60];
  assign shiftLeftOnePos[60] = \input[59] ;
  assign \input[59]  = \input  [59];
  assign shiftLeftOnePos[59] = \input[58] ;
  assign \input[58]  = \input  [58];
  assign shiftLeftOnePos[58] = \input[57] ;
  assign \input[57]  = \input  [57];
  assign shiftLeftOnePos[57] = \input[56] ;
  assign \input[56]  = \input  [56];
  assign shiftLeftOnePos[56] = \input[55] ;
  assign \input[55]  = \input  [55];
  assign shiftLeftOnePos[55] = \input[54] ;
  assign \input[54]  = \input  [54];
  assign shiftLeftOnePos[54] = \input[53] ;
  assign \input[53]  = \input  [53];
  assign shiftLeftOnePos[53] = \input[52] ;
  assign \input[52]  = \input  [52];
  assign shiftLeftOnePos[52] = \input[51] ;
  assign \input[51]  = \input  [51];
  assign shiftLeftOnePos[51] = \input[50] ;
  assign \input[50]  = \input  [50];
  assign shiftLeftOnePos[50] = \input[49] ;
  assign \input[49]  = \input  [49];
  assign shiftLeftOnePos[49] = \input[48] ;
  assign \input[48]  = \input  [48];
  assign shiftLeftOnePos[48] = \input[47] ;
  assign \input[47]  = \input  [47];
  assign shiftLeftOnePos[47] = \input[46] ;
  assign \input[46]  = \input  [46];
  assign shiftLeftOnePos[46] = \input[45] ;
  assign \input[45]  = \input  [45];
  assign shiftLeftOnePos[45] = \input[44] ;
  assign \input[44]  = \input  [44];
  assign shiftLeftOnePos[44] = \input[43] ;
  assign \input[43]  = \input  [43];
  assign shiftLeftOnePos[43] = \input[42] ;
  assign \input[42]  = \input  [42];
  assign shiftLeftOnePos[42] = \input[41] ;
  assign \input[41]  = \input  [41];
  assign shiftLeftOnePos[41] = \input[40] ;
  assign \input[40]  = \input  [40];
  assign shiftLeftOnePos[40] = \input[39] ;
  assign \input[39]  = \input  [39];
  assign shiftLeftOnePos[39] = \input[38] ;
  assign \input[38]  = \input  [38];
  assign shiftLeftOnePos[38] = \input[37] ;
  assign \input[37]  = \input  [37];
  assign shiftLeftOnePos[37] = \input[36] ;
  assign \input[36]  = \input  [36];
  assign shiftLeftOnePos[36] = \input[35] ;
  assign \input[35]  = \input  [35];
  assign shiftLeftOnePos[35] = \input[34] ;
  assign \input[34]  = \input  [34];
  assign shiftLeftOnePos[34] = \input[33] ;
  assign \input[33]  = \input  [33];
  assign shiftLeftOnePos[33] = \input[32] ;
  assign \input[32]  = \input  [32];
  assign shiftLeftOnePos[32] = \input[31] ;
  assign \input[31]  = \input  [31];
  assign shiftLeftOnePos[31] = \input[30] ;
  assign \input[30]  = \input  [30];
  assign shiftLeftOnePos[30] = \input[29] ;
  assign \input[29]  = \input  [29];
  assign shiftLeftOnePos[29] = \input[28] ;
  assign \input[28]  = \input  [28];
  assign shiftLeftOnePos[28] = \input[27] ;
  assign \input[27]  = \input  [27];
  assign shiftLeftOnePos[27] = \input[26] ;
  assign \input[26]  = \input  [26];
  assign shiftLeftOnePos[26] = \input[25] ;
  assign \input[25]  = \input  [25];
  assign shiftLeftOnePos[25] = \input[24] ;
  assign \input[24]  = \input  [24];
  assign shiftLeftOnePos[24] = \input[23] ;
  assign \input[23]  = \input  [23];
  assign shiftLeftOnePos[23] = \input[22] ;
  assign \input[22]  = \input  [22];
  assign shiftLeftOnePos[22] = \input[21] ;
  assign \input[21]  = \input  [21];
  assign shiftLeftOnePos[21] = \input[20] ;
  assign \input[20]  = \input  [20];
  assign shiftLeftOnePos[20] = \input[19] ;
  assign \input[19]  = \input  [19];
  assign shiftLeftOnePos[19] = \input[18] ;
  assign \input[18]  = \input  [18];
  assign shiftLeftOnePos[18] = \input[17] ;
  assign \input[17]  = \input  [17];
  assign shiftLeftOnePos[17] = \input[16] ;
  assign \input[16]  = \input  [16];
  assign shiftLeftOnePos[16] = \input[15] ;
  assign \input[15]  = \input  [15];
  assign shiftLeftOnePos[15] = \input[14] ;
  assign \input[14]  = \input  [14];
  assign shiftLeftOnePos[14] = \input[13] ;
  assign \input[13]  = \input  [13];
  assign shiftLeftOnePos[13] = \input[12] ;
  assign \input[12]  = \input  [12];
  assign shiftLeftOnePos[12] = \input[11] ;
  assign \input[11]  = \input  [11];
  assign shiftLeftOnePos[11] = \input[10] ;
  assign \input[10]  = \input  [10];
  assign shiftLeftOnePos[10] = \input[9] ;
  assign \input[9]  = \input  [9];
  assign shiftLeftOnePos[9] = \input[8] ;
  assign \input[8]  = \input  [8];
  assign shiftLeftOnePos[8] = \input[7] ;
  assign \input[7]  = \input  [7];
  assign shiftLeftOnePos[7] = \input[6] ;
  assign \input[6]  = \input  [6];
  assign shiftLeftOnePos[6] = \input[5] ;
  assign \input[5]  = \input  [5];
  assign shiftLeftOnePos[5] = \input[4] ;
  assign \input[4]  = \input  [4];
  assign shiftLeftOnePos[4] = \input[3] ;
  assign \input[3]  = \input  [3];
  assign shiftLeftOnePos[3] = \input[2] ;
  assign \input[2]  = \input  [2];
  assign shiftLeftOnePos[2] = \input[1] ;
  assign \input[1]  = \input  [1];
  assign shiftLeftOnePos[1] = \input[0] ;
  assign \input[0]  = \input  [0];

endmodule


module shifter_N64_13 ( \input , shiftLeftOnePos );
  input [63:0] \input ;
  output [63:0] shiftLeftOnePos;
  wire   \input[62] , \input[61] , \input[60] , \input[59] , \input[58] ,
         \input[57] , \input[56] , \input[55] , \input[54] , \input[53] ,
         \input[52] , \input[51] , \input[50] , \input[49] , \input[48] ,
         \input[47] , \input[46] , \input[45] , \input[44] , \input[43] ,
         \input[42] , \input[41] , \input[40] , \input[39] , \input[38] ,
         \input[37] , \input[36] , \input[35] , \input[34] , \input[33] ,
         \input[32] , \input[31] , \input[30] , \input[29] , \input[28] ,
         \input[27] , \input[26] , \input[25] , \input[24] , \input[23] ,
         \input[22] , \input[21] , \input[20] , \input[19] , \input[18] ,
         \input[17] , \input[16] , \input[15] , \input[14] , \input[13] ,
         \input[12] , \input[11] , \input[10] , \input[9] , \input[8] ,
         \input[7] , \input[6] , \input[5] , \input[4] , \input[3] ,
         \input[2] , \input[1] , \input[0] ;
  assign shiftLeftOnePos[0] = 1'b0;
  assign shiftLeftOnePos[63] = \input[62] ;
  assign \input[62]  = \input  [62];
  assign shiftLeftOnePos[62] = \input[61] ;
  assign \input[61]  = \input  [61];
  assign shiftLeftOnePos[61] = \input[60] ;
  assign \input[60]  = \input  [60];
  assign shiftLeftOnePos[60] = \input[59] ;
  assign \input[59]  = \input  [59];
  assign shiftLeftOnePos[59] = \input[58] ;
  assign \input[58]  = \input  [58];
  assign shiftLeftOnePos[58] = \input[57] ;
  assign \input[57]  = \input  [57];
  assign shiftLeftOnePos[57] = \input[56] ;
  assign \input[56]  = \input  [56];
  assign shiftLeftOnePos[56] = \input[55] ;
  assign \input[55]  = \input  [55];
  assign shiftLeftOnePos[55] = \input[54] ;
  assign \input[54]  = \input  [54];
  assign shiftLeftOnePos[54] = \input[53] ;
  assign \input[53]  = \input  [53];
  assign shiftLeftOnePos[53] = \input[52] ;
  assign \input[52]  = \input  [52];
  assign shiftLeftOnePos[52] = \input[51] ;
  assign \input[51]  = \input  [51];
  assign shiftLeftOnePos[51] = \input[50] ;
  assign \input[50]  = \input  [50];
  assign shiftLeftOnePos[50] = \input[49] ;
  assign \input[49]  = \input  [49];
  assign shiftLeftOnePos[49] = \input[48] ;
  assign \input[48]  = \input  [48];
  assign shiftLeftOnePos[48] = \input[47] ;
  assign \input[47]  = \input  [47];
  assign shiftLeftOnePos[47] = \input[46] ;
  assign \input[46]  = \input  [46];
  assign shiftLeftOnePos[46] = \input[45] ;
  assign \input[45]  = \input  [45];
  assign shiftLeftOnePos[45] = \input[44] ;
  assign \input[44]  = \input  [44];
  assign shiftLeftOnePos[44] = \input[43] ;
  assign \input[43]  = \input  [43];
  assign shiftLeftOnePos[43] = \input[42] ;
  assign \input[42]  = \input  [42];
  assign shiftLeftOnePos[42] = \input[41] ;
  assign \input[41]  = \input  [41];
  assign shiftLeftOnePos[41] = \input[40] ;
  assign \input[40]  = \input  [40];
  assign shiftLeftOnePos[40] = \input[39] ;
  assign \input[39]  = \input  [39];
  assign shiftLeftOnePos[39] = \input[38] ;
  assign \input[38]  = \input  [38];
  assign shiftLeftOnePos[38] = \input[37] ;
  assign \input[37]  = \input  [37];
  assign shiftLeftOnePos[37] = \input[36] ;
  assign \input[36]  = \input  [36];
  assign shiftLeftOnePos[36] = \input[35] ;
  assign \input[35]  = \input  [35];
  assign shiftLeftOnePos[35] = \input[34] ;
  assign \input[34]  = \input  [34];
  assign shiftLeftOnePos[34] = \input[33] ;
  assign \input[33]  = \input  [33];
  assign shiftLeftOnePos[33] = \input[32] ;
  assign \input[32]  = \input  [32];
  assign shiftLeftOnePos[32] = \input[31] ;
  assign \input[31]  = \input  [31];
  assign shiftLeftOnePos[31] = \input[30] ;
  assign \input[30]  = \input  [30];
  assign shiftLeftOnePos[30] = \input[29] ;
  assign \input[29]  = \input  [29];
  assign shiftLeftOnePos[29] = \input[28] ;
  assign \input[28]  = \input  [28];
  assign shiftLeftOnePos[28] = \input[27] ;
  assign \input[27]  = \input  [27];
  assign shiftLeftOnePos[27] = \input[26] ;
  assign \input[26]  = \input  [26];
  assign shiftLeftOnePos[26] = \input[25] ;
  assign \input[25]  = \input  [25];
  assign shiftLeftOnePos[25] = \input[24] ;
  assign \input[24]  = \input  [24];
  assign shiftLeftOnePos[24] = \input[23] ;
  assign \input[23]  = \input  [23];
  assign shiftLeftOnePos[23] = \input[22] ;
  assign \input[22]  = \input  [22];
  assign shiftLeftOnePos[22] = \input[21] ;
  assign \input[21]  = \input  [21];
  assign shiftLeftOnePos[21] = \input[20] ;
  assign \input[20]  = \input  [20];
  assign shiftLeftOnePos[20] = \input[19] ;
  assign \input[19]  = \input  [19];
  assign shiftLeftOnePos[19] = \input[18] ;
  assign \input[18]  = \input  [18];
  assign shiftLeftOnePos[18] = \input[17] ;
  assign \input[17]  = \input  [17];
  assign shiftLeftOnePos[17] = \input[16] ;
  assign \input[16]  = \input  [16];
  assign shiftLeftOnePos[16] = \input[15] ;
  assign \input[15]  = \input  [15];
  assign shiftLeftOnePos[15] = \input[14] ;
  assign \input[14]  = \input  [14];
  assign shiftLeftOnePos[14] = \input[13] ;
  assign \input[13]  = \input  [13];
  assign shiftLeftOnePos[13] = \input[12] ;
  assign \input[12]  = \input  [12];
  assign shiftLeftOnePos[12] = \input[11] ;
  assign \input[11]  = \input  [11];
  assign shiftLeftOnePos[11] = \input[10] ;
  assign \input[10]  = \input  [10];
  assign shiftLeftOnePos[10] = \input[9] ;
  assign \input[9]  = \input  [9];
  assign shiftLeftOnePos[9] = \input[8] ;
  assign \input[8]  = \input  [8];
  assign shiftLeftOnePos[8] = \input[7] ;
  assign \input[7]  = \input  [7];
  assign shiftLeftOnePos[7] = \input[6] ;
  assign \input[6]  = \input  [6];
  assign shiftLeftOnePos[6] = \input[5] ;
  assign \input[5]  = \input  [5];
  assign shiftLeftOnePos[5] = \input[4] ;
  assign \input[4]  = \input  [4];
  assign shiftLeftOnePos[4] = \input[3] ;
  assign \input[3]  = \input  [3];
  assign shiftLeftOnePos[3] = \input[2] ;
  assign \input[2]  = \input  [2];
  assign shiftLeftOnePos[2] = \input[1] ;
  assign \input[1]  = \input  [1];
  assign shiftLeftOnePos[1] = \input[0] ;
  assign \input[0]  = \input  [0];

endmodule


module complementer_N64_14_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n190, n191, n192, n193, n194, n196, n197, n198, n199, n200,
         n202, n203, n204, n206, n207, n208, n210, n211, n212, n213, n214,
         n216, n217, n218, n220, n221, n222, n224, n225, n226, n228, n229,
         n230, n232, n233, n234, n235, n237, n238, n239, n241, n242, n243,
         n245, n246, n247, n248, n249, n250, n251, n189, n195, n201, n205,
         n209, n215, n219, n223, n227, n231, n236, n240, n244;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U81 ( .A(n190), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U82 ( .A(n192), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U83 ( .A(n193), .B(B[6]), .Z(DIFF[6]) );
  XOR2_X1 U85 ( .A(n196), .B(B[62]), .Z(DIFF[62]) );
  XOR2_X1 U86 ( .A(n194), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U87 ( .A(n198), .B(B[59]), .Z(DIFF[59]) );
  XOR2_X1 U89 ( .A(n200), .B(B[57]), .Z(DIFF[57]) );
  XOR2_X1 U90 ( .A(n202), .B(B[55]), .Z(DIFF[55]) );
  XOR2_X1 U92 ( .A(n204), .B(B[53]), .Z(DIFF[53]) );
  XOR2_X1 U93 ( .A(n206), .B(B[51]), .Z(DIFF[51]) );
  XOR2_X1 U95 ( .A(n208), .B(B[49]), .Z(DIFF[49]) );
  XOR2_X1 U96 ( .A(n212), .B(B[47]), .Z(DIFF[47]) );
  XOR2_X1 U98 ( .A(n214), .B(B[45]), .Z(DIFF[45]) );
  XOR2_X1 U99 ( .A(n216), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U101 ( .A(n218), .B(B[41]), .Z(DIFF[41]) );
  XOR2_X1 U102 ( .A(n211), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U103 ( .A(n220), .B(B[39]), .Z(DIFF[39]) );
  XOR2_X1 U105 ( .A(n222), .B(B[37]), .Z(DIFF[37]) );
  XOR2_X1 U106 ( .A(n224), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U108 ( .A(n226), .B(B[33]), .Z(DIFF[33]) );
  XOR2_X1 U109 ( .A(n228), .B(B[31]), .Z(DIFF[31]) );
  XOR2_X1 U111 ( .A(n230), .B(B[29]), .Z(DIFF[29]) );
  XOR2_X1 U112 ( .A(n233), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U114 ( .A(n235), .B(B[25]), .Z(DIFF[25]) );
  XOR2_X1 U115 ( .A(n237), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U117 ( .A(n239), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U118 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U119 ( .A(n241), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U121 ( .A(n243), .B(B[17]), .Z(DIFF[17]) );
  XOR2_X1 U122 ( .A(n245), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U123 ( .A(n248), .B(B[14]), .Z(DIFF[14]) );
  XOR2_X1 U124 ( .A(n247), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U125 ( .A(n249), .B(B[11]), .Z(DIFF[11]) );
  XOR2_X1 U126 ( .A(n251), .B(B[10]), .Z(DIFF[10]) );
  XOR2_X1 U1 ( .A(n197), .B(n244), .Z(DIFF[61]) );
  NAND2_X1 U2 ( .A1(n197), .A2(n244), .ZN(n196) );
  NOR3_X1 U3 ( .A1(B[59]), .A2(B[60]), .A3(n198), .ZN(n197) );
  XNOR2_X1 U4 ( .A(n189), .B(B[54]), .ZN(DIFF[54]) );
  NOR2_X1 U5 ( .A1(n204), .A2(B[53]), .ZN(n189) );
  XNOR2_X1 U6 ( .A(B[56]), .B(n203), .ZN(DIFF[56]) );
  NOR2_X1 U7 ( .A1(B[55]), .A2(n202), .ZN(n203) );
  XNOR2_X1 U8 ( .A(B[60]), .B(n199), .ZN(DIFF[60]) );
  NOR2_X1 U9 ( .A1(B[59]), .A2(n198), .ZN(n199) );
  OR3_X1 U10 ( .A1(B[53]), .A2(B[54]), .A3(n204), .ZN(n202) );
  OR3_X1 U11 ( .A1(B[55]), .A2(B[56]), .A3(n202), .ZN(n200) );
  XNOR2_X1 U12 ( .A(B[52]), .B(n207), .ZN(DIFF[52]) );
  NOR2_X1 U13 ( .A1(B[51]), .A2(n206), .ZN(n207) );
  OR3_X1 U14 ( .A1(B[49]), .A2(B[50]), .A3(n208), .ZN(n206) );
  XNOR2_X1 U15 ( .A(n195), .B(B[50]), .ZN(DIFF[50]) );
  NOR2_X1 U16 ( .A1(n208), .A2(B[49]), .ZN(n195) );
  XNOR2_X1 U17 ( .A(n201), .B(B[63]), .ZN(DIFF[63]) );
  NOR2_X1 U18 ( .A1(n196), .A2(B[62]), .ZN(n201) );
  OR3_X1 U19 ( .A1(B[57]), .A2(B[58]), .A3(n200), .ZN(n198) );
  OR3_X1 U20 ( .A1(B[51]), .A2(B[52]), .A3(n206), .ZN(n204) );
  XNOR2_X1 U21 ( .A(n205), .B(B[58]), .ZN(DIFF[58]) );
  NOR2_X1 U22 ( .A1(n200), .A2(B[57]), .ZN(n205) );
  OR3_X1 U23 ( .A1(B[25]), .A2(B[26]), .A3(n235), .ZN(n233) );
  XNOR2_X1 U24 ( .A(n209), .B(B[26]), .ZN(DIFF[26]) );
  NOR2_X1 U25 ( .A1(n235), .A2(B[25]), .ZN(n209) );
  XNOR2_X1 U26 ( .A(B[44]), .B(n217), .ZN(DIFF[44]) );
  NOR2_X1 U27 ( .A1(B[43]), .A2(n216), .ZN(n217) );
  XNOR2_X1 U28 ( .A(B[40]), .B(n221), .ZN(DIFF[40]) );
  NOR2_X1 U29 ( .A1(B[39]), .A2(n220), .ZN(n221) );
  XNOR2_X1 U30 ( .A(B[36]), .B(n225), .ZN(DIFF[36]) );
  NOR2_X1 U31 ( .A1(B[35]), .A2(n224), .ZN(n225) );
  XNOR2_X1 U32 ( .A(B[32]), .B(n229), .ZN(DIFF[32]) );
  NOR2_X1 U33 ( .A1(B[31]), .A2(n228), .ZN(n229) );
  XNOR2_X1 U34 ( .A(B[28]), .B(n234), .ZN(DIFF[28]) );
  NOR2_X1 U35 ( .A1(B[27]), .A2(n233), .ZN(n234) );
  XNOR2_X1 U36 ( .A(B[48]), .B(n213), .ZN(DIFF[48]) );
  NOR2_X1 U37 ( .A1(B[47]), .A2(n212), .ZN(n213) );
  OR3_X1 U38 ( .A1(B[29]), .A2(B[30]), .A3(n230), .ZN(n228) );
  OR3_X1 U39 ( .A1(B[33]), .A2(B[34]), .A3(n226), .ZN(n224) );
  OR3_X1 U40 ( .A1(B[37]), .A2(B[38]), .A3(n222), .ZN(n220) );
  OR3_X1 U41 ( .A1(B[41]), .A2(B[42]), .A3(n218), .ZN(n216) );
  OR3_X1 U42 ( .A1(B[45]), .A2(B[46]), .A3(n214), .ZN(n212) );
  OR3_X1 U43 ( .A1(B[27]), .A2(B[28]), .A3(n233), .ZN(n230) );
  OR3_X1 U44 ( .A1(B[31]), .A2(B[32]), .A3(n228), .ZN(n226) );
  OR3_X1 U45 ( .A1(B[35]), .A2(B[36]), .A3(n224), .ZN(n222) );
  OR3_X1 U46 ( .A1(B[39]), .A2(B[40]), .A3(n220), .ZN(n218) );
  OR3_X1 U47 ( .A1(B[43]), .A2(B[44]), .A3(n216), .ZN(n214) );
  OR3_X1 U48 ( .A1(B[47]), .A2(B[48]), .A3(n212), .ZN(n208) );
  XNOR2_X1 U49 ( .A(n215), .B(B[46]), .ZN(DIFF[46]) );
  NOR2_X1 U50 ( .A1(n214), .A2(B[45]), .ZN(n215) );
  XNOR2_X1 U51 ( .A(n219), .B(B[42]), .ZN(DIFF[42]) );
  NOR2_X1 U52 ( .A1(n218), .A2(B[41]), .ZN(n219) );
  XNOR2_X1 U53 ( .A(n223), .B(B[38]), .ZN(DIFF[38]) );
  NOR2_X1 U54 ( .A1(n222), .A2(B[37]), .ZN(n223) );
  XNOR2_X1 U55 ( .A(n227), .B(B[34]), .ZN(DIFF[34]) );
  NOR2_X1 U56 ( .A1(n226), .A2(B[33]), .ZN(n227) );
  XNOR2_X1 U57 ( .A(n231), .B(B[30]), .ZN(DIFF[30]) );
  NOR2_X1 U58 ( .A1(n230), .A2(B[29]), .ZN(n231) );
  XNOR2_X1 U59 ( .A(B[24]), .B(n238), .ZN(DIFF[24]) );
  NOR2_X1 U60 ( .A1(B[23]), .A2(n237), .ZN(n238) );
  OR3_X1 U61 ( .A1(B[23]), .A2(B[24]), .A3(n237), .ZN(n235) );
  XNOR2_X1 U62 ( .A(n236), .B(B[22]), .ZN(DIFF[22]) );
  NOR2_X1 U63 ( .A1(n239), .A2(B[21]), .ZN(n236) );
  OR3_X1 U64 ( .A1(B[21]), .A2(B[22]), .A3(n239), .ZN(n237) );
  XNOR2_X1 U65 ( .A(B[20]), .B(n242), .ZN(DIFF[20]) );
  NOR2_X1 U66 ( .A1(B[19]), .A2(n241), .ZN(n242) );
  OR3_X1 U67 ( .A1(B[19]), .A2(B[20]), .A3(n241), .ZN(n239) );
  XNOR2_X1 U68 ( .A(n240), .B(B[18]), .ZN(DIFF[18]) );
  NOR2_X1 U69 ( .A1(n243), .A2(B[17]), .ZN(n240) );
  OR3_X1 U70 ( .A1(B[17]), .A2(B[18]), .A3(n243), .ZN(n241) );
  NOR2_X1 U71 ( .A1(B[15]), .A2(n245), .ZN(n246) );
  NOR2_X1 U72 ( .A1(B[11]), .A2(n249), .ZN(n250) );
  NOR2_X1 U73 ( .A1(B[7]), .A2(n192), .ZN(n191) );
  NOR2_X1 U74 ( .A1(B[3]), .A2(n211), .ZN(n210) );
  OR3_X1 U75 ( .A1(B[13]), .A2(B[14]), .A3(n247), .ZN(n245) );
  OR3_X1 U76 ( .A1(B[10]), .A2(B[9]), .A3(n190), .ZN(n249) );
  OR3_X1 U77 ( .A1(B[5]), .A2(B[6]), .A3(n194), .ZN(n192) );
  OR3_X1 U78 ( .A1(B[15]), .A2(B[16]), .A3(n245), .ZN(n243) );
  OR3_X1 U79 ( .A1(B[11]), .A2(B[12]), .A3(n249), .ZN(n247) );
  OR3_X1 U80 ( .A1(B[7]), .A2(B[8]), .A3(n192), .ZN(n190) );
  OR3_X1 U84 ( .A1(B[3]), .A2(B[4]), .A3(n211), .ZN(n194) );
  XNOR2_X1 U88 ( .A(B[16]), .B(n246), .ZN(DIFF[16]) );
  XNOR2_X1 U91 ( .A(B[12]), .B(n250), .ZN(DIFF[12]) );
  XNOR2_X1 U94 ( .A(B[8]), .B(n191), .ZN(DIFF[8]) );
  XNOR2_X1 U97 ( .A(B[4]), .B(n210), .ZN(DIFF[4]) );
  XNOR2_X1 U100 ( .A(B[2]), .B(n232), .ZN(DIFF[2]) );
  OR2_X1 U104 ( .A1(n247), .A2(B[13]), .ZN(n248) );
  OR2_X1 U107 ( .A1(n190), .A2(B[9]), .ZN(n251) );
  OR2_X1 U110 ( .A1(n194), .A2(B[5]), .ZN(n193) );
  OR3_X1 U113 ( .A1(B[1]), .A2(B[2]), .A3(\B[0] ), .ZN(n211) );
  NOR2_X1 U116 ( .A1(\B[0] ), .A2(B[1]), .ZN(n232) );
  INV_X1 U120 ( .A(B[61]), .ZN(n244) );
endmodule


module complementer_N64_14 ( \input , complement2 );
  input [63:0] \input ;
  output [63:0] complement2;


  complementer_N64_14_DW01_sub_0 sub_add_31_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(\input ), .CI(1'b0), .DIFF(complement2) );
endmodule


module complementer_N64_13_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n190, n191, n192, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n249, n250, n189, n193, n248, n251;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U81 ( .A(n190), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U82 ( .A(n192), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U84 ( .A(n195), .B(B[63]), .Z(DIFF[63]) );
  XOR2_X1 U85 ( .A(n196), .B(B[62]), .Z(DIFF[62]) );
  XOR2_X1 U86 ( .A(n194), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U87 ( .A(n198), .B(B[59]), .Z(DIFF[59]) );
  XOR2_X1 U88 ( .A(n201), .B(B[58]), .Z(DIFF[58]) );
  XOR2_X1 U89 ( .A(n200), .B(B[57]), .Z(DIFF[57]) );
  XOR2_X1 U90 ( .A(n202), .B(B[55]), .Z(DIFF[55]) );
  XOR2_X1 U91 ( .A(n205), .B(B[54]), .Z(DIFF[54]) );
  XOR2_X1 U92 ( .A(n204), .B(B[53]), .Z(DIFF[53]) );
  XOR2_X1 U93 ( .A(n206), .B(B[51]), .Z(DIFF[51]) );
  XOR2_X1 U94 ( .A(n209), .B(B[50]), .Z(DIFF[50]) );
  XOR2_X1 U95 ( .A(n208), .B(B[49]), .Z(DIFF[49]) );
  XOR2_X1 U96 ( .A(n212), .B(B[47]), .Z(DIFF[47]) );
  XOR2_X1 U97 ( .A(n215), .B(B[46]), .Z(DIFF[46]) );
  XOR2_X1 U98 ( .A(n214), .B(B[45]), .Z(DIFF[45]) );
  XOR2_X1 U99 ( .A(n216), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U100 ( .A(n219), .B(B[42]), .Z(DIFF[42]) );
  XOR2_X1 U101 ( .A(n218), .B(B[41]), .Z(DIFF[41]) );
  XOR2_X1 U102 ( .A(n211), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U103 ( .A(n220), .B(B[39]), .Z(DIFF[39]) );
  XOR2_X1 U104 ( .A(n223), .B(B[38]), .Z(DIFF[38]) );
  XOR2_X1 U105 ( .A(n222), .B(B[37]), .Z(DIFF[37]) );
  XOR2_X1 U106 ( .A(n224), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U107 ( .A(n227), .B(B[34]), .Z(DIFF[34]) );
  XOR2_X1 U108 ( .A(n226), .B(B[33]), .Z(DIFF[33]) );
  XOR2_X1 U109 ( .A(n228), .B(B[31]), .Z(DIFF[31]) );
  XOR2_X1 U110 ( .A(n231), .B(B[30]), .Z(DIFF[30]) );
  XOR2_X1 U111 ( .A(n230), .B(B[29]), .Z(DIFF[29]) );
  XOR2_X1 U112 ( .A(n233), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U113 ( .A(n236), .B(B[26]), .Z(DIFF[26]) );
  XOR2_X1 U114 ( .A(n235), .B(B[25]), .Z(DIFF[25]) );
  XOR2_X1 U115 ( .A(n237), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U116 ( .A(n240), .B(B[22]), .Z(DIFF[22]) );
  XOR2_X1 U117 ( .A(n239), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U118 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U119 ( .A(n241), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U120 ( .A(n244), .B(B[18]), .Z(DIFF[18]) );
  XOR2_X1 U121 ( .A(n243), .B(B[17]), .Z(DIFF[17]) );
  XOR2_X1 U122 ( .A(n245), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U124 ( .A(n247), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U125 ( .A(n249), .B(B[11]), .Z(DIFF[11]) );
  NAND2_X1 U1 ( .A1(n197), .A2(n251), .ZN(n196) );
  NOR3_X1 U2 ( .A1(B[59]), .A2(B[60]), .A3(n198), .ZN(n197) );
  NOR2_X1 U3 ( .A1(B[55]), .A2(n202), .ZN(n203) );
  NOR2_X1 U4 ( .A1(B[59]), .A2(n198), .ZN(n199) );
  OR3_X1 U5 ( .A1(B[57]), .A2(B[58]), .A3(n200), .ZN(n198) );
  OR3_X1 U6 ( .A1(B[53]), .A2(B[54]), .A3(n204), .ZN(n202) );
  OR3_X1 U7 ( .A1(B[55]), .A2(B[56]), .A3(n202), .ZN(n200) );
  OR2_X1 U8 ( .A1(n200), .A2(B[57]), .ZN(n201) );
  OR2_X1 U9 ( .A1(n204), .A2(B[53]), .ZN(n205) );
  OR2_X1 U10 ( .A1(n196), .A2(B[62]), .ZN(n195) );
  NOR2_X1 U11 ( .A1(B[51]), .A2(n206), .ZN(n207) );
  OR3_X1 U12 ( .A1(B[51]), .A2(B[52]), .A3(n206), .ZN(n204) );
  NOR2_X1 U13 ( .A1(B[47]), .A2(n212), .ZN(n213) );
  NOR2_X1 U14 ( .A1(B[43]), .A2(n216), .ZN(n217) );
  NOR2_X1 U15 ( .A1(B[39]), .A2(n220), .ZN(n221) );
  NOR2_X1 U16 ( .A1(B[35]), .A2(n224), .ZN(n225) );
  NOR2_X1 U17 ( .A1(B[31]), .A2(n228), .ZN(n229) );
  NOR2_X1 U18 ( .A1(B[27]), .A2(n233), .ZN(n234) );
  OR3_X1 U19 ( .A1(B[45]), .A2(B[46]), .A3(n214), .ZN(n212) );
  OR3_X1 U20 ( .A1(B[41]), .A2(B[42]), .A3(n218), .ZN(n216) );
  OR3_X1 U21 ( .A1(B[37]), .A2(B[38]), .A3(n222), .ZN(n220) );
  OR3_X1 U22 ( .A1(B[33]), .A2(B[34]), .A3(n226), .ZN(n224) );
  OR3_X1 U23 ( .A1(B[29]), .A2(B[30]), .A3(n230), .ZN(n228) );
  OR3_X1 U24 ( .A1(B[25]), .A2(B[26]), .A3(n235), .ZN(n233) );
  OR3_X1 U25 ( .A1(B[47]), .A2(B[48]), .A3(n212), .ZN(n208) );
  OR3_X1 U26 ( .A1(B[43]), .A2(B[44]), .A3(n216), .ZN(n214) );
  OR3_X1 U27 ( .A1(B[39]), .A2(B[40]), .A3(n220), .ZN(n218) );
  OR3_X1 U28 ( .A1(B[35]), .A2(B[36]), .A3(n224), .ZN(n222) );
  OR3_X1 U29 ( .A1(B[31]), .A2(B[32]), .A3(n228), .ZN(n226) );
  OR3_X1 U30 ( .A1(B[27]), .A2(B[28]), .A3(n233), .ZN(n230) );
  OR2_X1 U31 ( .A1(n214), .A2(B[45]), .ZN(n215) );
  OR2_X1 U32 ( .A1(n218), .A2(B[41]), .ZN(n219) );
  OR2_X1 U33 ( .A1(n222), .A2(B[37]), .ZN(n223) );
  OR2_X1 U34 ( .A1(n226), .A2(B[33]), .ZN(n227) );
  OR2_X1 U35 ( .A1(n230), .A2(B[29]), .ZN(n231) );
  OR2_X1 U36 ( .A1(n235), .A2(B[25]), .ZN(n236) );
  OR3_X1 U37 ( .A1(B[49]), .A2(B[50]), .A3(n208), .ZN(n206) );
  OR2_X1 U38 ( .A1(n208), .A2(B[49]), .ZN(n209) );
  NOR2_X1 U39 ( .A1(B[23]), .A2(n237), .ZN(n238) );
  XNOR2_X1 U40 ( .A(B[24]), .B(n238), .ZN(DIFF[24]) );
  OR3_X1 U41 ( .A1(B[23]), .A2(B[24]), .A3(n237), .ZN(n235) );
  XNOR2_X1 U42 ( .A(B[52]), .B(n207), .ZN(DIFF[52]) );
  XNOR2_X1 U43 ( .A(B[48]), .B(n213), .ZN(DIFF[48]) );
  XNOR2_X1 U44 ( .A(B[44]), .B(n217), .ZN(DIFF[44]) );
  XNOR2_X1 U45 ( .A(B[40]), .B(n221), .ZN(DIFF[40]) );
  XNOR2_X1 U46 ( .A(B[36]), .B(n225), .ZN(DIFF[36]) );
  XNOR2_X1 U47 ( .A(B[32]), .B(n229), .ZN(DIFF[32]) );
  XNOR2_X1 U48 ( .A(B[28]), .B(n234), .ZN(DIFF[28]) );
  XNOR2_X1 U49 ( .A(B[56]), .B(n203), .ZN(DIFF[56]) );
  XNOR2_X1 U50 ( .A(n197), .B(B[61]), .ZN(DIFF[61]) );
  XNOR2_X1 U51 ( .A(B[60]), .B(n199), .ZN(DIFF[60]) );
  XNOR2_X1 U52 ( .A(B[20]), .B(n242), .ZN(DIFF[20]) );
  OR3_X1 U53 ( .A1(B[21]), .A2(B[22]), .A3(n239), .ZN(n237) );
  OR2_X1 U54 ( .A1(n239), .A2(B[21]), .ZN(n240) );
  NOR2_X1 U55 ( .A1(B[19]), .A2(n241), .ZN(n242) );
  OR3_X1 U56 ( .A1(B[19]), .A2(B[20]), .A3(n241), .ZN(n239) );
  XNOR2_X1 U57 ( .A(n189), .B(B[14]), .ZN(DIFF[14]) );
  NOR2_X1 U58 ( .A1(n247), .A2(B[13]), .ZN(n189) );
  XNOR2_X1 U59 ( .A(n193), .B(B[10]), .ZN(DIFF[10]) );
  NOR2_X1 U60 ( .A1(n190), .A2(B[9]), .ZN(n193) );
  XNOR2_X1 U61 ( .A(n248), .B(B[6]), .ZN(DIFF[6]) );
  NOR2_X1 U62 ( .A1(n194), .A2(B[5]), .ZN(n248) );
  XNOR2_X1 U63 ( .A(B[16]), .B(n246), .ZN(DIFF[16]) );
  NOR2_X1 U64 ( .A1(B[15]), .A2(n245), .ZN(n246) );
  XNOR2_X1 U65 ( .A(B[12]), .B(n250), .ZN(DIFF[12]) );
  NOR2_X1 U66 ( .A1(B[11]), .A2(n249), .ZN(n250) );
  XNOR2_X1 U67 ( .A(B[8]), .B(n191), .ZN(DIFF[8]) );
  NOR2_X1 U68 ( .A1(B[7]), .A2(n192), .ZN(n191) );
  XNOR2_X1 U69 ( .A(B[2]), .B(n232), .ZN(DIFF[2]) );
  NOR2_X1 U70 ( .A1(\B[0] ), .A2(B[1]), .ZN(n232) );
  XNOR2_X1 U71 ( .A(B[4]), .B(n210), .ZN(DIFF[4]) );
  NOR2_X1 U72 ( .A1(B[3]), .A2(n211), .ZN(n210) );
  OR3_X1 U73 ( .A1(B[5]), .A2(B[6]), .A3(n194), .ZN(n192) );
  OR3_X1 U74 ( .A1(B[10]), .A2(B[9]), .A3(n190), .ZN(n249) );
  OR3_X1 U75 ( .A1(B[13]), .A2(B[14]), .A3(n247), .ZN(n245) );
  OR3_X1 U76 ( .A1(B[17]), .A2(B[18]), .A3(n243), .ZN(n241) );
  OR3_X1 U77 ( .A1(B[7]), .A2(B[8]), .A3(n192), .ZN(n190) );
  OR3_X1 U78 ( .A1(B[11]), .A2(B[12]), .A3(n249), .ZN(n247) );
  OR3_X1 U79 ( .A1(B[15]), .A2(B[16]), .A3(n245), .ZN(n243) );
  OR3_X1 U80 ( .A1(B[3]), .A2(B[4]), .A3(n211), .ZN(n194) );
  OR2_X1 U83 ( .A1(n243), .A2(B[17]), .ZN(n244) );
  OR3_X1 U123 ( .A1(B[1]), .A2(B[2]), .A3(\B[0] ), .ZN(n211) );
  INV_X1 U126 ( .A(B[61]), .ZN(n251) );
endmodule


module complementer_N64_13 ( \input , complement2 );
  input [63:0] \input ;
  output [63:0] complement2;


  complementer_N64_13_DW01_sub_0 sub_add_31_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(\input ), .CI(1'b0), .DIFF(complement2) );
endmodule


module ShiftnCompl_N64_7 ( plusA, plus2A_out, minus2A_out, plus4A_out, 
        minus4A_out );
  input [63:0] plusA;
  output [63:0] plus2A_out;
  output [63:0] minus2A_out;
  output [63:0] plus4A_out;
  output [63:0] minus4A_out;
  wire   n7, n8, n2, n9, n10;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign plus2A_out[0] = 1'b0;
  assign plus2A_out[51] = n2;
  assign plus4A_out[0] = 1'b0;

  shifter_N64_14 shifter_1 ( .\input (plusA), .shiftLeftOnePos({
        plus2A_out[63:59], n7, plus2A_out[57:54], n8, plus2A_out[52], n2, 
        plus2A_out[50:1], SYNOPSYS_UNCONNECTED__0}) );
  shifter_N64_13 shifter_2 ( .\input ({plus2A_out[63:52], n2, plus2A_out[50:1], 
        1'b0}), .shiftLeftOnePos({plus4A_out[63:59], n9, plus4A_out[57:54], 
        n10, plus4A_out[52:1], SYNOPSYS_UNCONNECTED__1}) );
  complementer_N64_14 complementer_1 ( .\input ({plus2A_out[63:52], n2, 
        plus2A_out[50:1], 1'b0}), .complement2(minus2A_out) );
  complementer_N64_13 complementer_2 ( .\input ({plus4A_out[63:1], 1'b0}), 
        .complement2(minus4A_out) );
  BUF_X1 U1 ( .A(n10), .Z(plus4A_out[53]) );
  BUF_X1 U4 ( .A(n8), .Z(plus2A_out[53]) );
  BUF_X1 U5 ( .A(n9), .Z(plus4A_out[58]) );
  BUF_X1 U6 ( .A(n7), .Z(plus2A_out[58]) );
endmodule


module MUX_GENERIC_N64_RADIX3_7 ( plusA, minusA, plus2A, minus2A, SEL, Y );
  input [63:0] plusA;
  input [63:0] minusA;
  input [63:0] plus2A;
  input [63:0] minus2A;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502;
  tri   [63:0] Y;

  TBUF_X1 \Y_tri[55]  ( .A(n446), .EN(n301), .Z(Y[55]) );
  TBUF_X1 \Y_tri[56]  ( .A(n445), .EN(n301), .Z(Y[56]) );
  TBUF_X1 \Y_tri[57]  ( .A(n444), .EN(n301), .Z(Y[57]) );
  TBUF_X1 \Y_tri[58]  ( .A(n443), .EN(n301), .Z(Y[58]) );
  TBUF_X1 \Y_tri[59]  ( .A(n442), .EN(n301), .Z(Y[59]) );
  TBUF_X1 \Y_tri[60]  ( .A(n441), .EN(n301), .Z(Y[60]) );
  TBUF_X1 \Y_tri[61]  ( .A(n440), .EN(n301), .Z(Y[61]) );
  TBUF_X1 \Y_tri[62]  ( .A(n439), .EN(n301), .Z(Y[62]) );
  TBUF_X1 \Y_tri[63]  ( .A(n438), .EN(n301), .Z(Y[63]) );
  TBUF_X1 \Y_tri[53]  ( .A(n448), .EN(n300), .Z(Y[53]) );
  TBUF_X1 \Y_tri[54]  ( .A(n447), .EN(n300), .Z(Y[54]) );
  TBUF_X1 \Y_tri[28]  ( .A(n473), .EN(n298), .Z(Y[28]) );
  TBUF_X1 \Y_tri[29]  ( .A(n472), .EN(n298), .Z(Y[29]) );
  TBUF_X1 \Y_tri[30]  ( .A(n471), .EN(n298), .Z(Y[30]) );
  TBUF_X1 \Y_tri[31]  ( .A(n470), .EN(n298), .Z(Y[31]) );
  TBUF_X1 \Y_tri[32]  ( .A(n469), .EN(n298), .Z(Y[32]) );
  TBUF_X1 \Y_tri[33]  ( .A(n468), .EN(n299), .Z(Y[33]) );
  TBUF_X1 \Y_tri[34]  ( .A(n467), .EN(n299), .Z(Y[34]) );
  TBUF_X1 \Y_tri[35]  ( .A(n466), .EN(n299), .Z(Y[35]) );
  TBUF_X1 \Y_tri[36]  ( .A(n465), .EN(n299), .Z(Y[36]) );
  TBUF_X1 \Y_tri[37]  ( .A(n464), .EN(n299), .Z(Y[37]) );
  TBUF_X1 \Y_tri[38]  ( .A(n463), .EN(n299), .Z(Y[38]) );
  TBUF_X1 \Y_tri[39]  ( .A(n462), .EN(n299), .Z(Y[39]) );
  TBUF_X1 \Y_tri[40]  ( .A(n461), .EN(n299), .Z(Y[40]) );
  TBUF_X1 \Y_tri[41]  ( .A(n460), .EN(n299), .Z(Y[41]) );
  TBUF_X1 \Y_tri[42]  ( .A(n459), .EN(n299), .Z(Y[42]) );
  TBUF_X1 \Y_tri[43]  ( .A(n458), .EN(n299), .Z(Y[43]) );
  TBUF_X1 \Y_tri[44]  ( .A(n457), .EN(n300), .Z(Y[44]) );
  TBUF_X1 \Y_tri[45]  ( .A(n456), .EN(n300), .Z(Y[45]) );
  TBUF_X1 \Y_tri[46]  ( .A(n455), .EN(n300), .Z(Y[46]) );
  TBUF_X1 \Y_tri[47]  ( .A(n454), .EN(n300), .Z(Y[47]) );
  TBUF_X1 \Y_tri[48]  ( .A(n453), .EN(n300), .Z(Y[48]) );
  TBUF_X1 \Y_tri[49]  ( .A(n452), .EN(n300), .Z(Y[49]) );
  TBUF_X1 \Y_tri[50]  ( .A(n451), .EN(n300), .Z(Y[50]) );
  TBUF_X1 \Y_tri[51]  ( .A(n450), .EN(n300), .Z(Y[51]) );
  TBUF_X1 \Y_tri[52]  ( .A(n449), .EN(n300), .Z(Y[52]) );
  TBUF_X1 \Y_tri[10]  ( .A(n491), .EN(n296), .Z(Y[10]) );
  TBUF_X1 \Y_tri[12]  ( .A(n489), .EN(n297), .Z(Y[12]) );
  TBUF_X1 \Y_tri[13]  ( .A(n488), .EN(n297), .Z(Y[13]) );
  TBUF_X1 \Y_tri[14]  ( .A(n487), .EN(n297), .Z(Y[14]) );
  TBUF_X1 \Y_tri[15]  ( .A(n486), .EN(n297), .Z(Y[15]) );
  TBUF_X1 \Y_tri[16]  ( .A(n485), .EN(n297), .Z(Y[16]) );
  TBUF_X1 \Y_tri[18]  ( .A(n483), .EN(n297), .Z(Y[18]) );
  TBUF_X1 \Y_tri[19]  ( .A(n482), .EN(n297), .Z(Y[19]) );
  TBUF_X1 \Y_tri[20]  ( .A(n481), .EN(n297), .Z(Y[20]) );
  TBUF_X1 \Y_tri[21]  ( .A(n480), .EN(n297), .Z(Y[21]) );
  TBUF_X1 \Y_tri[22]  ( .A(n479), .EN(n298), .Z(Y[22]) );
  TBUF_X1 \Y_tri[23]  ( .A(n478), .EN(n298), .Z(Y[23]) );
  TBUF_X1 \Y_tri[24]  ( .A(n477), .EN(n298), .Z(Y[24]) );
  TBUF_X1 \Y_tri[25]  ( .A(n476), .EN(n298), .Z(Y[25]) );
  TBUF_X1 \Y_tri[26]  ( .A(n475), .EN(n298), .Z(Y[26]) );
  TBUF_X1 \Y_tri[27]  ( .A(n474), .EN(n298), .Z(Y[27]) );
  TBUF_X1 \Y_tri[9]  ( .A(n492), .EN(n296), .Z(Y[9]) );
  TBUF_X1 \Y_tri[11]  ( .A(n490), .EN(n297), .Z(Y[11]) );
  TBUF_X1 \Y_tri[0]  ( .A(n502), .EN(n296), .Z(Y[0]) );
  TBUF_X1 \Y_tri[1]  ( .A(n501), .EN(n296), .Z(Y[1]) );
  TBUF_X1 \Y_tri[2]  ( .A(n500), .EN(n296), .Z(Y[2]) );
  TBUF_X1 \Y_tri[3]  ( .A(n499), .EN(n296), .Z(Y[3]) );
  TBUF_X1 \Y_tri[4]  ( .A(n498), .EN(n296), .Z(Y[4]) );
  TBUF_X1 \Y_tri[5]  ( .A(n497), .EN(n296), .Z(Y[5]) );
  TBUF_X1 \Y_tri[6]  ( .A(n496), .EN(n296), .Z(Y[6]) );
  TBUF_X1 \Y_tri[7]  ( .A(n495), .EN(n296), .Z(Y[7]) );
  TBUF_X1 \Y_tri[8]  ( .A(n494), .EN(n296), .Z(Y[8]) );
  TBUF_X1 \Y_tri[17]  ( .A(n484), .EN(n297), .Z(Y[17]) );
  NAND2_X1 U2 ( .A1(n351), .A2(n350), .ZN(n479) );
  AOI22_X1 U3 ( .A1(plusA[22]), .A2(n279), .B1(plus2A[22]), .B2(n273), .ZN(
        n351) );
  AOI22_X1 U4 ( .A1(minus2A[22]), .A2(n291), .B1(minusA[22]), .B2(n285), .ZN(
        n350) );
  NAND2_X1 U5 ( .A1(n357), .A2(n356), .ZN(n476) );
  AOI22_X1 U6 ( .A1(plusA[25]), .A2(n280), .B1(plus2A[25]), .B2(n274), .ZN(
        n357) );
  AOI22_X1 U7 ( .A1(minus2A[25]), .A2(n292), .B1(minusA[25]), .B2(n286), .ZN(
        n356) );
  NAND2_X1 U8 ( .A1(n361), .A2(n360), .ZN(n474) );
  AOI22_X1 U9 ( .A1(plusA[27]), .A2(n280), .B1(plus2A[27]), .B2(n274), .ZN(
        n361) );
  AOI22_X1 U10 ( .A1(minus2A[27]), .A2(n292), .B1(minusA[27]), .B2(n286), .ZN(
        n360) );
  NAND2_X1 U11 ( .A1(n353), .A2(n352), .ZN(n478) );
  AOI22_X1 U12 ( .A1(plusA[23]), .A2(n279), .B1(plus2A[23]), .B2(n273), .ZN(
        n353) );
  AOI22_X1 U13 ( .A1(minus2A[23]), .A2(n291), .B1(minusA[23]), .B2(n285), .ZN(
        n352) );
  NAND2_X1 U14 ( .A1(n359), .A2(n358), .ZN(n475) );
  AOI22_X1 U15 ( .A1(plusA[26]), .A2(n280), .B1(plus2A[26]), .B2(n274), .ZN(
        n359) );
  AOI22_X1 U16 ( .A1(minus2A[26]), .A2(n292), .B1(minusA[26]), .B2(n286), .ZN(
        n358) );
  NAND2_X1 U17 ( .A1(n355), .A2(n354), .ZN(n477) );
  AOI22_X1 U18 ( .A1(plusA[24]), .A2(n280), .B1(plus2A[24]), .B2(n274), .ZN(
        n355) );
  AOI22_X1 U19 ( .A1(minus2A[24]), .A2(n292), .B1(minusA[24]), .B2(n286), .ZN(
        n354) );
  NAND2_X1 U20 ( .A1(n407), .A2(n406), .ZN(n451) );
  AOI22_X1 U21 ( .A1(plusA[50]), .A2(n282), .B1(plus2A[50]), .B2(n276), .ZN(
        n407) );
  AOI22_X1 U22 ( .A1(minus2A[50]), .A2(n294), .B1(minusA[50]), .B2(n288), .ZN(
        n406) );
  NAND2_X1 U23 ( .A1(n397), .A2(n396), .ZN(n456) );
  AOI22_X1 U24 ( .A1(plusA[45]), .A2(n281), .B1(plus2A[45]), .B2(n275), .ZN(
        n397) );
  AOI22_X1 U25 ( .A1(minus2A[45]), .A2(n293), .B1(minusA[45]), .B2(n287), .ZN(
        n396) );
  NAND2_X1 U26 ( .A1(n389), .A2(n388), .ZN(n460) );
  AOI22_X1 U27 ( .A1(plusA[41]), .A2(n281), .B1(plus2A[41]), .B2(n275), .ZN(
        n389) );
  AOI22_X1 U28 ( .A1(minus2A[41]), .A2(n293), .B1(minusA[41]), .B2(n287), .ZN(
        n388) );
  NAND2_X1 U29 ( .A1(n381), .A2(n380), .ZN(n464) );
  AOI22_X1 U30 ( .A1(plusA[37]), .A2(n281), .B1(plus2A[37]), .B2(n275), .ZN(
        n381) );
  AOI22_X1 U31 ( .A1(minus2A[37]), .A2(n293), .B1(minusA[37]), .B2(n287), .ZN(
        n380) );
  NAND2_X1 U32 ( .A1(n373), .A2(n372), .ZN(n468) );
  AOI22_X1 U33 ( .A1(plusA[33]), .A2(n280), .B1(plus2A[33]), .B2(n274), .ZN(
        n373) );
  AOI22_X1 U34 ( .A1(minus2A[33]), .A2(n292), .B1(minusA[33]), .B2(n286), .ZN(
        n372) );
  NAND2_X1 U35 ( .A1(n365), .A2(n364), .ZN(n472) );
  AOI22_X1 U36 ( .A1(plusA[29]), .A2(n280), .B1(plus2A[29]), .B2(n274), .ZN(
        n365) );
  AOI22_X1 U37 ( .A1(minus2A[29]), .A2(n292), .B1(minusA[29]), .B2(n286), .ZN(
        n364) );
  NAND2_X1 U38 ( .A1(n401), .A2(n400), .ZN(n454) );
  AOI22_X1 U39 ( .A1(plusA[47]), .A2(n281), .B1(plus2A[47]), .B2(n275), .ZN(
        n401) );
  AOI22_X1 U40 ( .A1(minus2A[47]), .A2(n293), .B1(minusA[47]), .B2(n287), .ZN(
        n400) );
  NAND2_X1 U41 ( .A1(n393), .A2(n392), .ZN(n458) );
  AOI22_X1 U42 ( .A1(plusA[43]), .A2(n281), .B1(plus2A[43]), .B2(n275), .ZN(
        n393) );
  AOI22_X1 U43 ( .A1(minus2A[43]), .A2(n293), .B1(minusA[43]), .B2(n287), .ZN(
        n392) );
  NAND2_X1 U44 ( .A1(n385), .A2(n384), .ZN(n462) );
  AOI22_X1 U45 ( .A1(plusA[39]), .A2(n281), .B1(plus2A[39]), .B2(n275), .ZN(
        n385) );
  AOI22_X1 U46 ( .A1(minus2A[39]), .A2(n293), .B1(minusA[39]), .B2(n287), .ZN(
        n384) );
  NAND2_X1 U47 ( .A1(n377), .A2(n376), .ZN(n466) );
  AOI22_X1 U48 ( .A1(plusA[35]), .A2(n280), .B1(plus2A[35]), .B2(n274), .ZN(
        n377) );
  AOI22_X1 U49 ( .A1(minus2A[35]), .A2(n292), .B1(minusA[35]), .B2(n286), .ZN(
        n376) );
  NAND2_X1 U50 ( .A1(n369), .A2(n368), .ZN(n470) );
  AOI22_X1 U51 ( .A1(plusA[31]), .A2(n280), .B1(plus2A[31]), .B2(n274), .ZN(
        n369) );
  AOI22_X1 U52 ( .A1(minus2A[31]), .A2(n292), .B1(minusA[31]), .B2(n286), .ZN(
        n368) );
  NAND2_X1 U53 ( .A1(n409), .A2(n408), .ZN(n450) );
  AOI22_X1 U54 ( .A1(plusA[51]), .A2(n282), .B1(plus2A[51]), .B2(n276), .ZN(
        n409) );
  AOI22_X1 U55 ( .A1(minus2A[51]), .A2(n294), .B1(minusA[51]), .B2(n288), .ZN(
        n408) );
  NAND2_X1 U56 ( .A1(n411), .A2(n410), .ZN(n449) );
  AOI22_X1 U57 ( .A1(plusA[52]), .A2(n282), .B1(plus2A[52]), .B2(n276), .ZN(
        n411) );
  AOI22_X1 U58 ( .A1(minus2A[52]), .A2(n294), .B1(minusA[52]), .B2(n288), .ZN(
        n410) );
  NAND2_X1 U59 ( .A1(n399), .A2(n398), .ZN(n455) );
  AOI22_X1 U60 ( .A1(plusA[46]), .A2(n281), .B1(plus2A[46]), .B2(n275), .ZN(
        n399) );
  AOI22_X1 U61 ( .A1(minus2A[46]), .A2(n293), .B1(minusA[46]), .B2(n287), .ZN(
        n398) );
  NAND2_X1 U62 ( .A1(n391), .A2(n390), .ZN(n459) );
  AOI22_X1 U63 ( .A1(plusA[42]), .A2(n281), .B1(plus2A[42]), .B2(n275), .ZN(
        n391) );
  AOI22_X1 U64 ( .A1(minus2A[42]), .A2(n293), .B1(minusA[42]), .B2(n287), .ZN(
        n390) );
  NAND2_X1 U65 ( .A1(n383), .A2(n382), .ZN(n463) );
  AOI22_X1 U66 ( .A1(plusA[38]), .A2(n281), .B1(plus2A[38]), .B2(n275), .ZN(
        n383) );
  AOI22_X1 U67 ( .A1(minus2A[38]), .A2(n293), .B1(minusA[38]), .B2(n287), .ZN(
        n382) );
  NAND2_X1 U68 ( .A1(n375), .A2(n374), .ZN(n467) );
  AOI22_X1 U69 ( .A1(plusA[34]), .A2(n280), .B1(plus2A[34]), .B2(n274), .ZN(
        n375) );
  AOI22_X1 U70 ( .A1(minus2A[34]), .A2(n292), .B1(minusA[34]), .B2(n286), .ZN(
        n374) );
  NAND2_X1 U71 ( .A1(n367), .A2(n366), .ZN(n471) );
  AOI22_X1 U72 ( .A1(plusA[30]), .A2(n280), .B1(plus2A[30]), .B2(n274), .ZN(
        n367) );
  AOI22_X1 U73 ( .A1(minus2A[30]), .A2(n292), .B1(minusA[30]), .B2(n286), .ZN(
        n366) );
  NAND2_X1 U74 ( .A1(n405), .A2(n404), .ZN(n452) );
  AOI22_X1 U75 ( .A1(plusA[49]), .A2(n282), .B1(plus2A[49]), .B2(n276), .ZN(
        n405) );
  AOI22_X1 U76 ( .A1(minus2A[49]), .A2(n294), .B1(minusA[49]), .B2(n288), .ZN(
        n404) );
  NAND2_X1 U77 ( .A1(n403), .A2(n402), .ZN(n453) );
  AOI22_X1 U78 ( .A1(plusA[48]), .A2(n282), .B1(plus2A[48]), .B2(n276), .ZN(
        n403) );
  AOI22_X1 U79 ( .A1(minus2A[48]), .A2(n294), .B1(minusA[48]), .B2(n288), .ZN(
        n402) );
  NAND2_X1 U80 ( .A1(n395), .A2(n394), .ZN(n457) );
  AOI22_X1 U81 ( .A1(plusA[44]), .A2(n281), .B1(plus2A[44]), .B2(n275), .ZN(
        n395) );
  AOI22_X1 U82 ( .A1(minus2A[44]), .A2(n293), .B1(minusA[44]), .B2(n287), .ZN(
        n394) );
  NAND2_X1 U83 ( .A1(n387), .A2(n386), .ZN(n461) );
  AOI22_X1 U84 ( .A1(plusA[40]), .A2(n281), .B1(plus2A[40]), .B2(n275), .ZN(
        n387) );
  AOI22_X1 U85 ( .A1(minus2A[40]), .A2(n293), .B1(minusA[40]), .B2(n287), .ZN(
        n386) );
  NAND2_X1 U86 ( .A1(n379), .A2(n378), .ZN(n465) );
  AOI22_X1 U87 ( .A1(plusA[36]), .A2(n281), .B1(plus2A[36]), .B2(n275), .ZN(
        n379) );
  AOI22_X1 U88 ( .A1(minus2A[36]), .A2(n293), .B1(minusA[36]), .B2(n287), .ZN(
        n378) );
  NAND2_X1 U89 ( .A1(n371), .A2(n370), .ZN(n469) );
  AOI22_X1 U90 ( .A1(plusA[32]), .A2(n280), .B1(plus2A[32]), .B2(n274), .ZN(
        n371) );
  AOI22_X1 U91 ( .A1(minus2A[32]), .A2(n292), .B1(minusA[32]), .B2(n286), .ZN(
        n370) );
  NAND2_X1 U92 ( .A1(n363), .A2(n362), .ZN(n473) );
  AOI22_X1 U93 ( .A1(plusA[28]), .A2(n280), .B1(plus2A[28]), .B2(n274), .ZN(
        n363) );
  AOI22_X1 U94 ( .A1(minus2A[28]), .A2(n292), .B1(minusA[28]), .B2(n286), .ZN(
        n362) );
  NAND2_X1 U95 ( .A1(n419), .A2(n418), .ZN(n445) );
  AOI22_X1 U96 ( .A1(plusA[56]), .A2(n282), .B1(plus2A[56]), .B2(n276), .ZN(
        n419) );
  AOI22_X1 U97 ( .A1(minus2A[56]), .A2(n294), .B1(minusA[56]), .B2(n288), .ZN(
        n418) );
  NAND2_X1 U98 ( .A1(n415), .A2(n414), .ZN(n447) );
  AOI22_X1 U99 ( .A1(plusA[54]), .A2(n282), .B1(plus2A[54]), .B2(n276), .ZN(
        n415) );
  AOI22_X1 U100 ( .A1(minus2A[54]), .A2(n294), .B1(minusA[54]), .B2(n288), 
        .ZN(n414) );
  NAND2_X1 U101 ( .A1(n421), .A2(n420), .ZN(n444) );
  AOI22_X1 U102 ( .A1(plusA[57]), .A2(n282), .B1(plus2A[57]), .B2(n276), .ZN(
        n421) );
  AOI22_X1 U103 ( .A1(minus2A[57]), .A2(n294), .B1(minusA[57]), .B2(n288), 
        .ZN(n420) );
  NAND2_X1 U104 ( .A1(n417), .A2(n416), .ZN(n446) );
  AOI22_X1 U105 ( .A1(plusA[55]), .A2(n282), .B1(plus2A[55]), .B2(n276), .ZN(
        n417) );
  AOI22_X1 U106 ( .A1(minus2A[55]), .A2(n294), .B1(minusA[55]), .B2(n288), 
        .ZN(n416) );
  NAND2_X1 U107 ( .A1(n413), .A2(n412), .ZN(n448) );
  AOI22_X1 U108 ( .A1(plusA[53]), .A2(n282), .B1(plus2A[53]), .B2(n276), .ZN(
        n413) );
  AOI22_X1 U109 ( .A1(minus2A[53]), .A2(n294), .B1(minusA[53]), .B2(n288), 
        .ZN(n412) );
  NAND2_X1 U110 ( .A1(n437), .A2(n436), .ZN(n438) );
  AOI22_X1 U111 ( .A1(plusA[63]), .A2(n283), .B1(plus2A[63]), .B2(n277), .ZN(
        n437) );
  AOI22_X1 U112 ( .A1(minus2A[63]), .A2(n295), .B1(minusA[63]), .B2(n289), 
        .ZN(n436) );
  NAND2_X1 U113 ( .A1(n431), .A2(n430), .ZN(n439) );
  AOI22_X1 U114 ( .A1(plusA[62]), .A2(n283), .B1(plus2A[62]), .B2(n277), .ZN(
        n431) );
  AOI22_X1 U115 ( .A1(minus2A[62]), .A2(n295), .B1(minusA[62]), .B2(n289), 
        .ZN(n430) );
  NAND2_X1 U116 ( .A1(n429), .A2(n428), .ZN(n440) );
  AOI22_X1 U117 ( .A1(plusA[61]), .A2(n283), .B1(plus2A[61]), .B2(n277), .ZN(
        n429) );
  AOI22_X1 U118 ( .A1(minus2A[61]), .A2(n295), .B1(minusA[61]), .B2(n289), 
        .ZN(n428) );
  NAND2_X1 U119 ( .A1(n427), .A2(n426), .ZN(n441) );
  AOI22_X1 U120 ( .A1(plusA[60]), .A2(n283), .B1(plus2A[60]), .B2(n277), .ZN(
        n427) );
  AOI22_X1 U121 ( .A1(minus2A[60]), .A2(n295), .B1(minusA[60]), .B2(n289), 
        .ZN(n426) );
  NAND2_X1 U122 ( .A1(n425), .A2(n424), .ZN(n442) );
  AOI22_X1 U123 ( .A1(plusA[59]), .A2(n282), .B1(plus2A[59]), .B2(n276), .ZN(
        n425) );
  AOI22_X1 U124 ( .A1(minus2A[59]), .A2(n294), .B1(minusA[59]), .B2(n288), 
        .ZN(n424) );
  NAND2_X1 U125 ( .A1(n423), .A2(n422), .ZN(n443) );
  AOI22_X1 U126 ( .A1(plusA[58]), .A2(n282), .B1(plus2A[58]), .B2(n276), .ZN(
        n423) );
  AOI22_X1 U127 ( .A1(minus2A[58]), .A2(n294), .B1(minusA[58]), .B2(n288), 
        .ZN(n422) );
  BUF_X1 U128 ( .A(n493), .Z(n296) );
  BUF_X1 U129 ( .A(n433), .Z(n279) );
  BUF_X1 U130 ( .A(n434), .Z(n285) );
  BUF_X1 U131 ( .A(n432), .Z(n273) );
  BUF_X1 U132 ( .A(n493), .Z(n297) );
  NAND2_X1 U133 ( .A1(n349), .A2(n348), .ZN(n480) );
  AOI22_X1 U134 ( .A1(plusA[21]), .A2(n279), .B1(plus2A[21]), .B2(n273), .ZN(
        n349) );
  AOI22_X1 U135 ( .A1(minus2A[21]), .A2(n291), .B1(minusA[21]), .B2(n285), 
        .ZN(n348) );
  NAND2_X1 U136 ( .A1(n347), .A2(n346), .ZN(n481) );
  AOI22_X1 U137 ( .A1(plusA[20]), .A2(n279), .B1(plus2A[20]), .B2(n273), .ZN(
        n347) );
  AOI22_X1 U138 ( .A1(minus2A[20]), .A2(n291), .B1(minusA[20]), .B2(n285), 
        .ZN(n346) );
  BUF_X1 U139 ( .A(n433), .Z(n280) );
  BUF_X1 U140 ( .A(n435), .Z(n292) );
  BUF_X1 U141 ( .A(n435), .Z(n291) );
  BUF_X1 U142 ( .A(n434), .Z(n286) );
  BUF_X1 U143 ( .A(n432), .Z(n274) );
  BUF_X1 U144 ( .A(n493), .Z(n298) );
  BUF_X1 U145 ( .A(n433), .Z(n281) );
  BUF_X1 U146 ( .A(n435), .Z(n293) );
  BUF_X1 U147 ( .A(n434), .Z(n287) );
  BUF_X1 U148 ( .A(n432), .Z(n275) );
  BUF_X1 U149 ( .A(n493), .Z(n299) );
  BUF_X1 U150 ( .A(n433), .Z(n282) );
  BUF_X1 U151 ( .A(n435), .Z(n294) );
  BUF_X1 U152 ( .A(n434), .Z(n288) );
  BUF_X1 U153 ( .A(n432), .Z(n276) );
  BUF_X1 U154 ( .A(n493), .Z(n300) );
  BUF_X1 U155 ( .A(n493), .Z(n301) );
  BUF_X1 U156 ( .A(n433), .Z(n278) );
  BUF_X1 U157 ( .A(n435), .Z(n290) );
  BUF_X1 U158 ( .A(n434), .Z(n284) );
  BUF_X1 U159 ( .A(n432), .Z(n272) );
  NOR2_X1 U160 ( .A1(n323), .A2(n304), .ZN(n493) );
  INV_X1 U161 ( .A(SEL[2]), .ZN(n304) );
  NOR2_X1 U162 ( .A1(SEL[1]), .A2(SEL[0]), .ZN(n323) );
  NOR3_X1 U163 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n302), .ZN(n434) );
  NOR3_X1 U164 ( .A1(SEL[1]), .A2(SEL[2]), .A3(n303), .ZN(n433) );
  NOR3_X1 U165 ( .A1(n302), .A2(SEL[2]), .A3(n303), .ZN(n432) );
  NAND2_X1 U166 ( .A1(n345), .A2(n344), .ZN(n482) );
  AOI22_X1 U167 ( .A1(plusA[19]), .A2(n279), .B1(plus2A[19]), .B2(n273), .ZN(
        n345) );
  AOI22_X1 U168 ( .A1(minus2A[19]), .A2(n291), .B1(minusA[19]), .B2(n285), 
        .ZN(n344) );
  INV_X1 U169 ( .A(SEL[1]), .ZN(n302) );
  INV_X1 U170 ( .A(SEL[0]), .ZN(n303) );
  AND2_X1 U171 ( .A1(SEL[2]), .A2(n323), .ZN(n435) );
  NAND2_X1 U172 ( .A1(n343), .A2(n342), .ZN(n483) );
  AOI22_X1 U173 ( .A1(plusA[18]), .A2(n279), .B1(plus2A[18]), .B2(n273), .ZN(
        n343) );
  AOI22_X1 U174 ( .A1(minus2A[18]), .A2(n291), .B1(minusA[18]), .B2(n285), 
        .ZN(n342) );
  NAND2_X1 U175 ( .A1(n341), .A2(n340), .ZN(n484) );
  AOI22_X1 U176 ( .A1(plusA[17]), .A2(n279), .B1(plus2A[17]), .B2(n273), .ZN(
        n341) );
  AOI22_X1 U177 ( .A1(minus2A[17]), .A2(n291), .B1(minusA[17]), .B2(n285), 
        .ZN(n340) );
  NAND2_X1 U178 ( .A1(n337), .A2(n336), .ZN(n486) );
  AOI22_X1 U179 ( .A1(plusA[15]), .A2(n279), .B1(plus2A[15]), .B2(n273), .ZN(
        n337) );
  AOI22_X1 U180 ( .A1(minus2A[15]), .A2(n291), .B1(minusA[15]), .B2(n285), 
        .ZN(n336) );
  NAND2_X1 U181 ( .A1(n335), .A2(n334), .ZN(n487) );
  AOI22_X1 U182 ( .A1(plusA[14]), .A2(n279), .B1(plus2A[14]), .B2(n273), .ZN(
        n335) );
  AOI22_X1 U183 ( .A1(minus2A[14]), .A2(n291), .B1(minusA[14]), .B2(n285), 
        .ZN(n334) );
  NAND2_X1 U184 ( .A1(n333), .A2(n332), .ZN(n488) );
  AOI22_X1 U185 ( .A1(plusA[13]), .A2(n279), .B1(plus2A[13]), .B2(n273), .ZN(
        n333) );
  AOI22_X1 U186 ( .A1(minus2A[13]), .A2(n291), .B1(minusA[13]), .B2(n285), 
        .ZN(n332) );
  NAND2_X1 U187 ( .A1(n329), .A2(n328), .ZN(n490) );
  AOI22_X1 U188 ( .A1(plusA[11]), .A2(n278), .B1(plus2A[11]), .B2(n272), .ZN(
        n329) );
  AOI22_X1 U189 ( .A1(minus2A[11]), .A2(n290), .B1(minusA[11]), .B2(n284), 
        .ZN(n328) );
  NAND2_X1 U190 ( .A1(n327), .A2(n326), .ZN(n491) );
  AOI22_X1 U191 ( .A1(plusA[10]), .A2(n278), .B1(plus2A[10]), .B2(n272), .ZN(
        n327) );
  AOI22_X1 U192 ( .A1(minus2A[10]), .A2(n290), .B1(minusA[10]), .B2(n284), 
        .ZN(n326) );
  NAND2_X1 U193 ( .A1(n325), .A2(n324), .ZN(n492) );
  AOI22_X1 U194 ( .A1(plusA[9]), .A2(n278), .B1(plus2A[9]), .B2(n272), .ZN(
        n325) );
  AOI22_X1 U195 ( .A1(minus2A[9]), .A2(n290), .B1(minusA[9]), .B2(n284), .ZN(
        n324) );
  NAND2_X1 U196 ( .A1(n320), .A2(n319), .ZN(n495) );
  AOI22_X1 U197 ( .A1(plusA[7]), .A2(n278), .B1(plus2A[7]), .B2(n272), .ZN(
        n320) );
  AOI22_X1 U198 ( .A1(minus2A[7]), .A2(n290), .B1(minusA[7]), .B2(n284), .ZN(
        n319) );
  NAND2_X1 U199 ( .A1(n318), .A2(n317), .ZN(n496) );
  AOI22_X1 U200 ( .A1(plusA[6]), .A2(n278), .B1(plus2A[6]), .B2(n272), .ZN(
        n318) );
  AOI22_X1 U201 ( .A1(minus2A[6]), .A2(n290), .B1(minusA[6]), .B2(n284), .ZN(
        n317) );
  NAND2_X1 U202 ( .A1(n316), .A2(n315), .ZN(n497) );
  AOI22_X1 U203 ( .A1(plusA[5]), .A2(n278), .B1(plus2A[5]), .B2(n272), .ZN(
        n316) );
  AOI22_X1 U204 ( .A1(minus2A[5]), .A2(n290), .B1(minusA[5]), .B2(n284), .ZN(
        n315) );
  NAND2_X1 U205 ( .A1(n312), .A2(n311), .ZN(n499) );
  AOI22_X1 U206 ( .A1(plusA[3]), .A2(n278), .B1(plus2A[3]), .B2(n272), .ZN(
        n312) );
  AOI22_X1 U207 ( .A1(minus2A[3]), .A2(n290), .B1(minusA[3]), .B2(n284), .ZN(
        n311) );
  NAND2_X1 U208 ( .A1(n339), .A2(n338), .ZN(n485) );
  AOI22_X1 U209 ( .A1(plusA[16]), .A2(n279), .B1(plus2A[16]), .B2(n273), .ZN(
        n339) );
  AOI22_X1 U210 ( .A1(minus2A[16]), .A2(n291), .B1(minusA[16]), .B2(n285), 
        .ZN(n338) );
  NAND2_X1 U211 ( .A1(n331), .A2(n330), .ZN(n489) );
  AOI22_X1 U212 ( .A1(plusA[12]), .A2(n279), .B1(plus2A[12]), .B2(n273), .ZN(
        n331) );
  AOI22_X1 U213 ( .A1(minus2A[12]), .A2(n291), .B1(minusA[12]), .B2(n285), 
        .ZN(n330) );
  NAND2_X1 U214 ( .A1(n322), .A2(n321), .ZN(n494) );
  AOI22_X1 U215 ( .A1(plusA[8]), .A2(n278), .B1(plus2A[8]), .B2(n272), .ZN(
        n322) );
  AOI22_X1 U216 ( .A1(minus2A[8]), .A2(n290), .B1(minusA[8]), .B2(n284), .ZN(
        n321) );
  NAND2_X1 U217 ( .A1(n314), .A2(n313), .ZN(n498) );
  AOI22_X1 U218 ( .A1(plusA[4]), .A2(n278), .B1(plus2A[4]), .B2(n272), .ZN(
        n314) );
  AOI22_X1 U219 ( .A1(minus2A[4]), .A2(n290), .B1(minusA[4]), .B2(n284), .ZN(
        n313) );
  NAND2_X1 U220 ( .A1(n310), .A2(n309), .ZN(n500) );
  AOI22_X1 U221 ( .A1(plusA[2]), .A2(n278), .B1(plus2A[2]), .B2(n272), .ZN(
        n310) );
  AOI22_X1 U222 ( .A1(minus2A[2]), .A2(n290), .B1(minusA[2]), .B2(n284), .ZN(
        n309) );
  NAND2_X1 U223 ( .A1(n308), .A2(n307), .ZN(n501) );
  AOI22_X1 U224 ( .A1(plusA[1]), .A2(n278), .B1(plus2A[1]), .B2(n272), .ZN(
        n308) );
  AOI22_X1 U225 ( .A1(minus2A[1]), .A2(n290), .B1(minusA[1]), .B2(n284), .ZN(
        n307) );
  NAND2_X1 U226 ( .A1(n306), .A2(n305), .ZN(n502) );
  AOI22_X1 U227 ( .A1(plusA[0]), .A2(n278), .B1(plus2A[0]), .B2(n272), .ZN(
        n306) );
  AOI22_X1 U228 ( .A1(minus2A[0]), .A2(n290), .B1(minusA[0]), .B2(n284), .ZN(
        n305) );
  CLKBUF_X1 U229 ( .A(n432), .Z(n277) );
  CLKBUF_X1 U230 ( .A(n433), .Z(n283) );
  CLKBUF_X1 U231 ( .A(n434), .Z(n289) );
  CLKBUF_X1 U232 ( .A(n435), .Z(n295) );
endmodule


module FA_448 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_447 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_446 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_445 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_444 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_443 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_442 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_441 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_440 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_439 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(n5), .B(Ci), .Z(S) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_438 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_437 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_436 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_435 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_434 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_433 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_432 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_431 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  AOI22_X1 U4 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
  INV_X1 U5 ( .A(n7), .ZN(Co) );
endmodule


module FA_430 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_429 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_428 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_427 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_426 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_425 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_424 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_423 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_422 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_421 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_420 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_419 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_418 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_417 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_416 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_415 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_414 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_413 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_412 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_411 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_410 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_409 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_408 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_407 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_406 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_405 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_404 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_403 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_402 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_401 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_400 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_399 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_398 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_397 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_396 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_395 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_394 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_393 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_392 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_391 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_390 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_389 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_388 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_387 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_386 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_385 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N64_7 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Ci;
  output Co;

  wire   [63:1] CTMP;
  tri   [63:0] A;

  FA_448 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_447 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_446 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_445 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(CTMP[4]) );
  FA_444 FAI_5 ( .A(A[4]), .B(B[4]), .Ci(CTMP[4]), .S(S[4]), .Co(CTMP[5]) );
  FA_443 FAI_6 ( .A(A[5]), .B(B[5]), .Ci(CTMP[5]), .S(S[5]), .Co(CTMP[6]) );
  FA_442 FAI_7 ( .A(A[6]), .B(B[6]), .Ci(CTMP[6]), .S(S[6]), .Co(CTMP[7]) );
  FA_441 FAI_8 ( .A(A[7]), .B(B[7]), .Ci(CTMP[7]), .S(S[7]), .Co(CTMP[8]) );
  FA_440 FAI_9 ( .A(A[8]), .B(B[8]), .Ci(CTMP[8]), .S(S[8]), .Co(CTMP[9]) );
  FA_439 FAI_10 ( .A(A[9]), .B(B[9]), .Ci(CTMP[9]), .S(S[9]), .Co(CTMP[10]) );
  FA_438 FAI_11 ( .A(A[10]), .B(B[10]), .Ci(CTMP[10]), .S(S[10]), .Co(CTMP[11]) );
  FA_437 FAI_12 ( .A(A[11]), .B(B[11]), .Ci(CTMP[11]), .S(S[11]), .Co(CTMP[12]) );
  FA_436 FAI_13 ( .A(A[12]), .B(B[12]), .Ci(CTMP[12]), .S(S[12]), .Co(CTMP[13]) );
  FA_435 FAI_14 ( .A(A[13]), .B(B[13]), .Ci(CTMP[13]), .S(S[13]), .Co(CTMP[14]) );
  FA_434 FAI_15 ( .A(A[14]), .B(B[14]), .Ci(CTMP[14]), .S(S[14]), .Co(CTMP[15]) );
  FA_433 FAI_16 ( .A(A[15]), .B(B[15]), .Ci(CTMP[15]), .S(S[15]), .Co(CTMP[16]) );
  FA_432 FAI_17 ( .A(A[16]), .B(B[16]), .Ci(CTMP[16]), .S(S[16]), .Co(CTMP[17]) );
  FA_431 FAI_18 ( .A(A[17]), .B(B[17]), .Ci(CTMP[17]), .S(S[17]), .Co(CTMP[18]) );
  FA_430 FAI_19 ( .A(A[18]), .B(B[18]), .Ci(CTMP[18]), .S(S[18]), .Co(CTMP[19]) );
  FA_429 FAI_20 ( .A(A[19]), .B(B[19]), .Ci(CTMP[19]), .S(S[19]), .Co(CTMP[20]) );
  FA_428 FAI_21 ( .A(A[20]), .B(B[20]), .Ci(CTMP[20]), .S(S[20]), .Co(CTMP[21]) );
  FA_427 FAI_22 ( .A(A[21]), .B(B[21]), .Ci(CTMP[21]), .S(S[21]), .Co(CTMP[22]) );
  FA_426 FAI_23 ( .A(A[22]), .B(B[22]), .Ci(CTMP[22]), .S(S[22]), .Co(CTMP[23]) );
  FA_425 FAI_24 ( .A(A[23]), .B(B[23]), .Ci(CTMP[23]), .S(S[23]), .Co(CTMP[24]) );
  FA_424 FAI_25 ( .A(A[24]), .B(B[24]), .Ci(CTMP[24]), .S(S[24]), .Co(CTMP[25]) );
  FA_423 FAI_26 ( .A(A[25]), .B(B[25]), .Ci(CTMP[25]), .S(S[25]), .Co(CTMP[26]) );
  FA_422 FAI_27 ( .A(A[26]), .B(B[26]), .Ci(CTMP[26]), .S(S[26]), .Co(CTMP[27]) );
  FA_421 FAI_28 ( .A(A[27]), .B(B[27]), .Ci(CTMP[27]), .S(S[27]), .Co(CTMP[28]) );
  FA_420 FAI_29 ( .A(A[28]), .B(B[28]), .Ci(CTMP[28]), .S(S[28]), .Co(CTMP[29]) );
  FA_419 FAI_30 ( .A(A[29]), .B(B[29]), .Ci(CTMP[29]), .S(S[29]), .Co(CTMP[30]) );
  FA_418 FAI_31 ( .A(A[30]), .B(B[30]), .Ci(CTMP[30]), .S(S[30]), .Co(CTMP[31]) );
  FA_417 FAI_32 ( .A(A[31]), .B(B[31]), .Ci(CTMP[31]), .S(S[31]), .Co(CTMP[32]) );
  FA_416 FAI_33 ( .A(A[32]), .B(B[32]), .Ci(CTMP[32]), .S(S[32]), .Co(CTMP[33]) );
  FA_415 FAI_34 ( .A(A[33]), .B(B[33]), .Ci(CTMP[33]), .S(S[33]), .Co(CTMP[34]) );
  FA_414 FAI_35 ( .A(A[34]), .B(B[34]), .Ci(CTMP[34]), .S(S[34]), .Co(CTMP[35]) );
  FA_413 FAI_36 ( .A(A[35]), .B(B[35]), .Ci(CTMP[35]), .S(S[35]), .Co(CTMP[36]) );
  FA_412 FAI_37 ( .A(A[36]), .B(B[36]), .Ci(CTMP[36]), .S(S[36]), .Co(CTMP[37]) );
  FA_411 FAI_38 ( .A(A[37]), .B(B[37]), .Ci(CTMP[37]), .S(S[37]), .Co(CTMP[38]) );
  FA_410 FAI_39 ( .A(A[38]), .B(B[38]), .Ci(CTMP[38]), .S(S[38]), .Co(CTMP[39]) );
  FA_409 FAI_40 ( .A(A[39]), .B(B[39]), .Ci(CTMP[39]), .S(S[39]), .Co(CTMP[40]) );
  FA_408 FAI_41 ( .A(A[40]), .B(B[40]), .Ci(CTMP[40]), .S(S[40]), .Co(CTMP[41]) );
  FA_407 FAI_42 ( .A(A[41]), .B(B[41]), .Ci(CTMP[41]), .S(S[41]), .Co(CTMP[42]) );
  FA_406 FAI_43 ( .A(A[42]), .B(B[42]), .Ci(CTMP[42]), .S(S[42]), .Co(CTMP[43]) );
  FA_405 FAI_44 ( .A(A[43]), .B(B[43]), .Ci(CTMP[43]), .S(S[43]), .Co(CTMP[44]) );
  FA_404 FAI_45 ( .A(A[44]), .B(B[44]), .Ci(CTMP[44]), .S(S[44]), .Co(CTMP[45]) );
  FA_403 FAI_46 ( .A(A[45]), .B(B[45]), .Ci(CTMP[45]), .S(S[45]), .Co(CTMP[46]) );
  FA_402 FAI_47 ( .A(A[46]), .B(B[46]), .Ci(CTMP[46]), .S(S[46]), .Co(CTMP[47]) );
  FA_401 FAI_48 ( .A(A[47]), .B(B[47]), .Ci(CTMP[47]), .S(S[47]), .Co(CTMP[48]) );
  FA_400 FAI_49 ( .A(A[48]), .B(B[48]), .Ci(CTMP[48]), .S(S[48]), .Co(CTMP[49]) );
  FA_399 FAI_50 ( .A(A[49]), .B(B[49]), .Ci(CTMP[49]), .S(S[49]), .Co(CTMP[50]) );
  FA_398 FAI_51 ( .A(A[50]), .B(B[50]), .Ci(CTMP[50]), .S(S[50]), .Co(CTMP[51]) );
  FA_397 FAI_52 ( .A(A[51]), .B(B[51]), .Ci(CTMP[51]), .S(S[51]), .Co(CTMP[52]) );
  FA_396 FAI_53 ( .A(A[52]), .B(B[52]), .Ci(CTMP[52]), .S(S[52]), .Co(CTMP[53]) );
  FA_395 FAI_54 ( .A(A[53]), .B(B[53]), .Ci(CTMP[53]), .S(S[53]), .Co(CTMP[54]) );
  FA_394 FAI_55 ( .A(A[54]), .B(B[54]), .Ci(CTMP[54]), .S(S[54]), .Co(CTMP[55]) );
  FA_393 FAI_56 ( .A(A[55]), .B(B[55]), .Ci(CTMP[55]), .S(S[55]), .Co(CTMP[56]) );
  FA_392 FAI_57 ( .A(A[56]), .B(B[56]), .Ci(CTMP[56]), .S(S[56]), .Co(CTMP[57]) );
  FA_391 FAI_58 ( .A(A[57]), .B(B[57]), .Ci(CTMP[57]), .S(S[57]), .Co(CTMP[58]) );
  FA_390 FAI_59 ( .A(A[58]), .B(B[58]), .Ci(CTMP[58]), .S(S[58]), .Co(CTMP[59]) );
  FA_389 FAI_60 ( .A(A[59]), .B(B[59]), .Ci(CTMP[59]), .S(S[59]), .Co(CTMP[60]) );
  FA_388 FAI_61 ( .A(A[60]), .B(B[60]), .Ci(CTMP[60]), .S(S[60]), .Co(CTMP[61]) );
  FA_387 FAI_62 ( .A(A[61]), .B(B[61]), .Ci(CTMP[61]), .S(S[61]), .Co(CTMP[62]) );
  FA_386 FAI_63 ( .A(A[62]), .B(B[62]), .Ci(CTMP[62]), .S(S[62]), .Co(CTMP[63]) );
  FA_385 FAI_64 ( .A(A[63]), .B(B[63]), .Ci(CTMP[63]), .S(S[63]), .Co(Co) );
endmodule


module booth_mul_row_N64_RADIX3_7 ( prevA, prevSum, encoderIn, nextA, nextSum
 );
  input [63:0] prevA;
  input [63:0] prevSum;
  input [2:0] encoderIn;
  output [63:0] nextA;
  output [63:0] nextSum;
  wire   n4, n5;
  wire   [2:0] encoder_to_mux;
  wire   [63:0] plus2A_s;
  wire   [63:0] minus2A_s;
  wire   [63:0] minus4A_s;
  tri   [63:0] mux_to_adder;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign nextA[51] = n4;
  assign nextA[50] = n5;
  assign nextA[0] = 1'b0;

  encoder_N64_RADIX3_7 encoder_1 ( .X(encoderIn), .Z(encoder_to_mux) );
  ShiftnCompl_N64_7 ShiftnCompl_1 ( .plusA(prevA), .plus2A_out({plus2A_s[63:1], 
        SYNOPSYS_UNCONNECTED__0}), .minus2A_out(minus2A_s), .plus4A_out({
        nextA[63:52], n4, n5, nextA[49:1], SYNOPSYS_UNCONNECTED__1}), 
        .minus4A_out(minus4A_s) );
  MUX_GENERIC_N64_RADIX3_7 mux_1 ( .plusA({plus2A_s[63:1], 1'b0}), .minusA(
        minus2A_s), .plus2A({nextA[63:52], n4, n5, nextA[49:1], 1'b0}), 
        .minus2A(minus4A_s), .SEL(encoder_to_mux), .Y(mux_to_adder) );
  RCA_N64_7 rca_1 ( .A(mux_to_adder), .B(prevSum), .Ci(1'b0), .S(nextSum) );
endmodule


module encoder_N64_RADIX3_6 ( X, Z );
  input [2:0] X;
  output [2:0] Z;
  wire   n5, n7, n8;

  OAI22_X1 U1 ( .A1(n8), .A2(n5), .B1(X[2]), .B2(n7), .ZN(Z[1]) );
  INV_X1 U2 ( .A(X[2]), .ZN(n5) );
  AOI21_X1 U3 ( .B1(n8), .B2(n7), .A(X[2]), .ZN(Z[0]) );
  OAI21_X1 U4 ( .B1(X[1]), .B2(X[0]), .A(n7), .ZN(n8) );
  AND3_X1 U5 ( .A1(X[2]), .A2(n7), .A3(n8), .ZN(Z[2]) );
  NAND2_X1 U6 ( .A1(X[1]), .A2(X[0]), .ZN(n7) );
endmodule


module shifter_N64_12 ( \input , shiftLeftOnePos );
  input [63:0] \input ;
  output [63:0] shiftLeftOnePos;
  wire   \input[62] , \input[61] , \input[60] , \input[59] , \input[58] ,
         \input[57] , \input[56] , \input[55] , \input[54] , \input[53] ,
         \input[52] , \input[51] , \input[50] , \input[49] , \input[48] ,
         \input[47] , \input[46] , \input[45] , \input[44] , \input[43] ,
         \input[42] , \input[41] , \input[40] , \input[39] , \input[38] ,
         \input[37] , \input[36] , \input[35] , \input[34] , \input[33] ,
         \input[32] , \input[31] , \input[30] , \input[29] , \input[28] ,
         \input[27] , \input[26] , \input[25] , \input[24] , \input[23] ,
         \input[22] , \input[21] , \input[20] , \input[19] , \input[18] ,
         \input[17] , \input[16] , \input[15] , \input[14] , \input[13] ,
         \input[12] , \input[11] , \input[10] , \input[9] , \input[8] ,
         \input[7] , \input[6] , \input[5] , \input[4] , \input[3] ,
         \input[2] , \input[1] , \input[0] ;
  assign shiftLeftOnePos[0] = 1'b0;
  assign shiftLeftOnePos[63] = \input[62] ;
  assign \input[62]  = \input  [62];
  assign shiftLeftOnePos[62] = \input[61] ;
  assign \input[61]  = \input  [61];
  assign shiftLeftOnePos[61] = \input[60] ;
  assign \input[60]  = \input  [60];
  assign shiftLeftOnePos[60] = \input[59] ;
  assign \input[59]  = \input  [59];
  assign shiftLeftOnePos[59] = \input[58] ;
  assign \input[58]  = \input  [58];
  assign shiftLeftOnePos[58] = \input[57] ;
  assign \input[57]  = \input  [57];
  assign shiftLeftOnePos[57] = \input[56] ;
  assign \input[56]  = \input  [56];
  assign shiftLeftOnePos[56] = \input[55] ;
  assign \input[55]  = \input  [55];
  assign shiftLeftOnePos[55] = \input[54] ;
  assign \input[54]  = \input  [54];
  assign shiftLeftOnePos[54] = \input[53] ;
  assign \input[53]  = \input  [53];
  assign shiftLeftOnePos[53] = \input[52] ;
  assign \input[52]  = \input  [52];
  assign shiftLeftOnePos[52] = \input[51] ;
  assign \input[51]  = \input  [51];
  assign shiftLeftOnePos[51] = \input[50] ;
  assign \input[50]  = \input  [50];
  assign shiftLeftOnePos[50] = \input[49] ;
  assign \input[49]  = \input  [49];
  assign shiftLeftOnePos[49] = \input[48] ;
  assign \input[48]  = \input  [48];
  assign shiftLeftOnePos[48] = \input[47] ;
  assign \input[47]  = \input  [47];
  assign shiftLeftOnePos[47] = \input[46] ;
  assign \input[46]  = \input  [46];
  assign shiftLeftOnePos[46] = \input[45] ;
  assign \input[45]  = \input  [45];
  assign shiftLeftOnePos[45] = \input[44] ;
  assign \input[44]  = \input  [44];
  assign shiftLeftOnePos[44] = \input[43] ;
  assign \input[43]  = \input  [43];
  assign shiftLeftOnePos[43] = \input[42] ;
  assign \input[42]  = \input  [42];
  assign shiftLeftOnePos[42] = \input[41] ;
  assign \input[41]  = \input  [41];
  assign shiftLeftOnePos[41] = \input[40] ;
  assign \input[40]  = \input  [40];
  assign shiftLeftOnePos[40] = \input[39] ;
  assign \input[39]  = \input  [39];
  assign shiftLeftOnePos[39] = \input[38] ;
  assign \input[38]  = \input  [38];
  assign shiftLeftOnePos[38] = \input[37] ;
  assign \input[37]  = \input  [37];
  assign shiftLeftOnePos[37] = \input[36] ;
  assign \input[36]  = \input  [36];
  assign shiftLeftOnePos[36] = \input[35] ;
  assign \input[35]  = \input  [35];
  assign shiftLeftOnePos[35] = \input[34] ;
  assign \input[34]  = \input  [34];
  assign shiftLeftOnePos[34] = \input[33] ;
  assign \input[33]  = \input  [33];
  assign shiftLeftOnePos[33] = \input[32] ;
  assign \input[32]  = \input  [32];
  assign shiftLeftOnePos[32] = \input[31] ;
  assign \input[31]  = \input  [31];
  assign shiftLeftOnePos[31] = \input[30] ;
  assign \input[30]  = \input  [30];
  assign shiftLeftOnePos[30] = \input[29] ;
  assign \input[29]  = \input  [29];
  assign shiftLeftOnePos[29] = \input[28] ;
  assign \input[28]  = \input  [28];
  assign shiftLeftOnePos[28] = \input[27] ;
  assign \input[27]  = \input  [27];
  assign shiftLeftOnePos[27] = \input[26] ;
  assign \input[26]  = \input  [26];
  assign shiftLeftOnePos[26] = \input[25] ;
  assign \input[25]  = \input  [25];
  assign shiftLeftOnePos[25] = \input[24] ;
  assign \input[24]  = \input  [24];
  assign shiftLeftOnePos[24] = \input[23] ;
  assign \input[23]  = \input  [23];
  assign shiftLeftOnePos[23] = \input[22] ;
  assign \input[22]  = \input  [22];
  assign shiftLeftOnePos[22] = \input[21] ;
  assign \input[21]  = \input  [21];
  assign shiftLeftOnePos[21] = \input[20] ;
  assign \input[20]  = \input  [20];
  assign shiftLeftOnePos[20] = \input[19] ;
  assign \input[19]  = \input  [19];
  assign shiftLeftOnePos[19] = \input[18] ;
  assign \input[18]  = \input  [18];
  assign shiftLeftOnePos[18] = \input[17] ;
  assign \input[17]  = \input  [17];
  assign shiftLeftOnePos[17] = \input[16] ;
  assign \input[16]  = \input  [16];
  assign shiftLeftOnePos[16] = \input[15] ;
  assign \input[15]  = \input  [15];
  assign shiftLeftOnePos[15] = \input[14] ;
  assign \input[14]  = \input  [14];
  assign shiftLeftOnePos[14] = \input[13] ;
  assign \input[13]  = \input  [13];
  assign shiftLeftOnePos[13] = \input[12] ;
  assign \input[12]  = \input  [12];
  assign shiftLeftOnePos[12] = \input[11] ;
  assign \input[11]  = \input  [11];
  assign shiftLeftOnePos[11] = \input[10] ;
  assign \input[10]  = \input  [10];
  assign shiftLeftOnePos[10] = \input[9] ;
  assign \input[9]  = \input  [9];
  assign shiftLeftOnePos[9] = \input[8] ;
  assign \input[8]  = \input  [8];
  assign shiftLeftOnePos[8] = \input[7] ;
  assign \input[7]  = \input  [7];
  assign shiftLeftOnePos[7] = \input[6] ;
  assign \input[6]  = \input  [6];
  assign shiftLeftOnePos[6] = \input[5] ;
  assign \input[5]  = \input  [5];
  assign shiftLeftOnePos[5] = \input[4] ;
  assign \input[4]  = \input  [4];
  assign shiftLeftOnePos[4] = \input[3] ;
  assign \input[3]  = \input  [3];
  assign shiftLeftOnePos[3] = \input[2] ;
  assign \input[2]  = \input  [2];
  assign shiftLeftOnePos[2] = \input[1] ;
  assign \input[1]  = \input  [1];
  assign shiftLeftOnePos[1] = \input[0] ;
  assign \input[0]  = \input  [0];

endmodule


module shifter_N64_11 ( \input , shiftLeftOnePos );
  input [63:0] \input ;
  output [63:0] shiftLeftOnePos;
  wire   \input[62] , \input[61] , \input[60] , \input[59] , \input[58] ,
         \input[57] , \input[56] , \input[55] , \input[54] , \input[53] ,
         \input[52] , \input[51] , \input[50] , \input[49] , \input[48] ,
         \input[47] , \input[46] , \input[45] , \input[44] , \input[43] ,
         \input[42] , \input[41] , \input[40] , \input[39] , \input[38] ,
         \input[37] , \input[36] , \input[35] , \input[34] , \input[33] ,
         \input[32] , \input[31] , \input[30] , \input[29] , \input[28] ,
         \input[27] , \input[26] , \input[25] , \input[24] , \input[23] ,
         \input[22] , \input[21] , \input[20] , \input[19] , \input[18] ,
         \input[17] , \input[16] , \input[15] , \input[14] , \input[13] ,
         \input[12] , \input[11] , \input[10] , \input[9] , \input[8] ,
         \input[7] , \input[6] , \input[5] , \input[4] , \input[3] ,
         \input[2] , \input[1] , \input[0] ;
  assign shiftLeftOnePos[0] = 1'b0;
  assign shiftLeftOnePos[63] = \input[62] ;
  assign \input[62]  = \input  [62];
  assign shiftLeftOnePos[62] = \input[61] ;
  assign \input[61]  = \input  [61];
  assign shiftLeftOnePos[61] = \input[60] ;
  assign \input[60]  = \input  [60];
  assign shiftLeftOnePos[60] = \input[59] ;
  assign \input[59]  = \input  [59];
  assign shiftLeftOnePos[59] = \input[58] ;
  assign \input[58]  = \input  [58];
  assign shiftLeftOnePos[58] = \input[57] ;
  assign \input[57]  = \input  [57];
  assign shiftLeftOnePos[57] = \input[56] ;
  assign \input[56]  = \input  [56];
  assign shiftLeftOnePos[56] = \input[55] ;
  assign \input[55]  = \input  [55];
  assign shiftLeftOnePos[55] = \input[54] ;
  assign \input[54]  = \input  [54];
  assign shiftLeftOnePos[54] = \input[53] ;
  assign \input[53]  = \input  [53];
  assign shiftLeftOnePos[53] = \input[52] ;
  assign \input[52]  = \input  [52];
  assign shiftLeftOnePos[52] = \input[51] ;
  assign \input[51]  = \input  [51];
  assign shiftLeftOnePos[51] = \input[50] ;
  assign \input[50]  = \input  [50];
  assign shiftLeftOnePos[50] = \input[49] ;
  assign \input[49]  = \input  [49];
  assign shiftLeftOnePos[49] = \input[48] ;
  assign \input[48]  = \input  [48];
  assign shiftLeftOnePos[48] = \input[47] ;
  assign \input[47]  = \input  [47];
  assign shiftLeftOnePos[47] = \input[46] ;
  assign \input[46]  = \input  [46];
  assign shiftLeftOnePos[46] = \input[45] ;
  assign \input[45]  = \input  [45];
  assign shiftLeftOnePos[45] = \input[44] ;
  assign \input[44]  = \input  [44];
  assign shiftLeftOnePos[44] = \input[43] ;
  assign \input[43]  = \input  [43];
  assign shiftLeftOnePos[43] = \input[42] ;
  assign \input[42]  = \input  [42];
  assign shiftLeftOnePos[42] = \input[41] ;
  assign \input[41]  = \input  [41];
  assign shiftLeftOnePos[41] = \input[40] ;
  assign \input[40]  = \input  [40];
  assign shiftLeftOnePos[40] = \input[39] ;
  assign \input[39]  = \input  [39];
  assign shiftLeftOnePos[39] = \input[38] ;
  assign \input[38]  = \input  [38];
  assign shiftLeftOnePos[38] = \input[37] ;
  assign \input[37]  = \input  [37];
  assign shiftLeftOnePos[37] = \input[36] ;
  assign \input[36]  = \input  [36];
  assign shiftLeftOnePos[36] = \input[35] ;
  assign \input[35]  = \input  [35];
  assign shiftLeftOnePos[35] = \input[34] ;
  assign \input[34]  = \input  [34];
  assign shiftLeftOnePos[34] = \input[33] ;
  assign \input[33]  = \input  [33];
  assign shiftLeftOnePos[33] = \input[32] ;
  assign \input[32]  = \input  [32];
  assign shiftLeftOnePos[32] = \input[31] ;
  assign \input[31]  = \input  [31];
  assign shiftLeftOnePos[31] = \input[30] ;
  assign \input[30]  = \input  [30];
  assign shiftLeftOnePos[30] = \input[29] ;
  assign \input[29]  = \input  [29];
  assign shiftLeftOnePos[29] = \input[28] ;
  assign \input[28]  = \input  [28];
  assign shiftLeftOnePos[28] = \input[27] ;
  assign \input[27]  = \input  [27];
  assign shiftLeftOnePos[27] = \input[26] ;
  assign \input[26]  = \input  [26];
  assign shiftLeftOnePos[26] = \input[25] ;
  assign \input[25]  = \input  [25];
  assign shiftLeftOnePos[25] = \input[24] ;
  assign \input[24]  = \input  [24];
  assign shiftLeftOnePos[24] = \input[23] ;
  assign \input[23]  = \input  [23];
  assign shiftLeftOnePos[23] = \input[22] ;
  assign \input[22]  = \input  [22];
  assign shiftLeftOnePos[22] = \input[21] ;
  assign \input[21]  = \input  [21];
  assign shiftLeftOnePos[21] = \input[20] ;
  assign \input[20]  = \input  [20];
  assign shiftLeftOnePos[20] = \input[19] ;
  assign \input[19]  = \input  [19];
  assign shiftLeftOnePos[19] = \input[18] ;
  assign \input[18]  = \input  [18];
  assign shiftLeftOnePos[18] = \input[17] ;
  assign \input[17]  = \input  [17];
  assign shiftLeftOnePos[17] = \input[16] ;
  assign \input[16]  = \input  [16];
  assign shiftLeftOnePos[16] = \input[15] ;
  assign \input[15]  = \input  [15];
  assign shiftLeftOnePos[15] = \input[14] ;
  assign \input[14]  = \input  [14];
  assign shiftLeftOnePos[14] = \input[13] ;
  assign \input[13]  = \input  [13];
  assign shiftLeftOnePos[13] = \input[12] ;
  assign \input[12]  = \input  [12];
  assign shiftLeftOnePos[12] = \input[11] ;
  assign \input[11]  = \input  [11];
  assign shiftLeftOnePos[11] = \input[10] ;
  assign \input[10]  = \input  [10];
  assign shiftLeftOnePos[10] = \input[9] ;
  assign \input[9]  = \input  [9];
  assign shiftLeftOnePos[9] = \input[8] ;
  assign \input[8]  = \input  [8];
  assign shiftLeftOnePos[8] = \input[7] ;
  assign \input[7]  = \input  [7];
  assign shiftLeftOnePos[7] = \input[6] ;
  assign \input[6]  = \input  [6];
  assign shiftLeftOnePos[6] = \input[5] ;
  assign \input[5]  = \input  [5];
  assign shiftLeftOnePos[5] = \input[4] ;
  assign \input[4]  = \input  [4];
  assign shiftLeftOnePos[4] = \input[3] ;
  assign \input[3]  = \input  [3];
  assign shiftLeftOnePos[3] = \input[2] ;
  assign \input[2]  = \input  [2];
  assign shiftLeftOnePos[2] = \input[1] ;
  assign \input[1]  = \input  [1];
  assign shiftLeftOnePos[1] = \input[0] ;
  assign \input[0]  = \input  [0];

endmodule


module complementer_N64_12_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n190, n191, n192, n193, n194, n196, n197, n198, n199, n200,
         n202, n203, n204, n206, n207, n208, n210, n211, n212, n213, n214,
         n216, n217, n218, n220, n221, n222, n224, n225, n226, n228, n229,
         n230, n232, n233, n234, n235, n237, n238, n239, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n189, n195, n201,
         n205, n209, n215, n219, n223, n227, n231, n236, n240;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U81 ( .A(n190), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U82 ( .A(n192), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U83 ( .A(n193), .B(B[6]), .Z(DIFF[6]) );
  XOR2_X1 U85 ( .A(n196), .B(B[62]), .Z(DIFF[62]) );
  XOR2_X1 U86 ( .A(n194), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U87 ( .A(n198), .B(B[59]), .Z(DIFF[59]) );
  XOR2_X1 U89 ( .A(n200), .B(B[57]), .Z(DIFF[57]) );
  XOR2_X1 U90 ( .A(n202), .B(B[55]), .Z(DIFF[55]) );
  XOR2_X1 U92 ( .A(n204), .B(B[53]), .Z(DIFF[53]) );
  XOR2_X1 U93 ( .A(n206), .B(B[51]), .Z(DIFF[51]) );
  XOR2_X1 U95 ( .A(n208), .B(B[49]), .Z(DIFF[49]) );
  XOR2_X1 U96 ( .A(n212), .B(B[47]), .Z(DIFF[47]) );
  XOR2_X1 U98 ( .A(n214), .B(B[45]), .Z(DIFF[45]) );
  XOR2_X1 U99 ( .A(n216), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U101 ( .A(n218), .B(B[41]), .Z(DIFF[41]) );
  XOR2_X1 U102 ( .A(n211), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U103 ( .A(n220), .B(B[39]), .Z(DIFF[39]) );
  XOR2_X1 U105 ( .A(n222), .B(B[37]), .Z(DIFF[37]) );
  XOR2_X1 U106 ( .A(n224), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U108 ( .A(n226), .B(B[33]), .Z(DIFF[33]) );
  XOR2_X1 U109 ( .A(n228), .B(B[31]), .Z(DIFF[31]) );
  XOR2_X1 U111 ( .A(n230), .B(B[29]), .Z(DIFF[29]) );
  XOR2_X1 U112 ( .A(n233), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U114 ( .A(n235), .B(B[25]), .Z(DIFF[25]) );
  XOR2_X1 U115 ( .A(n237), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U117 ( .A(n239), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U118 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U119 ( .A(n241), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U120 ( .A(n244), .B(B[18]), .Z(DIFF[18]) );
  XOR2_X1 U121 ( .A(n243), .B(B[17]), .Z(DIFF[17]) );
  XOR2_X1 U122 ( .A(n245), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U123 ( .A(n248), .B(B[14]), .Z(DIFF[14]) );
  XOR2_X1 U124 ( .A(n247), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U125 ( .A(n249), .B(B[11]), .Z(DIFF[11]) );
  XOR2_X1 U126 ( .A(n251), .B(B[10]), .Z(DIFF[10]) );
  XOR2_X1 U1 ( .A(n197), .B(n240), .Z(DIFF[61]) );
  NAND2_X1 U2 ( .A1(n197), .A2(n240), .ZN(n196) );
  NOR3_X1 U3 ( .A1(B[59]), .A2(B[60]), .A3(n198), .ZN(n197) );
  XNOR2_X1 U4 ( .A(n189), .B(B[63]), .ZN(DIFF[63]) );
  NOR2_X1 U5 ( .A1(n196), .A2(B[62]), .ZN(n189) );
  XNOR2_X1 U6 ( .A(B[56]), .B(n203), .ZN(DIFF[56]) );
  NOR2_X1 U7 ( .A1(B[55]), .A2(n202), .ZN(n203) );
  XNOR2_X1 U8 ( .A(B[60]), .B(n199), .ZN(DIFF[60]) );
  NOR2_X1 U9 ( .A1(B[59]), .A2(n198), .ZN(n199) );
  OR3_X1 U10 ( .A1(B[57]), .A2(B[58]), .A3(n200), .ZN(n198) );
  OR3_X1 U11 ( .A1(B[53]), .A2(B[54]), .A3(n204), .ZN(n202) );
  OR3_X1 U12 ( .A1(B[55]), .A2(B[56]), .A3(n202), .ZN(n200) );
  XNOR2_X1 U13 ( .A(n195), .B(B[58]), .ZN(DIFF[58]) );
  NOR2_X1 U14 ( .A1(n200), .A2(B[57]), .ZN(n195) );
  XNOR2_X1 U15 ( .A(n201), .B(B[54]), .ZN(DIFF[54]) );
  NOR2_X1 U16 ( .A1(n204), .A2(B[53]), .ZN(n201) );
  XNOR2_X1 U17 ( .A(B[52]), .B(n207), .ZN(DIFF[52]) );
  NOR2_X1 U18 ( .A1(B[51]), .A2(n206), .ZN(n207) );
  OR3_X1 U19 ( .A1(B[51]), .A2(B[52]), .A3(n206), .ZN(n204) );
  XNOR2_X1 U20 ( .A(n205), .B(B[30]), .ZN(DIFF[30]) );
  NOR2_X1 U21 ( .A1(n230), .A2(B[29]), .ZN(n205) );
  XNOR2_X1 U22 ( .A(B[44]), .B(n217), .ZN(DIFF[44]) );
  NOR2_X1 U23 ( .A1(B[43]), .A2(n216), .ZN(n217) );
  XNOR2_X1 U24 ( .A(B[40]), .B(n221), .ZN(DIFF[40]) );
  NOR2_X1 U25 ( .A1(B[39]), .A2(n220), .ZN(n221) );
  XNOR2_X1 U26 ( .A(B[36]), .B(n225), .ZN(DIFF[36]) );
  NOR2_X1 U27 ( .A1(B[35]), .A2(n224), .ZN(n225) );
  XNOR2_X1 U28 ( .A(B[32]), .B(n229), .ZN(DIFF[32]) );
  NOR2_X1 U29 ( .A1(B[31]), .A2(n228), .ZN(n229) );
  XNOR2_X1 U30 ( .A(B[28]), .B(n234), .ZN(DIFF[28]) );
  NOR2_X1 U31 ( .A1(B[27]), .A2(n233), .ZN(n234) );
  OR3_X1 U32 ( .A1(B[29]), .A2(B[30]), .A3(n230), .ZN(n228) );
  OR3_X1 U33 ( .A1(B[33]), .A2(B[34]), .A3(n226), .ZN(n224) );
  OR3_X1 U34 ( .A1(B[37]), .A2(B[38]), .A3(n222), .ZN(n220) );
  OR3_X1 U35 ( .A1(B[41]), .A2(B[42]), .A3(n218), .ZN(n216) );
  OR3_X1 U36 ( .A1(B[27]), .A2(B[28]), .A3(n233), .ZN(n230) );
  OR3_X1 U37 ( .A1(B[31]), .A2(B[32]), .A3(n228), .ZN(n226) );
  OR3_X1 U38 ( .A1(B[35]), .A2(B[36]), .A3(n224), .ZN(n222) );
  OR3_X1 U39 ( .A1(B[39]), .A2(B[40]), .A3(n220), .ZN(n218) );
  XNOR2_X1 U40 ( .A(n209), .B(B[42]), .ZN(DIFF[42]) );
  NOR2_X1 U41 ( .A1(n218), .A2(B[41]), .ZN(n209) );
  XNOR2_X1 U42 ( .A(n215), .B(B[38]), .ZN(DIFF[38]) );
  NOR2_X1 U43 ( .A1(n222), .A2(B[37]), .ZN(n215) );
  XNOR2_X1 U44 ( .A(n219), .B(B[34]), .ZN(DIFF[34]) );
  NOR2_X1 U45 ( .A1(n226), .A2(B[33]), .ZN(n219) );
  XNOR2_X1 U46 ( .A(n223), .B(B[46]), .ZN(DIFF[46]) );
  NOR2_X1 U47 ( .A1(n214), .A2(B[45]), .ZN(n223) );
  XNOR2_X1 U48 ( .A(B[48]), .B(n213), .ZN(DIFF[48]) );
  NOR2_X1 U49 ( .A1(B[47]), .A2(n212), .ZN(n213) );
  OR3_X1 U50 ( .A1(B[45]), .A2(B[46]), .A3(n214), .ZN(n212) );
  OR3_X1 U51 ( .A1(B[49]), .A2(B[50]), .A3(n208), .ZN(n206) );
  OR3_X1 U52 ( .A1(B[43]), .A2(B[44]), .A3(n216), .ZN(n214) );
  OR3_X1 U53 ( .A1(B[47]), .A2(B[48]), .A3(n212), .ZN(n208) );
  XNOR2_X1 U54 ( .A(n227), .B(B[50]), .ZN(DIFF[50]) );
  NOR2_X1 U55 ( .A1(n208), .A2(B[49]), .ZN(n227) );
  OR3_X1 U56 ( .A1(B[25]), .A2(B[26]), .A3(n235), .ZN(n233) );
  XNOR2_X1 U57 ( .A(n231), .B(B[26]), .ZN(DIFF[26]) );
  NOR2_X1 U58 ( .A1(n235), .A2(B[25]), .ZN(n231) );
  XNOR2_X1 U59 ( .A(B[24]), .B(n238), .ZN(DIFF[24]) );
  NOR2_X1 U60 ( .A1(B[23]), .A2(n237), .ZN(n238) );
  OR3_X1 U61 ( .A1(B[23]), .A2(B[24]), .A3(n237), .ZN(n235) );
  XNOR2_X1 U62 ( .A(n236), .B(B[22]), .ZN(DIFF[22]) );
  NOR2_X1 U63 ( .A1(n239), .A2(B[21]), .ZN(n236) );
  OR3_X1 U64 ( .A1(B[21]), .A2(B[22]), .A3(n239), .ZN(n237) );
  OR3_X1 U65 ( .A1(B[19]), .A2(B[20]), .A3(n241), .ZN(n239) );
  XNOR2_X1 U66 ( .A(B[20]), .B(n242), .ZN(DIFF[20]) );
  NOR2_X1 U67 ( .A1(B[19]), .A2(n241), .ZN(n242) );
  NOR2_X1 U68 ( .A1(B[15]), .A2(n245), .ZN(n246) );
  NOR2_X1 U69 ( .A1(B[11]), .A2(n249), .ZN(n250) );
  NOR2_X1 U70 ( .A1(B[7]), .A2(n192), .ZN(n191) );
  NOR2_X1 U71 ( .A1(B[3]), .A2(n211), .ZN(n210) );
  OR3_X1 U72 ( .A1(B[17]), .A2(B[18]), .A3(n243), .ZN(n241) );
  OR3_X1 U73 ( .A1(B[13]), .A2(B[14]), .A3(n247), .ZN(n245) );
  OR3_X1 U74 ( .A1(B[10]), .A2(B[9]), .A3(n190), .ZN(n249) );
  OR3_X1 U75 ( .A1(B[5]), .A2(B[6]), .A3(n194), .ZN(n192) );
  OR3_X1 U76 ( .A1(B[15]), .A2(B[16]), .A3(n245), .ZN(n243) );
  OR3_X1 U77 ( .A1(B[11]), .A2(B[12]), .A3(n249), .ZN(n247) );
  OR3_X1 U78 ( .A1(B[7]), .A2(B[8]), .A3(n192), .ZN(n190) );
  OR3_X1 U79 ( .A1(B[3]), .A2(B[4]), .A3(n211), .ZN(n194) );
  XNOR2_X1 U80 ( .A(B[16]), .B(n246), .ZN(DIFF[16]) );
  XNOR2_X1 U84 ( .A(B[12]), .B(n250), .ZN(DIFF[12]) );
  XNOR2_X1 U88 ( .A(B[8]), .B(n191), .ZN(DIFF[8]) );
  XNOR2_X1 U91 ( .A(B[4]), .B(n210), .ZN(DIFF[4]) );
  XNOR2_X1 U94 ( .A(B[2]), .B(n232), .ZN(DIFF[2]) );
  OR2_X1 U97 ( .A1(n243), .A2(B[17]), .ZN(n244) );
  OR2_X1 U100 ( .A1(n247), .A2(B[13]), .ZN(n248) );
  OR2_X1 U104 ( .A1(n190), .A2(B[9]), .ZN(n251) );
  OR2_X1 U107 ( .A1(n194), .A2(B[5]), .ZN(n193) );
  OR3_X1 U110 ( .A1(B[1]), .A2(B[2]), .A3(\B[0] ), .ZN(n211) );
  NOR2_X1 U113 ( .A1(\B[0] ), .A2(B[1]), .ZN(n232) );
  INV_X1 U116 ( .A(B[61]), .ZN(n240) );
endmodule


module complementer_N64_12 ( \input , complement2 );
  input [63:0] \input ;
  output [63:0] complement2;


  complementer_N64_12_DW01_sub_0 sub_add_31_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(\input ), .CI(1'b0), .DIFF(complement2) );
endmodule


module complementer_N64_11_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n190, n191, n192, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n245,
         n246, n247, n249, n250, n189, n193, n244, n248, n251;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U81 ( .A(n190), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U82 ( .A(n192), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U84 ( .A(n195), .B(B[63]), .Z(DIFF[63]) );
  XOR2_X1 U85 ( .A(n196), .B(B[62]), .Z(DIFF[62]) );
  XOR2_X1 U86 ( .A(n194), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U87 ( .A(n198), .B(B[59]), .Z(DIFF[59]) );
  XOR2_X1 U88 ( .A(n201), .B(B[58]), .Z(DIFF[58]) );
  XOR2_X1 U89 ( .A(n200), .B(B[57]), .Z(DIFF[57]) );
  XOR2_X1 U90 ( .A(n202), .B(B[55]), .Z(DIFF[55]) );
  XOR2_X1 U91 ( .A(n205), .B(B[54]), .Z(DIFF[54]) );
  XOR2_X1 U92 ( .A(n204), .B(B[53]), .Z(DIFF[53]) );
  XOR2_X1 U93 ( .A(n206), .B(B[51]), .Z(DIFF[51]) );
  XOR2_X1 U94 ( .A(n209), .B(B[50]), .Z(DIFF[50]) );
  XOR2_X1 U95 ( .A(n208), .B(B[49]), .Z(DIFF[49]) );
  XOR2_X1 U96 ( .A(n212), .B(B[47]), .Z(DIFF[47]) );
  XOR2_X1 U97 ( .A(n215), .B(B[46]), .Z(DIFF[46]) );
  XOR2_X1 U98 ( .A(n214), .B(B[45]), .Z(DIFF[45]) );
  XOR2_X1 U99 ( .A(n216), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U100 ( .A(n219), .B(B[42]), .Z(DIFF[42]) );
  XOR2_X1 U101 ( .A(n218), .B(B[41]), .Z(DIFF[41]) );
  XOR2_X1 U102 ( .A(n211), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U103 ( .A(n220), .B(B[39]), .Z(DIFF[39]) );
  XOR2_X1 U104 ( .A(n223), .B(B[38]), .Z(DIFF[38]) );
  XOR2_X1 U105 ( .A(n222), .B(B[37]), .Z(DIFF[37]) );
  XOR2_X1 U106 ( .A(n224), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U107 ( .A(n227), .B(B[34]), .Z(DIFF[34]) );
  XOR2_X1 U108 ( .A(n226), .B(B[33]), .Z(DIFF[33]) );
  XOR2_X1 U109 ( .A(n228), .B(B[31]), .Z(DIFF[31]) );
  XOR2_X1 U110 ( .A(n231), .B(B[30]), .Z(DIFF[30]) );
  XOR2_X1 U111 ( .A(n230), .B(B[29]), .Z(DIFF[29]) );
  XOR2_X1 U112 ( .A(n233), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U113 ( .A(n236), .B(B[26]), .Z(DIFF[26]) );
  XOR2_X1 U114 ( .A(n235), .B(B[25]), .Z(DIFF[25]) );
  XOR2_X1 U115 ( .A(n237), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U116 ( .A(n240), .B(B[22]), .Z(DIFF[22]) );
  XOR2_X1 U117 ( .A(n239), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U118 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U119 ( .A(n241), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U121 ( .A(n243), .B(B[17]), .Z(DIFF[17]) );
  XOR2_X1 U122 ( .A(n245), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U124 ( .A(n247), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U125 ( .A(n249), .B(B[11]), .Z(DIFF[11]) );
  NOR2_X1 U1 ( .A1(B[59]), .A2(n198), .ZN(n199) );
  NAND2_X1 U2 ( .A1(n197), .A2(n251), .ZN(n196) );
  NOR3_X1 U3 ( .A1(B[59]), .A2(B[60]), .A3(n198), .ZN(n197) );
  NOR2_X1 U4 ( .A1(B[55]), .A2(n202), .ZN(n203) );
  OR3_X1 U5 ( .A1(B[57]), .A2(B[58]), .A3(n200), .ZN(n198) );
  OR3_X1 U6 ( .A1(B[53]), .A2(B[54]), .A3(n204), .ZN(n202) );
  OR3_X1 U7 ( .A1(B[55]), .A2(B[56]), .A3(n202), .ZN(n200) );
  OR2_X1 U8 ( .A1(n200), .A2(B[57]), .ZN(n201) );
  OR2_X1 U9 ( .A1(n204), .A2(B[53]), .ZN(n205) );
  OR2_X1 U10 ( .A1(n196), .A2(B[62]), .ZN(n195) );
  NOR2_X1 U11 ( .A1(B[51]), .A2(n206), .ZN(n207) );
  OR3_X1 U12 ( .A1(B[51]), .A2(B[52]), .A3(n206), .ZN(n204) );
  NOR2_X1 U13 ( .A1(B[39]), .A2(n220), .ZN(n221) );
  NOR2_X1 U14 ( .A1(B[35]), .A2(n224), .ZN(n225) );
  NOR2_X1 U15 ( .A1(B[31]), .A2(n228), .ZN(n229) );
  NOR2_X1 U16 ( .A1(B[27]), .A2(n233), .ZN(n234) );
  OR3_X1 U17 ( .A1(B[37]), .A2(B[38]), .A3(n222), .ZN(n220) );
  OR3_X1 U18 ( .A1(B[33]), .A2(B[34]), .A3(n226), .ZN(n224) );
  OR3_X1 U19 ( .A1(B[29]), .A2(B[30]), .A3(n230), .ZN(n228) );
  OR3_X1 U20 ( .A1(B[39]), .A2(B[40]), .A3(n220), .ZN(n218) );
  OR3_X1 U21 ( .A1(B[35]), .A2(B[36]), .A3(n224), .ZN(n222) );
  OR3_X1 U22 ( .A1(B[31]), .A2(B[32]), .A3(n228), .ZN(n226) );
  OR3_X1 U23 ( .A1(B[27]), .A2(B[28]), .A3(n233), .ZN(n230) );
  OR2_X1 U24 ( .A1(n222), .A2(B[37]), .ZN(n223) );
  OR2_X1 U25 ( .A1(n226), .A2(B[33]), .ZN(n227) );
  OR2_X1 U26 ( .A1(n230), .A2(B[29]), .ZN(n231) );
  NOR2_X1 U27 ( .A1(B[47]), .A2(n212), .ZN(n213) );
  NOR2_X1 U28 ( .A1(B[43]), .A2(n216), .ZN(n217) );
  OR3_X1 U29 ( .A1(B[49]), .A2(B[50]), .A3(n208), .ZN(n206) );
  OR3_X1 U30 ( .A1(B[45]), .A2(B[46]), .A3(n214), .ZN(n212) );
  OR3_X1 U31 ( .A1(B[41]), .A2(B[42]), .A3(n218), .ZN(n216) );
  OR3_X1 U32 ( .A1(B[47]), .A2(B[48]), .A3(n212), .ZN(n208) );
  OR3_X1 U33 ( .A1(B[43]), .A2(B[44]), .A3(n216), .ZN(n214) );
  OR2_X1 U34 ( .A1(n208), .A2(B[49]), .ZN(n209) );
  OR2_X1 U35 ( .A1(n214), .A2(B[45]), .ZN(n215) );
  OR2_X1 U36 ( .A1(n218), .A2(B[41]), .ZN(n219) );
  OR3_X1 U37 ( .A1(B[25]), .A2(B[26]), .A3(n235), .ZN(n233) );
  XNOR2_X1 U38 ( .A(B[44]), .B(n217), .ZN(DIFF[44]) );
  XNOR2_X1 U39 ( .A(B[40]), .B(n221), .ZN(DIFF[40]) );
  XNOR2_X1 U40 ( .A(B[36]), .B(n225), .ZN(DIFF[36]) );
  XNOR2_X1 U41 ( .A(B[32]), .B(n229), .ZN(DIFF[32]) );
  XNOR2_X1 U42 ( .A(B[28]), .B(n234), .ZN(DIFF[28]) );
  XNOR2_X1 U43 ( .A(B[24]), .B(n238), .ZN(DIFF[24]) );
  OR2_X1 U44 ( .A1(n235), .A2(B[25]), .ZN(n236) );
  XNOR2_X1 U45 ( .A(B[56]), .B(n203), .ZN(DIFF[56]) );
  XNOR2_X1 U46 ( .A(B[52]), .B(n207), .ZN(DIFF[52]) );
  XNOR2_X1 U47 ( .A(B[48]), .B(n213), .ZN(DIFF[48]) );
  XNOR2_X1 U48 ( .A(n197), .B(B[61]), .ZN(DIFF[61]) );
  XNOR2_X1 U49 ( .A(B[60]), .B(n199), .ZN(DIFF[60]) );
  NOR2_X1 U50 ( .A1(B[23]), .A2(n237), .ZN(n238) );
  OR3_X1 U51 ( .A1(B[23]), .A2(B[24]), .A3(n237), .ZN(n235) );
  OR3_X1 U52 ( .A1(B[21]), .A2(B[22]), .A3(n239), .ZN(n237) );
  OR2_X1 U53 ( .A1(n239), .A2(B[21]), .ZN(n240) );
  XNOR2_X1 U54 ( .A(B[20]), .B(n242), .ZN(DIFF[20]) );
  XNOR2_X1 U55 ( .A(n189), .B(B[18]), .ZN(DIFF[18]) );
  NOR2_X1 U56 ( .A1(n243), .A2(B[17]), .ZN(n189) );
  XNOR2_X1 U57 ( .A(n193), .B(B[14]), .ZN(DIFF[14]) );
  NOR2_X1 U58 ( .A1(n247), .A2(B[13]), .ZN(n193) );
  XNOR2_X1 U59 ( .A(n244), .B(B[10]), .ZN(DIFF[10]) );
  NOR2_X1 U60 ( .A1(n190), .A2(B[9]), .ZN(n244) );
  XNOR2_X1 U61 ( .A(n248), .B(B[6]), .ZN(DIFF[6]) );
  NOR2_X1 U62 ( .A1(n194), .A2(B[5]), .ZN(n248) );
  NOR2_X1 U63 ( .A1(B[19]), .A2(n241), .ZN(n242) );
  XNOR2_X1 U64 ( .A(B[16]), .B(n246), .ZN(DIFF[16]) );
  NOR2_X1 U65 ( .A1(B[15]), .A2(n245), .ZN(n246) );
  XNOR2_X1 U66 ( .A(B[12]), .B(n250), .ZN(DIFF[12]) );
  NOR2_X1 U67 ( .A1(B[11]), .A2(n249), .ZN(n250) );
  XNOR2_X1 U68 ( .A(B[8]), .B(n191), .ZN(DIFF[8]) );
  NOR2_X1 U69 ( .A1(B[7]), .A2(n192), .ZN(n191) );
  XNOR2_X1 U70 ( .A(B[2]), .B(n232), .ZN(DIFF[2]) );
  NOR2_X1 U71 ( .A1(\B[0] ), .A2(B[1]), .ZN(n232) );
  XNOR2_X1 U72 ( .A(B[4]), .B(n210), .ZN(DIFF[4]) );
  NOR2_X1 U73 ( .A1(B[3]), .A2(n211), .ZN(n210) );
  OR3_X1 U74 ( .A1(B[5]), .A2(B[6]), .A3(n194), .ZN(n192) );
  OR3_X1 U75 ( .A1(B[10]), .A2(B[9]), .A3(n190), .ZN(n249) );
  OR3_X1 U76 ( .A1(B[13]), .A2(B[14]), .A3(n247), .ZN(n245) );
  OR3_X1 U77 ( .A1(B[17]), .A2(B[18]), .A3(n243), .ZN(n241) );
  OR3_X1 U78 ( .A1(B[7]), .A2(B[8]), .A3(n192), .ZN(n190) );
  OR3_X1 U79 ( .A1(B[11]), .A2(B[12]), .A3(n249), .ZN(n247) );
  OR3_X1 U80 ( .A1(B[15]), .A2(B[16]), .A3(n245), .ZN(n243) );
  OR3_X1 U83 ( .A1(B[19]), .A2(B[20]), .A3(n241), .ZN(n239) );
  OR3_X1 U120 ( .A1(B[3]), .A2(B[4]), .A3(n211), .ZN(n194) );
  OR3_X1 U123 ( .A1(B[1]), .A2(B[2]), .A3(\B[0] ), .ZN(n211) );
  INV_X1 U126 ( .A(B[61]), .ZN(n251) );
endmodule


module complementer_N64_11 ( \input , complement2 );
  input [63:0] \input ;
  output [63:0] complement2;


  complementer_N64_11_DW01_sub_0 sub_add_31_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(\input ), .CI(1'b0), .DIFF(complement2) );
endmodule


module ShiftnCompl_N64_6 ( plusA, plus2A_out, minus2A_out, plus4A_out, 
        minus4A_out );
  input [63:0] plusA;
  output [63:0] plus2A_out;
  output [63:0] minus2A_out;
  output [63:0] plus4A_out;
  output [63:0] minus4A_out;
  wire   n7, n8, n9, n10, n11, n12;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign plus2A_out[0] = 1'b0;
  assign plus4A_out[0] = 1'b0;

  shifter_N64_12 shifter_1 ( .\input (plusA), .shiftLeftOnePos({
        plus2A_out[63:59], n7, plus2A_out[57:54], n8, plus2A_out[52:1], 
        SYNOPSYS_UNCONNECTED__0}) );
  shifter_N64_11 shifter_2 ( .\input ({plus2A_out[63:1], 1'b0}), 
        .shiftLeftOnePos({plus4A_out[63:59], n9, plus4A_out[57:54], n10, n11, 
        n12, plus4A_out[50:1], SYNOPSYS_UNCONNECTED__1}) );
  complementer_N64_12 complementer_1 ( .\input ({plus2A_out[63:1], 1'b0}), 
        .complement2(minus2A_out) );
  complementer_N64_11 complementer_2 ( .\input ({plus4A_out[63:1], 1'b0}), 
        .complement2(minus4A_out) );
  BUF_X1 U3 ( .A(n12), .Z(plus4A_out[51]) );
  BUF_X1 U4 ( .A(n8), .Z(plus2A_out[53]) );
  BUF_X1 U5 ( .A(n10), .Z(plus4A_out[53]) );
  BUF_X1 U6 ( .A(n11), .Z(plus4A_out[52]) );
  BUF_X1 U7 ( .A(n9), .Z(plus4A_out[58]) );
  BUF_X1 U8 ( .A(n7), .Z(plus2A_out[58]) );
endmodule


module MUX_GENERIC_N64_RADIX3_6 ( plusA, minusA, plus2A, minus2A, SEL, Y );
  input [63:0] plusA;
  input [63:0] minusA;
  input [63:0] plus2A;
  input [63:0] minus2A;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502;
  tri   [63:0] Y;

  TBUF_X1 \Y_tri[55]  ( .A(n446), .EN(n301), .Z(Y[55]) );
  TBUF_X1 \Y_tri[56]  ( .A(n445), .EN(n301), .Z(Y[56]) );
  TBUF_X1 \Y_tri[57]  ( .A(n444), .EN(n301), .Z(Y[57]) );
  TBUF_X1 \Y_tri[58]  ( .A(n443), .EN(n301), .Z(Y[58]) );
  TBUF_X1 \Y_tri[59]  ( .A(n442), .EN(n301), .Z(Y[59]) );
  TBUF_X1 \Y_tri[60]  ( .A(n441), .EN(n301), .Z(Y[60]) );
  TBUF_X1 \Y_tri[61]  ( .A(n440), .EN(n301), .Z(Y[61]) );
  TBUF_X1 \Y_tri[62]  ( .A(n439), .EN(n301), .Z(Y[62]) );
  TBUF_X1 \Y_tri[63]  ( .A(n438), .EN(n301), .Z(Y[63]) );
  TBUF_X1 \Y_tri[45]  ( .A(n456), .EN(n300), .Z(Y[45]) );
  TBUF_X1 \Y_tri[46]  ( .A(n455), .EN(n300), .Z(Y[46]) );
  TBUF_X1 \Y_tri[47]  ( .A(n454), .EN(n300), .Z(Y[47]) );
  TBUF_X1 \Y_tri[48]  ( .A(n453), .EN(n300), .Z(Y[48]) );
  TBUF_X1 \Y_tri[49]  ( .A(n452), .EN(n300), .Z(Y[49]) );
  TBUF_X1 \Y_tri[50]  ( .A(n451), .EN(n300), .Z(Y[50]) );
  TBUF_X1 \Y_tri[51]  ( .A(n450), .EN(n300), .Z(Y[51]) );
  TBUF_X1 \Y_tri[52]  ( .A(n449), .EN(n300), .Z(Y[52]) );
  TBUF_X1 \Y_tri[53]  ( .A(n448), .EN(n300), .Z(Y[53]) );
  TBUF_X1 \Y_tri[54]  ( .A(n447), .EN(n300), .Z(Y[54]) );
  TBUF_X1 \Y_tri[17]  ( .A(n484), .EN(n297), .Z(Y[17]) );
  TBUF_X1 \Y_tri[18]  ( .A(n483), .EN(n297), .Z(Y[18]) );
  TBUF_X1 \Y_tri[19]  ( .A(n482), .EN(n297), .Z(Y[19]) );
  TBUF_X1 \Y_tri[20]  ( .A(n481), .EN(n297), .Z(Y[20]) );
  TBUF_X1 \Y_tri[21]  ( .A(n480), .EN(n297), .Z(Y[21]) );
  TBUF_X1 \Y_tri[22]  ( .A(n479), .EN(n298), .Z(Y[22]) );
  TBUF_X1 \Y_tri[23]  ( .A(n478), .EN(n298), .Z(Y[23]) );
  TBUF_X1 \Y_tri[24]  ( .A(n477), .EN(n298), .Z(Y[24]) );
  TBUF_X1 \Y_tri[25]  ( .A(n476), .EN(n298), .Z(Y[25]) );
  TBUF_X1 \Y_tri[26]  ( .A(n475), .EN(n298), .Z(Y[26]) );
  TBUF_X1 \Y_tri[27]  ( .A(n474), .EN(n298), .Z(Y[27]) );
  TBUF_X1 \Y_tri[28]  ( .A(n473), .EN(n298), .Z(Y[28]) );
  TBUF_X1 \Y_tri[29]  ( .A(n472), .EN(n298), .Z(Y[29]) );
  TBUF_X1 \Y_tri[30]  ( .A(n471), .EN(n298), .Z(Y[30]) );
  TBUF_X1 \Y_tri[31]  ( .A(n470), .EN(n298), .Z(Y[31]) );
  TBUF_X1 \Y_tri[32]  ( .A(n469), .EN(n298), .Z(Y[32]) );
  TBUF_X1 \Y_tri[33]  ( .A(n468), .EN(n299), .Z(Y[33]) );
  TBUF_X1 \Y_tri[34]  ( .A(n467), .EN(n299), .Z(Y[34]) );
  TBUF_X1 \Y_tri[35]  ( .A(n466), .EN(n299), .Z(Y[35]) );
  TBUF_X1 \Y_tri[36]  ( .A(n465), .EN(n299), .Z(Y[36]) );
  TBUF_X1 \Y_tri[37]  ( .A(n464), .EN(n299), .Z(Y[37]) );
  TBUF_X1 \Y_tri[38]  ( .A(n463), .EN(n299), .Z(Y[38]) );
  TBUF_X1 \Y_tri[39]  ( .A(n462), .EN(n299), .Z(Y[39]) );
  TBUF_X1 \Y_tri[40]  ( .A(n461), .EN(n299), .Z(Y[40]) );
  TBUF_X1 \Y_tri[41]  ( .A(n460), .EN(n299), .Z(Y[41]) );
  TBUF_X1 \Y_tri[42]  ( .A(n459), .EN(n299), .Z(Y[42]) );
  TBUF_X1 \Y_tri[43]  ( .A(n458), .EN(n299), .Z(Y[43]) );
  TBUF_X1 \Y_tri[44]  ( .A(n457), .EN(n300), .Z(Y[44]) );
  TBUF_X1 \Y_tri[7]  ( .A(n495), .EN(n296), .Z(Y[7]) );
  TBUF_X1 \Y_tri[8]  ( .A(n494), .EN(n296), .Z(Y[8]) );
  TBUF_X1 \Y_tri[10]  ( .A(n491), .EN(n296), .Z(Y[10]) );
  TBUF_X1 \Y_tri[11]  ( .A(n490), .EN(n297), .Z(Y[11]) );
  TBUF_X1 \Y_tri[12]  ( .A(n489), .EN(n297), .Z(Y[12]) );
  TBUF_X1 \Y_tri[13]  ( .A(n488), .EN(n297), .Z(Y[13]) );
  TBUF_X1 \Y_tri[14]  ( .A(n487), .EN(n297), .Z(Y[14]) );
  TBUF_X1 \Y_tri[15]  ( .A(n486), .EN(n297), .Z(Y[15]) );
  TBUF_X1 \Y_tri[16]  ( .A(n485), .EN(n297), .Z(Y[16]) );
  TBUF_X1 \Y_tri[0]  ( .A(n502), .EN(n296), .Z(Y[0]) );
  TBUF_X1 \Y_tri[1]  ( .A(n501), .EN(n296), .Z(Y[1]) );
  TBUF_X1 \Y_tri[2]  ( .A(n500), .EN(n296), .Z(Y[2]) );
  TBUF_X1 \Y_tri[3]  ( .A(n499), .EN(n296), .Z(Y[3]) );
  TBUF_X1 \Y_tri[4]  ( .A(n498), .EN(n296), .Z(Y[4]) );
  TBUF_X1 \Y_tri[5]  ( .A(n497), .EN(n296), .Z(Y[5]) );
  TBUF_X1 \Y_tri[6]  ( .A(n496), .EN(n296), .Z(Y[6]) );
  TBUF_X1 \Y_tri[9]  ( .A(n492), .EN(n296), .Z(Y[9]) );
  NAND2_X1 U2 ( .A1(n393), .A2(n392), .ZN(n458) );
  AOI22_X1 U3 ( .A1(plusA[43]), .A2(n281), .B1(plus2A[43]), .B2(n275), .ZN(
        n393) );
  AOI22_X1 U4 ( .A1(minus2A[43]), .A2(n293), .B1(minusA[43]), .B2(n287), .ZN(
        n392) );
  NAND2_X1 U5 ( .A1(n385), .A2(n384), .ZN(n462) );
  AOI22_X1 U6 ( .A1(plusA[39]), .A2(n281), .B1(plus2A[39]), .B2(n275), .ZN(
        n385) );
  AOI22_X1 U7 ( .A1(minus2A[39]), .A2(n293), .B1(minusA[39]), .B2(n287), .ZN(
        n384) );
  NAND2_X1 U8 ( .A1(n377), .A2(n376), .ZN(n466) );
  AOI22_X1 U9 ( .A1(plusA[35]), .A2(n280), .B1(plus2A[35]), .B2(n274), .ZN(
        n377) );
  AOI22_X1 U10 ( .A1(minus2A[35]), .A2(n292), .B1(minusA[35]), .B2(n286), .ZN(
        n376) );
  NAND2_X1 U11 ( .A1(n369), .A2(n368), .ZN(n470) );
  AOI22_X1 U12 ( .A1(plusA[31]), .A2(n280), .B1(plus2A[31]), .B2(n274), .ZN(
        n369) );
  AOI22_X1 U13 ( .A1(minus2A[31]), .A2(n292), .B1(minusA[31]), .B2(n286), .ZN(
        n368) );
  NAND2_X1 U14 ( .A1(n361), .A2(n360), .ZN(n474) );
  AOI22_X1 U15 ( .A1(plusA[27]), .A2(n280), .B1(plus2A[27]), .B2(n274), .ZN(
        n361) );
  AOI22_X1 U16 ( .A1(minus2A[27]), .A2(n292), .B1(minusA[27]), .B2(n286), .ZN(
        n360) );
  NAND2_X1 U17 ( .A1(n389), .A2(n388), .ZN(n460) );
  AOI22_X1 U18 ( .A1(plusA[41]), .A2(n281), .B1(plus2A[41]), .B2(n275), .ZN(
        n389) );
  AOI22_X1 U19 ( .A1(minus2A[41]), .A2(n293), .B1(minusA[41]), .B2(n287), .ZN(
        n388) );
  NAND2_X1 U20 ( .A1(n381), .A2(n380), .ZN(n464) );
  AOI22_X1 U21 ( .A1(plusA[37]), .A2(n281), .B1(plus2A[37]), .B2(n275), .ZN(
        n381) );
  AOI22_X1 U22 ( .A1(minus2A[37]), .A2(n293), .B1(minusA[37]), .B2(n287), .ZN(
        n380) );
  NAND2_X1 U23 ( .A1(n373), .A2(n372), .ZN(n468) );
  AOI22_X1 U24 ( .A1(plusA[33]), .A2(n280), .B1(plus2A[33]), .B2(n274), .ZN(
        n373) );
  AOI22_X1 U25 ( .A1(minus2A[33]), .A2(n292), .B1(minusA[33]), .B2(n286), .ZN(
        n372) );
  NAND2_X1 U26 ( .A1(n365), .A2(n364), .ZN(n472) );
  AOI22_X1 U27 ( .A1(plusA[29]), .A2(n280), .B1(plus2A[29]), .B2(n274), .ZN(
        n365) );
  AOI22_X1 U28 ( .A1(minus2A[29]), .A2(n292), .B1(minusA[29]), .B2(n286), .ZN(
        n364) );
  NAND2_X1 U29 ( .A1(n357), .A2(n356), .ZN(n476) );
  AOI22_X1 U30 ( .A1(plusA[25]), .A2(n280), .B1(plus2A[25]), .B2(n274), .ZN(
        n357) );
  AOI22_X1 U31 ( .A1(minus2A[25]), .A2(n292), .B1(minusA[25]), .B2(n286), .ZN(
        n356) );
  NAND2_X1 U32 ( .A1(n395), .A2(n394), .ZN(n457) );
  AOI22_X1 U33 ( .A1(plusA[44]), .A2(n281), .B1(plus2A[44]), .B2(n275), .ZN(
        n395) );
  AOI22_X1 U34 ( .A1(minus2A[44]), .A2(n293), .B1(minusA[44]), .B2(n287), .ZN(
        n394) );
  NAND2_X1 U35 ( .A1(n387), .A2(n386), .ZN(n461) );
  AOI22_X1 U36 ( .A1(plusA[40]), .A2(n281), .B1(plus2A[40]), .B2(n275), .ZN(
        n387) );
  AOI22_X1 U37 ( .A1(minus2A[40]), .A2(n293), .B1(minusA[40]), .B2(n287), .ZN(
        n386) );
  NAND2_X1 U38 ( .A1(n379), .A2(n378), .ZN(n465) );
  AOI22_X1 U39 ( .A1(plusA[36]), .A2(n281), .B1(plus2A[36]), .B2(n275), .ZN(
        n379) );
  AOI22_X1 U40 ( .A1(minus2A[36]), .A2(n293), .B1(minusA[36]), .B2(n287), .ZN(
        n378) );
  NAND2_X1 U41 ( .A1(n371), .A2(n370), .ZN(n469) );
  AOI22_X1 U42 ( .A1(plusA[32]), .A2(n280), .B1(plus2A[32]), .B2(n274), .ZN(
        n371) );
  AOI22_X1 U43 ( .A1(minus2A[32]), .A2(n292), .B1(minusA[32]), .B2(n286), .ZN(
        n370) );
  NAND2_X1 U44 ( .A1(n363), .A2(n362), .ZN(n473) );
  AOI22_X1 U45 ( .A1(plusA[28]), .A2(n280), .B1(plus2A[28]), .B2(n274), .ZN(
        n363) );
  AOI22_X1 U46 ( .A1(minus2A[28]), .A2(n292), .B1(minusA[28]), .B2(n286), .ZN(
        n362) );
  NAND2_X1 U47 ( .A1(n355), .A2(n354), .ZN(n477) );
  AOI22_X1 U48 ( .A1(plusA[24]), .A2(n280), .B1(plus2A[24]), .B2(n274), .ZN(
        n355) );
  AOI22_X1 U49 ( .A1(minus2A[24]), .A2(n292), .B1(minusA[24]), .B2(n286), .ZN(
        n354) );
  NAND2_X1 U50 ( .A1(n391), .A2(n390), .ZN(n459) );
  AOI22_X1 U51 ( .A1(plusA[42]), .A2(n281), .B1(plus2A[42]), .B2(n275), .ZN(
        n391) );
  AOI22_X1 U52 ( .A1(minus2A[42]), .A2(n293), .B1(minusA[42]), .B2(n287), .ZN(
        n390) );
  NAND2_X1 U53 ( .A1(n383), .A2(n382), .ZN(n463) );
  AOI22_X1 U54 ( .A1(plusA[38]), .A2(n281), .B1(plus2A[38]), .B2(n275), .ZN(
        n383) );
  AOI22_X1 U55 ( .A1(minus2A[38]), .A2(n293), .B1(minusA[38]), .B2(n287), .ZN(
        n382) );
  NAND2_X1 U56 ( .A1(n375), .A2(n374), .ZN(n467) );
  AOI22_X1 U57 ( .A1(plusA[34]), .A2(n280), .B1(plus2A[34]), .B2(n274), .ZN(
        n375) );
  AOI22_X1 U58 ( .A1(minus2A[34]), .A2(n292), .B1(minusA[34]), .B2(n286), .ZN(
        n374) );
  NAND2_X1 U59 ( .A1(n367), .A2(n366), .ZN(n471) );
  AOI22_X1 U60 ( .A1(plusA[30]), .A2(n280), .B1(plus2A[30]), .B2(n274), .ZN(
        n367) );
  AOI22_X1 U61 ( .A1(minus2A[30]), .A2(n292), .B1(minusA[30]), .B2(n286), .ZN(
        n366) );
  NAND2_X1 U62 ( .A1(n359), .A2(n358), .ZN(n475) );
  AOI22_X1 U63 ( .A1(plusA[26]), .A2(n280), .B1(plus2A[26]), .B2(n274), .ZN(
        n359) );
  AOI22_X1 U64 ( .A1(minus2A[26]), .A2(n292), .B1(minusA[26]), .B2(n286), .ZN(
        n358) );
  NAND2_X1 U65 ( .A1(n437), .A2(n436), .ZN(n438) );
  AOI22_X1 U66 ( .A1(plusA[63]), .A2(n283), .B1(plus2A[63]), .B2(n277), .ZN(
        n437) );
  AOI22_X1 U67 ( .A1(minus2A[63]), .A2(n295), .B1(minusA[63]), .B2(n289), .ZN(
        n436) );
  NAND2_X1 U68 ( .A1(n409), .A2(n408), .ZN(n450) );
  AOI22_X1 U69 ( .A1(plusA[51]), .A2(n282), .B1(plus2A[51]), .B2(n276), .ZN(
        n409) );
  AOI22_X1 U70 ( .A1(minus2A[51]), .A2(n294), .B1(minusA[51]), .B2(n288), .ZN(
        n408) );
  NAND2_X1 U71 ( .A1(n401), .A2(n400), .ZN(n454) );
  AOI22_X1 U72 ( .A1(plusA[47]), .A2(n281), .B1(plus2A[47]), .B2(n275), .ZN(
        n401) );
  AOI22_X1 U73 ( .A1(minus2A[47]), .A2(n293), .B1(minusA[47]), .B2(n287), .ZN(
        n400) );
  NAND2_X1 U74 ( .A1(n419), .A2(n418), .ZN(n445) );
  AOI22_X1 U75 ( .A1(plusA[56]), .A2(n282), .B1(plus2A[56]), .B2(n276), .ZN(
        n419) );
  AOI22_X1 U76 ( .A1(minus2A[56]), .A2(n294), .B1(minusA[56]), .B2(n288), .ZN(
        n418) );
  NAND2_X1 U77 ( .A1(n415), .A2(n414), .ZN(n447) );
  AOI22_X1 U78 ( .A1(plusA[54]), .A2(n282), .B1(plus2A[54]), .B2(n276), .ZN(
        n415) );
  AOI22_X1 U79 ( .A1(minus2A[54]), .A2(n294), .B1(minusA[54]), .B2(n288), .ZN(
        n414) );
  NAND2_X1 U80 ( .A1(n421), .A2(n420), .ZN(n444) );
  AOI22_X1 U81 ( .A1(plusA[57]), .A2(n282), .B1(plus2A[57]), .B2(n276), .ZN(
        n421) );
  AOI22_X1 U82 ( .A1(minus2A[57]), .A2(n294), .B1(minusA[57]), .B2(n288), .ZN(
        n420) );
  NAND2_X1 U83 ( .A1(n417), .A2(n416), .ZN(n446) );
  AOI22_X1 U84 ( .A1(plusA[55]), .A2(n282), .B1(plus2A[55]), .B2(n276), .ZN(
        n417) );
  AOI22_X1 U85 ( .A1(minus2A[55]), .A2(n294), .B1(minusA[55]), .B2(n288), .ZN(
        n416) );
  NAND2_X1 U86 ( .A1(n413), .A2(n412), .ZN(n448) );
  AOI22_X1 U87 ( .A1(plusA[53]), .A2(n282), .B1(plus2A[53]), .B2(n276), .ZN(
        n413) );
  AOI22_X1 U88 ( .A1(minus2A[53]), .A2(n294), .B1(minusA[53]), .B2(n288), .ZN(
        n412) );
  NAND2_X1 U89 ( .A1(n405), .A2(n404), .ZN(n452) );
  AOI22_X1 U90 ( .A1(plusA[49]), .A2(n282), .B1(plus2A[49]), .B2(n276), .ZN(
        n405) );
  AOI22_X1 U91 ( .A1(minus2A[49]), .A2(n294), .B1(minusA[49]), .B2(n288), .ZN(
        n404) );
  NAND2_X1 U92 ( .A1(n397), .A2(n396), .ZN(n456) );
  AOI22_X1 U93 ( .A1(plusA[45]), .A2(n281), .B1(plus2A[45]), .B2(n275), .ZN(
        n397) );
  AOI22_X1 U94 ( .A1(minus2A[45]), .A2(n293), .B1(minusA[45]), .B2(n287), .ZN(
        n396) );
  NAND2_X1 U95 ( .A1(n411), .A2(n410), .ZN(n449) );
  AOI22_X1 U96 ( .A1(plusA[52]), .A2(n282), .B1(plus2A[52]), .B2(n276), .ZN(
        n411) );
  AOI22_X1 U97 ( .A1(minus2A[52]), .A2(n294), .B1(minusA[52]), .B2(n288), .ZN(
        n410) );
  NAND2_X1 U98 ( .A1(n403), .A2(n402), .ZN(n453) );
  AOI22_X1 U99 ( .A1(plusA[48]), .A2(n282), .B1(plus2A[48]), .B2(n276), .ZN(
        n403) );
  AOI22_X1 U100 ( .A1(minus2A[48]), .A2(n294), .B1(minusA[48]), .B2(n288), 
        .ZN(n402) );
  NAND2_X1 U101 ( .A1(n407), .A2(n406), .ZN(n451) );
  AOI22_X1 U102 ( .A1(plusA[50]), .A2(n282), .B1(plus2A[50]), .B2(n276), .ZN(
        n407) );
  AOI22_X1 U103 ( .A1(minus2A[50]), .A2(n294), .B1(minusA[50]), .B2(n288), 
        .ZN(n406) );
  NAND2_X1 U104 ( .A1(n399), .A2(n398), .ZN(n455) );
  AOI22_X1 U105 ( .A1(plusA[46]), .A2(n281), .B1(plus2A[46]), .B2(n275), .ZN(
        n399) );
  AOI22_X1 U106 ( .A1(minus2A[46]), .A2(n293), .B1(minusA[46]), .B2(n287), 
        .ZN(n398) );
  NAND2_X1 U107 ( .A1(n431), .A2(n430), .ZN(n439) );
  AOI22_X1 U108 ( .A1(plusA[62]), .A2(n283), .B1(plus2A[62]), .B2(n277), .ZN(
        n431) );
  AOI22_X1 U109 ( .A1(minus2A[62]), .A2(n295), .B1(minusA[62]), .B2(n289), 
        .ZN(n430) );
  NAND2_X1 U110 ( .A1(n429), .A2(n428), .ZN(n440) );
  AOI22_X1 U111 ( .A1(plusA[61]), .A2(n283), .B1(plus2A[61]), .B2(n277), .ZN(
        n429) );
  AOI22_X1 U112 ( .A1(minus2A[61]), .A2(n295), .B1(minusA[61]), .B2(n289), 
        .ZN(n428) );
  NAND2_X1 U113 ( .A1(n427), .A2(n426), .ZN(n441) );
  AOI22_X1 U114 ( .A1(plusA[60]), .A2(n283), .B1(plus2A[60]), .B2(n277), .ZN(
        n427) );
  AOI22_X1 U115 ( .A1(minus2A[60]), .A2(n295), .B1(minusA[60]), .B2(n289), 
        .ZN(n426) );
  NAND2_X1 U116 ( .A1(n425), .A2(n424), .ZN(n442) );
  AOI22_X1 U117 ( .A1(plusA[59]), .A2(n282), .B1(plus2A[59]), .B2(n276), .ZN(
        n425) );
  AOI22_X1 U118 ( .A1(minus2A[59]), .A2(n294), .B1(minusA[59]), .B2(n288), 
        .ZN(n424) );
  NAND2_X1 U119 ( .A1(n423), .A2(n422), .ZN(n443) );
  AOI22_X1 U120 ( .A1(plusA[58]), .A2(n282), .B1(plus2A[58]), .B2(n276), .ZN(
        n423) );
  AOI22_X1 U121 ( .A1(minus2A[58]), .A2(n294), .B1(minusA[58]), .B2(n288), 
        .ZN(n422) );
  BUF_X1 U122 ( .A(n493), .Z(n296) );
  BUF_X1 U123 ( .A(n493), .Z(n297) );
  BUF_X1 U124 ( .A(n433), .Z(n280) );
  BUF_X1 U125 ( .A(n433), .Z(n279) );
  BUF_X1 U126 ( .A(n435), .Z(n292) );
  BUF_X1 U127 ( .A(n435), .Z(n291) );
  BUF_X1 U128 ( .A(n434), .Z(n286) );
  BUF_X1 U129 ( .A(n432), .Z(n274) );
  BUF_X1 U130 ( .A(n434), .Z(n285) );
  BUF_X1 U131 ( .A(n432), .Z(n273) );
  BUF_X1 U132 ( .A(n493), .Z(n298) );
  NAND2_X1 U133 ( .A1(n353), .A2(n352), .ZN(n478) );
  AOI22_X1 U134 ( .A1(plusA[23]), .A2(n279), .B1(plus2A[23]), .B2(n273), .ZN(
        n353) );
  AOI22_X1 U135 ( .A1(minus2A[23]), .A2(n291), .B1(minusA[23]), .B2(n285), 
        .ZN(n352) );
  NAND2_X1 U136 ( .A1(n351), .A2(n350), .ZN(n479) );
  AOI22_X1 U137 ( .A1(plusA[22]), .A2(n279), .B1(plus2A[22]), .B2(n273), .ZN(
        n351) );
  AOI22_X1 U138 ( .A1(minus2A[22]), .A2(n291), .B1(minusA[22]), .B2(n285), 
        .ZN(n350) );
  BUF_X1 U139 ( .A(n433), .Z(n281) );
  BUF_X1 U140 ( .A(n435), .Z(n293) );
  BUF_X1 U141 ( .A(n434), .Z(n287) );
  BUF_X1 U142 ( .A(n432), .Z(n275) );
  BUF_X1 U143 ( .A(n493), .Z(n299) );
  BUF_X1 U144 ( .A(n433), .Z(n282) );
  BUF_X1 U145 ( .A(n435), .Z(n294) );
  BUF_X1 U146 ( .A(n434), .Z(n288) );
  BUF_X1 U147 ( .A(n432), .Z(n276) );
  BUF_X1 U148 ( .A(n493), .Z(n300) );
  BUF_X1 U149 ( .A(n493), .Z(n301) );
  BUF_X1 U150 ( .A(n433), .Z(n278) );
  BUF_X1 U151 ( .A(n435), .Z(n290) );
  BUF_X1 U152 ( .A(n434), .Z(n284) );
  BUF_X1 U153 ( .A(n432), .Z(n272) );
  NOR2_X1 U154 ( .A1(n323), .A2(n304), .ZN(n493) );
  INV_X1 U155 ( .A(SEL[2]), .ZN(n304) );
  NOR2_X1 U156 ( .A1(SEL[1]), .A2(SEL[0]), .ZN(n323) );
  NOR3_X1 U157 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n302), .ZN(n434) );
  NOR3_X1 U158 ( .A1(SEL[1]), .A2(SEL[2]), .A3(n303), .ZN(n433) );
  NOR3_X1 U159 ( .A1(n302), .A2(SEL[2]), .A3(n303), .ZN(n432) );
  AND2_X1 U160 ( .A1(SEL[2]), .A2(n323), .ZN(n435) );
  INV_X1 U161 ( .A(SEL[1]), .ZN(n302) );
  INV_X1 U162 ( .A(SEL[0]), .ZN(n303) );
  NAND2_X1 U163 ( .A1(n349), .A2(n348), .ZN(n480) );
  AOI22_X1 U164 ( .A1(plusA[21]), .A2(n279), .B1(plus2A[21]), .B2(n273), .ZN(
        n349) );
  AOI22_X1 U165 ( .A1(minus2A[21]), .A2(n291), .B1(minusA[21]), .B2(n285), 
        .ZN(n348) );
  NAND2_X1 U166 ( .A1(n347), .A2(n346), .ZN(n481) );
  AOI22_X1 U167 ( .A1(plusA[20]), .A2(n279), .B1(plus2A[20]), .B2(n273), .ZN(
        n347) );
  AOI22_X1 U168 ( .A1(minus2A[20]), .A2(n291), .B1(minusA[20]), .B2(n285), 
        .ZN(n346) );
  NAND2_X1 U169 ( .A1(n345), .A2(n344), .ZN(n482) );
  AOI22_X1 U170 ( .A1(plusA[19]), .A2(n279), .B1(plus2A[19]), .B2(n273), .ZN(
        n345) );
  AOI22_X1 U171 ( .A1(minus2A[19]), .A2(n291), .B1(minusA[19]), .B2(n285), 
        .ZN(n344) );
  NAND2_X1 U172 ( .A1(n343), .A2(n342), .ZN(n483) );
  AOI22_X1 U173 ( .A1(plusA[18]), .A2(n279), .B1(plus2A[18]), .B2(n273), .ZN(
        n343) );
  AOI22_X1 U174 ( .A1(minus2A[18]), .A2(n291), .B1(minusA[18]), .B2(n285), 
        .ZN(n342) );
  NAND2_X1 U175 ( .A1(n341), .A2(n340), .ZN(n484) );
  AOI22_X1 U176 ( .A1(plusA[17]), .A2(n279), .B1(plus2A[17]), .B2(n273), .ZN(
        n341) );
  AOI22_X1 U177 ( .A1(minus2A[17]), .A2(n291), .B1(minusA[17]), .B2(n285), 
        .ZN(n340) );
  NAND2_X1 U178 ( .A1(n337), .A2(n336), .ZN(n486) );
  AOI22_X1 U179 ( .A1(plusA[15]), .A2(n279), .B1(plus2A[15]), .B2(n273), .ZN(
        n337) );
  AOI22_X1 U180 ( .A1(minus2A[15]), .A2(n291), .B1(minusA[15]), .B2(n285), 
        .ZN(n336) );
  NAND2_X1 U181 ( .A1(n335), .A2(n334), .ZN(n487) );
  AOI22_X1 U182 ( .A1(plusA[14]), .A2(n279), .B1(plus2A[14]), .B2(n273), .ZN(
        n335) );
  AOI22_X1 U183 ( .A1(minus2A[14]), .A2(n291), .B1(minusA[14]), .B2(n285), 
        .ZN(n334) );
  NAND2_X1 U184 ( .A1(n333), .A2(n332), .ZN(n488) );
  AOI22_X1 U185 ( .A1(plusA[13]), .A2(n279), .B1(plus2A[13]), .B2(n273), .ZN(
        n333) );
  AOI22_X1 U186 ( .A1(minus2A[13]), .A2(n291), .B1(minusA[13]), .B2(n285), 
        .ZN(n332) );
  NAND2_X1 U187 ( .A1(n329), .A2(n328), .ZN(n490) );
  AOI22_X1 U188 ( .A1(plusA[11]), .A2(n278), .B1(plus2A[11]), .B2(n272), .ZN(
        n329) );
  AOI22_X1 U189 ( .A1(minus2A[11]), .A2(n290), .B1(minusA[11]), .B2(n284), 
        .ZN(n328) );
  NAND2_X1 U190 ( .A1(n327), .A2(n326), .ZN(n491) );
  AOI22_X1 U191 ( .A1(plusA[10]), .A2(n278), .B1(plus2A[10]), .B2(n272), .ZN(
        n327) );
  AOI22_X1 U192 ( .A1(minus2A[10]), .A2(n290), .B1(minusA[10]), .B2(n284), 
        .ZN(n326) );
  NAND2_X1 U193 ( .A1(n325), .A2(n324), .ZN(n492) );
  AOI22_X1 U194 ( .A1(plusA[9]), .A2(n278), .B1(plus2A[9]), .B2(n272), .ZN(
        n325) );
  AOI22_X1 U195 ( .A1(minus2A[9]), .A2(n290), .B1(minusA[9]), .B2(n284), .ZN(
        n324) );
  NAND2_X1 U196 ( .A1(n320), .A2(n319), .ZN(n495) );
  AOI22_X1 U197 ( .A1(plusA[7]), .A2(n278), .B1(plus2A[7]), .B2(n272), .ZN(
        n320) );
  AOI22_X1 U198 ( .A1(minus2A[7]), .A2(n290), .B1(minusA[7]), .B2(n284), .ZN(
        n319) );
  NAND2_X1 U199 ( .A1(n318), .A2(n317), .ZN(n496) );
  AOI22_X1 U200 ( .A1(plusA[6]), .A2(n278), .B1(plus2A[6]), .B2(n272), .ZN(
        n318) );
  AOI22_X1 U201 ( .A1(minus2A[6]), .A2(n290), .B1(minusA[6]), .B2(n284), .ZN(
        n317) );
  NAND2_X1 U202 ( .A1(n316), .A2(n315), .ZN(n497) );
  AOI22_X1 U203 ( .A1(plusA[5]), .A2(n278), .B1(plus2A[5]), .B2(n272), .ZN(
        n316) );
  AOI22_X1 U204 ( .A1(minus2A[5]), .A2(n290), .B1(minusA[5]), .B2(n284), .ZN(
        n315) );
  NAND2_X1 U205 ( .A1(n312), .A2(n311), .ZN(n499) );
  AOI22_X1 U206 ( .A1(plusA[3]), .A2(n278), .B1(plus2A[3]), .B2(n272), .ZN(
        n312) );
  AOI22_X1 U207 ( .A1(minus2A[3]), .A2(n290), .B1(minusA[3]), .B2(n284), .ZN(
        n311) );
  NAND2_X1 U208 ( .A1(n339), .A2(n338), .ZN(n485) );
  AOI22_X1 U209 ( .A1(plusA[16]), .A2(n279), .B1(plus2A[16]), .B2(n273), .ZN(
        n339) );
  AOI22_X1 U210 ( .A1(minus2A[16]), .A2(n291), .B1(minusA[16]), .B2(n285), 
        .ZN(n338) );
  NAND2_X1 U211 ( .A1(n331), .A2(n330), .ZN(n489) );
  AOI22_X1 U212 ( .A1(plusA[12]), .A2(n279), .B1(plus2A[12]), .B2(n273), .ZN(
        n331) );
  AOI22_X1 U213 ( .A1(minus2A[12]), .A2(n291), .B1(minusA[12]), .B2(n285), 
        .ZN(n330) );
  NAND2_X1 U214 ( .A1(n322), .A2(n321), .ZN(n494) );
  AOI22_X1 U215 ( .A1(plusA[8]), .A2(n278), .B1(plus2A[8]), .B2(n272), .ZN(
        n322) );
  AOI22_X1 U216 ( .A1(minus2A[8]), .A2(n290), .B1(minusA[8]), .B2(n284), .ZN(
        n321) );
  NAND2_X1 U217 ( .A1(n314), .A2(n313), .ZN(n498) );
  AOI22_X1 U218 ( .A1(plusA[4]), .A2(n278), .B1(plus2A[4]), .B2(n272), .ZN(
        n314) );
  AOI22_X1 U219 ( .A1(minus2A[4]), .A2(n290), .B1(minusA[4]), .B2(n284), .ZN(
        n313) );
  NAND2_X1 U220 ( .A1(n310), .A2(n309), .ZN(n500) );
  AOI22_X1 U221 ( .A1(plusA[2]), .A2(n278), .B1(plus2A[2]), .B2(n272), .ZN(
        n310) );
  AOI22_X1 U222 ( .A1(minus2A[2]), .A2(n290), .B1(minusA[2]), .B2(n284), .ZN(
        n309) );
  NAND2_X1 U223 ( .A1(n308), .A2(n307), .ZN(n501) );
  AOI22_X1 U224 ( .A1(plusA[1]), .A2(n278), .B1(plus2A[1]), .B2(n272), .ZN(
        n308) );
  AOI22_X1 U225 ( .A1(minus2A[1]), .A2(n290), .B1(minusA[1]), .B2(n284), .ZN(
        n307) );
  NAND2_X1 U226 ( .A1(n306), .A2(n305), .ZN(n502) );
  AOI22_X1 U227 ( .A1(plusA[0]), .A2(n278), .B1(plus2A[0]), .B2(n272), .ZN(
        n306) );
  AOI22_X1 U228 ( .A1(minus2A[0]), .A2(n290), .B1(minusA[0]), .B2(n284), .ZN(
        n305) );
  CLKBUF_X1 U229 ( .A(n432), .Z(n277) );
  CLKBUF_X1 U230 ( .A(n433), .Z(n283) );
  CLKBUF_X1 U231 ( .A(n434), .Z(n289) );
  CLKBUF_X1 U232 ( .A(n435), .Z(n295) );
endmodule


module FA_384 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_383 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_382 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_381 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_380 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_379 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_378 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_377 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_376 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_375 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_374 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_373 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_372 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_371 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_370 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_369 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_368 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_367 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_366 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_365 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_364 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_363 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_362 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_361 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_360 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_359 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_358 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_357 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_356 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_355 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_354 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_353 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_352 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_351 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_350 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_349 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_348 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_347 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_346 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_345 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_344 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_343 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_342 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_341 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_340 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_339 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_338 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_337 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_336 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_335 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_334 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_333 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_332 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_331 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_330 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_329 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_328 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_327 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_326 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_325 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_324 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_323 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_322 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_321 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N64_6 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Ci;
  output Co;

  wire   [63:1] CTMP;
  tri   [63:0] A;

  FA_384 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_383 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_382 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_381 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(CTMP[4]) );
  FA_380 FAI_5 ( .A(A[4]), .B(B[4]), .Ci(CTMP[4]), .S(S[4]), .Co(CTMP[5]) );
  FA_379 FAI_6 ( .A(A[5]), .B(B[5]), .Ci(CTMP[5]), .S(S[5]), .Co(CTMP[6]) );
  FA_378 FAI_7 ( .A(A[6]), .B(B[6]), .Ci(CTMP[6]), .S(S[6]), .Co(CTMP[7]) );
  FA_377 FAI_8 ( .A(A[7]), .B(B[7]), .Ci(CTMP[7]), .S(S[7]), .Co(CTMP[8]) );
  FA_376 FAI_9 ( .A(A[8]), .B(B[8]), .Ci(CTMP[8]), .S(S[8]), .Co(CTMP[9]) );
  FA_375 FAI_10 ( .A(A[9]), .B(B[9]), .Ci(CTMP[9]), .S(S[9]), .Co(CTMP[10]) );
  FA_374 FAI_11 ( .A(A[10]), .B(B[10]), .Ci(CTMP[10]), .S(S[10]), .Co(CTMP[11]) );
  FA_373 FAI_12 ( .A(A[11]), .B(B[11]), .Ci(CTMP[11]), .S(S[11]), .Co(CTMP[12]) );
  FA_372 FAI_13 ( .A(A[12]), .B(B[12]), .Ci(CTMP[12]), .S(S[12]), .Co(CTMP[13]) );
  FA_371 FAI_14 ( .A(A[13]), .B(B[13]), .Ci(CTMP[13]), .S(S[13]), .Co(CTMP[14]) );
  FA_370 FAI_15 ( .A(A[14]), .B(B[14]), .Ci(CTMP[14]), .S(S[14]), .Co(CTMP[15]) );
  FA_369 FAI_16 ( .A(A[15]), .B(B[15]), .Ci(CTMP[15]), .S(S[15]), .Co(CTMP[16]) );
  FA_368 FAI_17 ( .A(A[16]), .B(B[16]), .Ci(CTMP[16]), .S(S[16]), .Co(CTMP[17]) );
  FA_367 FAI_18 ( .A(A[17]), .B(B[17]), .Ci(CTMP[17]), .S(S[17]), .Co(CTMP[18]) );
  FA_366 FAI_19 ( .A(A[18]), .B(B[18]), .Ci(CTMP[18]), .S(S[18]), .Co(CTMP[19]) );
  FA_365 FAI_20 ( .A(A[19]), .B(B[19]), .Ci(CTMP[19]), .S(S[19]), .Co(CTMP[20]) );
  FA_364 FAI_21 ( .A(A[20]), .B(B[20]), .Ci(CTMP[20]), .S(S[20]), .Co(CTMP[21]) );
  FA_363 FAI_22 ( .A(A[21]), .B(B[21]), .Ci(CTMP[21]), .S(S[21]), .Co(CTMP[22]) );
  FA_362 FAI_23 ( .A(A[22]), .B(B[22]), .Ci(CTMP[22]), .S(S[22]), .Co(CTMP[23]) );
  FA_361 FAI_24 ( .A(A[23]), .B(B[23]), .Ci(CTMP[23]), .S(S[23]), .Co(CTMP[24]) );
  FA_360 FAI_25 ( .A(A[24]), .B(B[24]), .Ci(CTMP[24]), .S(S[24]), .Co(CTMP[25]) );
  FA_359 FAI_26 ( .A(A[25]), .B(B[25]), .Ci(CTMP[25]), .S(S[25]), .Co(CTMP[26]) );
  FA_358 FAI_27 ( .A(A[26]), .B(B[26]), .Ci(CTMP[26]), .S(S[26]), .Co(CTMP[27]) );
  FA_357 FAI_28 ( .A(A[27]), .B(B[27]), .Ci(CTMP[27]), .S(S[27]), .Co(CTMP[28]) );
  FA_356 FAI_29 ( .A(A[28]), .B(B[28]), .Ci(CTMP[28]), .S(S[28]), .Co(CTMP[29]) );
  FA_355 FAI_30 ( .A(A[29]), .B(B[29]), .Ci(CTMP[29]), .S(S[29]), .Co(CTMP[30]) );
  FA_354 FAI_31 ( .A(A[30]), .B(B[30]), .Ci(CTMP[30]), .S(S[30]), .Co(CTMP[31]) );
  FA_353 FAI_32 ( .A(A[31]), .B(B[31]), .Ci(CTMP[31]), .S(S[31]), .Co(CTMP[32]) );
  FA_352 FAI_33 ( .A(A[32]), .B(B[32]), .Ci(CTMP[32]), .S(S[32]), .Co(CTMP[33]) );
  FA_351 FAI_34 ( .A(A[33]), .B(B[33]), .Ci(CTMP[33]), .S(S[33]), .Co(CTMP[34]) );
  FA_350 FAI_35 ( .A(A[34]), .B(B[34]), .Ci(CTMP[34]), .S(S[34]), .Co(CTMP[35]) );
  FA_349 FAI_36 ( .A(A[35]), .B(B[35]), .Ci(CTMP[35]), .S(S[35]), .Co(CTMP[36]) );
  FA_348 FAI_37 ( .A(A[36]), .B(B[36]), .Ci(CTMP[36]), .S(S[36]), .Co(CTMP[37]) );
  FA_347 FAI_38 ( .A(A[37]), .B(B[37]), .Ci(CTMP[37]), .S(S[37]), .Co(CTMP[38]) );
  FA_346 FAI_39 ( .A(A[38]), .B(B[38]), .Ci(CTMP[38]), .S(S[38]), .Co(CTMP[39]) );
  FA_345 FAI_40 ( .A(A[39]), .B(B[39]), .Ci(CTMP[39]), .S(S[39]), .Co(CTMP[40]) );
  FA_344 FAI_41 ( .A(A[40]), .B(B[40]), .Ci(CTMP[40]), .S(S[40]), .Co(CTMP[41]) );
  FA_343 FAI_42 ( .A(A[41]), .B(B[41]), .Ci(CTMP[41]), .S(S[41]), .Co(CTMP[42]) );
  FA_342 FAI_43 ( .A(A[42]), .B(B[42]), .Ci(CTMP[42]), .S(S[42]), .Co(CTMP[43]) );
  FA_341 FAI_44 ( .A(A[43]), .B(B[43]), .Ci(CTMP[43]), .S(S[43]), .Co(CTMP[44]) );
  FA_340 FAI_45 ( .A(A[44]), .B(B[44]), .Ci(CTMP[44]), .S(S[44]), .Co(CTMP[45]) );
  FA_339 FAI_46 ( .A(A[45]), .B(B[45]), .Ci(CTMP[45]), .S(S[45]), .Co(CTMP[46]) );
  FA_338 FAI_47 ( .A(A[46]), .B(B[46]), .Ci(CTMP[46]), .S(S[46]), .Co(CTMP[47]) );
  FA_337 FAI_48 ( .A(A[47]), .B(B[47]), .Ci(CTMP[47]), .S(S[47]), .Co(CTMP[48]) );
  FA_336 FAI_49 ( .A(A[48]), .B(B[48]), .Ci(CTMP[48]), .S(S[48]), .Co(CTMP[49]) );
  FA_335 FAI_50 ( .A(A[49]), .B(B[49]), .Ci(CTMP[49]), .S(S[49]), .Co(CTMP[50]) );
  FA_334 FAI_51 ( .A(A[50]), .B(B[50]), .Ci(CTMP[50]), .S(S[50]), .Co(CTMP[51]) );
  FA_333 FAI_52 ( .A(A[51]), .B(B[51]), .Ci(CTMP[51]), .S(S[51]), .Co(CTMP[52]) );
  FA_332 FAI_53 ( .A(A[52]), .B(B[52]), .Ci(CTMP[52]), .S(S[52]), .Co(CTMP[53]) );
  FA_331 FAI_54 ( .A(A[53]), .B(B[53]), .Ci(CTMP[53]), .S(S[53]), .Co(CTMP[54]) );
  FA_330 FAI_55 ( .A(A[54]), .B(B[54]), .Ci(CTMP[54]), .S(S[54]), .Co(CTMP[55]) );
  FA_329 FAI_56 ( .A(A[55]), .B(B[55]), .Ci(CTMP[55]), .S(S[55]), .Co(CTMP[56]) );
  FA_328 FAI_57 ( .A(A[56]), .B(B[56]), .Ci(CTMP[56]), .S(S[56]), .Co(CTMP[57]) );
  FA_327 FAI_58 ( .A(A[57]), .B(B[57]), .Ci(CTMP[57]), .S(S[57]), .Co(CTMP[58]) );
  FA_326 FAI_59 ( .A(A[58]), .B(B[58]), .Ci(CTMP[58]), .S(S[58]), .Co(CTMP[59]) );
  FA_325 FAI_60 ( .A(A[59]), .B(B[59]), .Ci(CTMP[59]), .S(S[59]), .Co(CTMP[60]) );
  FA_324 FAI_61 ( .A(A[60]), .B(B[60]), .Ci(CTMP[60]), .S(S[60]), .Co(CTMP[61]) );
  FA_323 FAI_62 ( .A(A[61]), .B(B[61]), .Ci(CTMP[61]), .S(S[61]), .Co(CTMP[62]) );
  FA_322 FAI_63 ( .A(A[62]), .B(B[62]), .Ci(CTMP[62]), .S(S[62]), .Co(CTMP[63]) );
  FA_321 FAI_64 ( .A(A[63]), .B(B[63]), .Ci(CTMP[63]), .S(S[63]), .Co(Co) );
endmodule


module booth_mul_row_N64_RADIX3_6 ( prevA, prevSum, encoderIn, nextA, nextSum
 );
  input [63:0] prevA;
  input [63:0] prevSum;
  input [2:0] encoderIn;
  output [63:0] nextA;
  output [63:0] nextSum;

  wire   [2:0] encoder_to_mux;
  wire   [63:0] plus2A_s;
  wire   [63:0] minus2A_s;
  wire   [63:0] minus4A_s;
  tri   [63:0] mux_to_adder;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign nextA[0] = 1'b0;

  encoder_N64_RADIX3_6 encoder_1 ( .X(encoderIn), .Z(encoder_to_mux) );
  ShiftnCompl_N64_6 ShiftnCompl_1 ( .plusA(prevA), .plus2A_out({plus2A_s[63:1], 
        SYNOPSYS_UNCONNECTED__0}), .minus2A_out(minus2A_s), .plus4A_out({
        nextA[63:1], SYNOPSYS_UNCONNECTED__1}), .minus4A_out(minus4A_s) );
  MUX_GENERIC_N64_RADIX3_6 mux_1 ( .plusA({plus2A_s[63:1], 1'b0}), .minusA(
        minus2A_s), .plus2A({nextA[63:1], 1'b0}), .minus2A(minus4A_s), .SEL(
        encoder_to_mux), .Y(mux_to_adder) );
  RCA_N64_6 rca_1 ( .A(mux_to_adder), .B(prevSum), .Ci(1'b0), .S(nextSum) );
endmodule


module encoder_N64_RADIX3_5 ( X, Z );
  input [2:0] X;
  output [2:0] Z;
  wire   n5, n7, n8;

  OAI22_X1 U1 ( .A1(n8), .A2(n5), .B1(X[2]), .B2(n7), .ZN(Z[1]) );
  INV_X1 U2 ( .A(X[2]), .ZN(n5) );
  AOI21_X1 U3 ( .B1(n8), .B2(n7), .A(X[2]), .ZN(Z[0]) );
  OAI21_X1 U4 ( .B1(X[1]), .B2(X[0]), .A(n7), .ZN(n8) );
  AND3_X1 U5 ( .A1(X[2]), .A2(n7), .A3(n8), .ZN(Z[2]) );
  NAND2_X1 U6 ( .A1(X[1]), .A2(X[0]), .ZN(n7) );
endmodule


module shifter_N64_10 ( \input , shiftLeftOnePos );
  input [63:0] \input ;
  output [63:0] shiftLeftOnePos;
  wire   \input[62] , \input[61] , \input[60] , \input[59] , \input[58] ,
         \input[57] , \input[56] , \input[55] , \input[54] , \input[53] ,
         \input[52] , \input[51] , \input[50] , \input[49] , \input[48] ,
         \input[47] , \input[46] , \input[45] , \input[44] , \input[43] ,
         \input[42] , \input[41] , \input[40] , \input[39] , \input[38] ,
         \input[37] , \input[36] , \input[35] , \input[34] , \input[33] ,
         \input[32] , \input[31] , \input[30] , \input[29] , \input[28] ,
         \input[27] , \input[26] , \input[25] , \input[24] , \input[23] ,
         \input[22] , \input[21] , \input[20] , \input[19] , \input[18] ,
         \input[17] , \input[16] , \input[15] , \input[14] , \input[13] ,
         \input[12] , \input[11] , \input[10] , \input[9] , \input[8] ,
         \input[7] , \input[6] , \input[5] , \input[4] , \input[3] ,
         \input[2] , \input[1] , \input[0] ;
  assign shiftLeftOnePos[0] = 1'b0;
  assign shiftLeftOnePos[63] = \input[62] ;
  assign \input[62]  = \input  [62];
  assign shiftLeftOnePos[62] = \input[61] ;
  assign \input[61]  = \input  [61];
  assign shiftLeftOnePos[61] = \input[60] ;
  assign \input[60]  = \input  [60];
  assign shiftLeftOnePos[60] = \input[59] ;
  assign \input[59]  = \input  [59];
  assign shiftLeftOnePos[59] = \input[58] ;
  assign \input[58]  = \input  [58];
  assign shiftLeftOnePos[58] = \input[57] ;
  assign \input[57]  = \input  [57];
  assign shiftLeftOnePos[57] = \input[56] ;
  assign \input[56]  = \input  [56];
  assign shiftLeftOnePos[56] = \input[55] ;
  assign \input[55]  = \input  [55];
  assign shiftLeftOnePos[55] = \input[54] ;
  assign \input[54]  = \input  [54];
  assign shiftLeftOnePos[54] = \input[53] ;
  assign \input[53]  = \input  [53];
  assign shiftLeftOnePos[53] = \input[52] ;
  assign \input[52]  = \input  [52];
  assign shiftLeftOnePos[52] = \input[51] ;
  assign \input[51]  = \input  [51];
  assign shiftLeftOnePos[51] = \input[50] ;
  assign \input[50]  = \input  [50];
  assign shiftLeftOnePos[50] = \input[49] ;
  assign \input[49]  = \input  [49];
  assign shiftLeftOnePos[49] = \input[48] ;
  assign \input[48]  = \input  [48];
  assign shiftLeftOnePos[48] = \input[47] ;
  assign \input[47]  = \input  [47];
  assign shiftLeftOnePos[47] = \input[46] ;
  assign \input[46]  = \input  [46];
  assign shiftLeftOnePos[46] = \input[45] ;
  assign \input[45]  = \input  [45];
  assign shiftLeftOnePos[45] = \input[44] ;
  assign \input[44]  = \input  [44];
  assign shiftLeftOnePos[44] = \input[43] ;
  assign \input[43]  = \input  [43];
  assign shiftLeftOnePos[43] = \input[42] ;
  assign \input[42]  = \input  [42];
  assign shiftLeftOnePos[42] = \input[41] ;
  assign \input[41]  = \input  [41];
  assign shiftLeftOnePos[41] = \input[40] ;
  assign \input[40]  = \input  [40];
  assign shiftLeftOnePos[40] = \input[39] ;
  assign \input[39]  = \input  [39];
  assign shiftLeftOnePos[39] = \input[38] ;
  assign \input[38]  = \input  [38];
  assign shiftLeftOnePos[38] = \input[37] ;
  assign \input[37]  = \input  [37];
  assign shiftLeftOnePos[37] = \input[36] ;
  assign \input[36]  = \input  [36];
  assign shiftLeftOnePos[36] = \input[35] ;
  assign \input[35]  = \input  [35];
  assign shiftLeftOnePos[35] = \input[34] ;
  assign \input[34]  = \input  [34];
  assign shiftLeftOnePos[34] = \input[33] ;
  assign \input[33]  = \input  [33];
  assign shiftLeftOnePos[33] = \input[32] ;
  assign \input[32]  = \input  [32];
  assign shiftLeftOnePos[32] = \input[31] ;
  assign \input[31]  = \input  [31];
  assign shiftLeftOnePos[31] = \input[30] ;
  assign \input[30]  = \input  [30];
  assign shiftLeftOnePos[30] = \input[29] ;
  assign \input[29]  = \input  [29];
  assign shiftLeftOnePos[29] = \input[28] ;
  assign \input[28]  = \input  [28];
  assign shiftLeftOnePos[28] = \input[27] ;
  assign \input[27]  = \input  [27];
  assign shiftLeftOnePos[27] = \input[26] ;
  assign \input[26]  = \input  [26];
  assign shiftLeftOnePos[26] = \input[25] ;
  assign \input[25]  = \input  [25];
  assign shiftLeftOnePos[25] = \input[24] ;
  assign \input[24]  = \input  [24];
  assign shiftLeftOnePos[24] = \input[23] ;
  assign \input[23]  = \input  [23];
  assign shiftLeftOnePos[23] = \input[22] ;
  assign \input[22]  = \input  [22];
  assign shiftLeftOnePos[22] = \input[21] ;
  assign \input[21]  = \input  [21];
  assign shiftLeftOnePos[21] = \input[20] ;
  assign \input[20]  = \input  [20];
  assign shiftLeftOnePos[20] = \input[19] ;
  assign \input[19]  = \input  [19];
  assign shiftLeftOnePos[19] = \input[18] ;
  assign \input[18]  = \input  [18];
  assign shiftLeftOnePos[18] = \input[17] ;
  assign \input[17]  = \input  [17];
  assign shiftLeftOnePos[17] = \input[16] ;
  assign \input[16]  = \input  [16];
  assign shiftLeftOnePos[16] = \input[15] ;
  assign \input[15]  = \input  [15];
  assign shiftLeftOnePos[15] = \input[14] ;
  assign \input[14]  = \input  [14];
  assign shiftLeftOnePos[14] = \input[13] ;
  assign \input[13]  = \input  [13];
  assign shiftLeftOnePos[13] = \input[12] ;
  assign \input[12]  = \input  [12];
  assign shiftLeftOnePos[12] = \input[11] ;
  assign \input[11]  = \input  [11];
  assign shiftLeftOnePos[11] = \input[10] ;
  assign \input[10]  = \input  [10];
  assign shiftLeftOnePos[10] = \input[9] ;
  assign \input[9]  = \input  [9];
  assign shiftLeftOnePos[9] = \input[8] ;
  assign \input[8]  = \input  [8];
  assign shiftLeftOnePos[8] = \input[7] ;
  assign \input[7]  = \input  [7];
  assign shiftLeftOnePos[7] = \input[6] ;
  assign \input[6]  = \input  [6];
  assign shiftLeftOnePos[6] = \input[5] ;
  assign \input[5]  = \input  [5];
  assign shiftLeftOnePos[5] = \input[4] ;
  assign \input[4]  = \input  [4];
  assign shiftLeftOnePos[4] = \input[3] ;
  assign \input[3]  = \input  [3];
  assign shiftLeftOnePos[3] = \input[2] ;
  assign \input[2]  = \input  [2];
  assign shiftLeftOnePos[2] = \input[1] ;
  assign \input[1]  = \input  [1];
  assign shiftLeftOnePos[1] = \input[0] ;
  assign \input[0]  = \input  [0];

endmodule


module shifter_N64_9 ( \input , shiftLeftOnePos );
  input [63:0] \input ;
  output [63:0] shiftLeftOnePos;
  wire   \input[62] , \input[61] , \input[60] , \input[59] , \input[58] ,
         \input[57] , \input[56] , \input[55] , \input[54] , \input[53] ,
         \input[52] , \input[51] , \input[50] , \input[49] , \input[48] ,
         \input[47] , \input[46] , \input[45] , \input[44] , \input[43] ,
         \input[42] , \input[41] , \input[40] , \input[39] , \input[38] ,
         \input[37] , \input[36] , \input[35] , \input[34] , \input[33] ,
         \input[32] , \input[31] , \input[30] , \input[29] , \input[28] ,
         \input[27] , \input[26] , \input[25] , \input[24] , \input[23] ,
         \input[22] , \input[21] , \input[20] , \input[19] , \input[18] ,
         \input[17] , \input[16] , \input[15] , \input[14] , \input[13] ,
         \input[12] , \input[11] , \input[10] , \input[9] , \input[8] ,
         \input[7] , \input[6] , \input[5] , \input[4] , \input[3] ,
         \input[2] , \input[1] , \input[0] ;
  assign shiftLeftOnePos[0] = 1'b0;
  assign shiftLeftOnePos[63] = \input[62] ;
  assign \input[62]  = \input  [62];
  assign shiftLeftOnePos[62] = \input[61] ;
  assign \input[61]  = \input  [61];
  assign shiftLeftOnePos[61] = \input[60] ;
  assign \input[60]  = \input  [60];
  assign shiftLeftOnePos[60] = \input[59] ;
  assign \input[59]  = \input  [59];
  assign shiftLeftOnePos[59] = \input[58] ;
  assign \input[58]  = \input  [58];
  assign shiftLeftOnePos[58] = \input[57] ;
  assign \input[57]  = \input  [57];
  assign shiftLeftOnePos[57] = \input[56] ;
  assign \input[56]  = \input  [56];
  assign shiftLeftOnePos[56] = \input[55] ;
  assign \input[55]  = \input  [55];
  assign shiftLeftOnePos[55] = \input[54] ;
  assign \input[54]  = \input  [54];
  assign shiftLeftOnePos[54] = \input[53] ;
  assign \input[53]  = \input  [53];
  assign shiftLeftOnePos[53] = \input[52] ;
  assign \input[52]  = \input  [52];
  assign shiftLeftOnePos[52] = \input[51] ;
  assign \input[51]  = \input  [51];
  assign shiftLeftOnePos[51] = \input[50] ;
  assign \input[50]  = \input  [50];
  assign shiftLeftOnePos[50] = \input[49] ;
  assign \input[49]  = \input  [49];
  assign shiftLeftOnePos[49] = \input[48] ;
  assign \input[48]  = \input  [48];
  assign shiftLeftOnePos[48] = \input[47] ;
  assign \input[47]  = \input  [47];
  assign shiftLeftOnePos[47] = \input[46] ;
  assign \input[46]  = \input  [46];
  assign shiftLeftOnePos[46] = \input[45] ;
  assign \input[45]  = \input  [45];
  assign shiftLeftOnePos[45] = \input[44] ;
  assign \input[44]  = \input  [44];
  assign shiftLeftOnePos[44] = \input[43] ;
  assign \input[43]  = \input  [43];
  assign shiftLeftOnePos[43] = \input[42] ;
  assign \input[42]  = \input  [42];
  assign shiftLeftOnePos[42] = \input[41] ;
  assign \input[41]  = \input  [41];
  assign shiftLeftOnePos[41] = \input[40] ;
  assign \input[40]  = \input  [40];
  assign shiftLeftOnePos[40] = \input[39] ;
  assign \input[39]  = \input  [39];
  assign shiftLeftOnePos[39] = \input[38] ;
  assign \input[38]  = \input  [38];
  assign shiftLeftOnePos[38] = \input[37] ;
  assign \input[37]  = \input  [37];
  assign shiftLeftOnePos[37] = \input[36] ;
  assign \input[36]  = \input  [36];
  assign shiftLeftOnePos[36] = \input[35] ;
  assign \input[35]  = \input  [35];
  assign shiftLeftOnePos[35] = \input[34] ;
  assign \input[34]  = \input  [34];
  assign shiftLeftOnePos[34] = \input[33] ;
  assign \input[33]  = \input  [33];
  assign shiftLeftOnePos[33] = \input[32] ;
  assign \input[32]  = \input  [32];
  assign shiftLeftOnePos[32] = \input[31] ;
  assign \input[31]  = \input  [31];
  assign shiftLeftOnePos[31] = \input[30] ;
  assign \input[30]  = \input  [30];
  assign shiftLeftOnePos[30] = \input[29] ;
  assign \input[29]  = \input  [29];
  assign shiftLeftOnePos[29] = \input[28] ;
  assign \input[28]  = \input  [28];
  assign shiftLeftOnePos[28] = \input[27] ;
  assign \input[27]  = \input  [27];
  assign shiftLeftOnePos[27] = \input[26] ;
  assign \input[26]  = \input  [26];
  assign shiftLeftOnePos[26] = \input[25] ;
  assign \input[25]  = \input  [25];
  assign shiftLeftOnePos[25] = \input[24] ;
  assign \input[24]  = \input  [24];
  assign shiftLeftOnePos[24] = \input[23] ;
  assign \input[23]  = \input  [23];
  assign shiftLeftOnePos[23] = \input[22] ;
  assign \input[22]  = \input  [22];
  assign shiftLeftOnePos[22] = \input[21] ;
  assign \input[21]  = \input  [21];
  assign shiftLeftOnePos[21] = \input[20] ;
  assign \input[20]  = \input  [20];
  assign shiftLeftOnePos[20] = \input[19] ;
  assign \input[19]  = \input  [19];
  assign shiftLeftOnePos[19] = \input[18] ;
  assign \input[18]  = \input  [18];
  assign shiftLeftOnePos[18] = \input[17] ;
  assign \input[17]  = \input  [17];
  assign shiftLeftOnePos[17] = \input[16] ;
  assign \input[16]  = \input  [16];
  assign shiftLeftOnePos[16] = \input[15] ;
  assign \input[15]  = \input  [15];
  assign shiftLeftOnePos[15] = \input[14] ;
  assign \input[14]  = \input  [14];
  assign shiftLeftOnePos[14] = \input[13] ;
  assign \input[13]  = \input  [13];
  assign shiftLeftOnePos[13] = \input[12] ;
  assign \input[12]  = \input  [12];
  assign shiftLeftOnePos[12] = \input[11] ;
  assign \input[11]  = \input  [11];
  assign shiftLeftOnePos[11] = \input[10] ;
  assign \input[10]  = \input  [10];
  assign shiftLeftOnePos[10] = \input[9] ;
  assign \input[9]  = \input  [9];
  assign shiftLeftOnePos[9] = \input[8] ;
  assign \input[8]  = \input  [8];
  assign shiftLeftOnePos[8] = \input[7] ;
  assign \input[7]  = \input  [7];
  assign shiftLeftOnePos[7] = \input[6] ;
  assign \input[6]  = \input  [6];
  assign shiftLeftOnePos[6] = \input[5] ;
  assign \input[5]  = \input  [5];
  assign shiftLeftOnePos[5] = \input[4] ;
  assign \input[4]  = \input  [4];
  assign shiftLeftOnePos[4] = \input[3] ;
  assign \input[3]  = \input  [3];
  assign shiftLeftOnePos[3] = \input[2] ;
  assign \input[2]  = \input  [2];
  assign shiftLeftOnePos[2] = \input[1] ;
  assign \input[1]  = \input  [1];
  assign shiftLeftOnePos[1] = \input[0] ;
  assign \input[0]  = \input  [0];

endmodule


module complementer_N64_10_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n190, n191, n192, n193, n194, n196, n197, n198, n199, n200,
         n202, n203, n204, n206, n207, n208, n210, n211, n212, n213, n214,
         n216, n217, n218, n220, n221, n222, n224, n225, n226, n228, n229,
         n230, n232, n233, n234, n235, n237, n238, n239, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n189, n195, n201,
         n205, n209, n215, n219, n223, n227, n231, n236, n240;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U81 ( .A(n190), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U82 ( .A(n192), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U83 ( .A(n193), .B(B[6]), .Z(DIFF[6]) );
  XOR2_X1 U85 ( .A(n196), .B(B[62]), .Z(DIFF[62]) );
  XOR2_X1 U86 ( .A(n194), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U87 ( .A(n198), .B(B[59]), .Z(DIFF[59]) );
  XOR2_X1 U89 ( .A(n200), .B(B[57]), .Z(DIFF[57]) );
  XOR2_X1 U90 ( .A(n202), .B(B[55]), .Z(DIFF[55]) );
  XOR2_X1 U92 ( .A(n204), .B(B[53]), .Z(DIFF[53]) );
  XOR2_X1 U93 ( .A(n206), .B(B[51]), .Z(DIFF[51]) );
  XOR2_X1 U95 ( .A(n208), .B(B[49]), .Z(DIFF[49]) );
  XOR2_X1 U96 ( .A(n212), .B(B[47]), .Z(DIFF[47]) );
  XOR2_X1 U98 ( .A(n214), .B(B[45]), .Z(DIFF[45]) );
  XOR2_X1 U99 ( .A(n216), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U101 ( .A(n218), .B(B[41]), .Z(DIFF[41]) );
  XOR2_X1 U102 ( .A(n211), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U103 ( .A(n220), .B(B[39]), .Z(DIFF[39]) );
  XOR2_X1 U105 ( .A(n222), .B(B[37]), .Z(DIFF[37]) );
  XOR2_X1 U106 ( .A(n224), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U108 ( .A(n226), .B(B[33]), .Z(DIFF[33]) );
  XOR2_X1 U109 ( .A(n228), .B(B[31]), .Z(DIFF[31]) );
  XOR2_X1 U111 ( .A(n230), .B(B[29]), .Z(DIFF[29]) );
  XOR2_X1 U112 ( .A(n233), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U114 ( .A(n235), .B(B[25]), .Z(DIFF[25]) );
  XOR2_X1 U115 ( .A(n237), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U117 ( .A(n239), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U118 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U119 ( .A(n241), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U120 ( .A(n244), .B(B[18]), .Z(DIFF[18]) );
  XOR2_X1 U121 ( .A(n243), .B(B[17]), .Z(DIFF[17]) );
  XOR2_X1 U122 ( .A(n245), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U123 ( .A(n248), .B(B[14]), .Z(DIFF[14]) );
  XOR2_X1 U124 ( .A(n247), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U125 ( .A(n249), .B(B[11]), .Z(DIFF[11]) );
  XOR2_X1 U126 ( .A(n251), .B(B[10]), .Z(DIFF[10]) );
  NOR3_X1 U1 ( .A1(B[59]), .A2(B[60]), .A3(n198), .ZN(n197) );
  XNOR2_X1 U2 ( .A(B[60]), .B(n199), .ZN(DIFF[60]) );
  NOR2_X1 U3 ( .A1(B[59]), .A2(n198), .ZN(n199) );
  XOR2_X1 U4 ( .A(n197), .B(n240), .Z(DIFF[61]) );
  NAND2_X1 U5 ( .A1(n197), .A2(n240), .ZN(n196) );
  XNOR2_X1 U6 ( .A(n189), .B(B[63]), .ZN(DIFF[63]) );
  NOR2_X1 U7 ( .A1(n196), .A2(B[62]), .ZN(n189) );
  XNOR2_X1 U8 ( .A(B[56]), .B(n203), .ZN(DIFF[56]) );
  NOR2_X1 U9 ( .A1(B[55]), .A2(n202), .ZN(n203) );
  OR3_X1 U10 ( .A1(B[57]), .A2(B[58]), .A3(n200), .ZN(n198) );
  OR3_X1 U11 ( .A1(B[53]), .A2(B[54]), .A3(n204), .ZN(n202) );
  OR3_X1 U12 ( .A1(B[55]), .A2(B[56]), .A3(n202), .ZN(n200) );
  XNOR2_X1 U13 ( .A(n195), .B(B[58]), .ZN(DIFF[58]) );
  NOR2_X1 U14 ( .A1(n200), .A2(B[57]), .ZN(n195) );
  XNOR2_X1 U15 ( .A(n201), .B(B[54]), .ZN(DIFF[54]) );
  NOR2_X1 U16 ( .A1(n204), .A2(B[53]), .ZN(n201) );
  XNOR2_X1 U17 ( .A(B[40]), .B(n221), .ZN(DIFF[40]) );
  NOR2_X1 U18 ( .A1(B[39]), .A2(n220), .ZN(n221) );
  XNOR2_X1 U19 ( .A(B[36]), .B(n225), .ZN(DIFF[36]) );
  NOR2_X1 U20 ( .A1(B[35]), .A2(n224), .ZN(n225) );
  XNOR2_X1 U21 ( .A(B[32]), .B(n229), .ZN(DIFF[32]) );
  NOR2_X1 U22 ( .A1(B[31]), .A2(n228), .ZN(n229) );
  OR3_X1 U23 ( .A1(B[33]), .A2(B[34]), .A3(n226), .ZN(n224) );
  OR3_X1 U24 ( .A1(B[37]), .A2(B[38]), .A3(n222), .ZN(n220) );
  OR3_X1 U25 ( .A1(B[31]), .A2(B[32]), .A3(n228), .ZN(n226) );
  OR3_X1 U26 ( .A1(B[35]), .A2(B[36]), .A3(n224), .ZN(n222) );
  OR3_X1 U27 ( .A1(B[39]), .A2(B[40]), .A3(n220), .ZN(n218) );
  XNOR2_X1 U28 ( .A(n205), .B(B[38]), .ZN(DIFF[38]) );
  NOR2_X1 U29 ( .A1(n222), .A2(B[37]), .ZN(n205) );
  XNOR2_X1 U30 ( .A(n209), .B(B[34]), .ZN(DIFF[34]) );
  NOR2_X1 U31 ( .A1(n226), .A2(B[33]), .ZN(n209) );
  XNOR2_X1 U32 ( .A(B[52]), .B(n207), .ZN(DIFF[52]) );
  NOR2_X1 U33 ( .A1(B[51]), .A2(n206), .ZN(n207) );
  XNOR2_X1 U34 ( .A(B[48]), .B(n213), .ZN(DIFF[48]) );
  NOR2_X1 U35 ( .A1(B[47]), .A2(n212), .ZN(n213) );
  XNOR2_X1 U36 ( .A(B[44]), .B(n217), .ZN(DIFF[44]) );
  NOR2_X1 U37 ( .A1(B[43]), .A2(n216), .ZN(n217) );
  OR3_X1 U38 ( .A1(B[41]), .A2(B[42]), .A3(n218), .ZN(n216) );
  OR3_X1 U39 ( .A1(B[45]), .A2(B[46]), .A3(n214), .ZN(n212) );
  OR3_X1 U40 ( .A1(B[49]), .A2(B[50]), .A3(n208), .ZN(n206) );
  OR3_X1 U41 ( .A1(B[43]), .A2(B[44]), .A3(n216), .ZN(n214) );
  OR3_X1 U42 ( .A1(B[47]), .A2(B[48]), .A3(n212), .ZN(n208) );
  OR3_X1 U43 ( .A1(B[51]), .A2(B[52]), .A3(n206), .ZN(n204) );
  XNOR2_X1 U44 ( .A(n215), .B(B[50]), .ZN(DIFF[50]) );
  NOR2_X1 U45 ( .A1(n208), .A2(B[49]), .ZN(n215) );
  XNOR2_X1 U46 ( .A(n219), .B(B[46]), .ZN(DIFF[46]) );
  NOR2_X1 U47 ( .A1(n214), .A2(B[45]), .ZN(n219) );
  XNOR2_X1 U48 ( .A(n223), .B(B[42]), .ZN(DIFF[42]) );
  NOR2_X1 U49 ( .A1(n218), .A2(B[41]), .ZN(n223) );
  OR3_X1 U50 ( .A1(B[29]), .A2(B[30]), .A3(n230), .ZN(n228) );
  XNOR2_X1 U51 ( .A(n227), .B(B[30]), .ZN(DIFF[30]) );
  NOR2_X1 U52 ( .A1(n230), .A2(B[29]), .ZN(n227) );
  XNOR2_X1 U53 ( .A(B[28]), .B(n234), .ZN(DIFF[28]) );
  NOR2_X1 U54 ( .A1(B[27]), .A2(n233), .ZN(n234) );
  OR3_X1 U55 ( .A1(B[27]), .A2(B[28]), .A3(n233), .ZN(n230) );
  OR3_X1 U56 ( .A1(B[25]), .A2(B[26]), .A3(n235), .ZN(n233) );
  XNOR2_X1 U57 ( .A(n231), .B(B[26]), .ZN(DIFF[26]) );
  NOR2_X1 U58 ( .A1(n235), .A2(B[25]), .ZN(n231) );
  XNOR2_X1 U59 ( .A(B[24]), .B(n238), .ZN(DIFF[24]) );
  NOR2_X1 U60 ( .A1(B[23]), .A2(n237), .ZN(n238) );
  OR3_X1 U61 ( .A1(B[23]), .A2(B[24]), .A3(n237), .ZN(n235) );
  XNOR2_X1 U62 ( .A(n236), .B(B[22]), .ZN(DIFF[22]) );
  NOR2_X1 U63 ( .A1(n239), .A2(B[21]), .ZN(n236) );
  OR3_X1 U64 ( .A1(B[21]), .A2(B[22]), .A3(n239), .ZN(n237) );
  NOR2_X1 U65 ( .A1(B[19]), .A2(n241), .ZN(n242) );
  NOR2_X1 U66 ( .A1(B[15]), .A2(n245), .ZN(n246) );
  NOR2_X1 U67 ( .A1(B[11]), .A2(n249), .ZN(n250) );
  NOR2_X1 U68 ( .A1(B[7]), .A2(n192), .ZN(n191) );
  NOR2_X1 U69 ( .A1(B[3]), .A2(n211), .ZN(n210) );
  OR3_X1 U70 ( .A1(B[17]), .A2(B[18]), .A3(n243), .ZN(n241) );
  OR3_X1 U71 ( .A1(B[13]), .A2(B[14]), .A3(n247), .ZN(n245) );
  OR3_X1 U72 ( .A1(B[10]), .A2(B[9]), .A3(n190), .ZN(n249) );
  OR3_X1 U73 ( .A1(B[5]), .A2(B[6]), .A3(n194), .ZN(n192) );
  OR3_X1 U74 ( .A1(B[19]), .A2(B[20]), .A3(n241), .ZN(n239) );
  OR3_X1 U75 ( .A1(B[15]), .A2(B[16]), .A3(n245), .ZN(n243) );
  OR3_X1 U76 ( .A1(B[11]), .A2(B[12]), .A3(n249), .ZN(n247) );
  OR3_X1 U77 ( .A1(B[7]), .A2(B[8]), .A3(n192), .ZN(n190) );
  OR3_X1 U78 ( .A1(B[3]), .A2(B[4]), .A3(n211), .ZN(n194) );
  XNOR2_X1 U79 ( .A(B[20]), .B(n242), .ZN(DIFF[20]) );
  XNOR2_X1 U80 ( .A(B[16]), .B(n246), .ZN(DIFF[16]) );
  XNOR2_X1 U84 ( .A(B[12]), .B(n250), .ZN(DIFF[12]) );
  XNOR2_X1 U88 ( .A(B[8]), .B(n191), .ZN(DIFF[8]) );
  XNOR2_X1 U91 ( .A(B[4]), .B(n210), .ZN(DIFF[4]) );
  XNOR2_X1 U94 ( .A(B[2]), .B(n232), .ZN(DIFF[2]) );
  OR2_X1 U97 ( .A1(n243), .A2(B[17]), .ZN(n244) );
  OR2_X1 U100 ( .A1(n247), .A2(B[13]), .ZN(n248) );
  OR2_X1 U104 ( .A1(n190), .A2(B[9]), .ZN(n251) );
  OR2_X1 U107 ( .A1(n194), .A2(B[5]), .ZN(n193) );
  OR3_X1 U110 ( .A1(B[1]), .A2(B[2]), .A3(\B[0] ), .ZN(n211) );
  NOR2_X1 U113 ( .A1(\B[0] ), .A2(B[1]), .ZN(n232) );
  INV_X1 U116 ( .A(B[61]), .ZN(n240) );
endmodule


module complementer_N64_10 ( \input , complement2 );
  input [63:0] \input ;
  output [63:0] complement2;


  complementer_N64_10_DW01_sub_0 sub_add_31_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(\input ), .CI(1'b0), .DIFF(complement2) );
endmodule


module complementer_N64_9_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n190, n191, n192, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n245,
         n246, n247, n249, n250, n189, n193, n244, n248, n251;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U81 ( .A(n190), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U82 ( .A(n192), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U84 ( .A(n195), .B(B[63]), .Z(DIFF[63]) );
  XOR2_X1 U85 ( .A(n196), .B(B[62]), .Z(DIFF[62]) );
  XOR2_X1 U86 ( .A(n194), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U87 ( .A(n198), .B(B[59]), .Z(DIFF[59]) );
  XOR2_X1 U88 ( .A(n201), .B(B[58]), .Z(DIFF[58]) );
  XOR2_X1 U89 ( .A(n200), .B(B[57]), .Z(DIFF[57]) );
  XOR2_X1 U90 ( .A(n202), .B(B[55]), .Z(DIFF[55]) );
  XOR2_X1 U91 ( .A(n205), .B(B[54]), .Z(DIFF[54]) );
  XOR2_X1 U92 ( .A(n204), .B(B[53]), .Z(DIFF[53]) );
  XOR2_X1 U93 ( .A(n206), .B(B[51]), .Z(DIFF[51]) );
  XOR2_X1 U94 ( .A(n209), .B(B[50]), .Z(DIFF[50]) );
  XOR2_X1 U95 ( .A(n208), .B(B[49]), .Z(DIFF[49]) );
  XOR2_X1 U96 ( .A(n212), .B(B[47]), .Z(DIFF[47]) );
  XOR2_X1 U97 ( .A(n215), .B(B[46]), .Z(DIFF[46]) );
  XOR2_X1 U98 ( .A(n214), .B(B[45]), .Z(DIFF[45]) );
  XOR2_X1 U99 ( .A(n216), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U100 ( .A(n219), .B(B[42]), .Z(DIFF[42]) );
  XOR2_X1 U101 ( .A(n218), .B(B[41]), .Z(DIFF[41]) );
  XOR2_X1 U102 ( .A(n211), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U103 ( .A(n220), .B(B[39]), .Z(DIFF[39]) );
  XOR2_X1 U104 ( .A(n223), .B(B[38]), .Z(DIFF[38]) );
  XOR2_X1 U105 ( .A(n222), .B(B[37]), .Z(DIFF[37]) );
  XOR2_X1 U106 ( .A(n224), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U107 ( .A(n227), .B(B[34]), .Z(DIFF[34]) );
  XOR2_X1 U108 ( .A(n226), .B(B[33]), .Z(DIFF[33]) );
  XOR2_X1 U109 ( .A(n228), .B(B[31]), .Z(DIFF[31]) );
  XOR2_X1 U110 ( .A(n231), .B(B[30]), .Z(DIFF[30]) );
  XOR2_X1 U111 ( .A(n230), .B(B[29]), .Z(DIFF[29]) );
  XOR2_X1 U112 ( .A(n233), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U113 ( .A(n236), .B(B[26]), .Z(DIFF[26]) );
  XOR2_X1 U114 ( .A(n235), .B(B[25]), .Z(DIFF[25]) );
  XOR2_X1 U115 ( .A(n237), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U116 ( .A(n240), .B(B[22]), .Z(DIFF[22]) );
  XOR2_X1 U117 ( .A(n239), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U118 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U119 ( .A(n241), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U121 ( .A(n243), .B(B[17]), .Z(DIFF[17]) );
  XOR2_X1 U122 ( .A(n245), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U124 ( .A(n247), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U125 ( .A(n249), .B(B[11]), .Z(DIFF[11]) );
  NAND2_X1 U1 ( .A1(n197), .A2(n251), .ZN(n196) );
  NOR3_X1 U2 ( .A1(B[59]), .A2(B[60]), .A3(n198), .ZN(n197) );
  NOR2_X1 U3 ( .A1(B[59]), .A2(n198), .ZN(n199) );
  NOR2_X1 U4 ( .A1(B[55]), .A2(n202), .ZN(n203) );
  OR3_X1 U5 ( .A1(B[57]), .A2(B[58]), .A3(n200), .ZN(n198) );
  OR3_X1 U6 ( .A1(B[55]), .A2(B[56]), .A3(n202), .ZN(n200) );
  OR2_X1 U7 ( .A1(n200), .A2(B[57]), .ZN(n201) );
  OR2_X1 U8 ( .A1(n196), .A2(B[62]), .ZN(n195) );
  NOR2_X1 U9 ( .A1(B[35]), .A2(n224), .ZN(n225) );
  NOR2_X1 U10 ( .A1(B[31]), .A2(n228), .ZN(n229) );
  OR3_X1 U11 ( .A1(B[33]), .A2(B[34]), .A3(n226), .ZN(n224) );
  OR3_X1 U12 ( .A1(B[35]), .A2(B[36]), .A3(n224), .ZN(n222) );
  OR3_X1 U13 ( .A1(B[31]), .A2(B[32]), .A3(n228), .ZN(n226) );
  OR2_X1 U14 ( .A1(n222), .A2(B[37]), .ZN(n223) );
  OR2_X1 U15 ( .A1(n226), .A2(B[33]), .ZN(n227) );
  NOR2_X1 U16 ( .A1(B[51]), .A2(n206), .ZN(n207) );
  NOR2_X1 U17 ( .A1(B[47]), .A2(n212), .ZN(n213) );
  NOR2_X1 U18 ( .A1(B[43]), .A2(n216), .ZN(n217) );
  NOR2_X1 U19 ( .A1(B[39]), .A2(n220), .ZN(n221) );
  OR3_X1 U20 ( .A1(B[53]), .A2(B[54]), .A3(n204), .ZN(n202) );
  OR3_X1 U21 ( .A1(B[49]), .A2(B[50]), .A3(n208), .ZN(n206) );
  OR3_X1 U22 ( .A1(B[45]), .A2(B[46]), .A3(n214), .ZN(n212) );
  OR3_X1 U23 ( .A1(B[41]), .A2(B[42]), .A3(n218), .ZN(n216) );
  OR3_X1 U24 ( .A1(B[37]), .A2(B[38]), .A3(n222), .ZN(n220) );
  OR3_X1 U25 ( .A1(B[51]), .A2(B[52]), .A3(n206), .ZN(n204) );
  OR3_X1 U26 ( .A1(B[47]), .A2(B[48]), .A3(n212), .ZN(n208) );
  OR3_X1 U27 ( .A1(B[43]), .A2(B[44]), .A3(n216), .ZN(n214) );
  OR3_X1 U28 ( .A1(B[39]), .A2(B[40]), .A3(n220), .ZN(n218) );
  OR2_X1 U29 ( .A1(n204), .A2(B[53]), .ZN(n205) );
  OR2_X1 U30 ( .A1(n208), .A2(B[49]), .ZN(n209) );
  OR2_X1 U31 ( .A1(n214), .A2(B[45]), .ZN(n215) );
  OR2_X1 U32 ( .A1(n218), .A2(B[41]), .ZN(n219) );
  OR3_X1 U33 ( .A1(B[29]), .A2(B[30]), .A3(n230), .ZN(n228) );
  OR2_X1 U34 ( .A1(n230), .A2(B[29]), .ZN(n231) );
  NOR2_X1 U35 ( .A1(B[27]), .A2(n233), .ZN(n234) );
  OR3_X1 U36 ( .A1(B[27]), .A2(B[28]), .A3(n233), .ZN(n230) );
  XNOR2_X1 U37 ( .A(B[40]), .B(n221), .ZN(DIFF[40]) );
  XNOR2_X1 U38 ( .A(B[36]), .B(n225), .ZN(DIFF[36]) );
  XNOR2_X1 U39 ( .A(B[32]), .B(n229), .ZN(DIFF[32]) );
  XNOR2_X1 U40 ( .A(B[28]), .B(n234), .ZN(DIFF[28]) );
  XNOR2_X1 U41 ( .A(n197), .B(B[61]), .ZN(DIFF[61]) );
  XNOR2_X1 U42 ( .A(B[52]), .B(n207), .ZN(DIFF[52]) );
  XNOR2_X1 U43 ( .A(B[48]), .B(n213), .ZN(DIFF[48]) );
  XNOR2_X1 U44 ( .A(B[44]), .B(n217), .ZN(DIFF[44]) );
  XNOR2_X1 U45 ( .A(B[56]), .B(n203), .ZN(DIFF[56]) );
  XNOR2_X1 U46 ( .A(B[60]), .B(n199), .ZN(DIFF[60]) );
  OR3_X1 U47 ( .A1(B[25]), .A2(B[26]), .A3(n235), .ZN(n233) );
  XNOR2_X1 U48 ( .A(B[24]), .B(n238), .ZN(DIFF[24]) );
  OR2_X1 U49 ( .A1(n235), .A2(B[25]), .ZN(n236) );
  NOR2_X1 U50 ( .A1(B[23]), .A2(n237), .ZN(n238) );
  OR3_X1 U51 ( .A1(B[23]), .A2(B[24]), .A3(n237), .ZN(n235) );
  XNOR2_X1 U52 ( .A(n189), .B(B[18]), .ZN(DIFF[18]) );
  NOR2_X1 U53 ( .A1(n243), .A2(B[17]), .ZN(n189) );
  XNOR2_X1 U54 ( .A(n193), .B(B[14]), .ZN(DIFF[14]) );
  NOR2_X1 U55 ( .A1(n247), .A2(B[13]), .ZN(n193) );
  XNOR2_X1 U56 ( .A(n244), .B(B[6]), .ZN(DIFF[6]) );
  NOR2_X1 U57 ( .A1(n194), .A2(B[5]), .ZN(n244) );
  XNOR2_X1 U58 ( .A(n248), .B(B[10]), .ZN(DIFF[10]) );
  NOR2_X1 U59 ( .A1(n190), .A2(B[9]), .ZN(n248) );
  XNOR2_X1 U60 ( .A(B[20]), .B(n242), .ZN(DIFF[20]) );
  NOR2_X1 U61 ( .A1(B[19]), .A2(n241), .ZN(n242) );
  XNOR2_X1 U62 ( .A(B[16]), .B(n246), .ZN(DIFF[16]) );
  NOR2_X1 U63 ( .A1(B[15]), .A2(n245), .ZN(n246) );
  XNOR2_X1 U64 ( .A(B[12]), .B(n250), .ZN(DIFF[12]) );
  NOR2_X1 U65 ( .A1(B[11]), .A2(n249), .ZN(n250) );
  XNOR2_X1 U66 ( .A(B[8]), .B(n191), .ZN(DIFF[8]) );
  NOR2_X1 U67 ( .A1(B[7]), .A2(n192), .ZN(n191) );
  XNOR2_X1 U68 ( .A(B[2]), .B(n232), .ZN(DIFF[2]) );
  NOR2_X1 U69 ( .A1(\B[0] ), .A2(B[1]), .ZN(n232) );
  XNOR2_X1 U70 ( .A(B[4]), .B(n210), .ZN(DIFF[4]) );
  NOR2_X1 U71 ( .A1(B[3]), .A2(n211), .ZN(n210) );
  OR3_X1 U72 ( .A1(B[5]), .A2(B[6]), .A3(n194), .ZN(n192) );
  OR3_X1 U73 ( .A1(B[10]), .A2(B[9]), .A3(n190), .ZN(n249) );
  OR3_X1 U74 ( .A1(B[13]), .A2(B[14]), .A3(n247), .ZN(n245) );
  OR3_X1 U75 ( .A1(B[17]), .A2(B[18]), .A3(n243), .ZN(n241) );
  OR3_X1 U76 ( .A1(B[21]), .A2(B[22]), .A3(n239), .ZN(n237) );
  OR3_X1 U77 ( .A1(B[7]), .A2(B[8]), .A3(n192), .ZN(n190) );
  OR3_X1 U78 ( .A1(B[11]), .A2(B[12]), .A3(n249), .ZN(n247) );
  OR3_X1 U79 ( .A1(B[15]), .A2(B[16]), .A3(n245), .ZN(n243) );
  OR3_X1 U80 ( .A1(B[19]), .A2(B[20]), .A3(n241), .ZN(n239) );
  OR3_X1 U83 ( .A1(B[3]), .A2(B[4]), .A3(n211), .ZN(n194) );
  OR2_X1 U120 ( .A1(n239), .A2(B[21]), .ZN(n240) );
  OR3_X1 U123 ( .A1(B[1]), .A2(B[2]), .A3(\B[0] ), .ZN(n211) );
  INV_X1 U126 ( .A(B[61]), .ZN(n251) );
endmodule


module complementer_N64_9 ( \input , complement2 );
  input [63:0] \input ;
  output [63:0] complement2;


  complementer_N64_9_DW01_sub_0 sub_add_31_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(\input ), .CI(1'b0), .DIFF(complement2) );
endmodule


module ShiftnCompl_N64_5 ( plusA, plus2A_out, minus2A_out, plus4A_out, 
        minus4A_out );
  input [63:0] plusA;
  output [63:0] plus2A_out;
  output [63:0] minus2A_out;
  output [63:0] plus4A_out;
  output [63:0] minus4A_out;
  wire   n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign plus2A_out[0] = 1'b0;
  assign plus4A_out[0] = 1'b0;

  shifter_N64_10 shifter_1 ( .\input (plusA), .shiftLeftOnePos({
        plus2A_out[63:59], n33, plus2A_out[57:52], n34, n35, n36, n37, n38, 
        n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, 
        n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, 
        plus2A_out[21:1], SYNOPSYS_UNCONNECTED__0}) );
  shifter_N64_9 shifter_2 ( .\input ({plus2A_out[63:1], 1'b0}), 
        .shiftLeftOnePos({plus4A_out[63:59], n64, plus4A_out[57:1], 
        SYNOPSYS_UNCONNECTED__1}) );
  complementer_N64_10 complementer_1 ( .\input ({plus2A_out[63:1], 1'b0}), 
        .complement2(minus2A_out) );
  complementer_N64_9 complementer_2 ( .\input ({plus4A_out[63:1], 1'b0}), 
        .complement2(minus4A_out) );
  BUF_X1 U3 ( .A(n50), .Z(plus2A_out[35]) );
  BUF_X1 U4 ( .A(n54), .Z(plus2A_out[31]) );
  BUF_X1 U5 ( .A(n38), .Z(plus2A_out[47]) );
  BUF_X1 U6 ( .A(n42), .Z(plus2A_out[43]) );
  BUF_X1 U7 ( .A(n46), .Z(plus2A_out[39]) );
  BUF_X1 U8 ( .A(n34), .Z(plus2A_out[51]) );
  BUF_X1 U9 ( .A(n64), .Z(plus4A_out[58]) );
  BUF_X1 U10 ( .A(n33), .Z(plus2A_out[58]) );
  BUF_X1 U11 ( .A(n58), .Z(plus2A_out[27]) );
  BUF_X1 U12 ( .A(n62), .Z(plus2A_out[23]) );
  BUF_X1 U13 ( .A(n56), .Z(plus2A_out[29]) );
  BUF_X1 U14 ( .A(n60), .Z(plus2A_out[25]) );
  BUF_X1 U15 ( .A(n57), .Z(plus2A_out[28]) );
  BUF_X1 U16 ( .A(n61), .Z(plus2A_out[24]) );
  BUF_X1 U17 ( .A(n59), .Z(plus2A_out[26]) );
  BUF_X1 U18 ( .A(n63), .Z(plus2A_out[22]) );
  BUF_X1 U19 ( .A(n48), .Z(plus2A_out[37]) );
  BUF_X1 U20 ( .A(n52), .Z(plus2A_out[33]) );
  BUF_X1 U21 ( .A(n45), .Z(plus2A_out[40]) );
  BUF_X1 U22 ( .A(n49), .Z(plus2A_out[36]) );
  BUF_X1 U23 ( .A(n53), .Z(plus2A_out[32]) );
  BUF_X1 U24 ( .A(n47), .Z(plus2A_out[38]) );
  BUF_X1 U25 ( .A(n51), .Z(plus2A_out[34]) );
  BUF_X1 U26 ( .A(n55), .Z(plus2A_out[30]) );
  BUF_X1 U27 ( .A(n36), .Z(plus2A_out[49]) );
  BUF_X1 U28 ( .A(n40), .Z(plus2A_out[45]) );
  BUF_X1 U29 ( .A(n44), .Z(plus2A_out[41]) );
  BUF_X1 U30 ( .A(n37), .Z(plus2A_out[48]) );
  BUF_X1 U31 ( .A(n41), .Z(plus2A_out[44]) );
  BUF_X1 U32 ( .A(n35), .Z(plus2A_out[50]) );
  BUF_X1 U33 ( .A(n39), .Z(plus2A_out[46]) );
  BUF_X1 U34 ( .A(n43), .Z(plus2A_out[42]) );
endmodule


module MUX_GENERIC_N64_RADIX3_5 ( plusA, minusA, plus2A, minus2A, SEL, Y );
  input [63:0] plusA;
  input [63:0] minusA;
  input [63:0] plus2A;
  input [63:0] minus2A;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502;
  tri   [63:0] Y;

  TBUF_X1 \Y_tri[55]  ( .A(n446), .EN(n301), .Z(Y[55]) );
  TBUF_X1 \Y_tri[56]  ( .A(n445), .EN(n301), .Z(Y[56]) );
  TBUF_X1 \Y_tri[57]  ( .A(n444), .EN(n301), .Z(Y[57]) );
  TBUF_X1 \Y_tri[58]  ( .A(n443), .EN(n301), .Z(Y[58]) );
  TBUF_X1 \Y_tri[59]  ( .A(n442), .EN(n301), .Z(Y[59]) );
  TBUF_X1 \Y_tri[60]  ( .A(n441), .EN(n301), .Z(Y[60]) );
  TBUF_X1 \Y_tri[61]  ( .A(n440), .EN(n301), .Z(Y[61]) );
  TBUF_X1 \Y_tri[62]  ( .A(n439), .EN(n301), .Z(Y[62]) );
  TBUF_X1 \Y_tri[63]  ( .A(n438), .EN(n301), .Z(Y[63]) );
  TBUF_X1 \Y_tri[42]  ( .A(n459), .EN(n299), .Z(Y[42]) );
  TBUF_X1 \Y_tri[43]  ( .A(n458), .EN(n299), .Z(Y[43]) );
  TBUF_X1 \Y_tri[44]  ( .A(n457), .EN(n300), .Z(Y[44]) );
  TBUF_X1 \Y_tri[45]  ( .A(n456), .EN(n300), .Z(Y[45]) );
  TBUF_X1 \Y_tri[46]  ( .A(n455), .EN(n300), .Z(Y[46]) );
  TBUF_X1 \Y_tri[47]  ( .A(n454), .EN(n300), .Z(Y[47]) );
  TBUF_X1 \Y_tri[48]  ( .A(n453), .EN(n300), .Z(Y[48]) );
  TBUF_X1 \Y_tri[49]  ( .A(n452), .EN(n300), .Z(Y[49]) );
  TBUF_X1 \Y_tri[50]  ( .A(n451), .EN(n300), .Z(Y[50]) );
  TBUF_X1 \Y_tri[51]  ( .A(n450), .EN(n300), .Z(Y[51]) );
  TBUF_X1 \Y_tri[52]  ( .A(n449), .EN(n300), .Z(Y[52]) );
  TBUF_X1 \Y_tri[53]  ( .A(n448), .EN(n300), .Z(Y[53]) );
  TBUF_X1 \Y_tri[54]  ( .A(n447), .EN(n300), .Z(Y[54]) );
  TBUF_X1 \Y_tri[16]  ( .A(n485), .EN(n297), .Z(Y[16]) );
  TBUF_X1 \Y_tri[17]  ( .A(n484), .EN(n297), .Z(Y[17]) );
  TBUF_X1 \Y_tri[18]  ( .A(n483), .EN(n297), .Z(Y[18]) );
  TBUF_X1 \Y_tri[19]  ( .A(n482), .EN(n297), .Z(Y[19]) );
  TBUF_X1 \Y_tri[20]  ( .A(n481), .EN(n297), .Z(Y[20]) );
  TBUF_X1 \Y_tri[21]  ( .A(n480), .EN(n297), .Z(Y[21]) );
  TBUF_X1 \Y_tri[22]  ( .A(n479), .EN(n298), .Z(Y[22]) );
  TBUF_X1 \Y_tri[23]  ( .A(n478), .EN(n298), .Z(Y[23]) );
  TBUF_X1 \Y_tri[24]  ( .A(n477), .EN(n298), .Z(Y[24]) );
  TBUF_X1 \Y_tri[25]  ( .A(n476), .EN(n298), .Z(Y[25]) );
  TBUF_X1 \Y_tri[26]  ( .A(n475), .EN(n298), .Z(Y[26]) );
  TBUF_X1 \Y_tri[27]  ( .A(n474), .EN(n298), .Z(Y[27]) );
  TBUF_X1 \Y_tri[28]  ( .A(n473), .EN(n298), .Z(Y[28]) );
  TBUF_X1 \Y_tri[29]  ( .A(n472), .EN(n298), .Z(Y[29]) );
  TBUF_X1 \Y_tri[30]  ( .A(n471), .EN(n298), .Z(Y[30]) );
  TBUF_X1 \Y_tri[31]  ( .A(n470), .EN(n298), .Z(Y[31]) );
  TBUF_X1 \Y_tri[32]  ( .A(n469), .EN(n298), .Z(Y[32]) );
  TBUF_X1 \Y_tri[33]  ( .A(n468), .EN(n299), .Z(Y[33]) );
  TBUF_X1 \Y_tri[34]  ( .A(n467), .EN(n299), .Z(Y[34]) );
  TBUF_X1 \Y_tri[35]  ( .A(n466), .EN(n299), .Z(Y[35]) );
  TBUF_X1 \Y_tri[36]  ( .A(n465), .EN(n299), .Z(Y[36]) );
  TBUF_X1 \Y_tri[37]  ( .A(n464), .EN(n299), .Z(Y[37]) );
  TBUF_X1 \Y_tri[38]  ( .A(n463), .EN(n299), .Z(Y[38]) );
  TBUF_X1 \Y_tri[39]  ( .A(n462), .EN(n299), .Z(Y[39]) );
  TBUF_X1 \Y_tri[40]  ( .A(n461), .EN(n299), .Z(Y[40]) );
  TBUF_X1 \Y_tri[41]  ( .A(n460), .EN(n299), .Z(Y[41]) );
  TBUF_X1 \Y_tri[5]  ( .A(n497), .EN(n296), .Z(Y[5]) );
  TBUF_X1 \Y_tri[6]  ( .A(n496), .EN(n296), .Z(Y[6]) );
  TBUF_X1 \Y_tri[7]  ( .A(n495), .EN(n296), .Z(Y[7]) );
  TBUF_X1 \Y_tri[8]  ( .A(n494), .EN(n296), .Z(Y[8]) );
  TBUF_X1 \Y_tri[9]  ( .A(n492), .EN(n296), .Z(Y[9]) );
  TBUF_X1 \Y_tri[10]  ( .A(n491), .EN(n296), .Z(Y[10]) );
  TBUF_X1 \Y_tri[11]  ( .A(n490), .EN(n297), .Z(Y[11]) );
  TBUF_X1 \Y_tri[12]  ( .A(n489), .EN(n297), .Z(Y[12]) );
  TBUF_X1 \Y_tri[13]  ( .A(n488), .EN(n297), .Z(Y[13]) );
  TBUF_X1 \Y_tri[14]  ( .A(n487), .EN(n297), .Z(Y[14]) );
  TBUF_X1 \Y_tri[15]  ( .A(n486), .EN(n297), .Z(Y[15]) );
  TBUF_X1 \Y_tri[0]  ( .A(n502), .EN(n296), .Z(Y[0]) );
  TBUF_X1 \Y_tri[1]  ( .A(n501), .EN(n296), .Z(Y[1]) );
  TBUF_X1 \Y_tri[2]  ( .A(n500), .EN(n296), .Z(Y[2]) );
  TBUF_X1 \Y_tri[3]  ( .A(n499), .EN(n296), .Z(Y[3]) );
  TBUF_X1 \Y_tri[4]  ( .A(n498), .EN(n296), .Z(Y[4]) );
  NAND2_X1 U2 ( .A1(n387), .A2(n386), .ZN(n461) );
  AOI22_X1 U3 ( .A1(plusA[40]), .A2(n281), .B1(plus2A[40]), .B2(n275), .ZN(
        n387) );
  AOI22_X1 U4 ( .A1(minus2A[40]), .A2(n293), .B1(minusA[40]), .B2(n287), .ZN(
        n386) );
  NAND2_X1 U5 ( .A1(n379), .A2(n378), .ZN(n465) );
  AOI22_X1 U6 ( .A1(plusA[36]), .A2(n281), .B1(plus2A[36]), .B2(n275), .ZN(
        n379) );
  AOI22_X1 U7 ( .A1(minus2A[36]), .A2(n293), .B1(minusA[36]), .B2(n287), .ZN(
        n378) );
  NAND2_X1 U8 ( .A1(n371), .A2(n370), .ZN(n469) );
  AOI22_X1 U9 ( .A1(plusA[32]), .A2(n280), .B1(plus2A[32]), .B2(n274), .ZN(
        n371) );
  AOI22_X1 U10 ( .A1(minus2A[32]), .A2(n292), .B1(minusA[32]), .B2(n286), .ZN(
        n370) );
  NAND2_X1 U11 ( .A1(n363), .A2(n362), .ZN(n473) );
  AOI22_X1 U12 ( .A1(plusA[28]), .A2(n280), .B1(plus2A[28]), .B2(n274), .ZN(
        n363) );
  AOI22_X1 U13 ( .A1(minus2A[28]), .A2(n292), .B1(minusA[28]), .B2(n286), .ZN(
        n362) );
  NAND2_X1 U14 ( .A1(n383), .A2(n382), .ZN(n463) );
  AOI22_X1 U15 ( .A1(plusA[38]), .A2(n281), .B1(plus2A[38]), .B2(n275), .ZN(
        n383) );
  AOI22_X1 U16 ( .A1(minus2A[38]), .A2(n293), .B1(minusA[38]), .B2(n287), .ZN(
        n382) );
  NAND2_X1 U17 ( .A1(n375), .A2(n374), .ZN(n467) );
  AOI22_X1 U18 ( .A1(plusA[34]), .A2(n280), .B1(plus2A[34]), .B2(n274), .ZN(
        n375) );
  AOI22_X1 U19 ( .A1(minus2A[34]), .A2(n292), .B1(minusA[34]), .B2(n286), .ZN(
        n374) );
  NAND2_X1 U20 ( .A1(n367), .A2(n366), .ZN(n471) );
  AOI22_X1 U21 ( .A1(plusA[30]), .A2(n280), .B1(plus2A[30]), .B2(n274), .ZN(
        n367) );
  AOI22_X1 U22 ( .A1(minus2A[30]), .A2(n292), .B1(minusA[30]), .B2(n286), .ZN(
        n366) );
  NAND2_X1 U23 ( .A1(n359), .A2(n358), .ZN(n475) );
  AOI22_X1 U24 ( .A1(plusA[26]), .A2(n280), .B1(plus2A[26]), .B2(n274), .ZN(
        n359) );
  AOI22_X1 U25 ( .A1(minus2A[26]), .A2(n292), .B1(minusA[26]), .B2(n286), .ZN(
        n358) );
  NAND2_X1 U26 ( .A1(n389), .A2(n388), .ZN(n460) );
  AOI22_X1 U27 ( .A1(plusA[41]), .A2(n281), .B1(plus2A[41]), .B2(n275), .ZN(
        n389) );
  AOI22_X1 U28 ( .A1(minus2A[41]), .A2(n293), .B1(minusA[41]), .B2(n287), .ZN(
        n388) );
  NAND2_X1 U29 ( .A1(n381), .A2(n380), .ZN(n464) );
  AOI22_X1 U30 ( .A1(plusA[37]), .A2(n281), .B1(plus2A[37]), .B2(n275), .ZN(
        n381) );
  AOI22_X1 U31 ( .A1(minus2A[37]), .A2(n293), .B1(minusA[37]), .B2(n287), .ZN(
        n380) );
  NAND2_X1 U32 ( .A1(n373), .A2(n372), .ZN(n468) );
  AOI22_X1 U33 ( .A1(plusA[33]), .A2(n280), .B1(plus2A[33]), .B2(n274), .ZN(
        n373) );
  AOI22_X1 U34 ( .A1(minus2A[33]), .A2(n292), .B1(minusA[33]), .B2(n286), .ZN(
        n372) );
  NAND2_X1 U35 ( .A1(n365), .A2(n364), .ZN(n472) );
  AOI22_X1 U36 ( .A1(plusA[29]), .A2(n280), .B1(plus2A[29]), .B2(n274), .ZN(
        n365) );
  AOI22_X1 U37 ( .A1(minus2A[29]), .A2(n292), .B1(minusA[29]), .B2(n286), .ZN(
        n364) );
  NAND2_X1 U38 ( .A1(n385), .A2(n384), .ZN(n462) );
  AOI22_X1 U39 ( .A1(plusA[39]), .A2(n281), .B1(plus2A[39]), .B2(n275), .ZN(
        n385) );
  AOI22_X1 U40 ( .A1(minus2A[39]), .A2(n293), .B1(minusA[39]), .B2(n287), .ZN(
        n384) );
  NAND2_X1 U41 ( .A1(n377), .A2(n376), .ZN(n466) );
  AOI22_X1 U42 ( .A1(plusA[35]), .A2(n280), .B1(plus2A[35]), .B2(n274), .ZN(
        n377) );
  AOI22_X1 U43 ( .A1(minus2A[35]), .A2(n292), .B1(minusA[35]), .B2(n286), .ZN(
        n376) );
  NAND2_X1 U44 ( .A1(n369), .A2(n368), .ZN(n470) );
  AOI22_X1 U45 ( .A1(plusA[31]), .A2(n280), .B1(plus2A[31]), .B2(n274), .ZN(
        n369) );
  AOI22_X1 U46 ( .A1(minus2A[31]), .A2(n292), .B1(minusA[31]), .B2(n286), .ZN(
        n368) );
  NAND2_X1 U47 ( .A1(n361), .A2(n360), .ZN(n474) );
  AOI22_X1 U48 ( .A1(plusA[27]), .A2(n280), .B1(plus2A[27]), .B2(n274), .ZN(
        n361) );
  AOI22_X1 U49 ( .A1(minus2A[27]), .A2(n292), .B1(minusA[27]), .B2(n286), .ZN(
        n360) );
  NAND2_X1 U50 ( .A1(n429), .A2(n428), .ZN(n440) );
  AOI22_X1 U51 ( .A1(plusA[61]), .A2(n283), .B1(plus2A[61]), .B2(n277), .ZN(
        n429) );
  AOI22_X1 U52 ( .A1(minus2A[61]), .A2(n295), .B1(minusA[61]), .B2(n289), .ZN(
        n428) );
  NAND2_X1 U53 ( .A1(n411), .A2(n410), .ZN(n449) );
  AOI22_X1 U54 ( .A1(plusA[52]), .A2(n282), .B1(plus2A[52]), .B2(n276), .ZN(
        n411) );
  AOI22_X1 U55 ( .A1(minus2A[52]), .A2(n294), .B1(minusA[52]), .B2(n288), .ZN(
        n410) );
  NAND2_X1 U56 ( .A1(n403), .A2(n402), .ZN(n453) );
  AOI22_X1 U57 ( .A1(plusA[48]), .A2(n282), .B1(plus2A[48]), .B2(n276), .ZN(
        n403) );
  AOI22_X1 U58 ( .A1(minus2A[48]), .A2(n294), .B1(minusA[48]), .B2(n288), .ZN(
        n402) );
  NAND2_X1 U59 ( .A1(n395), .A2(n394), .ZN(n457) );
  AOI22_X1 U60 ( .A1(plusA[44]), .A2(n281), .B1(plus2A[44]), .B2(n275), .ZN(
        n395) );
  AOI22_X1 U61 ( .A1(minus2A[44]), .A2(n293), .B1(minusA[44]), .B2(n287), .ZN(
        n394) );
  NAND2_X1 U62 ( .A1(n413), .A2(n412), .ZN(n448) );
  AOI22_X1 U63 ( .A1(plusA[53]), .A2(n282), .B1(plus2A[53]), .B2(n276), .ZN(
        n413) );
  AOI22_X1 U64 ( .A1(minus2A[53]), .A2(n294), .B1(minusA[53]), .B2(n288), .ZN(
        n412) );
  NAND2_X1 U65 ( .A1(n419), .A2(n418), .ZN(n445) );
  AOI22_X1 U66 ( .A1(plusA[56]), .A2(n282), .B1(plus2A[56]), .B2(n276), .ZN(
        n419) );
  AOI22_X1 U67 ( .A1(minus2A[56]), .A2(n294), .B1(minusA[56]), .B2(n288), .ZN(
        n418) );
  NAND2_X1 U68 ( .A1(n407), .A2(n406), .ZN(n451) );
  AOI22_X1 U69 ( .A1(plusA[50]), .A2(n282), .B1(plus2A[50]), .B2(n276), .ZN(
        n407) );
  AOI22_X1 U70 ( .A1(minus2A[50]), .A2(n294), .B1(minusA[50]), .B2(n288), .ZN(
        n406) );
  NAND2_X1 U71 ( .A1(n399), .A2(n398), .ZN(n455) );
  AOI22_X1 U72 ( .A1(plusA[46]), .A2(n281), .B1(plus2A[46]), .B2(n275), .ZN(
        n399) );
  AOI22_X1 U73 ( .A1(minus2A[46]), .A2(n293), .B1(minusA[46]), .B2(n287), .ZN(
        n398) );
  NAND2_X1 U74 ( .A1(n391), .A2(n390), .ZN(n459) );
  AOI22_X1 U75 ( .A1(plusA[42]), .A2(n281), .B1(plus2A[42]), .B2(n275), .ZN(
        n391) );
  AOI22_X1 U76 ( .A1(minus2A[42]), .A2(n293), .B1(minusA[42]), .B2(n287), .ZN(
        n390) );
  NAND2_X1 U77 ( .A1(n421), .A2(n420), .ZN(n444) );
  AOI22_X1 U78 ( .A1(plusA[57]), .A2(n282), .B1(plus2A[57]), .B2(n276), .ZN(
        n421) );
  AOI22_X1 U79 ( .A1(minus2A[57]), .A2(n294), .B1(minusA[57]), .B2(n288), .ZN(
        n420) );
  NAND2_X1 U80 ( .A1(n417), .A2(n416), .ZN(n446) );
  AOI22_X1 U81 ( .A1(plusA[55]), .A2(n282), .B1(plus2A[55]), .B2(n276), .ZN(
        n417) );
  AOI22_X1 U82 ( .A1(minus2A[55]), .A2(n294), .B1(minusA[55]), .B2(n288), .ZN(
        n416) );
  NAND2_X1 U83 ( .A1(n405), .A2(n404), .ZN(n452) );
  AOI22_X1 U84 ( .A1(plusA[49]), .A2(n282), .B1(plus2A[49]), .B2(n276), .ZN(
        n405) );
  AOI22_X1 U85 ( .A1(minus2A[49]), .A2(n294), .B1(minusA[49]), .B2(n288), .ZN(
        n404) );
  NAND2_X1 U86 ( .A1(n397), .A2(n396), .ZN(n456) );
  AOI22_X1 U87 ( .A1(plusA[45]), .A2(n281), .B1(plus2A[45]), .B2(n275), .ZN(
        n397) );
  AOI22_X1 U88 ( .A1(minus2A[45]), .A2(n293), .B1(minusA[45]), .B2(n287), .ZN(
        n396) );
  NAND2_X1 U89 ( .A1(n415), .A2(n414), .ZN(n447) );
  AOI22_X1 U90 ( .A1(plusA[54]), .A2(n282), .B1(plus2A[54]), .B2(n276), .ZN(
        n415) );
  AOI22_X1 U91 ( .A1(minus2A[54]), .A2(n294), .B1(minusA[54]), .B2(n288), .ZN(
        n414) );
  NAND2_X1 U92 ( .A1(n409), .A2(n408), .ZN(n450) );
  AOI22_X1 U93 ( .A1(plusA[51]), .A2(n282), .B1(plus2A[51]), .B2(n276), .ZN(
        n409) );
  AOI22_X1 U94 ( .A1(minus2A[51]), .A2(n294), .B1(minusA[51]), .B2(n288), .ZN(
        n408) );
  NAND2_X1 U95 ( .A1(n401), .A2(n400), .ZN(n454) );
  AOI22_X1 U96 ( .A1(plusA[47]), .A2(n281), .B1(plus2A[47]), .B2(n275), .ZN(
        n401) );
  AOI22_X1 U97 ( .A1(minus2A[47]), .A2(n293), .B1(minusA[47]), .B2(n287), .ZN(
        n400) );
  NAND2_X1 U98 ( .A1(n393), .A2(n392), .ZN(n458) );
  AOI22_X1 U99 ( .A1(plusA[43]), .A2(n281), .B1(plus2A[43]), .B2(n275), .ZN(
        n393) );
  AOI22_X1 U100 ( .A1(minus2A[43]), .A2(n293), .B1(minusA[43]), .B2(n287), 
        .ZN(n392) );
  NAND2_X1 U101 ( .A1(n437), .A2(n436), .ZN(n438) );
  AOI22_X1 U102 ( .A1(plusA[63]), .A2(n283), .B1(plus2A[63]), .B2(n277), .ZN(
        n437) );
  AOI22_X1 U103 ( .A1(minus2A[63]), .A2(n295), .B1(minusA[63]), .B2(n289), 
        .ZN(n436) );
  NAND2_X1 U104 ( .A1(n431), .A2(n430), .ZN(n439) );
  AOI22_X1 U105 ( .A1(plusA[62]), .A2(n283), .B1(plus2A[62]), .B2(n277), .ZN(
        n431) );
  AOI22_X1 U106 ( .A1(minus2A[62]), .A2(n295), .B1(minusA[62]), .B2(n289), 
        .ZN(n430) );
  NAND2_X1 U107 ( .A1(n427), .A2(n426), .ZN(n441) );
  AOI22_X1 U108 ( .A1(plusA[60]), .A2(n283), .B1(plus2A[60]), .B2(n277), .ZN(
        n427) );
  AOI22_X1 U109 ( .A1(minus2A[60]), .A2(n295), .B1(minusA[60]), .B2(n289), 
        .ZN(n426) );
  NAND2_X1 U110 ( .A1(n425), .A2(n424), .ZN(n442) );
  AOI22_X1 U111 ( .A1(plusA[59]), .A2(n282), .B1(plus2A[59]), .B2(n276), .ZN(
        n425) );
  AOI22_X1 U112 ( .A1(minus2A[59]), .A2(n294), .B1(minusA[59]), .B2(n288), 
        .ZN(n424) );
  NAND2_X1 U113 ( .A1(n423), .A2(n422), .ZN(n443) );
  AOI22_X1 U114 ( .A1(plusA[58]), .A2(n282), .B1(plus2A[58]), .B2(n276), .ZN(
        n423) );
  AOI22_X1 U115 ( .A1(minus2A[58]), .A2(n294), .B1(minusA[58]), .B2(n288), 
        .ZN(n422) );
  BUF_X1 U116 ( .A(n493), .Z(n296) );
  BUF_X1 U117 ( .A(n493), .Z(n297) );
  BUF_X1 U118 ( .A(n433), .Z(n280) );
  BUF_X1 U119 ( .A(n433), .Z(n279) );
  BUF_X1 U120 ( .A(n435), .Z(n292) );
  BUF_X1 U121 ( .A(n435), .Z(n291) );
  BUF_X1 U122 ( .A(n434), .Z(n286) );
  BUF_X1 U123 ( .A(n432), .Z(n274) );
  BUF_X1 U124 ( .A(n434), .Z(n285) );
  BUF_X1 U125 ( .A(n432), .Z(n273) );
  BUF_X1 U126 ( .A(n493), .Z(n298) );
  NAND2_X1 U127 ( .A1(n355), .A2(n354), .ZN(n477) );
  AOI22_X1 U128 ( .A1(plusA[24]), .A2(n280), .B1(plus2A[24]), .B2(n274), .ZN(
        n355) );
  AOI22_X1 U129 ( .A1(minus2A[24]), .A2(n292), .B1(minusA[24]), .B2(n286), 
        .ZN(n354) );
  NAND2_X1 U130 ( .A1(n357), .A2(n356), .ZN(n476) );
  AOI22_X1 U131 ( .A1(plusA[25]), .A2(n280), .B1(plus2A[25]), .B2(n274), .ZN(
        n357) );
  AOI22_X1 U132 ( .A1(minus2A[25]), .A2(n292), .B1(minusA[25]), .B2(n286), 
        .ZN(n356) );
  BUF_X1 U133 ( .A(n433), .Z(n281) );
  BUF_X1 U134 ( .A(n435), .Z(n293) );
  BUF_X1 U135 ( .A(n434), .Z(n287) );
  BUF_X1 U136 ( .A(n432), .Z(n275) );
  BUF_X1 U137 ( .A(n493), .Z(n299) );
  BUF_X1 U138 ( .A(n493), .Z(n300) );
  BUF_X1 U139 ( .A(n433), .Z(n282) );
  BUF_X1 U140 ( .A(n435), .Z(n294) );
  BUF_X1 U141 ( .A(n434), .Z(n288) );
  BUF_X1 U142 ( .A(n432), .Z(n276) );
  BUF_X1 U143 ( .A(n493), .Z(n301) );
  BUF_X1 U144 ( .A(n433), .Z(n278) );
  BUF_X1 U145 ( .A(n435), .Z(n290) );
  BUF_X1 U146 ( .A(n434), .Z(n284) );
  BUF_X1 U147 ( .A(n432), .Z(n272) );
  NOR2_X1 U148 ( .A1(n323), .A2(n304), .ZN(n493) );
  INV_X1 U149 ( .A(SEL[2]), .ZN(n304) );
  NOR2_X1 U150 ( .A1(SEL[1]), .A2(SEL[0]), .ZN(n323) );
  NOR3_X1 U151 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n302), .ZN(n434) );
  NOR3_X1 U152 ( .A1(SEL[1]), .A2(SEL[2]), .A3(n303), .ZN(n433) );
  NOR3_X1 U153 ( .A1(n302), .A2(SEL[2]), .A3(n303), .ZN(n432) );
  AND2_X1 U154 ( .A1(SEL[2]), .A2(n323), .ZN(n435) );
  INV_X1 U155 ( .A(SEL[1]), .ZN(n302) );
  INV_X1 U156 ( .A(SEL[0]), .ZN(n303) );
  NAND2_X1 U157 ( .A1(n353), .A2(n352), .ZN(n478) );
  AOI22_X1 U158 ( .A1(plusA[23]), .A2(n279), .B1(plus2A[23]), .B2(n273), .ZN(
        n353) );
  AOI22_X1 U159 ( .A1(minus2A[23]), .A2(n291), .B1(minusA[23]), .B2(n285), 
        .ZN(n352) );
  NAND2_X1 U160 ( .A1(n351), .A2(n350), .ZN(n479) );
  AOI22_X1 U161 ( .A1(plusA[22]), .A2(n279), .B1(plus2A[22]), .B2(n273), .ZN(
        n351) );
  AOI22_X1 U162 ( .A1(minus2A[22]), .A2(n291), .B1(minusA[22]), .B2(n285), 
        .ZN(n350) );
  NAND2_X1 U163 ( .A1(n349), .A2(n348), .ZN(n480) );
  AOI22_X1 U164 ( .A1(plusA[21]), .A2(n279), .B1(plus2A[21]), .B2(n273), .ZN(
        n349) );
  AOI22_X1 U165 ( .A1(minus2A[21]), .A2(n291), .B1(minusA[21]), .B2(n285), 
        .ZN(n348) );
  NAND2_X1 U166 ( .A1(n345), .A2(n344), .ZN(n482) );
  AOI22_X1 U167 ( .A1(plusA[19]), .A2(n279), .B1(plus2A[19]), .B2(n273), .ZN(
        n345) );
  AOI22_X1 U168 ( .A1(minus2A[19]), .A2(n291), .B1(minusA[19]), .B2(n285), 
        .ZN(n344) );
  NAND2_X1 U169 ( .A1(n343), .A2(n342), .ZN(n483) );
  AOI22_X1 U170 ( .A1(plusA[18]), .A2(n279), .B1(plus2A[18]), .B2(n273), .ZN(
        n343) );
  AOI22_X1 U171 ( .A1(minus2A[18]), .A2(n291), .B1(minusA[18]), .B2(n285), 
        .ZN(n342) );
  NAND2_X1 U172 ( .A1(n341), .A2(n340), .ZN(n484) );
  AOI22_X1 U173 ( .A1(plusA[17]), .A2(n279), .B1(plus2A[17]), .B2(n273), .ZN(
        n341) );
  AOI22_X1 U174 ( .A1(minus2A[17]), .A2(n291), .B1(minusA[17]), .B2(n285), 
        .ZN(n340) );
  NAND2_X1 U175 ( .A1(n337), .A2(n336), .ZN(n486) );
  AOI22_X1 U176 ( .A1(plusA[15]), .A2(n279), .B1(plus2A[15]), .B2(n273), .ZN(
        n337) );
  AOI22_X1 U177 ( .A1(minus2A[15]), .A2(n291), .B1(minusA[15]), .B2(n285), 
        .ZN(n336) );
  NAND2_X1 U178 ( .A1(n335), .A2(n334), .ZN(n487) );
  AOI22_X1 U179 ( .A1(plusA[14]), .A2(n279), .B1(plus2A[14]), .B2(n273), .ZN(
        n335) );
  AOI22_X1 U180 ( .A1(minus2A[14]), .A2(n291), .B1(minusA[14]), .B2(n285), 
        .ZN(n334) );
  NAND2_X1 U181 ( .A1(n333), .A2(n332), .ZN(n488) );
  AOI22_X1 U182 ( .A1(plusA[13]), .A2(n279), .B1(plus2A[13]), .B2(n273), .ZN(
        n333) );
  AOI22_X1 U183 ( .A1(minus2A[13]), .A2(n291), .B1(minusA[13]), .B2(n285), 
        .ZN(n332) );
  NAND2_X1 U184 ( .A1(n329), .A2(n328), .ZN(n490) );
  AOI22_X1 U185 ( .A1(plusA[11]), .A2(n278), .B1(plus2A[11]), .B2(n272), .ZN(
        n329) );
  AOI22_X1 U186 ( .A1(minus2A[11]), .A2(n290), .B1(minusA[11]), .B2(n284), 
        .ZN(n328) );
  NAND2_X1 U187 ( .A1(n327), .A2(n326), .ZN(n491) );
  AOI22_X1 U188 ( .A1(plusA[10]), .A2(n278), .B1(plus2A[10]), .B2(n272), .ZN(
        n327) );
  AOI22_X1 U189 ( .A1(minus2A[10]), .A2(n290), .B1(minusA[10]), .B2(n284), 
        .ZN(n326) );
  NAND2_X1 U190 ( .A1(n325), .A2(n324), .ZN(n492) );
  AOI22_X1 U191 ( .A1(plusA[9]), .A2(n278), .B1(plus2A[9]), .B2(n272), .ZN(
        n325) );
  AOI22_X1 U192 ( .A1(minus2A[9]), .A2(n290), .B1(minusA[9]), .B2(n284), .ZN(
        n324) );
  NAND2_X1 U193 ( .A1(n320), .A2(n319), .ZN(n495) );
  AOI22_X1 U194 ( .A1(plusA[7]), .A2(n278), .B1(plus2A[7]), .B2(n272), .ZN(
        n320) );
  AOI22_X1 U195 ( .A1(minus2A[7]), .A2(n290), .B1(minusA[7]), .B2(n284), .ZN(
        n319) );
  NAND2_X1 U196 ( .A1(n318), .A2(n317), .ZN(n496) );
  AOI22_X1 U197 ( .A1(plusA[6]), .A2(n278), .B1(plus2A[6]), .B2(n272), .ZN(
        n318) );
  AOI22_X1 U198 ( .A1(minus2A[6]), .A2(n290), .B1(minusA[6]), .B2(n284), .ZN(
        n317) );
  NAND2_X1 U199 ( .A1(n316), .A2(n315), .ZN(n497) );
  AOI22_X1 U200 ( .A1(plusA[5]), .A2(n278), .B1(plus2A[5]), .B2(n272), .ZN(
        n316) );
  AOI22_X1 U201 ( .A1(minus2A[5]), .A2(n290), .B1(minusA[5]), .B2(n284), .ZN(
        n315) );
  NAND2_X1 U202 ( .A1(n312), .A2(n311), .ZN(n499) );
  AOI22_X1 U203 ( .A1(plusA[3]), .A2(n278), .B1(plus2A[3]), .B2(n272), .ZN(
        n312) );
  AOI22_X1 U204 ( .A1(minus2A[3]), .A2(n290), .B1(minusA[3]), .B2(n284), .ZN(
        n311) );
  NAND2_X1 U205 ( .A1(n347), .A2(n346), .ZN(n481) );
  AOI22_X1 U206 ( .A1(plusA[20]), .A2(n279), .B1(plus2A[20]), .B2(n273), .ZN(
        n347) );
  AOI22_X1 U207 ( .A1(minus2A[20]), .A2(n291), .B1(minusA[20]), .B2(n285), 
        .ZN(n346) );
  NAND2_X1 U208 ( .A1(n339), .A2(n338), .ZN(n485) );
  AOI22_X1 U209 ( .A1(plusA[16]), .A2(n279), .B1(plus2A[16]), .B2(n273), .ZN(
        n339) );
  AOI22_X1 U210 ( .A1(minus2A[16]), .A2(n291), .B1(minusA[16]), .B2(n285), 
        .ZN(n338) );
  NAND2_X1 U211 ( .A1(n331), .A2(n330), .ZN(n489) );
  AOI22_X1 U212 ( .A1(plusA[12]), .A2(n279), .B1(plus2A[12]), .B2(n273), .ZN(
        n331) );
  AOI22_X1 U213 ( .A1(minus2A[12]), .A2(n291), .B1(minusA[12]), .B2(n285), 
        .ZN(n330) );
  NAND2_X1 U214 ( .A1(n322), .A2(n321), .ZN(n494) );
  AOI22_X1 U215 ( .A1(plusA[8]), .A2(n278), .B1(plus2A[8]), .B2(n272), .ZN(
        n322) );
  AOI22_X1 U216 ( .A1(minus2A[8]), .A2(n290), .B1(minusA[8]), .B2(n284), .ZN(
        n321) );
  NAND2_X1 U217 ( .A1(n314), .A2(n313), .ZN(n498) );
  AOI22_X1 U218 ( .A1(plusA[4]), .A2(n278), .B1(plus2A[4]), .B2(n272), .ZN(
        n314) );
  AOI22_X1 U219 ( .A1(minus2A[4]), .A2(n290), .B1(minusA[4]), .B2(n284), .ZN(
        n313) );
  NAND2_X1 U220 ( .A1(n310), .A2(n309), .ZN(n500) );
  AOI22_X1 U221 ( .A1(plusA[2]), .A2(n278), .B1(plus2A[2]), .B2(n272), .ZN(
        n310) );
  AOI22_X1 U222 ( .A1(minus2A[2]), .A2(n290), .B1(minusA[2]), .B2(n284), .ZN(
        n309) );
  NAND2_X1 U223 ( .A1(n308), .A2(n307), .ZN(n501) );
  AOI22_X1 U224 ( .A1(plusA[1]), .A2(n278), .B1(plus2A[1]), .B2(n272), .ZN(
        n308) );
  AOI22_X1 U225 ( .A1(minus2A[1]), .A2(n290), .B1(minusA[1]), .B2(n284), .ZN(
        n307) );
  NAND2_X1 U226 ( .A1(n306), .A2(n305), .ZN(n502) );
  AOI22_X1 U227 ( .A1(plusA[0]), .A2(n278), .B1(plus2A[0]), .B2(n272), .ZN(
        n306) );
  AOI22_X1 U228 ( .A1(minus2A[0]), .A2(n290), .B1(minusA[0]), .B2(n284), .ZN(
        n305) );
  CLKBUF_X1 U229 ( .A(n432), .Z(n277) );
  CLKBUF_X1 U230 ( .A(n433), .Z(n283) );
  CLKBUF_X1 U231 ( .A(n434), .Z(n289) );
  CLKBUF_X1 U232 ( .A(n435), .Z(n295) );
endmodule


module FA_320 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_319 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_318 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_317 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_316 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  XOR2_X1 U1 ( .A(Ci), .B(n5), .Z(S) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_315 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_314 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_313 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_312 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_311 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_310 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_309 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_308 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_307 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_306 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_305 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_304 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_303 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_302 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_301 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_300 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_299 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_298 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_297 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_296 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_295 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_294 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_293 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_292 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_291 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_290 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_289 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_288 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_287 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_286 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_285 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_284 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_283 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_282 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_281 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_280 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_279 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_278 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_277 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_276 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_275 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_274 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_273 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_272 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_271 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_270 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_269 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_268 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_267 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_266 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_265 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_264 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_263 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_262 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_261 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_260 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_259 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_258 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_257 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N64_5 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Ci;
  output Co;

  wire   [63:1] CTMP;
  tri   [63:0] A;

  FA_320 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_319 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_318 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_317 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(CTMP[4]) );
  FA_316 FAI_5 ( .A(A[4]), .B(B[4]), .Ci(CTMP[4]), .S(S[4]), .Co(CTMP[5]) );
  FA_315 FAI_6 ( .A(A[5]), .B(B[5]), .Ci(CTMP[5]), .S(S[5]), .Co(CTMP[6]) );
  FA_314 FAI_7 ( .A(A[6]), .B(B[6]), .Ci(CTMP[6]), .S(S[6]), .Co(CTMP[7]) );
  FA_313 FAI_8 ( .A(A[7]), .B(B[7]), .Ci(CTMP[7]), .S(S[7]), .Co(CTMP[8]) );
  FA_312 FAI_9 ( .A(A[8]), .B(B[8]), .Ci(CTMP[8]), .S(S[8]), .Co(CTMP[9]) );
  FA_311 FAI_10 ( .A(A[9]), .B(B[9]), .Ci(CTMP[9]), .S(S[9]), .Co(CTMP[10]) );
  FA_310 FAI_11 ( .A(A[10]), .B(B[10]), .Ci(CTMP[10]), .S(S[10]), .Co(CTMP[11]) );
  FA_309 FAI_12 ( .A(A[11]), .B(B[11]), .Ci(CTMP[11]), .S(S[11]), .Co(CTMP[12]) );
  FA_308 FAI_13 ( .A(A[12]), .B(B[12]), .Ci(CTMP[12]), .S(S[12]), .Co(CTMP[13]) );
  FA_307 FAI_14 ( .A(A[13]), .B(B[13]), .Ci(CTMP[13]), .S(S[13]), .Co(CTMP[14]) );
  FA_306 FAI_15 ( .A(A[14]), .B(B[14]), .Ci(CTMP[14]), .S(S[14]), .Co(CTMP[15]) );
  FA_305 FAI_16 ( .A(A[15]), .B(B[15]), .Ci(CTMP[15]), .S(S[15]), .Co(CTMP[16]) );
  FA_304 FAI_17 ( .A(A[16]), .B(B[16]), .Ci(CTMP[16]), .S(S[16]), .Co(CTMP[17]) );
  FA_303 FAI_18 ( .A(A[17]), .B(B[17]), .Ci(CTMP[17]), .S(S[17]), .Co(CTMP[18]) );
  FA_302 FAI_19 ( .A(A[18]), .B(B[18]), .Ci(CTMP[18]), .S(S[18]), .Co(CTMP[19]) );
  FA_301 FAI_20 ( .A(A[19]), .B(B[19]), .Ci(CTMP[19]), .S(S[19]), .Co(CTMP[20]) );
  FA_300 FAI_21 ( .A(A[20]), .B(B[20]), .Ci(CTMP[20]), .S(S[20]), .Co(CTMP[21]) );
  FA_299 FAI_22 ( .A(A[21]), .B(B[21]), .Ci(CTMP[21]), .S(S[21]), .Co(CTMP[22]) );
  FA_298 FAI_23 ( .A(A[22]), .B(B[22]), .Ci(CTMP[22]), .S(S[22]), .Co(CTMP[23]) );
  FA_297 FAI_24 ( .A(A[23]), .B(B[23]), .Ci(CTMP[23]), .S(S[23]), .Co(CTMP[24]) );
  FA_296 FAI_25 ( .A(A[24]), .B(B[24]), .Ci(CTMP[24]), .S(S[24]), .Co(CTMP[25]) );
  FA_295 FAI_26 ( .A(A[25]), .B(B[25]), .Ci(CTMP[25]), .S(S[25]), .Co(CTMP[26]) );
  FA_294 FAI_27 ( .A(A[26]), .B(B[26]), .Ci(CTMP[26]), .S(S[26]), .Co(CTMP[27]) );
  FA_293 FAI_28 ( .A(A[27]), .B(B[27]), .Ci(CTMP[27]), .S(S[27]), .Co(CTMP[28]) );
  FA_292 FAI_29 ( .A(A[28]), .B(B[28]), .Ci(CTMP[28]), .S(S[28]), .Co(CTMP[29]) );
  FA_291 FAI_30 ( .A(A[29]), .B(B[29]), .Ci(CTMP[29]), .S(S[29]), .Co(CTMP[30]) );
  FA_290 FAI_31 ( .A(A[30]), .B(B[30]), .Ci(CTMP[30]), .S(S[30]), .Co(CTMP[31]) );
  FA_289 FAI_32 ( .A(A[31]), .B(B[31]), .Ci(CTMP[31]), .S(S[31]), .Co(CTMP[32]) );
  FA_288 FAI_33 ( .A(A[32]), .B(B[32]), .Ci(CTMP[32]), .S(S[32]), .Co(CTMP[33]) );
  FA_287 FAI_34 ( .A(A[33]), .B(B[33]), .Ci(CTMP[33]), .S(S[33]), .Co(CTMP[34]) );
  FA_286 FAI_35 ( .A(A[34]), .B(B[34]), .Ci(CTMP[34]), .S(S[34]), .Co(CTMP[35]) );
  FA_285 FAI_36 ( .A(A[35]), .B(B[35]), .Ci(CTMP[35]), .S(S[35]), .Co(CTMP[36]) );
  FA_284 FAI_37 ( .A(A[36]), .B(B[36]), .Ci(CTMP[36]), .S(S[36]), .Co(CTMP[37]) );
  FA_283 FAI_38 ( .A(A[37]), .B(B[37]), .Ci(CTMP[37]), .S(S[37]), .Co(CTMP[38]) );
  FA_282 FAI_39 ( .A(A[38]), .B(B[38]), .Ci(CTMP[38]), .S(S[38]), .Co(CTMP[39]) );
  FA_281 FAI_40 ( .A(A[39]), .B(B[39]), .Ci(CTMP[39]), .S(S[39]), .Co(CTMP[40]) );
  FA_280 FAI_41 ( .A(A[40]), .B(B[40]), .Ci(CTMP[40]), .S(S[40]), .Co(CTMP[41]) );
  FA_279 FAI_42 ( .A(A[41]), .B(B[41]), .Ci(CTMP[41]), .S(S[41]), .Co(CTMP[42]) );
  FA_278 FAI_43 ( .A(A[42]), .B(B[42]), .Ci(CTMP[42]), .S(S[42]), .Co(CTMP[43]) );
  FA_277 FAI_44 ( .A(A[43]), .B(B[43]), .Ci(CTMP[43]), .S(S[43]), .Co(CTMP[44]) );
  FA_276 FAI_45 ( .A(A[44]), .B(B[44]), .Ci(CTMP[44]), .S(S[44]), .Co(CTMP[45]) );
  FA_275 FAI_46 ( .A(A[45]), .B(B[45]), .Ci(CTMP[45]), .S(S[45]), .Co(CTMP[46]) );
  FA_274 FAI_47 ( .A(A[46]), .B(B[46]), .Ci(CTMP[46]), .S(S[46]), .Co(CTMP[47]) );
  FA_273 FAI_48 ( .A(A[47]), .B(B[47]), .Ci(CTMP[47]), .S(S[47]), .Co(CTMP[48]) );
  FA_272 FAI_49 ( .A(A[48]), .B(B[48]), .Ci(CTMP[48]), .S(S[48]), .Co(CTMP[49]) );
  FA_271 FAI_50 ( .A(A[49]), .B(B[49]), .Ci(CTMP[49]), .S(S[49]), .Co(CTMP[50]) );
  FA_270 FAI_51 ( .A(A[50]), .B(B[50]), .Ci(CTMP[50]), .S(S[50]), .Co(CTMP[51]) );
  FA_269 FAI_52 ( .A(A[51]), .B(B[51]), .Ci(CTMP[51]), .S(S[51]), .Co(CTMP[52]) );
  FA_268 FAI_53 ( .A(A[52]), .B(B[52]), .Ci(CTMP[52]), .S(S[52]), .Co(CTMP[53]) );
  FA_267 FAI_54 ( .A(A[53]), .B(B[53]), .Ci(CTMP[53]), .S(S[53]), .Co(CTMP[54]) );
  FA_266 FAI_55 ( .A(A[54]), .B(B[54]), .Ci(CTMP[54]), .S(S[54]), .Co(CTMP[55]) );
  FA_265 FAI_56 ( .A(A[55]), .B(B[55]), .Ci(CTMP[55]), .S(S[55]), .Co(CTMP[56]) );
  FA_264 FAI_57 ( .A(A[56]), .B(B[56]), .Ci(CTMP[56]), .S(S[56]), .Co(CTMP[57]) );
  FA_263 FAI_58 ( .A(A[57]), .B(B[57]), .Ci(CTMP[57]), .S(S[57]), .Co(CTMP[58]) );
  FA_262 FAI_59 ( .A(A[58]), .B(B[58]), .Ci(CTMP[58]), .S(S[58]), .Co(CTMP[59]) );
  FA_261 FAI_60 ( .A(A[59]), .B(B[59]), .Ci(CTMP[59]), .S(S[59]), .Co(CTMP[60]) );
  FA_260 FAI_61 ( .A(A[60]), .B(B[60]), .Ci(CTMP[60]), .S(S[60]), .Co(CTMP[61]) );
  FA_259 FAI_62 ( .A(A[61]), .B(B[61]), .Ci(CTMP[61]), .S(S[61]), .Co(CTMP[62]) );
  FA_258 FAI_63 ( .A(A[62]), .B(B[62]), .Ci(CTMP[62]), .S(S[62]), .Co(CTMP[63]) );
  FA_257 FAI_64 ( .A(A[63]), .B(B[63]), .Ci(CTMP[63]), .S(S[63]), .Co(Co) );
endmodule


module booth_mul_row_N64_RADIX3_5 ( prevA, prevSum, encoderIn, nextA, nextSum
 );
  input [63:0] prevA;
  input [63:0] prevSum;
  input [2:0] encoderIn;
  output [63:0] nextA;
  output [63:0] nextSum;

  wire   [2:0] encoder_to_mux;
  wire   [63:0] plus2A_s;
  wire   [63:0] minus2A_s;
  wire   [63:0] minus4A_s;
  tri   [63:0] mux_to_adder;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign nextA[0] = 1'b0;

  encoder_N64_RADIX3_5 encoder_1 ( .X(encoderIn), .Z(encoder_to_mux) );
  ShiftnCompl_N64_5 ShiftnCompl_1 ( .plusA(prevA), .plus2A_out({plus2A_s[63:1], 
        SYNOPSYS_UNCONNECTED__0}), .minus2A_out(minus2A_s), .plus4A_out({
        nextA[63:1], SYNOPSYS_UNCONNECTED__1}), .minus4A_out(minus4A_s) );
  MUX_GENERIC_N64_RADIX3_5 mux_1 ( .plusA({plus2A_s[63:1], 1'b0}), .minusA(
        minus2A_s), .plus2A({nextA[63:1], 1'b0}), .minus2A(minus4A_s), .SEL(
        encoder_to_mux), .Y(mux_to_adder) );
  RCA_N64_5 rca_1 ( .A(mux_to_adder), .B(prevSum), .Ci(1'b0), .S(nextSum) );
endmodule


module encoder_N64_RADIX3_4 ( X, Z );
  input [2:0] X;
  output [2:0] Z;
  wire   n5, n7, n8;

  OAI22_X1 U1 ( .A1(n8), .A2(n5), .B1(X[2]), .B2(n7), .ZN(Z[1]) );
  INV_X1 U2 ( .A(X[2]), .ZN(n5) );
  AOI21_X1 U3 ( .B1(n8), .B2(n7), .A(X[2]), .ZN(Z[0]) );
  OAI21_X1 U4 ( .B1(X[1]), .B2(X[0]), .A(n7), .ZN(n8) );
  AND3_X1 U5 ( .A1(X[2]), .A2(n7), .A3(n8), .ZN(Z[2]) );
  NAND2_X1 U6 ( .A1(X[1]), .A2(X[0]), .ZN(n7) );
endmodule


module shifter_N64_8 ( \input , shiftLeftOnePos );
  input [63:0] \input ;
  output [63:0] shiftLeftOnePos;
  wire   \input[62] , \input[61] , \input[60] , \input[59] , \input[58] ,
         \input[57] , \input[56] , \input[55] , \input[54] , \input[53] ,
         \input[52] , \input[51] , \input[50] , \input[49] , \input[48] ,
         \input[47] , \input[46] , \input[45] , \input[44] , \input[43] ,
         \input[42] , \input[41] , \input[40] , \input[39] , \input[38] ,
         \input[37] , \input[36] , \input[35] , \input[34] , \input[33] ,
         \input[32] , \input[31] , \input[30] , \input[29] , \input[28] ,
         \input[27] , \input[26] , \input[25] , \input[24] , \input[23] ,
         \input[22] , \input[21] , \input[20] , \input[19] , \input[18] ,
         \input[17] , \input[16] , \input[15] , \input[14] , \input[13] ,
         \input[12] , \input[11] , \input[10] , \input[9] , \input[8] ,
         \input[7] , \input[6] , \input[5] , \input[4] , \input[3] ,
         \input[2] , \input[1] , \input[0] ;
  assign shiftLeftOnePos[0] = 1'b0;
  assign shiftLeftOnePos[63] = \input[62] ;
  assign \input[62]  = \input  [62];
  assign shiftLeftOnePos[62] = \input[61] ;
  assign \input[61]  = \input  [61];
  assign shiftLeftOnePos[61] = \input[60] ;
  assign \input[60]  = \input  [60];
  assign shiftLeftOnePos[60] = \input[59] ;
  assign \input[59]  = \input  [59];
  assign shiftLeftOnePos[59] = \input[58] ;
  assign \input[58]  = \input  [58];
  assign shiftLeftOnePos[58] = \input[57] ;
  assign \input[57]  = \input  [57];
  assign shiftLeftOnePos[57] = \input[56] ;
  assign \input[56]  = \input  [56];
  assign shiftLeftOnePos[56] = \input[55] ;
  assign \input[55]  = \input  [55];
  assign shiftLeftOnePos[55] = \input[54] ;
  assign \input[54]  = \input  [54];
  assign shiftLeftOnePos[54] = \input[53] ;
  assign \input[53]  = \input  [53];
  assign shiftLeftOnePos[53] = \input[52] ;
  assign \input[52]  = \input  [52];
  assign shiftLeftOnePos[52] = \input[51] ;
  assign \input[51]  = \input  [51];
  assign shiftLeftOnePos[51] = \input[50] ;
  assign \input[50]  = \input  [50];
  assign shiftLeftOnePos[50] = \input[49] ;
  assign \input[49]  = \input  [49];
  assign shiftLeftOnePos[49] = \input[48] ;
  assign \input[48]  = \input  [48];
  assign shiftLeftOnePos[48] = \input[47] ;
  assign \input[47]  = \input  [47];
  assign shiftLeftOnePos[47] = \input[46] ;
  assign \input[46]  = \input  [46];
  assign shiftLeftOnePos[46] = \input[45] ;
  assign \input[45]  = \input  [45];
  assign shiftLeftOnePos[45] = \input[44] ;
  assign \input[44]  = \input  [44];
  assign shiftLeftOnePos[44] = \input[43] ;
  assign \input[43]  = \input  [43];
  assign shiftLeftOnePos[43] = \input[42] ;
  assign \input[42]  = \input  [42];
  assign shiftLeftOnePos[42] = \input[41] ;
  assign \input[41]  = \input  [41];
  assign shiftLeftOnePos[41] = \input[40] ;
  assign \input[40]  = \input  [40];
  assign shiftLeftOnePos[40] = \input[39] ;
  assign \input[39]  = \input  [39];
  assign shiftLeftOnePos[39] = \input[38] ;
  assign \input[38]  = \input  [38];
  assign shiftLeftOnePos[38] = \input[37] ;
  assign \input[37]  = \input  [37];
  assign shiftLeftOnePos[37] = \input[36] ;
  assign \input[36]  = \input  [36];
  assign shiftLeftOnePos[36] = \input[35] ;
  assign \input[35]  = \input  [35];
  assign shiftLeftOnePos[35] = \input[34] ;
  assign \input[34]  = \input  [34];
  assign shiftLeftOnePos[34] = \input[33] ;
  assign \input[33]  = \input  [33];
  assign shiftLeftOnePos[33] = \input[32] ;
  assign \input[32]  = \input  [32];
  assign shiftLeftOnePos[32] = \input[31] ;
  assign \input[31]  = \input  [31];
  assign shiftLeftOnePos[31] = \input[30] ;
  assign \input[30]  = \input  [30];
  assign shiftLeftOnePos[30] = \input[29] ;
  assign \input[29]  = \input  [29];
  assign shiftLeftOnePos[29] = \input[28] ;
  assign \input[28]  = \input  [28];
  assign shiftLeftOnePos[28] = \input[27] ;
  assign \input[27]  = \input  [27];
  assign shiftLeftOnePos[27] = \input[26] ;
  assign \input[26]  = \input  [26];
  assign shiftLeftOnePos[26] = \input[25] ;
  assign \input[25]  = \input  [25];
  assign shiftLeftOnePos[25] = \input[24] ;
  assign \input[24]  = \input  [24];
  assign shiftLeftOnePos[24] = \input[23] ;
  assign \input[23]  = \input  [23];
  assign shiftLeftOnePos[23] = \input[22] ;
  assign \input[22]  = \input  [22];
  assign shiftLeftOnePos[22] = \input[21] ;
  assign \input[21]  = \input  [21];
  assign shiftLeftOnePos[21] = \input[20] ;
  assign \input[20]  = \input  [20];
  assign shiftLeftOnePos[20] = \input[19] ;
  assign \input[19]  = \input  [19];
  assign shiftLeftOnePos[19] = \input[18] ;
  assign \input[18]  = \input  [18];
  assign shiftLeftOnePos[18] = \input[17] ;
  assign \input[17]  = \input  [17];
  assign shiftLeftOnePos[17] = \input[16] ;
  assign \input[16]  = \input  [16];
  assign shiftLeftOnePos[16] = \input[15] ;
  assign \input[15]  = \input  [15];
  assign shiftLeftOnePos[15] = \input[14] ;
  assign \input[14]  = \input  [14];
  assign shiftLeftOnePos[14] = \input[13] ;
  assign \input[13]  = \input  [13];
  assign shiftLeftOnePos[13] = \input[12] ;
  assign \input[12]  = \input  [12];
  assign shiftLeftOnePos[12] = \input[11] ;
  assign \input[11]  = \input  [11];
  assign shiftLeftOnePos[11] = \input[10] ;
  assign \input[10]  = \input  [10];
  assign shiftLeftOnePos[10] = \input[9] ;
  assign \input[9]  = \input  [9];
  assign shiftLeftOnePos[9] = \input[8] ;
  assign \input[8]  = \input  [8];
  assign shiftLeftOnePos[8] = \input[7] ;
  assign \input[7]  = \input  [7];
  assign shiftLeftOnePos[7] = \input[6] ;
  assign \input[6]  = \input  [6];
  assign shiftLeftOnePos[6] = \input[5] ;
  assign \input[5]  = \input  [5];
  assign shiftLeftOnePos[5] = \input[4] ;
  assign \input[4]  = \input  [4];
  assign shiftLeftOnePos[4] = \input[3] ;
  assign \input[3]  = \input  [3];
  assign shiftLeftOnePos[3] = \input[2] ;
  assign \input[2]  = \input  [2];
  assign shiftLeftOnePos[2] = \input[1] ;
  assign \input[1]  = \input  [1];
  assign shiftLeftOnePos[1] = \input[0] ;
  assign \input[0]  = \input  [0];

endmodule


module shifter_N64_7 ( \input , shiftLeftOnePos );
  input [63:0] \input ;
  output [63:0] shiftLeftOnePos;
  wire   \input[62] , \input[61] , \input[60] , \input[59] , \input[58] ,
         \input[57] , \input[56] , \input[55] , \input[54] , \input[53] ,
         \input[52] , \input[51] , \input[50] , \input[49] , \input[48] ,
         \input[47] , \input[46] , \input[45] , \input[44] , \input[43] ,
         \input[42] , \input[41] , \input[40] , \input[39] , \input[38] ,
         \input[37] , \input[36] , \input[35] , \input[34] , \input[33] ,
         \input[32] , \input[31] , \input[30] , \input[29] , \input[28] ,
         \input[27] , \input[26] , \input[25] , \input[24] , \input[23] ,
         \input[22] , \input[21] , \input[20] , \input[19] , \input[18] ,
         \input[17] , \input[16] , \input[15] , \input[14] , \input[13] ,
         \input[12] , \input[11] , \input[10] , \input[9] , \input[8] ,
         \input[7] , \input[6] , \input[5] , \input[4] , \input[3] ,
         \input[2] , \input[1] , \input[0] ;
  assign shiftLeftOnePos[0] = 1'b0;
  assign shiftLeftOnePos[63] = \input[62] ;
  assign \input[62]  = \input  [62];
  assign shiftLeftOnePos[62] = \input[61] ;
  assign \input[61]  = \input  [61];
  assign shiftLeftOnePos[61] = \input[60] ;
  assign \input[60]  = \input  [60];
  assign shiftLeftOnePos[60] = \input[59] ;
  assign \input[59]  = \input  [59];
  assign shiftLeftOnePos[59] = \input[58] ;
  assign \input[58]  = \input  [58];
  assign shiftLeftOnePos[58] = \input[57] ;
  assign \input[57]  = \input  [57];
  assign shiftLeftOnePos[57] = \input[56] ;
  assign \input[56]  = \input  [56];
  assign shiftLeftOnePos[56] = \input[55] ;
  assign \input[55]  = \input  [55];
  assign shiftLeftOnePos[55] = \input[54] ;
  assign \input[54]  = \input  [54];
  assign shiftLeftOnePos[54] = \input[53] ;
  assign \input[53]  = \input  [53];
  assign shiftLeftOnePos[53] = \input[52] ;
  assign \input[52]  = \input  [52];
  assign shiftLeftOnePos[52] = \input[51] ;
  assign \input[51]  = \input  [51];
  assign shiftLeftOnePos[51] = \input[50] ;
  assign \input[50]  = \input  [50];
  assign shiftLeftOnePos[50] = \input[49] ;
  assign \input[49]  = \input  [49];
  assign shiftLeftOnePos[49] = \input[48] ;
  assign \input[48]  = \input  [48];
  assign shiftLeftOnePos[48] = \input[47] ;
  assign \input[47]  = \input  [47];
  assign shiftLeftOnePos[47] = \input[46] ;
  assign \input[46]  = \input  [46];
  assign shiftLeftOnePos[46] = \input[45] ;
  assign \input[45]  = \input  [45];
  assign shiftLeftOnePos[45] = \input[44] ;
  assign \input[44]  = \input  [44];
  assign shiftLeftOnePos[44] = \input[43] ;
  assign \input[43]  = \input  [43];
  assign shiftLeftOnePos[43] = \input[42] ;
  assign \input[42]  = \input  [42];
  assign shiftLeftOnePos[42] = \input[41] ;
  assign \input[41]  = \input  [41];
  assign shiftLeftOnePos[41] = \input[40] ;
  assign \input[40]  = \input  [40];
  assign shiftLeftOnePos[40] = \input[39] ;
  assign \input[39]  = \input  [39];
  assign shiftLeftOnePos[39] = \input[38] ;
  assign \input[38]  = \input  [38];
  assign shiftLeftOnePos[38] = \input[37] ;
  assign \input[37]  = \input  [37];
  assign shiftLeftOnePos[37] = \input[36] ;
  assign \input[36]  = \input  [36];
  assign shiftLeftOnePos[36] = \input[35] ;
  assign \input[35]  = \input  [35];
  assign shiftLeftOnePos[35] = \input[34] ;
  assign \input[34]  = \input  [34];
  assign shiftLeftOnePos[34] = \input[33] ;
  assign \input[33]  = \input  [33];
  assign shiftLeftOnePos[33] = \input[32] ;
  assign \input[32]  = \input  [32];
  assign shiftLeftOnePos[32] = \input[31] ;
  assign \input[31]  = \input  [31];
  assign shiftLeftOnePos[31] = \input[30] ;
  assign \input[30]  = \input  [30];
  assign shiftLeftOnePos[30] = \input[29] ;
  assign \input[29]  = \input  [29];
  assign shiftLeftOnePos[29] = \input[28] ;
  assign \input[28]  = \input  [28];
  assign shiftLeftOnePos[28] = \input[27] ;
  assign \input[27]  = \input  [27];
  assign shiftLeftOnePos[27] = \input[26] ;
  assign \input[26]  = \input  [26];
  assign shiftLeftOnePos[26] = \input[25] ;
  assign \input[25]  = \input  [25];
  assign shiftLeftOnePos[25] = \input[24] ;
  assign \input[24]  = \input  [24];
  assign shiftLeftOnePos[24] = \input[23] ;
  assign \input[23]  = \input  [23];
  assign shiftLeftOnePos[23] = \input[22] ;
  assign \input[22]  = \input  [22];
  assign shiftLeftOnePos[22] = \input[21] ;
  assign \input[21]  = \input  [21];
  assign shiftLeftOnePos[21] = \input[20] ;
  assign \input[20]  = \input  [20];
  assign shiftLeftOnePos[20] = \input[19] ;
  assign \input[19]  = \input  [19];
  assign shiftLeftOnePos[19] = \input[18] ;
  assign \input[18]  = \input  [18];
  assign shiftLeftOnePos[18] = \input[17] ;
  assign \input[17]  = \input  [17];
  assign shiftLeftOnePos[17] = \input[16] ;
  assign \input[16]  = \input  [16];
  assign shiftLeftOnePos[16] = \input[15] ;
  assign \input[15]  = \input  [15];
  assign shiftLeftOnePos[15] = \input[14] ;
  assign \input[14]  = \input  [14];
  assign shiftLeftOnePos[14] = \input[13] ;
  assign \input[13]  = \input  [13];
  assign shiftLeftOnePos[13] = \input[12] ;
  assign \input[12]  = \input  [12];
  assign shiftLeftOnePos[12] = \input[11] ;
  assign \input[11]  = \input  [11];
  assign shiftLeftOnePos[11] = \input[10] ;
  assign \input[10]  = \input  [10];
  assign shiftLeftOnePos[10] = \input[9] ;
  assign \input[9]  = \input  [9];
  assign shiftLeftOnePos[9] = \input[8] ;
  assign \input[8]  = \input  [8];
  assign shiftLeftOnePos[8] = \input[7] ;
  assign \input[7]  = \input  [7];
  assign shiftLeftOnePos[7] = \input[6] ;
  assign \input[6]  = \input  [6];
  assign shiftLeftOnePos[6] = \input[5] ;
  assign \input[5]  = \input  [5];
  assign shiftLeftOnePos[5] = \input[4] ;
  assign \input[4]  = \input  [4];
  assign shiftLeftOnePos[4] = \input[3] ;
  assign \input[3]  = \input  [3];
  assign shiftLeftOnePos[3] = \input[2] ;
  assign \input[2]  = \input  [2];
  assign shiftLeftOnePos[2] = \input[1] ;
  assign \input[1]  = \input  [1];
  assign shiftLeftOnePos[1] = \input[0] ;
  assign \input[0]  = \input  [0];

endmodule


module complementer_N64_8_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n190, n191, n192, n193, n194, n196, n197, n198, n199, n200,
         n202, n203, n204, n206, n207, n208, n210, n211, n212, n213, n214,
         n216, n217, n218, n220, n221, n222, n224, n225, n226, n228, n229,
         n230, n232, n233, n234, n235, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n189, n195,
         n201, n205, n209, n215, n219, n223, n227, n231, n236;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U81 ( .A(n190), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U82 ( .A(n192), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U83 ( .A(n193), .B(B[6]), .Z(DIFF[6]) );
  XOR2_X1 U85 ( .A(n196), .B(B[62]), .Z(DIFF[62]) );
  XOR2_X1 U86 ( .A(n194), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U87 ( .A(n198), .B(B[59]), .Z(DIFF[59]) );
  XOR2_X1 U89 ( .A(n200), .B(B[57]), .Z(DIFF[57]) );
  XOR2_X1 U90 ( .A(n202), .B(B[55]), .Z(DIFF[55]) );
  XOR2_X1 U92 ( .A(n204), .B(B[53]), .Z(DIFF[53]) );
  XOR2_X1 U93 ( .A(n206), .B(B[51]), .Z(DIFF[51]) );
  XOR2_X1 U95 ( .A(n208), .B(B[49]), .Z(DIFF[49]) );
  XOR2_X1 U96 ( .A(n212), .B(B[47]), .Z(DIFF[47]) );
  XOR2_X1 U98 ( .A(n214), .B(B[45]), .Z(DIFF[45]) );
  XOR2_X1 U99 ( .A(n216), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U101 ( .A(n218), .B(B[41]), .Z(DIFF[41]) );
  XOR2_X1 U102 ( .A(n211), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U103 ( .A(n220), .B(B[39]), .Z(DIFF[39]) );
  XOR2_X1 U105 ( .A(n222), .B(B[37]), .Z(DIFF[37]) );
  XOR2_X1 U106 ( .A(n224), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U108 ( .A(n226), .B(B[33]), .Z(DIFF[33]) );
  XOR2_X1 U109 ( .A(n228), .B(B[31]), .Z(DIFF[31]) );
  XOR2_X1 U111 ( .A(n230), .B(B[29]), .Z(DIFF[29]) );
  XOR2_X1 U112 ( .A(n233), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U114 ( .A(n235), .B(B[25]), .Z(DIFF[25]) );
  XOR2_X1 U115 ( .A(n237), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U116 ( .A(n240), .B(B[22]), .Z(DIFF[22]) );
  XOR2_X1 U117 ( .A(n239), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U118 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U119 ( .A(n241), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U120 ( .A(n244), .B(B[18]), .Z(DIFF[18]) );
  XOR2_X1 U121 ( .A(n243), .B(B[17]), .Z(DIFF[17]) );
  XOR2_X1 U122 ( .A(n245), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U123 ( .A(n248), .B(B[14]), .Z(DIFF[14]) );
  XOR2_X1 U124 ( .A(n247), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U125 ( .A(n249), .B(B[11]), .Z(DIFF[11]) );
  XOR2_X1 U126 ( .A(n251), .B(B[10]), .Z(DIFF[10]) );
  XOR2_X1 U1 ( .A(n197), .B(n236), .Z(DIFF[61]) );
  NAND2_X1 U2 ( .A1(n197), .A2(n236), .ZN(n196) );
  XNOR2_X1 U3 ( .A(n189), .B(B[58]), .ZN(DIFF[58]) );
  NOR2_X1 U4 ( .A1(n200), .A2(B[57]), .ZN(n189) );
  NOR3_X1 U5 ( .A1(B[59]), .A2(B[60]), .A3(n198), .ZN(n197) );
  XNOR2_X1 U6 ( .A(B[60]), .B(n199), .ZN(DIFF[60]) );
  NOR2_X1 U7 ( .A1(B[59]), .A2(n198), .ZN(n199) );
  OR3_X1 U8 ( .A1(B[57]), .A2(B[58]), .A3(n200), .ZN(n198) );
  XNOR2_X1 U9 ( .A(B[56]), .B(n203), .ZN(DIFF[56]) );
  NOR2_X1 U10 ( .A1(B[55]), .A2(n202), .ZN(n203) );
  OR3_X1 U11 ( .A1(B[55]), .A2(B[56]), .A3(n202), .ZN(n200) );
  XNOR2_X1 U12 ( .A(n195), .B(B[63]), .ZN(DIFF[63]) );
  NOR2_X1 U13 ( .A1(n196), .A2(B[62]), .ZN(n195) );
  OR3_X1 U14 ( .A1(B[33]), .A2(B[34]), .A3(n226), .ZN(n224) );
  OR3_X1 U15 ( .A1(B[35]), .A2(B[36]), .A3(n224), .ZN(n222) );
  XNOR2_X1 U16 ( .A(n201), .B(B[34]), .ZN(DIFF[34]) );
  NOR2_X1 U17 ( .A1(n226), .A2(B[33]), .ZN(n201) );
  XNOR2_X1 U18 ( .A(n205), .B(B[50]), .ZN(DIFF[50]) );
  NOR2_X1 U19 ( .A1(n208), .A2(B[49]), .ZN(n205) );
  XNOR2_X1 U20 ( .A(n209), .B(B[42]), .ZN(DIFF[42]) );
  NOR2_X1 U21 ( .A1(n218), .A2(B[41]), .ZN(n209) );
  XNOR2_X1 U22 ( .A(B[52]), .B(n207), .ZN(DIFF[52]) );
  NOR2_X1 U23 ( .A1(B[51]), .A2(n206), .ZN(n207) );
  XNOR2_X1 U24 ( .A(B[48]), .B(n213), .ZN(DIFF[48]) );
  NOR2_X1 U25 ( .A1(B[47]), .A2(n212), .ZN(n213) );
  XNOR2_X1 U26 ( .A(B[44]), .B(n217), .ZN(DIFF[44]) );
  NOR2_X1 U27 ( .A1(B[43]), .A2(n216), .ZN(n217) );
  XNOR2_X1 U28 ( .A(B[40]), .B(n221), .ZN(DIFF[40]) );
  NOR2_X1 U29 ( .A1(B[39]), .A2(n220), .ZN(n221) );
  XNOR2_X1 U30 ( .A(B[36]), .B(n225), .ZN(DIFF[36]) );
  NOR2_X1 U31 ( .A1(B[35]), .A2(n224), .ZN(n225) );
  OR3_X1 U32 ( .A1(B[37]), .A2(B[38]), .A3(n222), .ZN(n220) );
  OR3_X1 U33 ( .A1(B[41]), .A2(B[42]), .A3(n218), .ZN(n216) );
  OR3_X1 U34 ( .A1(B[45]), .A2(B[46]), .A3(n214), .ZN(n212) );
  OR3_X1 U35 ( .A1(B[49]), .A2(B[50]), .A3(n208), .ZN(n206) );
  OR3_X1 U36 ( .A1(B[53]), .A2(B[54]), .A3(n204), .ZN(n202) );
  OR3_X1 U37 ( .A1(B[39]), .A2(B[40]), .A3(n220), .ZN(n218) );
  OR3_X1 U38 ( .A1(B[43]), .A2(B[44]), .A3(n216), .ZN(n214) );
  OR3_X1 U39 ( .A1(B[47]), .A2(B[48]), .A3(n212), .ZN(n208) );
  OR3_X1 U40 ( .A1(B[51]), .A2(B[52]), .A3(n206), .ZN(n204) );
  XNOR2_X1 U41 ( .A(n215), .B(B[54]), .ZN(DIFF[54]) );
  NOR2_X1 U42 ( .A1(n204), .A2(B[53]), .ZN(n215) );
  XNOR2_X1 U43 ( .A(n219), .B(B[46]), .ZN(DIFF[46]) );
  NOR2_X1 U44 ( .A1(n214), .A2(B[45]), .ZN(n219) );
  XNOR2_X1 U45 ( .A(n223), .B(B[38]), .ZN(DIFF[38]) );
  NOR2_X1 U46 ( .A1(n222), .A2(B[37]), .ZN(n223) );
  XNOR2_X1 U47 ( .A(B[32]), .B(n229), .ZN(DIFF[32]) );
  NOR2_X1 U48 ( .A1(B[31]), .A2(n228), .ZN(n229) );
  OR3_X1 U49 ( .A1(B[31]), .A2(B[32]), .A3(n228), .ZN(n226) );
  OR3_X1 U50 ( .A1(B[29]), .A2(B[30]), .A3(n230), .ZN(n228) );
  XNOR2_X1 U51 ( .A(n227), .B(B[30]), .ZN(DIFF[30]) );
  NOR2_X1 U52 ( .A1(n230), .A2(B[29]), .ZN(n227) );
  XNOR2_X1 U53 ( .A(B[28]), .B(n234), .ZN(DIFF[28]) );
  NOR2_X1 U54 ( .A1(B[27]), .A2(n233), .ZN(n234) );
  OR3_X1 U55 ( .A1(B[27]), .A2(B[28]), .A3(n233), .ZN(n230) );
  OR3_X1 U56 ( .A1(B[25]), .A2(B[26]), .A3(n235), .ZN(n233) );
  XNOR2_X1 U57 ( .A(n231), .B(B[26]), .ZN(DIFF[26]) );
  NOR2_X1 U58 ( .A1(n235), .A2(B[25]), .ZN(n231) );
  OR3_X1 U59 ( .A1(B[23]), .A2(B[24]), .A3(n237), .ZN(n235) );
  XNOR2_X1 U60 ( .A(B[24]), .B(n238), .ZN(DIFF[24]) );
  NOR2_X1 U61 ( .A1(B[23]), .A2(n237), .ZN(n238) );
  NOR2_X1 U62 ( .A1(B[19]), .A2(n241), .ZN(n242) );
  NOR2_X1 U63 ( .A1(B[15]), .A2(n245), .ZN(n246) );
  NOR2_X1 U64 ( .A1(B[11]), .A2(n249), .ZN(n250) );
  NOR2_X1 U65 ( .A1(B[7]), .A2(n192), .ZN(n191) );
  NOR2_X1 U66 ( .A1(B[3]), .A2(n211), .ZN(n210) );
  OR3_X1 U67 ( .A1(B[21]), .A2(B[22]), .A3(n239), .ZN(n237) );
  OR3_X1 U68 ( .A1(B[17]), .A2(B[18]), .A3(n243), .ZN(n241) );
  OR3_X1 U69 ( .A1(B[13]), .A2(B[14]), .A3(n247), .ZN(n245) );
  OR3_X1 U70 ( .A1(B[10]), .A2(B[9]), .A3(n190), .ZN(n249) );
  OR3_X1 U71 ( .A1(B[5]), .A2(B[6]), .A3(n194), .ZN(n192) );
  OR3_X1 U72 ( .A1(B[19]), .A2(B[20]), .A3(n241), .ZN(n239) );
  OR3_X1 U73 ( .A1(B[15]), .A2(B[16]), .A3(n245), .ZN(n243) );
  OR3_X1 U74 ( .A1(B[11]), .A2(B[12]), .A3(n249), .ZN(n247) );
  OR3_X1 U75 ( .A1(B[7]), .A2(B[8]), .A3(n192), .ZN(n190) );
  OR3_X1 U76 ( .A1(B[3]), .A2(B[4]), .A3(n211), .ZN(n194) );
  XNOR2_X1 U77 ( .A(B[20]), .B(n242), .ZN(DIFF[20]) );
  XNOR2_X1 U78 ( .A(B[16]), .B(n246), .ZN(DIFF[16]) );
  XNOR2_X1 U79 ( .A(B[12]), .B(n250), .ZN(DIFF[12]) );
  XNOR2_X1 U80 ( .A(B[8]), .B(n191), .ZN(DIFF[8]) );
  XNOR2_X1 U84 ( .A(B[4]), .B(n210), .ZN(DIFF[4]) );
  XNOR2_X1 U88 ( .A(B[2]), .B(n232), .ZN(DIFF[2]) );
  OR2_X1 U91 ( .A1(n239), .A2(B[21]), .ZN(n240) );
  OR2_X1 U94 ( .A1(n243), .A2(B[17]), .ZN(n244) );
  OR2_X1 U97 ( .A1(n247), .A2(B[13]), .ZN(n248) );
  OR2_X1 U100 ( .A1(n190), .A2(B[9]), .ZN(n251) );
  OR2_X1 U104 ( .A1(n194), .A2(B[5]), .ZN(n193) );
  OR3_X1 U107 ( .A1(B[1]), .A2(B[2]), .A3(\B[0] ), .ZN(n211) );
  NOR2_X1 U110 ( .A1(\B[0] ), .A2(B[1]), .ZN(n232) );
  INV_X1 U113 ( .A(B[61]), .ZN(n236) );
endmodule


module complementer_N64_8 ( \input , complement2 );
  input [63:0] \input ;
  output [63:0] complement2;


  complementer_N64_8_DW01_sub_0 sub_add_31_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(\input ), .CI(1'b0), .DIFF(complement2) );
endmodule


module complementer_N64_7_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n190, n191, n192, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n241, n242, n243, n245, n246,
         n247, n249, n250, n189, n193, n240, n244, n248, n251;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U81 ( .A(n190), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U82 ( .A(n192), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U84 ( .A(n195), .B(B[63]), .Z(DIFF[63]) );
  XOR2_X1 U85 ( .A(n196), .B(B[62]), .Z(DIFF[62]) );
  XOR2_X1 U86 ( .A(n194), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U87 ( .A(n198), .B(B[59]), .Z(DIFF[59]) );
  XOR2_X1 U88 ( .A(n201), .B(B[58]), .Z(DIFF[58]) );
  XOR2_X1 U89 ( .A(n200), .B(B[57]), .Z(DIFF[57]) );
  XOR2_X1 U90 ( .A(n202), .B(B[55]), .Z(DIFF[55]) );
  XOR2_X1 U91 ( .A(n205), .B(B[54]), .Z(DIFF[54]) );
  XOR2_X1 U92 ( .A(n204), .B(B[53]), .Z(DIFF[53]) );
  XOR2_X1 U93 ( .A(n206), .B(B[51]), .Z(DIFF[51]) );
  XOR2_X1 U94 ( .A(n209), .B(B[50]), .Z(DIFF[50]) );
  XOR2_X1 U95 ( .A(n208), .B(B[49]), .Z(DIFF[49]) );
  XOR2_X1 U96 ( .A(n212), .B(B[47]), .Z(DIFF[47]) );
  XOR2_X1 U97 ( .A(n215), .B(B[46]), .Z(DIFF[46]) );
  XOR2_X1 U98 ( .A(n214), .B(B[45]), .Z(DIFF[45]) );
  XOR2_X1 U99 ( .A(n216), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U100 ( .A(n219), .B(B[42]), .Z(DIFF[42]) );
  XOR2_X1 U101 ( .A(n218), .B(B[41]), .Z(DIFF[41]) );
  XOR2_X1 U102 ( .A(n211), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U103 ( .A(n220), .B(B[39]), .Z(DIFF[39]) );
  XOR2_X1 U104 ( .A(n223), .B(B[38]), .Z(DIFF[38]) );
  XOR2_X1 U105 ( .A(n222), .B(B[37]), .Z(DIFF[37]) );
  XOR2_X1 U106 ( .A(n224), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U107 ( .A(n227), .B(B[34]), .Z(DIFF[34]) );
  XOR2_X1 U108 ( .A(n226), .B(B[33]), .Z(DIFF[33]) );
  XOR2_X1 U109 ( .A(n228), .B(B[31]), .Z(DIFF[31]) );
  XOR2_X1 U110 ( .A(n231), .B(B[30]), .Z(DIFF[30]) );
  XOR2_X1 U111 ( .A(n230), .B(B[29]), .Z(DIFF[29]) );
  XOR2_X1 U112 ( .A(n233), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U113 ( .A(n236), .B(B[26]), .Z(DIFF[26]) );
  XOR2_X1 U114 ( .A(n235), .B(B[25]), .Z(DIFF[25]) );
  XOR2_X1 U115 ( .A(n237), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U117 ( .A(n239), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U118 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U119 ( .A(n241), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U121 ( .A(n243), .B(B[17]), .Z(DIFF[17]) );
  XOR2_X1 U122 ( .A(n245), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U124 ( .A(n247), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U125 ( .A(n249), .B(B[11]), .Z(DIFF[11]) );
  NAND2_X1 U1 ( .A1(n197), .A2(n251), .ZN(n196) );
  NOR3_X1 U2 ( .A1(B[59]), .A2(B[60]), .A3(n198), .ZN(n197) );
  NOR2_X1 U3 ( .A1(B[59]), .A2(n198), .ZN(n199) );
  OR2_X1 U4 ( .A1(n196), .A2(B[62]), .ZN(n195) );
  OR3_X1 U5 ( .A1(B[57]), .A2(B[58]), .A3(n200), .ZN(n198) );
  OR2_X1 U6 ( .A1(n200), .A2(B[57]), .ZN(n201) );
  OR3_X1 U7 ( .A1(B[33]), .A2(B[34]), .A3(n226), .ZN(n224) );
  OR3_X1 U8 ( .A1(B[35]), .A2(B[36]), .A3(n224), .ZN(n222) );
  NOR2_X1 U9 ( .A1(B[51]), .A2(n206), .ZN(n207) );
  NOR2_X1 U10 ( .A1(B[47]), .A2(n212), .ZN(n213) );
  NOR2_X1 U11 ( .A1(B[43]), .A2(n216), .ZN(n217) );
  NOR2_X1 U12 ( .A1(B[39]), .A2(n220), .ZN(n221) );
  NOR2_X1 U13 ( .A1(B[35]), .A2(n224), .ZN(n225) );
  OR3_X1 U14 ( .A1(B[53]), .A2(B[54]), .A3(n204), .ZN(n202) );
  OR3_X1 U15 ( .A1(B[49]), .A2(B[50]), .A3(n208), .ZN(n206) );
  OR3_X1 U16 ( .A1(B[45]), .A2(B[46]), .A3(n214), .ZN(n212) );
  OR3_X1 U17 ( .A1(B[41]), .A2(B[42]), .A3(n218), .ZN(n216) );
  OR3_X1 U18 ( .A1(B[37]), .A2(B[38]), .A3(n222), .ZN(n220) );
  OR3_X1 U19 ( .A1(B[51]), .A2(B[52]), .A3(n206), .ZN(n204) );
  OR3_X1 U20 ( .A1(B[47]), .A2(B[48]), .A3(n212), .ZN(n208) );
  OR3_X1 U21 ( .A1(B[43]), .A2(B[44]), .A3(n216), .ZN(n214) );
  OR3_X1 U22 ( .A1(B[39]), .A2(B[40]), .A3(n220), .ZN(n218) );
  OR2_X1 U23 ( .A1(n204), .A2(B[53]), .ZN(n205) );
  OR2_X1 U24 ( .A1(n208), .A2(B[49]), .ZN(n209) );
  OR2_X1 U25 ( .A1(n214), .A2(B[45]), .ZN(n215) );
  OR2_X1 U26 ( .A1(n218), .A2(B[41]), .ZN(n219) );
  OR2_X1 U27 ( .A1(n222), .A2(B[37]), .ZN(n223) );
  OR2_X1 U28 ( .A1(n226), .A2(B[33]), .ZN(n227) );
  NOR2_X1 U29 ( .A1(B[55]), .A2(n202), .ZN(n203) );
  OR3_X1 U30 ( .A1(B[55]), .A2(B[56]), .A3(n202), .ZN(n200) );
  OR3_X1 U31 ( .A1(B[31]), .A2(B[32]), .A3(n228), .ZN(n226) );
  NOR2_X1 U32 ( .A1(B[31]), .A2(n228), .ZN(n229) );
  OR3_X1 U33 ( .A1(B[29]), .A2(B[30]), .A3(n230), .ZN(n228) );
  XNOR2_X1 U34 ( .A(B[32]), .B(n229), .ZN(DIFF[32]) );
  XNOR2_X1 U35 ( .A(B[28]), .B(n234), .ZN(DIFF[28]) );
  OR2_X1 U36 ( .A1(n230), .A2(B[29]), .ZN(n231) );
  XNOR2_X1 U37 ( .A(B[52]), .B(n207), .ZN(DIFF[52]) );
  XNOR2_X1 U38 ( .A(B[48]), .B(n213), .ZN(DIFF[48]) );
  XNOR2_X1 U39 ( .A(B[44]), .B(n217), .ZN(DIFF[44]) );
  XNOR2_X1 U40 ( .A(B[40]), .B(n221), .ZN(DIFF[40]) );
  XNOR2_X1 U41 ( .A(B[36]), .B(n225), .ZN(DIFF[36]) );
  XNOR2_X1 U42 ( .A(B[56]), .B(n203), .ZN(DIFF[56]) );
  XNOR2_X1 U43 ( .A(n197), .B(B[61]), .ZN(DIFF[61]) );
  XNOR2_X1 U44 ( .A(B[60]), .B(n199), .ZN(DIFF[60]) );
  NOR2_X1 U45 ( .A1(B[27]), .A2(n233), .ZN(n234) );
  OR3_X1 U46 ( .A1(B[27]), .A2(B[28]), .A3(n233), .ZN(n230) );
  OR3_X1 U47 ( .A1(B[25]), .A2(B[26]), .A3(n235), .ZN(n233) );
  OR2_X1 U48 ( .A1(n235), .A2(B[25]), .ZN(n236) );
  XNOR2_X1 U49 ( .A(B[24]), .B(n238), .ZN(DIFF[24]) );
  XNOR2_X1 U50 ( .A(n189), .B(B[22]), .ZN(DIFF[22]) );
  NOR2_X1 U51 ( .A1(n239), .A2(B[21]), .ZN(n189) );
  XNOR2_X1 U52 ( .A(n193), .B(B[18]), .ZN(DIFF[18]) );
  NOR2_X1 U53 ( .A1(n243), .A2(B[17]), .ZN(n193) );
  XNOR2_X1 U54 ( .A(n240), .B(B[14]), .ZN(DIFF[14]) );
  NOR2_X1 U55 ( .A1(n247), .A2(B[13]), .ZN(n240) );
  XNOR2_X1 U56 ( .A(n244), .B(B[10]), .ZN(DIFF[10]) );
  NOR2_X1 U57 ( .A1(n190), .A2(B[9]), .ZN(n244) );
  XNOR2_X1 U58 ( .A(n248), .B(B[6]), .ZN(DIFF[6]) );
  NOR2_X1 U59 ( .A1(n194), .A2(B[5]), .ZN(n248) );
  NOR2_X1 U60 ( .A1(B[23]), .A2(n237), .ZN(n238) );
  XNOR2_X1 U61 ( .A(B[20]), .B(n242), .ZN(DIFF[20]) );
  NOR2_X1 U62 ( .A1(B[19]), .A2(n241), .ZN(n242) );
  XNOR2_X1 U63 ( .A(B[16]), .B(n246), .ZN(DIFF[16]) );
  NOR2_X1 U64 ( .A1(B[15]), .A2(n245), .ZN(n246) );
  XNOR2_X1 U65 ( .A(B[12]), .B(n250), .ZN(DIFF[12]) );
  NOR2_X1 U66 ( .A1(B[11]), .A2(n249), .ZN(n250) );
  XNOR2_X1 U67 ( .A(B[8]), .B(n191), .ZN(DIFF[8]) );
  NOR2_X1 U68 ( .A1(B[7]), .A2(n192), .ZN(n191) );
  XNOR2_X1 U69 ( .A(B[2]), .B(n232), .ZN(DIFF[2]) );
  NOR2_X1 U70 ( .A1(\B[0] ), .A2(B[1]), .ZN(n232) );
  XNOR2_X1 U71 ( .A(B[4]), .B(n210), .ZN(DIFF[4]) );
  NOR2_X1 U72 ( .A1(B[3]), .A2(n211), .ZN(n210) );
  OR3_X1 U73 ( .A1(B[5]), .A2(B[6]), .A3(n194), .ZN(n192) );
  OR3_X1 U74 ( .A1(B[10]), .A2(B[9]), .A3(n190), .ZN(n249) );
  OR3_X1 U75 ( .A1(B[13]), .A2(B[14]), .A3(n247), .ZN(n245) );
  OR3_X1 U76 ( .A1(B[17]), .A2(B[18]), .A3(n243), .ZN(n241) );
  OR3_X1 U77 ( .A1(B[21]), .A2(B[22]), .A3(n239), .ZN(n237) );
  OR3_X1 U78 ( .A1(B[7]), .A2(B[8]), .A3(n192), .ZN(n190) );
  OR3_X1 U79 ( .A1(B[11]), .A2(B[12]), .A3(n249), .ZN(n247) );
  OR3_X1 U80 ( .A1(B[15]), .A2(B[16]), .A3(n245), .ZN(n243) );
  OR3_X1 U83 ( .A1(B[19]), .A2(B[20]), .A3(n241), .ZN(n239) );
  OR3_X1 U116 ( .A1(B[23]), .A2(B[24]), .A3(n237), .ZN(n235) );
  OR3_X1 U120 ( .A1(B[3]), .A2(B[4]), .A3(n211), .ZN(n194) );
  OR3_X1 U123 ( .A1(B[1]), .A2(B[2]), .A3(\B[0] ), .ZN(n211) );
  INV_X1 U126 ( .A(B[61]), .ZN(n251) );
endmodule


module complementer_N64_7 ( \input , complement2 );
  input [63:0] \input ;
  output [63:0] complement2;


  complementer_N64_7_DW01_sub_0 sub_add_31_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(\input ), .CI(1'b0), .DIFF(complement2) );
endmodule


module ShiftnCompl_N64_4 ( plusA, plus2A_out, minus2A_out, plus4A_out, 
        minus4A_out );
  input [63:0] plusA;
  output [63:0] plus2A_out;
  output [63:0] minus2A_out;
  output [63:0] plus4A_out;
  output [63:0] minus4A_out;
  wire   n3, n4;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign plus2A_out[0] = 1'b0;
  assign plus4A_out[0] = 1'b0;

  shifter_N64_8 shifter_1 ( .\input (plusA), .shiftLeftOnePos({
        plus2A_out[63:59], n3, plus2A_out[57:1], SYNOPSYS_UNCONNECTED__0}) );
  shifter_N64_7 shifter_2 ( .\input ({plus2A_out[63:1], 1'b0}), 
        .shiftLeftOnePos({plus4A_out[63:59], n4, plus4A_out[57:1], 
        SYNOPSYS_UNCONNECTED__1}) );
  complementer_N64_8 complementer_1 ( .\input ({plus2A_out[63:1], 1'b0}), 
        .complement2(minus2A_out) );
  complementer_N64_7 complementer_2 ( .\input ({plus4A_out[63:1], 1'b0}), 
        .complement2(minus4A_out) );
  BUF_X1 U3 ( .A(n4), .Z(plus4A_out[58]) );
  BUF_X1 U4 ( .A(n3), .Z(plus2A_out[58]) );
endmodule


module MUX_GENERIC_N64_RADIX3_4 ( plusA, minusA, plus2A, minus2A, SEL, Y );
  input [63:0] plusA;
  input [63:0] minusA;
  input [63:0] plus2A;
  input [63:0] minus2A;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502;
  tri   [63:0] Y;

  TBUF_X1 \Y_tri[59]  ( .A(n442), .EN(n301), .Z(Y[59]) );
  TBUF_X1 \Y_tri[60]  ( .A(n441), .EN(n301), .Z(Y[60]) );
  TBUF_X1 \Y_tri[61]  ( .A(n440), .EN(n301), .Z(Y[61]) );
  TBUF_X1 \Y_tri[62]  ( .A(n439), .EN(n301), .Z(Y[62]) );
  TBUF_X1 \Y_tri[63]  ( .A(n438), .EN(n301), .Z(Y[63]) );
  TBUF_X1 \Y_tri[55]  ( .A(n446), .EN(n301), .Z(Y[55]) );
  TBUF_X1 \Y_tri[56]  ( .A(n445), .EN(n301), .Z(Y[56]) );
  TBUF_X1 \Y_tri[57]  ( .A(n444), .EN(n301), .Z(Y[57]) );
  TBUF_X1 \Y_tri[58]  ( .A(n443), .EN(n301), .Z(Y[58]) );
  TBUF_X1 \Y_tri[35]  ( .A(n466), .EN(n299), .Z(Y[35]) );
  TBUF_X1 \Y_tri[36]  ( .A(n465), .EN(n299), .Z(Y[36]) );
  TBUF_X1 \Y_tri[38]  ( .A(n463), .EN(n299), .Z(Y[38]) );
  TBUF_X1 \Y_tri[39]  ( .A(n462), .EN(n299), .Z(Y[39]) );
  TBUF_X1 \Y_tri[40]  ( .A(n461), .EN(n299), .Z(Y[40]) );
  TBUF_X1 \Y_tri[41]  ( .A(n460), .EN(n299), .Z(Y[41]) );
  TBUF_X1 \Y_tri[42]  ( .A(n459), .EN(n299), .Z(Y[42]) );
  TBUF_X1 \Y_tri[43]  ( .A(n458), .EN(n299), .Z(Y[43]) );
  TBUF_X1 \Y_tri[44]  ( .A(n457), .EN(n300), .Z(Y[44]) );
  TBUF_X1 \Y_tri[45]  ( .A(n456), .EN(n300), .Z(Y[45]) );
  TBUF_X1 \Y_tri[46]  ( .A(n455), .EN(n300), .Z(Y[46]) );
  TBUF_X1 \Y_tri[47]  ( .A(n454), .EN(n300), .Z(Y[47]) );
  TBUF_X1 \Y_tri[48]  ( .A(n453), .EN(n300), .Z(Y[48]) );
  TBUF_X1 \Y_tri[49]  ( .A(n452), .EN(n300), .Z(Y[49]) );
  TBUF_X1 \Y_tri[50]  ( .A(n451), .EN(n300), .Z(Y[50]) );
  TBUF_X1 \Y_tri[51]  ( .A(n450), .EN(n300), .Z(Y[51]) );
  TBUF_X1 \Y_tri[52]  ( .A(n449), .EN(n300), .Z(Y[52]) );
  TBUF_X1 \Y_tri[53]  ( .A(n448), .EN(n300), .Z(Y[53]) );
  TBUF_X1 \Y_tri[54]  ( .A(n447), .EN(n300), .Z(Y[54]) );
  TBUF_X1 \Y_tri[14]  ( .A(n487), .EN(n297), .Z(Y[14]) );
  TBUF_X1 \Y_tri[15]  ( .A(n486), .EN(n297), .Z(Y[15]) );
  TBUF_X1 \Y_tri[16]  ( .A(n485), .EN(n297), .Z(Y[16]) );
  TBUF_X1 \Y_tri[17]  ( .A(n484), .EN(n297), .Z(Y[17]) );
  TBUF_X1 \Y_tri[18]  ( .A(n483), .EN(n297), .Z(Y[18]) );
  TBUF_X1 \Y_tri[19]  ( .A(n482), .EN(n297), .Z(Y[19]) );
  TBUF_X1 \Y_tri[20]  ( .A(n481), .EN(n297), .Z(Y[20]) );
  TBUF_X1 \Y_tri[21]  ( .A(n480), .EN(n297), .Z(Y[21]) );
  TBUF_X1 \Y_tri[22]  ( .A(n479), .EN(n298), .Z(Y[22]) );
  TBUF_X1 \Y_tri[23]  ( .A(n478), .EN(n298), .Z(Y[23]) );
  TBUF_X1 \Y_tri[24]  ( .A(n477), .EN(n298), .Z(Y[24]) );
  TBUF_X1 \Y_tri[25]  ( .A(n476), .EN(n298), .Z(Y[25]) );
  TBUF_X1 \Y_tri[26]  ( .A(n475), .EN(n298), .Z(Y[26]) );
  TBUF_X1 \Y_tri[27]  ( .A(n474), .EN(n298), .Z(Y[27]) );
  TBUF_X1 \Y_tri[28]  ( .A(n473), .EN(n298), .Z(Y[28]) );
  TBUF_X1 \Y_tri[29]  ( .A(n472), .EN(n298), .Z(Y[29]) );
  TBUF_X1 \Y_tri[30]  ( .A(n471), .EN(n298), .Z(Y[30]) );
  TBUF_X1 \Y_tri[31]  ( .A(n470), .EN(n298), .Z(Y[31]) );
  TBUF_X1 \Y_tri[32]  ( .A(n469), .EN(n298), .Z(Y[32]) );
  TBUF_X1 \Y_tri[33]  ( .A(n468), .EN(n299), .Z(Y[33]) );
  TBUF_X1 \Y_tri[34]  ( .A(n467), .EN(n299), .Z(Y[34]) );
  TBUF_X1 \Y_tri[3]  ( .A(n499), .EN(n296), .Z(Y[3]) );
  TBUF_X1 \Y_tri[4]  ( .A(n498), .EN(n296), .Z(Y[4]) );
  TBUF_X1 \Y_tri[5]  ( .A(n497), .EN(n296), .Z(Y[5]) );
  TBUF_X1 \Y_tri[6]  ( .A(n496), .EN(n296), .Z(Y[6]) );
  TBUF_X1 \Y_tri[7]  ( .A(n495), .EN(n296), .Z(Y[7]) );
  TBUF_X1 \Y_tri[8]  ( .A(n494), .EN(n296), .Z(Y[8]) );
  TBUF_X1 \Y_tri[9]  ( .A(n492), .EN(n296), .Z(Y[9]) );
  TBUF_X1 \Y_tri[10]  ( .A(n491), .EN(n296), .Z(Y[10]) );
  TBUF_X1 \Y_tri[11]  ( .A(n490), .EN(n297), .Z(Y[11]) );
  TBUF_X1 \Y_tri[12]  ( .A(n489), .EN(n297), .Z(Y[12]) );
  TBUF_X1 \Y_tri[13]  ( .A(n488), .EN(n297), .Z(Y[13]) );
  TBUF_X1 \Y_tri[0]  ( .A(n502), .EN(n296), .Z(Y[0]) );
  TBUF_X1 \Y_tri[1]  ( .A(n501), .EN(n296), .Z(Y[1]) );
  TBUF_X1 \Y_tri[2]  ( .A(n500), .EN(n296), .Z(Y[2]) );
  TBUF_X1 \Y_tri[37]  ( .A(n464), .EN(n299), .Z(Y[37]) );
  NAND2_X1 U2 ( .A1(n375), .A2(n374), .ZN(n467) );
  AOI22_X1 U3 ( .A1(plusA[34]), .A2(n280), .B1(plus2A[34]), .B2(n274), .ZN(
        n375) );
  AOI22_X1 U4 ( .A1(minus2A[34]), .A2(n292), .B1(minusA[34]), .B2(n286), .ZN(
        n374) );
  NAND2_X1 U5 ( .A1(n367), .A2(n366), .ZN(n471) );
  AOI22_X1 U6 ( .A1(plusA[30]), .A2(n280), .B1(plus2A[30]), .B2(n274), .ZN(
        n367) );
  AOI22_X1 U7 ( .A1(minus2A[30]), .A2(n292), .B1(minusA[30]), .B2(n286), .ZN(
        n366) );
  NAND2_X1 U8 ( .A1(n371), .A2(n370), .ZN(n469) );
  AOI22_X1 U9 ( .A1(plusA[32]), .A2(n280), .B1(plus2A[32]), .B2(n274), .ZN(
        n371) );
  AOI22_X1 U10 ( .A1(minus2A[32]), .A2(n292), .B1(minusA[32]), .B2(n286), .ZN(
        n370) );
  NAND2_X1 U11 ( .A1(n363), .A2(n362), .ZN(n473) );
  AOI22_X1 U12 ( .A1(plusA[28]), .A2(n280), .B1(plus2A[28]), .B2(n274), .ZN(
        n363) );
  AOI22_X1 U13 ( .A1(minus2A[28]), .A2(n292), .B1(minusA[28]), .B2(n286), .ZN(
        n362) );
  NAND2_X1 U14 ( .A1(n369), .A2(n368), .ZN(n470) );
  AOI22_X1 U15 ( .A1(plusA[31]), .A2(n280), .B1(plus2A[31]), .B2(n274), .ZN(
        n369) );
  AOI22_X1 U16 ( .A1(minus2A[31]), .A2(n292), .B1(minusA[31]), .B2(n286), .ZN(
        n368) );
  NAND2_X1 U17 ( .A1(n381), .A2(n380), .ZN(n464) );
  AOI22_X1 U18 ( .A1(plusA[37]), .A2(n281), .B1(plus2A[37]), .B2(n275), .ZN(
        n381) );
  AOI22_X1 U19 ( .A1(minus2A[37]), .A2(n293), .B1(minusA[37]), .B2(n287), .ZN(
        n380) );
  NAND2_X1 U20 ( .A1(n373), .A2(n372), .ZN(n468) );
  AOI22_X1 U21 ( .A1(plusA[33]), .A2(n280), .B1(plus2A[33]), .B2(n274), .ZN(
        n373) );
  AOI22_X1 U22 ( .A1(minus2A[33]), .A2(n292), .B1(minusA[33]), .B2(n286), .ZN(
        n372) );
  NAND2_X1 U23 ( .A1(n365), .A2(n364), .ZN(n472) );
  AOI22_X1 U24 ( .A1(plusA[29]), .A2(n280), .B1(plus2A[29]), .B2(n274), .ZN(
        n365) );
  AOI22_X1 U25 ( .A1(minus2A[29]), .A2(n292), .B1(minusA[29]), .B2(n286), .ZN(
        n364) );
  NAND2_X1 U26 ( .A1(n415), .A2(n414), .ZN(n447) );
  AOI22_X1 U27 ( .A1(plusA[54]), .A2(n282), .B1(plus2A[54]), .B2(n276), .ZN(
        n415) );
  AOI22_X1 U28 ( .A1(minus2A[54]), .A2(n294), .B1(minusA[54]), .B2(n288), .ZN(
        n414) );
  NAND2_X1 U29 ( .A1(n407), .A2(n406), .ZN(n451) );
  AOI22_X1 U30 ( .A1(plusA[50]), .A2(n282), .B1(plus2A[50]), .B2(n276), .ZN(
        n407) );
  AOI22_X1 U31 ( .A1(minus2A[50]), .A2(n294), .B1(minusA[50]), .B2(n288), .ZN(
        n406) );
  NAND2_X1 U32 ( .A1(n399), .A2(n398), .ZN(n455) );
  AOI22_X1 U33 ( .A1(plusA[46]), .A2(n281), .B1(plus2A[46]), .B2(n275), .ZN(
        n399) );
  AOI22_X1 U34 ( .A1(minus2A[46]), .A2(n293), .B1(minusA[46]), .B2(n287), .ZN(
        n398) );
  NAND2_X1 U35 ( .A1(n391), .A2(n390), .ZN(n459) );
  AOI22_X1 U36 ( .A1(plusA[42]), .A2(n281), .B1(plus2A[42]), .B2(n275), .ZN(
        n391) );
  AOI22_X1 U37 ( .A1(minus2A[42]), .A2(n293), .B1(minusA[42]), .B2(n287), .ZN(
        n390) );
  NAND2_X1 U38 ( .A1(n383), .A2(n382), .ZN(n463) );
  AOI22_X1 U39 ( .A1(plusA[38]), .A2(n281), .B1(plus2A[38]), .B2(n275), .ZN(
        n383) );
  AOI22_X1 U40 ( .A1(minus2A[38]), .A2(n293), .B1(minusA[38]), .B2(n287), .ZN(
        n382) );
  NAND2_X1 U41 ( .A1(n417), .A2(n416), .ZN(n446) );
  AOI22_X1 U42 ( .A1(plusA[55]), .A2(n282), .B1(plus2A[55]), .B2(n276), .ZN(
        n417) );
  AOI22_X1 U43 ( .A1(minus2A[55]), .A2(n294), .B1(minusA[55]), .B2(n288), .ZN(
        n416) );
  NAND2_X1 U44 ( .A1(n411), .A2(n410), .ZN(n449) );
  AOI22_X1 U45 ( .A1(plusA[52]), .A2(n282), .B1(plus2A[52]), .B2(n276), .ZN(
        n411) );
  AOI22_X1 U46 ( .A1(minus2A[52]), .A2(n294), .B1(minusA[52]), .B2(n288), .ZN(
        n410) );
  NAND2_X1 U47 ( .A1(n403), .A2(n402), .ZN(n453) );
  AOI22_X1 U48 ( .A1(plusA[48]), .A2(n282), .B1(plus2A[48]), .B2(n276), .ZN(
        n403) );
  AOI22_X1 U49 ( .A1(minus2A[48]), .A2(n294), .B1(minusA[48]), .B2(n288), .ZN(
        n402) );
  NAND2_X1 U50 ( .A1(n395), .A2(n394), .ZN(n457) );
  AOI22_X1 U51 ( .A1(plusA[44]), .A2(n281), .B1(plus2A[44]), .B2(n275), .ZN(
        n395) );
  AOI22_X1 U52 ( .A1(minus2A[44]), .A2(n293), .B1(minusA[44]), .B2(n287), .ZN(
        n394) );
  NAND2_X1 U53 ( .A1(n387), .A2(n386), .ZN(n461) );
  AOI22_X1 U54 ( .A1(plusA[40]), .A2(n281), .B1(plus2A[40]), .B2(n275), .ZN(
        n387) );
  AOI22_X1 U55 ( .A1(minus2A[40]), .A2(n293), .B1(minusA[40]), .B2(n287), .ZN(
        n386) );
  NAND2_X1 U56 ( .A1(n379), .A2(n378), .ZN(n465) );
  AOI22_X1 U57 ( .A1(plusA[36]), .A2(n281), .B1(plus2A[36]), .B2(n275), .ZN(
        n379) );
  AOI22_X1 U58 ( .A1(minus2A[36]), .A2(n293), .B1(minusA[36]), .B2(n287), .ZN(
        n378) );
  NAND2_X1 U59 ( .A1(n421), .A2(n420), .ZN(n444) );
  AOI22_X1 U60 ( .A1(plusA[57]), .A2(n282), .B1(plus2A[57]), .B2(n276), .ZN(
        n421) );
  AOI22_X1 U61 ( .A1(minus2A[57]), .A2(n294), .B1(minusA[57]), .B2(n288), .ZN(
        n420) );
  NAND2_X1 U62 ( .A1(n409), .A2(n408), .ZN(n450) );
  AOI22_X1 U63 ( .A1(plusA[51]), .A2(n282), .B1(plus2A[51]), .B2(n276), .ZN(
        n409) );
  AOI22_X1 U64 ( .A1(minus2A[51]), .A2(n294), .B1(minusA[51]), .B2(n288), .ZN(
        n408) );
  NAND2_X1 U65 ( .A1(n401), .A2(n400), .ZN(n454) );
  AOI22_X1 U66 ( .A1(plusA[47]), .A2(n281), .B1(plus2A[47]), .B2(n275), .ZN(
        n401) );
  AOI22_X1 U67 ( .A1(minus2A[47]), .A2(n293), .B1(minusA[47]), .B2(n287), .ZN(
        n400) );
  NAND2_X1 U68 ( .A1(n393), .A2(n392), .ZN(n458) );
  AOI22_X1 U69 ( .A1(plusA[43]), .A2(n281), .B1(plus2A[43]), .B2(n275), .ZN(
        n393) );
  AOI22_X1 U70 ( .A1(minus2A[43]), .A2(n293), .B1(minusA[43]), .B2(n287), .ZN(
        n392) );
  NAND2_X1 U71 ( .A1(n385), .A2(n384), .ZN(n462) );
  AOI22_X1 U72 ( .A1(plusA[39]), .A2(n281), .B1(plus2A[39]), .B2(n275), .ZN(
        n385) );
  AOI22_X1 U73 ( .A1(minus2A[39]), .A2(n293), .B1(minusA[39]), .B2(n287), .ZN(
        n384) );
  NAND2_X1 U74 ( .A1(n377), .A2(n376), .ZN(n466) );
  AOI22_X1 U75 ( .A1(plusA[35]), .A2(n280), .B1(plus2A[35]), .B2(n274), .ZN(
        n377) );
  AOI22_X1 U76 ( .A1(minus2A[35]), .A2(n292), .B1(minusA[35]), .B2(n286), .ZN(
        n376) );
  NAND2_X1 U77 ( .A1(n419), .A2(n418), .ZN(n445) );
  AOI22_X1 U78 ( .A1(plusA[56]), .A2(n282), .B1(plus2A[56]), .B2(n276), .ZN(
        n419) );
  AOI22_X1 U79 ( .A1(minus2A[56]), .A2(n294), .B1(minusA[56]), .B2(n288), .ZN(
        n418) );
  NAND2_X1 U80 ( .A1(n413), .A2(n412), .ZN(n448) );
  AOI22_X1 U81 ( .A1(plusA[53]), .A2(n282), .B1(plus2A[53]), .B2(n276), .ZN(
        n413) );
  AOI22_X1 U82 ( .A1(minus2A[53]), .A2(n294), .B1(minusA[53]), .B2(n288), .ZN(
        n412) );
  NAND2_X1 U83 ( .A1(n405), .A2(n404), .ZN(n452) );
  AOI22_X1 U84 ( .A1(plusA[49]), .A2(n282), .B1(plus2A[49]), .B2(n276), .ZN(
        n405) );
  AOI22_X1 U85 ( .A1(minus2A[49]), .A2(n294), .B1(minusA[49]), .B2(n288), .ZN(
        n404) );
  NAND2_X1 U86 ( .A1(n397), .A2(n396), .ZN(n456) );
  AOI22_X1 U87 ( .A1(plusA[45]), .A2(n281), .B1(plus2A[45]), .B2(n275), .ZN(
        n397) );
  AOI22_X1 U88 ( .A1(minus2A[45]), .A2(n293), .B1(minusA[45]), .B2(n287), .ZN(
        n396) );
  NAND2_X1 U89 ( .A1(n389), .A2(n388), .ZN(n460) );
  AOI22_X1 U90 ( .A1(plusA[41]), .A2(n281), .B1(plus2A[41]), .B2(n275), .ZN(
        n389) );
  AOI22_X1 U91 ( .A1(minus2A[41]), .A2(n293), .B1(minusA[41]), .B2(n287), .ZN(
        n388) );
  NAND2_X1 U92 ( .A1(n423), .A2(n422), .ZN(n443) );
  AOI22_X1 U93 ( .A1(plusA[58]), .A2(n282), .B1(plus2A[58]), .B2(n276), .ZN(
        n423) );
  AOI22_X1 U94 ( .A1(minus2A[58]), .A2(n294), .B1(minusA[58]), .B2(n288), .ZN(
        n422) );
  NAND2_X1 U95 ( .A1(n437), .A2(n436), .ZN(n438) );
  AOI22_X1 U96 ( .A1(plusA[63]), .A2(n283), .B1(plus2A[63]), .B2(n277), .ZN(
        n437) );
  AOI22_X1 U97 ( .A1(minus2A[63]), .A2(n295), .B1(minusA[63]), .B2(n289), .ZN(
        n436) );
  NAND2_X1 U98 ( .A1(n429), .A2(n428), .ZN(n440) );
  AOI22_X1 U99 ( .A1(plusA[61]), .A2(n283), .B1(plus2A[61]), .B2(n277), .ZN(
        n429) );
  AOI22_X1 U100 ( .A1(minus2A[61]), .A2(n295), .B1(minusA[61]), .B2(n289), 
        .ZN(n428) );
  NAND2_X1 U101 ( .A1(n427), .A2(n426), .ZN(n441) );
  AOI22_X1 U102 ( .A1(plusA[60]), .A2(n283), .B1(plus2A[60]), .B2(n277), .ZN(
        n427) );
  AOI22_X1 U103 ( .A1(minus2A[60]), .A2(n295), .B1(minusA[60]), .B2(n289), 
        .ZN(n426) );
  NAND2_X1 U104 ( .A1(n431), .A2(n430), .ZN(n439) );
  AOI22_X1 U105 ( .A1(plusA[62]), .A2(n283), .B1(plus2A[62]), .B2(n277), .ZN(
        n431) );
  AOI22_X1 U106 ( .A1(minus2A[62]), .A2(n295), .B1(minusA[62]), .B2(n289), 
        .ZN(n430) );
  NAND2_X1 U107 ( .A1(n425), .A2(n424), .ZN(n442) );
  AOI22_X1 U108 ( .A1(plusA[59]), .A2(n282), .B1(plus2A[59]), .B2(n276), .ZN(
        n425) );
  AOI22_X1 U109 ( .A1(minus2A[59]), .A2(n294), .B1(minusA[59]), .B2(n288), 
        .ZN(n424) );
  BUF_X1 U110 ( .A(n493), .Z(n296) );
  BUF_X1 U111 ( .A(n493), .Z(n297) );
  BUF_X1 U112 ( .A(n493), .Z(n298) );
  NAND2_X1 U113 ( .A1(n359), .A2(n358), .ZN(n475) );
  AOI22_X1 U114 ( .A1(plusA[26]), .A2(n280), .B1(plus2A[26]), .B2(n274), .ZN(
        n359) );
  AOI22_X1 U115 ( .A1(minus2A[26]), .A2(n292), .B1(minusA[26]), .B2(n286), 
        .ZN(n358) );
  NAND2_X1 U116 ( .A1(n361), .A2(n360), .ZN(n474) );
  AOI22_X1 U117 ( .A1(plusA[27]), .A2(n280), .B1(plus2A[27]), .B2(n274), .ZN(
        n361) );
  AOI22_X1 U118 ( .A1(minus2A[27]), .A2(n292), .B1(minusA[27]), .B2(n286), 
        .ZN(n360) );
  BUF_X1 U119 ( .A(n433), .Z(n281) );
  BUF_X1 U120 ( .A(n433), .Z(n280) );
  BUF_X1 U121 ( .A(n435), .Z(n293) );
  BUF_X1 U122 ( .A(n435), .Z(n292) );
  BUF_X1 U123 ( .A(n434), .Z(n287) );
  BUF_X1 U124 ( .A(n432), .Z(n275) );
  BUF_X1 U125 ( .A(n434), .Z(n286) );
  BUF_X1 U126 ( .A(n432), .Z(n274) );
  BUF_X1 U127 ( .A(n493), .Z(n299) );
  BUF_X1 U128 ( .A(n493), .Z(n300) );
  BUF_X1 U129 ( .A(n433), .Z(n282) );
  BUF_X1 U130 ( .A(n435), .Z(n294) );
  BUF_X1 U131 ( .A(n434), .Z(n288) );
  BUF_X1 U132 ( .A(n432), .Z(n276) );
  BUF_X1 U133 ( .A(n493), .Z(n301) );
  BUF_X1 U134 ( .A(n433), .Z(n279) );
  BUF_X1 U135 ( .A(n433), .Z(n278) );
  BUF_X1 U136 ( .A(n435), .Z(n291) );
  BUF_X1 U137 ( .A(n435), .Z(n290) );
  BUF_X1 U138 ( .A(n434), .Z(n285) );
  BUF_X1 U139 ( .A(n432), .Z(n273) );
  BUF_X1 U140 ( .A(n434), .Z(n284) );
  BUF_X1 U141 ( .A(n432), .Z(n272) );
  NOR2_X1 U142 ( .A1(n323), .A2(n304), .ZN(n493) );
  INV_X1 U143 ( .A(SEL[2]), .ZN(n304) );
  NOR2_X1 U144 ( .A1(SEL[1]), .A2(SEL[0]), .ZN(n323) );
  NAND2_X1 U145 ( .A1(n357), .A2(n356), .ZN(n476) );
  AOI22_X1 U146 ( .A1(plusA[25]), .A2(n280), .B1(plus2A[25]), .B2(n274), .ZN(
        n357) );
  AOI22_X1 U147 ( .A1(minus2A[25]), .A2(n292), .B1(minusA[25]), .B2(n286), 
        .ZN(n356) );
  NOR3_X1 U148 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n302), .ZN(n434) );
  NOR3_X1 U149 ( .A1(SEL[1]), .A2(SEL[2]), .A3(n303), .ZN(n433) );
  NOR3_X1 U150 ( .A1(n302), .A2(SEL[2]), .A3(n303), .ZN(n432) );
  AND2_X1 U151 ( .A1(SEL[2]), .A2(n323), .ZN(n435) );
  INV_X1 U152 ( .A(SEL[1]), .ZN(n302) );
  INV_X1 U153 ( .A(SEL[0]), .ZN(n303) );
  NAND2_X1 U154 ( .A1(n355), .A2(n354), .ZN(n477) );
  AOI22_X1 U155 ( .A1(plusA[24]), .A2(n280), .B1(plus2A[24]), .B2(n274), .ZN(
        n355) );
  AOI22_X1 U156 ( .A1(minus2A[24]), .A2(n292), .B1(minusA[24]), .B2(n286), 
        .ZN(n354) );
  NAND2_X1 U157 ( .A1(n353), .A2(n352), .ZN(n478) );
  AOI22_X1 U158 ( .A1(plusA[23]), .A2(n279), .B1(plus2A[23]), .B2(n273), .ZN(
        n353) );
  AOI22_X1 U159 ( .A1(minus2A[23]), .A2(n291), .B1(minusA[23]), .B2(n285), 
        .ZN(n352) );
  NAND2_X1 U160 ( .A1(n351), .A2(n350), .ZN(n479) );
  AOI22_X1 U161 ( .A1(plusA[22]), .A2(n279), .B1(plus2A[22]), .B2(n273), .ZN(
        n351) );
  AOI22_X1 U162 ( .A1(minus2A[22]), .A2(n291), .B1(minusA[22]), .B2(n285), 
        .ZN(n350) );
  NAND2_X1 U163 ( .A1(n349), .A2(n348), .ZN(n480) );
  AOI22_X1 U164 ( .A1(plusA[21]), .A2(n279), .B1(plus2A[21]), .B2(n273), .ZN(
        n349) );
  AOI22_X1 U165 ( .A1(minus2A[21]), .A2(n291), .B1(minusA[21]), .B2(n285), 
        .ZN(n348) );
  NAND2_X1 U166 ( .A1(n345), .A2(n344), .ZN(n482) );
  AOI22_X1 U167 ( .A1(plusA[19]), .A2(n279), .B1(plus2A[19]), .B2(n273), .ZN(
        n345) );
  AOI22_X1 U168 ( .A1(minus2A[19]), .A2(n291), .B1(minusA[19]), .B2(n285), 
        .ZN(n344) );
  NAND2_X1 U169 ( .A1(n343), .A2(n342), .ZN(n483) );
  AOI22_X1 U170 ( .A1(plusA[18]), .A2(n279), .B1(plus2A[18]), .B2(n273), .ZN(
        n343) );
  AOI22_X1 U171 ( .A1(minus2A[18]), .A2(n291), .B1(minusA[18]), .B2(n285), 
        .ZN(n342) );
  NAND2_X1 U172 ( .A1(n341), .A2(n340), .ZN(n484) );
  AOI22_X1 U173 ( .A1(plusA[17]), .A2(n279), .B1(plus2A[17]), .B2(n273), .ZN(
        n341) );
  AOI22_X1 U174 ( .A1(minus2A[17]), .A2(n291), .B1(minusA[17]), .B2(n285), 
        .ZN(n340) );
  NAND2_X1 U175 ( .A1(n337), .A2(n336), .ZN(n486) );
  AOI22_X1 U176 ( .A1(plusA[15]), .A2(n279), .B1(plus2A[15]), .B2(n273), .ZN(
        n337) );
  AOI22_X1 U177 ( .A1(minus2A[15]), .A2(n291), .B1(minusA[15]), .B2(n285), 
        .ZN(n336) );
  NAND2_X1 U178 ( .A1(n335), .A2(n334), .ZN(n487) );
  AOI22_X1 U179 ( .A1(plusA[14]), .A2(n279), .B1(plus2A[14]), .B2(n273), .ZN(
        n335) );
  AOI22_X1 U180 ( .A1(minus2A[14]), .A2(n291), .B1(minusA[14]), .B2(n285), 
        .ZN(n334) );
  NAND2_X1 U181 ( .A1(n333), .A2(n332), .ZN(n488) );
  AOI22_X1 U182 ( .A1(plusA[13]), .A2(n279), .B1(plus2A[13]), .B2(n273), .ZN(
        n333) );
  AOI22_X1 U183 ( .A1(minus2A[13]), .A2(n291), .B1(minusA[13]), .B2(n285), 
        .ZN(n332) );
  NAND2_X1 U184 ( .A1(n329), .A2(n328), .ZN(n490) );
  AOI22_X1 U185 ( .A1(plusA[11]), .A2(n278), .B1(plus2A[11]), .B2(n272), .ZN(
        n329) );
  AOI22_X1 U186 ( .A1(minus2A[11]), .A2(n290), .B1(minusA[11]), .B2(n284), 
        .ZN(n328) );
  NAND2_X1 U187 ( .A1(n327), .A2(n326), .ZN(n491) );
  AOI22_X1 U188 ( .A1(plusA[10]), .A2(n278), .B1(plus2A[10]), .B2(n272), .ZN(
        n327) );
  AOI22_X1 U189 ( .A1(minus2A[10]), .A2(n290), .B1(minusA[10]), .B2(n284), 
        .ZN(n326) );
  NAND2_X1 U190 ( .A1(n325), .A2(n324), .ZN(n492) );
  AOI22_X1 U191 ( .A1(plusA[9]), .A2(n278), .B1(plus2A[9]), .B2(n272), .ZN(
        n325) );
  AOI22_X1 U192 ( .A1(minus2A[9]), .A2(n290), .B1(minusA[9]), .B2(n284), .ZN(
        n324) );
  NAND2_X1 U193 ( .A1(n320), .A2(n319), .ZN(n495) );
  AOI22_X1 U194 ( .A1(plusA[7]), .A2(n278), .B1(plus2A[7]), .B2(n272), .ZN(
        n320) );
  AOI22_X1 U195 ( .A1(minus2A[7]), .A2(n290), .B1(minusA[7]), .B2(n284), .ZN(
        n319) );
  NAND2_X1 U196 ( .A1(n318), .A2(n317), .ZN(n496) );
  AOI22_X1 U197 ( .A1(plusA[6]), .A2(n278), .B1(plus2A[6]), .B2(n272), .ZN(
        n318) );
  AOI22_X1 U198 ( .A1(minus2A[6]), .A2(n290), .B1(minusA[6]), .B2(n284), .ZN(
        n317) );
  NAND2_X1 U199 ( .A1(n316), .A2(n315), .ZN(n497) );
  AOI22_X1 U200 ( .A1(plusA[5]), .A2(n278), .B1(plus2A[5]), .B2(n272), .ZN(
        n316) );
  AOI22_X1 U201 ( .A1(minus2A[5]), .A2(n290), .B1(minusA[5]), .B2(n284), .ZN(
        n315) );
  NAND2_X1 U202 ( .A1(n312), .A2(n311), .ZN(n499) );
  AOI22_X1 U203 ( .A1(plusA[3]), .A2(n278), .B1(plus2A[3]), .B2(n272), .ZN(
        n312) );
  AOI22_X1 U204 ( .A1(minus2A[3]), .A2(n290), .B1(minusA[3]), .B2(n284), .ZN(
        n311) );
  NAND2_X1 U205 ( .A1(n347), .A2(n346), .ZN(n481) );
  AOI22_X1 U206 ( .A1(plusA[20]), .A2(n279), .B1(plus2A[20]), .B2(n273), .ZN(
        n347) );
  AOI22_X1 U207 ( .A1(minus2A[20]), .A2(n291), .B1(minusA[20]), .B2(n285), 
        .ZN(n346) );
  NAND2_X1 U208 ( .A1(n339), .A2(n338), .ZN(n485) );
  AOI22_X1 U209 ( .A1(plusA[16]), .A2(n279), .B1(plus2A[16]), .B2(n273), .ZN(
        n339) );
  AOI22_X1 U210 ( .A1(minus2A[16]), .A2(n291), .B1(minusA[16]), .B2(n285), 
        .ZN(n338) );
  NAND2_X1 U211 ( .A1(n331), .A2(n330), .ZN(n489) );
  AOI22_X1 U212 ( .A1(plusA[12]), .A2(n279), .B1(plus2A[12]), .B2(n273), .ZN(
        n331) );
  AOI22_X1 U213 ( .A1(minus2A[12]), .A2(n291), .B1(minusA[12]), .B2(n285), 
        .ZN(n330) );
  NAND2_X1 U214 ( .A1(n322), .A2(n321), .ZN(n494) );
  AOI22_X1 U215 ( .A1(plusA[8]), .A2(n278), .B1(plus2A[8]), .B2(n272), .ZN(
        n322) );
  AOI22_X1 U216 ( .A1(minus2A[8]), .A2(n290), .B1(minusA[8]), .B2(n284), .ZN(
        n321) );
  NAND2_X1 U217 ( .A1(n314), .A2(n313), .ZN(n498) );
  AOI22_X1 U218 ( .A1(plusA[4]), .A2(n278), .B1(plus2A[4]), .B2(n272), .ZN(
        n314) );
  AOI22_X1 U219 ( .A1(minus2A[4]), .A2(n290), .B1(minusA[4]), .B2(n284), .ZN(
        n313) );
  NAND2_X1 U220 ( .A1(n310), .A2(n309), .ZN(n500) );
  AOI22_X1 U221 ( .A1(plusA[2]), .A2(n278), .B1(plus2A[2]), .B2(n272), .ZN(
        n310) );
  AOI22_X1 U222 ( .A1(minus2A[2]), .A2(n290), .B1(minusA[2]), .B2(n284), .ZN(
        n309) );
  NAND2_X1 U223 ( .A1(n308), .A2(n307), .ZN(n501) );
  AOI22_X1 U224 ( .A1(plusA[1]), .A2(n278), .B1(plus2A[1]), .B2(n272), .ZN(
        n308) );
  AOI22_X1 U225 ( .A1(minus2A[1]), .A2(n290), .B1(minusA[1]), .B2(n284), .ZN(
        n307) );
  NAND2_X1 U226 ( .A1(n306), .A2(n305), .ZN(n502) );
  AOI22_X1 U227 ( .A1(plusA[0]), .A2(n278), .B1(plus2A[0]), .B2(n272), .ZN(
        n306) );
  AOI22_X1 U228 ( .A1(minus2A[0]), .A2(n290), .B1(minusA[0]), .B2(n284), .ZN(
        n305) );
  CLKBUF_X1 U229 ( .A(n432), .Z(n277) );
  CLKBUF_X1 U230 ( .A(n433), .Z(n283) );
  CLKBUF_X1 U231 ( .A(n434), .Z(n289) );
  CLKBUF_X1 U232 ( .A(n435), .Z(n295) );
endmodule


module FA_256 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_255 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_254 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_253 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_252 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_251 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_250 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_249 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_248 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_247 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_246 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_245 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_244 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_243 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_242 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_241 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_240 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_239 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_238 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_237 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_236 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_235 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_234 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_233 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_232 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_231 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_230 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_229 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_228 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_227 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_226 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_225 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_224 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_223 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_222 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_221 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_220 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_219 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_218 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_217 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_216 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_215 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_214 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_213 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_212 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_211 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_210 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_209 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_208 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_207 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_206 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_205 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_204 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_203 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_202 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_201 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_200 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_199 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_198 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_197 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_196 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_195 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_194 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_193 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N64_4 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Ci;
  output Co;

  wire   [63:1] CTMP;
  tri   [63:0] A;

  FA_256 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_255 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_254 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_253 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(CTMP[4]) );
  FA_252 FAI_5 ( .A(A[4]), .B(B[4]), .Ci(CTMP[4]), .S(S[4]), .Co(CTMP[5]) );
  FA_251 FAI_6 ( .A(A[5]), .B(B[5]), .Ci(CTMP[5]), .S(S[5]), .Co(CTMP[6]) );
  FA_250 FAI_7 ( .A(A[6]), .B(B[6]), .Ci(CTMP[6]), .S(S[6]), .Co(CTMP[7]) );
  FA_249 FAI_8 ( .A(A[7]), .B(B[7]), .Ci(CTMP[7]), .S(S[7]), .Co(CTMP[8]) );
  FA_248 FAI_9 ( .A(A[8]), .B(B[8]), .Ci(CTMP[8]), .S(S[8]), .Co(CTMP[9]) );
  FA_247 FAI_10 ( .A(A[9]), .B(B[9]), .Ci(CTMP[9]), .S(S[9]), .Co(CTMP[10]) );
  FA_246 FAI_11 ( .A(A[10]), .B(B[10]), .Ci(CTMP[10]), .S(S[10]), .Co(CTMP[11]) );
  FA_245 FAI_12 ( .A(A[11]), .B(B[11]), .Ci(CTMP[11]), .S(S[11]), .Co(CTMP[12]) );
  FA_244 FAI_13 ( .A(A[12]), .B(B[12]), .Ci(CTMP[12]), .S(S[12]), .Co(CTMP[13]) );
  FA_243 FAI_14 ( .A(A[13]), .B(B[13]), .Ci(CTMP[13]), .S(S[13]), .Co(CTMP[14]) );
  FA_242 FAI_15 ( .A(A[14]), .B(B[14]), .Ci(CTMP[14]), .S(S[14]), .Co(CTMP[15]) );
  FA_241 FAI_16 ( .A(A[15]), .B(B[15]), .Ci(CTMP[15]), .S(S[15]), .Co(CTMP[16]) );
  FA_240 FAI_17 ( .A(A[16]), .B(B[16]), .Ci(CTMP[16]), .S(S[16]), .Co(CTMP[17]) );
  FA_239 FAI_18 ( .A(A[17]), .B(B[17]), .Ci(CTMP[17]), .S(S[17]), .Co(CTMP[18]) );
  FA_238 FAI_19 ( .A(A[18]), .B(B[18]), .Ci(CTMP[18]), .S(S[18]), .Co(CTMP[19]) );
  FA_237 FAI_20 ( .A(A[19]), .B(B[19]), .Ci(CTMP[19]), .S(S[19]), .Co(CTMP[20]) );
  FA_236 FAI_21 ( .A(A[20]), .B(B[20]), .Ci(CTMP[20]), .S(S[20]), .Co(CTMP[21]) );
  FA_235 FAI_22 ( .A(A[21]), .B(B[21]), .Ci(CTMP[21]), .S(S[21]), .Co(CTMP[22]) );
  FA_234 FAI_23 ( .A(A[22]), .B(B[22]), .Ci(CTMP[22]), .S(S[22]), .Co(CTMP[23]) );
  FA_233 FAI_24 ( .A(A[23]), .B(B[23]), .Ci(CTMP[23]), .S(S[23]), .Co(CTMP[24]) );
  FA_232 FAI_25 ( .A(A[24]), .B(B[24]), .Ci(CTMP[24]), .S(S[24]), .Co(CTMP[25]) );
  FA_231 FAI_26 ( .A(A[25]), .B(B[25]), .Ci(CTMP[25]), .S(S[25]), .Co(CTMP[26]) );
  FA_230 FAI_27 ( .A(A[26]), .B(B[26]), .Ci(CTMP[26]), .S(S[26]), .Co(CTMP[27]) );
  FA_229 FAI_28 ( .A(A[27]), .B(B[27]), .Ci(CTMP[27]), .S(S[27]), .Co(CTMP[28]) );
  FA_228 FAI_29 ( .A(A[28]), .B(B[28]), .Ci(CTMP[28]), .S(S[28]), .Co(CTMP[29]) );
  FA_227 FAI_30 ( .A(A[29]), .B(B[29]), .Ci(CTMP[29]), .S(S[29]), .Co(CTMP[30]) );
  FA_226 FAI_31 ( .A(A[30]), .B(B[30]), .Ci(CTMP[30]), .S(S[30]), .Co(CTMP[31]) );
  FA_225 FAI_32 ( .A(A[31]), .B(B[31]), .Ci(CTMP[31]), .S(S[31]), .Co(CTMP[32]) );
  FA_224 FAI_33 ( .A(A[32]), .B(B[32]), .Ci(CTMP[32]), .S(S[32]), .Co(CTMP[33]) );
  FA_223 FAI_34 ( .A(A[33]), .B(B[33]), .Ci(CTMP[33]), .S(S[33]), .Co(CTMP[34]) );
  FA_222 FAI_35 ( .A(A[34]), .B(B[34]), .Ci(CTMP[34]), .S(S[34]), .Co(CTMP[35]) );
  FA_221 FAI_36 ( .A(A[35]), .B(B[35]), .Ci(CTMP[35]), .S(S[35]), .Co(CTMP[36]) );
  FA_220 FAI_37 ( .A(A[36]), .B(B[36]), .Ci(CTMP[36]), .S(S[36]), .Co(CTMP[37]) );
  FA_219 FAI_38 ( .A(A[37]), .B(B[37]), .Ci(CTMP[37]), .S(S[37]), .Co(CTMP[38]) );
  FA_218 FAI_39 ( .A(A[38]), .B(B[38]), .Ci(CTMP[38]), .S(S[38]), .Co(CTMP[39]) );
  FA_217 FAI_40 ( .A(A[39]), .B(B[39]), .Ci(CTMP[39]), .S(S[39]), .Co(CTMP[40]) );
  FA_216 FAI_41 ( .A(A[40]), .B(B[40]), .Ci(CTMP[40]), .S(S[40]), .Co(CTMP[41]) );
  FA_215 FAI_42 ( .A(A[41]), .B(B[41]), .Ci(CTMP[41]), .S(S[41]), .Co(CTMP[42]) );
  FA_214 FAI_43 ( .A(A[42]), .B(B[42]), .Ci(CTMP[42]), .S(S[42]), .Co(CTMP[43]) );
  FA_213 FAI_44 ( .A(A[43]), .B(B[43]), .Ci(CTMP[43]), .S(S[43]), .Co(CTMP[44]) );
  FA_212 FAI_45 ( .A(A[44]), .B(B[44]), .Ci(CTMP[44]), .S(S[44]), .Co(CTMP[45]) );
  FA_211 FAI_46 ( .A(A[45]), .B(B[45]), .Ci(CTMP[45]), .S(S[45]), .Co(CTMP[46]) );
  FA_210 FAI_47 ( .A(A[46]), .B(B[46]), .Ci(CTMP[46]), .S(S[46]), .Co(CTMP[47]) );
  FA_209 FAI_48 ( .A(A[47]), .B(B[47]), .Ci(CTMP[47]), .S(S[47]), .Co(CTMP[48]) );
  FA_208 FAI_49 ( .A(A[48]), .B(B[48]), .Ci(CTMP[48]), .S(S[48]), .Co(CTMP[49]) );
  FA_207 FAI_50 ( .A(A[49]), .B(B[49]), .Ci(CTMP[49]), .S(S[49]), .Co(CTMP[50]) );
  FA_206 FAI_51 ( .A(A[50]), .B(B[50]), .Ci(CTMP[50]), .S(S[50]), .Co(CTMP[51]) );
  FA_205 FAI_52 ( .A(A[51]), .B(B[51]), .Ci(CTMP[51]), .S(S[51]), .Co(CTMP[52]) );
  FA_204 FAI_53 ( .A(A[52]), .B(B[52]), .Ci(CTMP[52]), .S(S[52]), .Co(CTMP[53]) );
  FA_203 FAI_54 ( .A(A[53]), .B(B[53]), .Ci(CTMP[53]), .S(S[53]), .Co(CTMP[54]) );
  FA_202 FAI_55 ( .A(A[54]), .B(B[54]), .Ci(CTMP[54]), .S(S[54]), .Co(CTMP[55]) );
  FA_201 FAI_56 ( .A(A[55]), .B(B[55]), .Ci(CTMP[55]), .S(S[55]), .Co(CTMP[56]) );
  FA_200 FAI_57 ( .A(A[56]), .B(B[56]), .Ci(CTMP[56]), .S(S[56]), .Co(CTMP[57]) );
  FA_199 FAI_58 ( .A(A[57]), .B(B[57]), .Ci(CTMP[57]), .S(S[57]), .Co(CTMP[58]) );
  FA_198 FAI_59 ( .A(A[58]), .B(B[58]), .Ci(CTMP[58]), .S(S[58]), .Co(CTMP[59]) );
  FA_197 FAI_60 ( .A(A[59]), .B(B[59]), .Ci(CTMP[59]), .S(S[59]), .Co(CTMP[60]) );
  FA_196 FAI_61 ( .A(A[60]), .B(B[60]), .Ci(CTMP[60]), .S(S[60]), .Co(CTMP[61]) );
  FA_195 FAI_62 ( .A(A[61]), .B(B[61]), .Ci(CTMP[61]), .S(S[61]), .Co(CTMP[62]) );
  FA_194 FAI_63 ( .A(A[62]), .B(B[62]), .Ci(CTMP[62]), .S(S[62]), .Co(CTMP[63]) );
  FA_193 FAI_64 ( .A(A[63]), .B(B[63]), .Ci(CTMP[63]), .S(S[63]), .Co(Co) );
endmodule


module booth_mul_row_N64_RADIX3_4 ( prevA, prevSum, encoderIn, nextA, nextSum
 );
  input [63:0] prevA;
  input [63:0] prevSum;
  input [2:0] encoderIn;
  output [63:0] nextA;
  output [63:0] nextSum;

  wire   [2:0] encoder_to_mux;
  wire   [63:0] plus2A_s;
  wire   [63:0] minus2A_s;
  wire   [63:0] minus4A_s;
  tri   [63:0] mux_to_adder;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign nextA[0] = 1'b0;

  encoder_N64_RADIX3_4 encoder_1 ( .X(encoderIn), .Z(encoder_to_mux) );
  ShiftnCompl_N64_4 ShiftnCompl_1 ( .plusA(prevA), .plus2A_out({plus2A_s[63:1], 
        SYNOPSYS_UNCONNECTED__0}), .minus2A_out(minus2A_s), .plus4A_out({
        nextA[63:1], SYNOPSYS_UNCONNECTED__1}), .minus4A_out(minus4A_s) );
  MUX_GENERIC_N64_RADIX3_4 mux_1 ( .plusA({plus2A_s[63:1], 1'b0}), .minusA(
        minus2A_s), .plus2A({nextA[63:1], 1'b0}), .minus2A(minus4A_s), .SEL(
        encoder_to_mux), .Y(mux_to_adder) );
  RCA_N64_4 rca_1 ( .A(mux_to_adder), .B(prevSum), .Ci(1'b0), .S(nextSum) );
endmodule


module encoder_N64_RADIX3_3 ( X, Z );
  input [2:0] X;
  output [2:0] Z;
  wire   n5, n7, n8;

  OAI22_X1 U1 ( .A1(n8), .A2(n5), .B1(X[2]), .B2(n7), .ZN(Z[1]) );
  INV_X1 U2 ( .A(X[2]), .ZN(n5) );
  AOI21_X1 U3 ( .B1(n8), .B2(n7), .A(X[2]), .ZN(Z[0]) );
  OAI21_X1 U4 ( .B1(X[1]), .B2(X[0]), .A(n7), .ZN(n8) );
  AND3_X1 U5 ( .A1(X[2]), .A2(n7), .A3(n8), .ZN(Z[2]) );
  NAND2_X1 U6 ( .A1(X[1]), .A2(X[0]), .ZN(n7) );
endmodule


module shifter_N64_6 ( \input , shiftLeftOnePos );
  input [63:0] \input ;
  output [63:0] shiftLeftOnePos;
  wire   \input[62] , \input[61] , \input[60] , \input[59] , \input[58] ,
         \input[57] , \input[56] , \input[55] , \input[54] , \input[53] ,
         \input[52] , \input[51] , \input[50] , \input[49] , \input[48] ,
         \input[47] , \input[46] , \input[45] , \input[44] , \input[43] ,
         \input[42] , \input[41] , \input[40] , \input[39] , \input[38] ,
         \input[37] , \input[36] , \input[35] , \input[34] , \input[33] ,
         \input[32] , \input[31] , \input[30] , \input[29] , \input[28] ,
         \input[27] , \input[26] , \input[25] , \input[24] , \input[23] ,
         \input[22] , \input[21] , \input[20] , \input[19] , \input[18] ,
         \input[17] , \input[16] , \input[15] , \input[14] , \input[13] ,
         \input[12] , \input[11] , \input[10] , \input[9] , \input[8] ,
         \input[7] , \input[6] , \input[5] , \input[4] , \input[3] ,
         \input[2] , \input[1] , \input[0] ;
  assign shiftLeftOnePos[0] = 1'b0;
  assign shiftLeftOnePos[63] = \input[62] ;
  assign \input[62]  = \input  [62];
  assign shiftLeftOnePos[62] = \input[61] ;
  assign \input[61]  = \input  [61];
  assign shiftLeftOnePos[61] = \input[60] ;
  assign \input[60]  = \input  [60];
  assign shiftLeftOnePos[60] = \input[59] ;
  assign \input[59]  = \input  [59];
  assign shiftLeftOnePos[59] = \input[58] ;
  assign \input[58]  = \input  [58];
  assign shiftLeftOnePos[58] = \input[57] ;
  assign \input[57]  = \input  [57];
  assign shiftLeftOnePos[57] = \input[56] ;
  assign \input[56]  = \input  [56];
  assign shiftLeftOnePos[56] = \input[55] ;
  assign \input[55]  = \input  [55];
  assign shiftLeftOnePos[55] = \input[54] ;
  assign \input[54]  = \input  [54];
  assign shiftLeftOnePos[54] = \input[53] ;
  assign \input[53]  = \input  [53];
  assign shiftLeftOnePos[53] = \input[52] ;
  assign \input[52]  = \input  [52];
  assign shiftLeftOnePos[52] = \input[51] ;
  assign \input[51]  = \input  [51];
  assign shiftLeftOnePos[51] = \input[50] ;
  assign \input[50]  = \input  [50];
  assign shiftLeftOnePos[50] = \input[49] ;
  assign \input[49]  = \input  [49];
  assign shiftLeftOnePos[49] = \input[48] ;
  assign \input[48]  = \input  [48];
  assign shiftLeftOnePos[48] = \input[47] ;
  assign \input[47]  = \input  [47];
  assign shiftLeftOnePos[47] = \input[46] ;
  assign \input[46]  = \input  [46];
  assign shiftLeftOnePos[46] = \input[45] ;
  assign \input[45]  = \input  [45];
  assign shiftLeftOnePos[45] = \input[44] ;
  assign \input[44]  = \input  [44];
  assign shiftLeftOnePos[44] = \input[43] ;
  assign \input[43]  = \input  [43];
  assign shiftLeftOnePos[43] = \input[42] ;
  assign \input[42]  = \input  [42];
  assign shiftLeftOnePos[42] = \input[41] ;
  assign \input[41]  = \input  [41];
  assign shiftLeftOnePos[41] = \input[40] ;
  assign \input[40]  = \input  [40];
  assign shiftLeftOnePos[40] = \input[39] ;
  assign \input[39]  = \input  [39];
  assign shiftLeftOnePos[39] = \input[38] ;
  assign \input[38]  = \input  [38];
  assign shiftLeftOnePos[38] = \input[37] ;
  assign \input[37]  = \input  [37];
  assign shiftLeftOnePos[37] = \input[36] ;
  assign \input[36]  = \input  [36];
  assign shiftLeftOnePos[36] = \input[35] ;
  assign \input[35]  = \input  [35];
  assign shiftLeftOnePos[35] = \input[34] ;
  assign \input[34]  = \input  [34];
  assign shiftLeftOnePos[34] = \input[33] ;
  assign \input[33]  = \input  [33];
  assign shiftLeftOnePos[33] = \input[32] ;
  assign \input[32]  = \input  [32];
  assign shiftLeftOnePos[32] = \input[31] ;
  assign \input[31]  = \input  [31];
  assign shiftLeftOnePos[31] = \input[30] ;
  assign \input[30]  = \input  [30];
  assign shiftLeftOnePos[30] = \input[29] ;
  assign \input[29]  = \input  [29];
  assign shiftLeftOnePos[29] = \input[28] ;
  assign \input[28]  = \input  [28];
  assign shiftLeftOnePos[28] = \input[27] ;
  assign \input[27]  = \input  [27];
  assign shiftLeftOnePos[27] = \input[26] ;
  assign \input[26]  = \input  [26];
  assign shiftLeftOnePos[26] = \input[25] ;
  assign \input[25]  = \input  [25];
  assign shiftLeftOnePos[25] = \input[24] ;
  assign \input[24]  = \input  [24];
  assign shiftLeftOnePos[24] = \input[23] ;
  assign \input[23]  = \input  [23];
  assign shiftLeftOnePos[23] = \input[22] ;
  assign \input[22]  = \input  [22];
  assign shiftLeftOnePos[22] = \input[21] ;
  assign \input[21]  = \input  [21];
  assign shiftLeftOnePos[21] = \input[20] ;
  assign \input[20]  = \input  [20];
  assign shiftLeftOnePos[20] = \input[19] ;
  assign \input[19]  = \input  [19];
  assign shiftLeftOnePos[19] = \input[18] ;
  assign \input[18]  = \input  [18];
  assign shiftLeftOnePos[18] = \input[17] ;
  assign \input[17]  = \input  [17];
  assign shiftLeftOnePos[17] = \input[16] ;
  assign \input[16]  = \input  [16];
  assign shiftLeftOnePos[16] = \input[15] ;
  assign \input[15]  = \input  [15];
  assign shiftLeftOnePos[15] = \input[14] ;
  assign \input[14]  = \input  [14];
  assign shiftLeftOnePos[14] = \input[13] ;
  assign \input[13]  = \input  [13];
  assign shiftLeftOnePos[13] = \input[12] ;
  assign \input[12]  = \input  [12];
  assign shiftLeftOnePos[12] = \input[11] ;
  assign \input[11]  = \input  [11];
  assign shiftLeftOnePos[11] = \input[10] ;
  assign \input[10]  = \input  [10];
  assign shiftLeftOnePos[10] = \input[9] ;
  assign \input[9]  = \input  [9];
  assign shiftLeftOnePos[9] = \input[8] ;
  assign \input[8]  = \input  [8];
  assign shiftLeftOnePos[8] = \input[7] ;
  assign \input[7]  = \input  [7];
  assign shiftLeftOnePos[7] = \input[6] ;
  assign \input[6]  = \input  [6];
  assign shiftLeftOnePos[6] = \input[5] ;
  assign \input[5]  = \input  [5];
  assign shiftLeftOnePos[5] = \input[4] ;
  assign \input[4]  = \input  [4];
  assign shiftLeftOnePos[4] = \input[3] ;
  assign \input[3]  = \input  [3];
  assign shiftLeftOnePos[3] = \input[2] ;
  assign \input[2]  = \input  [2];
  assign shiftLeftOnePos[2] = \input[1] ;
  assign \input[1]  = \input  [1];
  assign shiftLeftOnePos[1] = \input[0] ;
  assign \input[0]  = \input  [0];

endmodule


module shifter_N64_5 ( \input , shiftLeftOnePos );
  input [63:0] \input ;
  output [63:0] shiftLeftOnePos;
  wire   \input[62] , \input[61] , \input[60] , \input[59] , \input[58] ,
         \input[57] , \input[56] , \input[55] , \input[54] , \input[53] ,
         \input[52] , \input[51] , \input[50] , \input[49] , \input[48] ,
         \input[47] , \input[46] , \input[45] , \input[44] , \input[43] ,
         \input[42] , \input[41] , \input[40] , \input[39] , \input[38] ,
         \input[37] , \input[36] , \input[35] , \input[34] , \input[33] ,
         \input[32] , \input[31] , \input[30] , \input[29] , \input[28] ,
         \input[27] , \input[26] , \input[25] , \input[24] , \input[23] ,
         \input[22] , \input[21] , \input[20] , \input[19] , \input[18] ,
         \input[17] , \input[16] , \input[15] , \input[14] , \input[13] ,
         \input[12] , \input[11] , \input[10] , \input[9] , \input[8] ,
         \input[7] , \input[6] , \input[5] , \input[4] , \input[3] ,
         \input[2] , \input[1] , \input[0] ;
  assign shiftLeftOnePos[0] = 1'b0;
  assign shiftLeftOnePos[63] = \input[62] ;
  assign \input[62]  = \input  [62];
  assign shiftLeftOnePos[62] = \input[61] ;
  assign \input[61]  = \input  [61];
  assign shiftLeftOnePos[61] = \input[60] ;
  assign \input[60]  = \input  [60];
  assign shiftLeftOnePos[60] = \input[59] ;
  assign \input[59]  = \input  [59];
  assign shiftLeftOnePos[59] = \input[58] ;
  assign \input[58]  = \input  [58];
  assign shiftLeftOnePos[58] = \input[57] ;
  assign \input[57]  = \input  [57];
  assign shiftLeftOnePos[57] = \input[56] ;
  assign \input[56]  = \input  [56];
  assign shiftLeftOnePos[56] = \input[55] ;
  assign \input[55]  = \input  [55];
  assign shiftLeftOnePos[55] = \input[54] ;
  assign \input[54]  = \input  [54];
  assign shiftLeftOnePos[54] = \input[53] ;
  assign \input[53]  = \input  [53];
  assign shiftLeftOnePos[53] = \input[52] ;
  assign \input[52]  = \input  [52];
  assign shiftLeftOnePos[52] = \input[51] ;
  assign \input[51]  = \input  [51];
  assign shiftLeftOnePos[51] = \input[50] ;
  assign \input[50]  = \input  [50];
  assign shiftLeftOnePos[50] = \input[49] ;
  assign \input[49]  = \input  [49];
  assign shiftLeftOnePos[49] = \input[48] ;
  assign \input[48]  = \input  [48];
  assign shiftLeftOnePos[48] = \input[47] ;
  assign \input[47]  = \input  [47];
  assign shiftLeftOnePos[47] = \input[46] ;
  assign \input[46]  = \input  [46];
  assign shiftLeftOnePos[46] = \input[45] ;
  assign \input[45]  = \input  [45];
  assign shiftLeftOnePos[45] = \input[44] ;
  assign \input[44]  = \input  [44];
  assign shiftLeftOnePos[44] = \input[43] ;
  assign \input[43]  = \input  [43];
  assign shiftLeftOnePos[43] = \input[42] ;
  assign \input[42]  = \input  [42];
  assign shiftLeftOnePos[42] = \input[41] ;
  assign \input[41]  = \input  [41];
  assign shiftLeftOnePos[41] = \input[40] ;
  assign \input[40]  = \input  [40];
  assign shiftLeftOnePos[40] = \input[39] ;
  assign \input[39]  = \input  [39];
  assign shiftLeftOnePos[39] = \input[38] ;
  assign \input[38]  = \input  [38];
  assign shiftLeftOnePos[38] = \input[37] ;
  assign \input[37]  = \input  [37];
  assign shiftLeftOnePos[37] = \input[36] ;
  assign \input[36]  = \input  [36];
  assign shiftLeftOnePos[36] = \input[35] ;
  assign \input[35]  = \input  [35];
  assign shiftLeftOnePos[35] = \input[34] ;
  assign \input[34]  = \input  [34];
  assign shiftLeftOnePos[34] = \input[33] ;
  assign \input[33]  = \input  [33];
  assign shiftLeftOnePos[33] = \input[32] ;
  assign \input[32]  = \input  [32];
  assign shiftLeftOnePos[32] = \input[31] ;
  assign \input[31]  = \input  [31];
  assign shiftLeftOnePos[31] = \input[30] ;
  assign \input[30]  = \input  [30];
  assign shiftLeftOnePos[30] = \input[29] ;
  assign \input[29]  = \input  [29];
  assign shiftLeftOnePos[29] = \input[28] ;
  assign \input[28]  = \input  [28];
  assign shiftLeftOnePos[28] = \input[27] ;
  assign \input[27]  = \input  [27];
  assign shiftLeftOnePos[27] = \input[26] ;
  assign \input[26]  = \input  [26];
  assign shiftLeftOnePos[26] = \input[25] ;
  assign \input[25]  = \input  [25];
  assign shiftLeftOnePos[25] = \input[24] ;
  assign \input[24]  = \input  [24];
  assign shiftLeftOnePos[24] = \input[23] ;
  assign \input[23]  = \input  [23];
  assign shiftLeftOnePos[23] = \input[22] ;
  assign \input[22]  = \input  [22];
  assign shiftLeftOnePos[22] = \input[21] ;
  assign \input[21]  = \input  [21];
  assign shiftLeftOnePos[21] = \input[20] ;
  assign \input[20]  = \input  [20];
  assign shiftLeftOnePos[20] = \input[19] ;
  assign \input[19]  = \input  [19];
  assign shiftLeftOnePos[19] = \input[18] ;
  assign \input[18]  = \input  [18];
  assign shiftLeftOnePos[18] = \input[17] ;
  assign \input[17]  = \input  [17];
  assign shiftLeftOnePos[17] = \input[16] ;
  assign \input[16]  = \input  [16];
  assign shiftLeftOnePos[16] = \input[15] ;
  assign \input[15]  = \input  [15];
  assign shiftLeftOnePos[15] = \input[14] ;
  assign \input[14]  = \input  [14];
  assign shiftLeftOnePos[14] = \input[13] ;
  assign \input[13]  = \input  [13];
  assign shiftLeftOnePos[13] = \input[12] ;
  assign \input[12]  = \input  [12];
  assign shiftLeftOnePos[12] = \input[11] ;
  assign \input[11]  = \input  [11];
  assign shiftLeftOnePos[11] = \input[10] ;
  assign \input[10]  = \input  [10];
  assign shiftLeftOnePos[10] = \input[9] ;
  assign \input[9]  = \input  [9];
  assign shiftLeftOnePos[9] = \input[8] ;
  assign \input[8]  = \input  [8];
  assign shiftLeftOnePos[8] = \input[7] ;
  assign \input[7]  = \input  [7];
  assign shiftLeftOnePos[7] = \input[6] ;
  assign \input[6]  = \input  [6];
  assign shiftLeftOnePos[6] = \input[5] ;
  assign \input[5]  = \input  [5];
  assign shiftLeftOnePos[5] = \input[4] ;
  assign \input[4]  = \input  [4];
  assign shiftLeftOnePos[4] = \input[3] ;
  assign \input[3]  = \input  [3];
  assign shiftLeftOnePos[3] = \input[2] ;
  assign \input[2]  = \input  [2];
  assign shiftLeftOnePos[2] = \input[1] ;
  assign \input[1]  = \input  [1];
  assign shiftLeftOnePos[1] = \input[0] ;
  assign \input[0]  = \input  [0];

endmodule


module complementer_N64_6_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n189, n236;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U81 ( .A(n190), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U82 ( .A(n192), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U83 ( .A(n193), .B(B[6]), .Z(DIFF[6]) );
  XOR2_X1 U84 ( .A(n195), .B(B[63]), .Z(DIFF[63]) );
  XOR2_X1 U85 ( .A(n196), .B(B[62]), .Z(DIFF[62]) );
  XOR2_X1 U86 ( .A(n194), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U87 ( .A(n198), .B(B[59]), .Z(DIFF[59]) );
  XOR2_X1 U88 ( .A(n201), .B(B[58]), .Z(DIFF[58]) );
  XOR2_X1 U89 ( .A(n200), .B(B[57]), .Z(DIFF[57]) );
  XOR2_X1 U90 ( .A(n202), .B(B[55]), .Z(DIFF[55]) );
  XOR2_X1 U91 ( .A(n205), .B(B[54]), .Z(DIFF[54]) );
  XOR2_X1 U92 ( .A(n204), .B(B[53]), .Z(DIFF[53]) );
  XOR2_X1 U93 ( .A(n206), .B(B[51]), .Z(DIFF[51]) );
  XOR2_X1 U94 ( .A(n209), .B(B[50]), .Z(DIFF[50]) );
  XOR2_X1 U95 ( .A(n208), .B(B[49]), .Z(DIFF[49]) );
  XOR2_X1 U96 ( .A(n212), .B(B[47]), .Z(DIFF[47]) );
  XOR2_X1 U97 ( .A(n215), .B(B[46]), .Z(DIFF[46]) );
  XOR2_X1 U98 ( .A(n214), .B(B[45]), .Z(DIFF[45]) );
  XOR2_X1 U99 ( .A(n216), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U100 ( .A(n219), .B(B[42]), .Z(DIFF[42]) );
  XOR2_X1 U101 ( .A(n218), .B(B[41]), .Z(DIFF[41]) );
  XOR2_X1 U102 ( .A(n211), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U103 ( .A(n220), .B(B[39]), .Z(DIFF[39]) );
  XOR2_X1 U104 ( .A(n223), .B(B[38]), .Z(DIFF[38]) );
  XOR2_X1 U105 ( .A(n222), .B(B[37]), .Z(DIFF[37]) );
  XOR2_X1 U106 ( .A(n224), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U107 ( .A(n227), .B(B[34]), .Z(DIFF[34]) );
  XOR2_X1 U108 ( .A(n226), .B(B[33]), .Z(DIFF[33]) );
  XOR2_X1 U109 ( .A(n228), .B(B[31]), .Z(DIFF[31]) );
  XOR2_X1 U110 ( .A(n231), .B(B[30]), .Z(DIFF[30]) );
  XOR2_X1 U111 ( .A(n230), .B(B[29]), .Z(DIFF[29]) );
  XOR2_X1 U112 ( .A(n233), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U114 ( .A(n235), .B(B[25]), .Z(DIFF[25]) );
  XOR2_X1 U115 ( .A(n237), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U116 ( .A(n240), .B(B[22]), .Z(DIFF[22]) );
  XOR2_X1 U117 ( .A(n239), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U118 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U119 ( .A(n241), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U120 ( .A(n244), .B(B[18]), .Z(DIFF[18]) );
  XOR2_X1 U121 ( .A(n243), .B(B[17]), .Z(DIFF[17]) );
  XOR2_X1 U122 ( .A(n245), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U123 ( .A(n248), .B(B[14]), .Z(DIFF[14]) );
  XOR2_X1 U124 ( .A(n247), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U125 ( .A(n249), .B(B[11]), .Z(DIFF[11]) );
  XOR2_X1 U126 ( .A(n251), .B(B[10]), .Z(DIFF[10]) );
  NAND2_X1 U1 ( .A1(n197), .A2(n236), .ZN(n196) );
  NOR3_X1 U2 ( .A1(B[59]), .A2(B[60]), .A3(n198), .ZN(n197) );
  NOR2_X1 U3 ( .A1(B[59]), .A2(n198), .ZN(n199) );
  OR2_X1 U4 ( .A1(n196), .A2(B[62]), .ZN(n195) );
  OR3_X1 U5 ( .A1(B[57]), .A2(B[58]), .A3(n200), .ZN(n198) );
  OR2_X1 U6 ( .A1(n200), .A2(B[57]), .ZN(n201) );
  NOR2_X1 U7 ( .A1(B[47]), .A2(n212), .ZN(n213) );
  NOR2_X1 U8 ( .A1(B[43]), .A2(n216), .ZN(n217) );
  NOR2_X1 U9 ( .A1(B[39]), .A2(n220), .ZN(n221) );
  NOR2_X1 U10 ( .A1(B[35]), .A2(n224), .ZN(n225) );
  OR3_X1 U11 ( .A1(B[49]), .A2(B[50]), .A3(n208), .ZN(n206) );
  OR3_X1 U12 ( .A1(B[45]), .A2(B[46]), .A3(n214), .ZN(n212) );
  OR3_X1 U13 ( .A1(B[41]), .A2(B[42]), .A3(n218), .ZN(n216) );
  OR3_X1 U14 ( .A1(B[37]), .A2(B[38]), .A3(n222), .ZN(n220) );
  OR3_X1 U15 ( .A1(B[47]), .A2(B[48]), .A3(n212), .ZN(n208) );
  OR3_X1 U16 ( .A1(B[43]), .A2(B[44]), .A3(n216), .ZN(n214) );
  OR3_X1 U17 ( .A1(B[39]), .A2(B[40]), .A3(n220), .ZN(n218) );
  OR3_X1 U18 ( .A1(B[35]), .A2(B[36]), .A3(n224), .ZN(n222) );
  OR2_X1 U19 ( .A1(n208), .A2(B[49]), .ZN(n209) );
  OR2_X1 U20 ( .A1(n214), .A2(B[45]), .ZN(n215) );
  OR2_X1 U21 ( .A1(n218), .A2(B[41]), .ZN(n219) );
  OR2_X1 U22 ( .A1(n222), .A2(B[37]), .ZN(n223) );
  NOR2_X1 U23 ( .A1(B[55]), .A2(n202), .ZN(n203) );
  NOR2_X1 U24 ( .A1(B[51]), .A2(n206), .ZN(n207) );
  OR3_X1 U25 ( .A1(B[53]), .A2(B[54]), .A3(n204), .ZN(n202) );
  OR3_X1 U26 ( .A1(B[55]), .A2(B[56]), .A3(n202), .ZN(n200) );
  OR3_X1 U27 ( .A1(B[51]), .A2(B[52]), .A3(n206), .ZN(n204) );
  OR2_X1 U28 ( .A1(n204), .A2(B[53]), .ZN(n205) );
  OR3_X1 U29 ( .A1(B[33]), .A2(B[34]), .A3(n226), .ZN(n224) );
  OR2_X1 U30 ( .A1(n226), .A2(B[33]), .ZN(n227) );
  NOR2_X1 U31 ( .A1(B[31]), .A2(n228), .ZN(n229) );
  OR3_X1 U32 ( .A1(B[31]), .A2(B[32]), .A3(n228), .ZN(n226) );
  XNOR2_X1 U33 ( .A(B[52]), .B(n207), .ZN(DIFF[52]) );
  XNOR2_X1 U34 ( .A(B[48]), .B(n213), .ZN(DIFF[48]) );
  XNOR2_X1 U35 ( .A(B[44]), .B(n217), .ZN(DIFF[44]) );
  XNOR2_X1 U36 ( .A(B[40]), .B(n221), .ZN(DIFF[40]) );
  XNOR2_X1 U37 ( .A(B[36]), .B(n225), .ZN(DIFF[36]) );
  XNOR2_X1 U38 ( .A(B[32]), .B(n229), .ZN(DIFF[32]) );
  XNOR2_X1 U39 ( .A(B[60]), .B(n199), .ZN(DIFF[60]) );
  XNOR2_X1 U40 ( .A(B[56]), .B(n203), .ZN(DIFF[56]) );
  XNOR2_X1 U41 ( .A(n197), .B(B[61]), .ZN(DIFF[61]) );
  OR3_X1 U42 ( .A1(B[29]), .A2(B[30]), .A3(n230), .ZN(n228) );
  XNOR2_X1 U43 ( .A(B[28]), .B(n234), .ZN(DIFF[28]) );
  OR2_X1 U44 ( .A1(n230), .A2(B[29]), .ZN(n231) );
  NOR2_X1 U45 ( .A1(B[27]), .A2(n233), .ZN(n234) );
  OR3_X1 U46 ( .A1(B[27]), .A2(B[28]), .A3(n233), .ZN(n230) );
  XNOR2_X1 U47 ( .A(n189), .B(B[26]), .ZN(DIFF[26]) );
  NOR2_X1 U48 ( .A1(n235), .A2(B[25]), .ZN(n189) );
  OR3_X1 U49 ( .A1(B[25]), .A2(B[26]), .A3(n235), .ZN(n233) );
  NOR2_X1 U50 ( .A1(B[23]), .A2(n237), .ZN(n238) );
  NOR2_X1 U51 ( .A1(B[19]), .A2(n241), .ZN(n242) );
  NOR2_X1 U52 ( .A1(B[15]), .A2(n245), .ZN(n246) );
  NOR2_X1 U53 ( .A1(B[11]), .A2(n249), .ZN(n250) );
  NOR2_X1 U54 ( .A1(B[7]), .A2(n192), .ZN(n191) );
  NOR2_X1 U55 ( .A1(B[3]), .A2(n211), .ZN(n210) );
  OR3_X1 U56 ( .A1(B[21]), .A2(B[22]), .A3(n239), .ZN(n237) );
  OR3_X1 U57 ( .A1(B[17]), .A2(B[18]), .A3(n243), .ZN(n241) );
  OR3_X1 U58 ( .A1(B[13]), .A2(B[14]), .A3(n247), .ZN(n245) );
  OR3_X1 U59 ( .A1(B[10]), .A2(B[9]), .A3(n190), .ZN(n249) );
  OR3_X1 U60 ( .A1(B[5]), .A2(B[6]), .A3(n194), .ZN(n192) );
  OR3_X1 U61 ( .A1(B[23]), .A2(B[24]), .A3(n237), .ZN(n235) );
  OR3_X1 U62 ( .A1(B[19]), .A2(B[20]), .A3(n241), .ZN(n239) );
  OR3_X1 U63 ( .A1(B[15]), .A2(B[16]), .A3(n245), .ZN(n243) );
  OR3_X1 U64 ( .A1(B[11]), .A2(B[12]), .A3(n249), .ZN(n247) );
  OR3_X1 U65 ( .A1(B[7]), .A2(B[8]), .A3(n192), .ZN(n190) );
  OR3_X1 U66 ( .A1(B[3]), .A2(B[4]), .A3(n211), .ZN(n194) );
  XNOR2_X1 U67 ( .A(B[24]), .B(n238), .ZN(DIFF[24]) );
  XNOR2_X1 U68 ( .A(B[20]), .B(n242), .ZN(DIFF[20]) );
  XNOR2_X1 U69 ( .A(B[16]), .B(n246), .ZN(DIFF[16]) );
  XNOR2_X1 U70 ( .A(B[12]), .B(n250), .ZN(DIFF[12]) );
  XNOR2_X1 U71 ( .A(B[8]), .B(n191), .ZN(DIFF[8]) );
  XNOR2_X1 U72 ( .A(B[4]), .B(n210), .ZN(DIFF[4]) );
  XNOR2_X1 U73 ( .A(B[2]), .B(n232), .ZN(DIFF[2]) );
  OR2_X1 U74 ( .A1(n239), .A2(B[21]), .ZN(n240) );
  OR2_X1 U75 ( .A1(n243), .A2(B[17]), .ZN(n244) );
  OR2_X1 U76 ( .A1(n247), .A2(B[13]), .ZN(n248) );
  OR2_X1 U77 ( .A1(n190), .A2(B[9]), .ZN(n251) );
  OR2_X1 U78 ( .A1(n194), .A2(B[5]), .ZN(n193) );
  OR3_X1 U79 ( .A1(B[1]), .A2(B[2]), .A3(\B[0] ), .ZN(n211) );
  NOR2_X1 U80 ( .A1(\B[0] ), .A2(B[1]), .ZN(n232) );
  INV_X1 U113 ( .A(B[61]), .ZN(n236) );
endmodule


module complementer_N64_6 ( \input , complement2 );
  input [63:0] \input ;
  output [63:0] complement2;


  complementer_N64_6_DW01_sub_0 sub_add_31_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(\input ), .CI(1'b0), .DIFF(complement2) );
endmodule


module complementer_N64_5_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n190, n191, n192, n194, n196, n197, n198, n199, n200, n202,
         n203, n204, n206, n207, n208, n210, n211, n212, n213, n214, n216,
         n217, n218, n220, n221, n222, n224, n225, n226, n228, n229, n230,
         n232, n233, n234, n235, n236, n237, n238, n239, n241, n242, n243,
         n245, n246, n247, n249, n250, n189, n193, n195, n201, n205, n209,
         n215, n219, n223, n227, n231, n240, n244, n248, n251;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U81 ( .A(n190), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U82 ( .A(n192), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U85 ( .A(n196), .B(B[62]), .Z(DIFF[62]) );
  XOR2_X1 U86 ( .A(n194), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U87 ( .A(n198), .B(B[59]), .Z(DIFF[59]) );
  XOR2_X1 U89 ( .A(n200), .B(B[57]), .Z(DIFF[57]) );
  XOR2_X1 U90 ( .A(n202), .B(B[55]), .Z(DIFF[55]) );
  XOR2_X1 U92 ( .A(n204), .B(B[53]), .Z(DIFF[53]) );
  XOR2_X1 U93 ( .A(n206), .B(B[51]), .Z(DIFF[51]) );
  XOR2_X1 U95 ( .A(n208), .B(B[49]), .Z(DIFF[49]) );
  XOR2_X1 U96 ( .A(n212), .B(B[47]), .Z(DIFF[47]) );
  XOR2_X1 U98 ( .A(n214), .B(B[45]), .Z(DIFF[45]) );
  XOR2_X1 U99 ( .A(n216), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U101 ( .A(n218), .B(B[41]), .Z(DIFF[41]) );
  XOR2_X1 U102 ( .A(n211), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U103 ( .A(n220), .B(B[39]), .Z(DIFF[39]) );
  XOR2_X1 U105 ( .A(n222), .B(B[37]), .Z(DIFF[37]) );
  XOR2_X1 U106 ( .A(n224), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U108 ( .A(n226), .B(B[33]), .Z(DIFF[33]) );
  XOR2_X1 U109 ( .A(n228), .B(B[31]), .Z(DIFF[31]) );
  XOR2_X1 U111 ( .A(n230), .B(B[29]), .Z(DIFF[29]) );
  XOR2_X1 U112 ( .A(n233), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U113 ( .A(n236), .B(B[26]), .Z(DIFF[26]) );
  XOR2_X1 U114 ( .A(n235), .B(B[25]), .Z(DIFF[25]) );
  XOR2_X1 U115 ( .A(n237), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U117 ( .A(n239), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U118 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U119 ( .A(n241), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U121 ( .A(n243), .B(B[17]), .Z(DIFF[17]) );
  XOR2_X1 U122 ( .A(n245), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U124 ( .A(n247), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U125 ( .A(n249), .B(B[11]), .Z(DIFF[11]) );
  XOR2_X1 U1 ( .A(n197), .B(n251), .Z(DIFF[61]) );
  NAND2_X1 U2 ( .A1(n197), .A2(n251), .ZN(n196) );
  NOR3_X1 U3 ( .A1(B[59]), .A2(B[60]), .A3(n198), .ZN(n197) );
  XNOR2_X1 U4 ( .A(n189), .B(B[63]), .ZN(DIFF[63]) );
  NOR2_X1 U5 ( .A1(n196), .A2(B[62]), .ZN(n189) );
  XNOR2_X1 U6 ( .A(B[60]), .B(n199), .ZN(DIFF[60]) );
  NOR2_X1 U7 ( .A1(B[59]), .A2(n198), .ZN(n199) );
  XNOR2_X1 U8 ( .A(B[52]), .B(n207), .ZN(DIFF[52]) );
  NOR2_X1 U9 ( .A1(B[51]), .A2(n206), .ZN(n207) );
  XNOR2_X1 U10 ( .A(B[48]), .B(n213), .ZN(DIFF[48]) );
  NOR2_X1 U11 ( .A1(B[47]), .A2(n212), .ZN(n213) );
  XNOR2_X1 U12 ( .A(B[44]), .B(n217), .ZN(DIFF[44]) );
  NOR2_X1 U13 ( .A1(B[43]), .A2(n216), .ZN(n217) );
  XNOR2_X1 U14 ( .A(B[40]), .B(n221), .ZN(DIFF[40]) );
  NOR2_X1 U15 ( .A1(B[39]), .A2(n220), .ZN(n221) );
  OR3_X1 U16 ( .A1(B[37]), .A2(B[38]), .A3(n222), .ZN(n220) );
  OR3_X1 U17 ( .A1(B[41]), .A2(B[42]), .A3(n218), .ZN(n216) );
  OR3_X1 U18 ( .A1(B[45]), .A2(B[46]), .A3(n214), .ZN(n212) );
  OR3_X1 U19 ( .A1(B[49]), .A2(B[50]), .A3(n208), .ZN(n206) );
  OR3_X1 U20 ( .A1(B[39]), .A2(B[40]), .A3(n220), .ZN(n218) );
  OR3_X1 U21 ( .A1(B[43]), .A2(B[44]), .A3(n216), .ZN(n214) );
  OR3_X1 U22 ( .A1(B[47]), .A2(B[48]), .A3(n212), .ZN(n208) );
  XNOR2_X1 U23 ( .A(n193), .B(B[50]), .ZN(DIFF[50]) );
  NOR2_X1 U24 ( .A1(n208), .A2(B[49]), .ZN(n193) );
  XNOR2_X1 U25 ( .A(n195), .B(B[46]), .ZN(DIFF[46]) );
  NOR2_X1 U26 ( .A1(n214), .A2(B[45]), .ZN(n195) );
  XNOR2_X1 U27 ( .A(n201), .B(B[42]), .ZN(DIFF[42]) );
  NOR2_X1 U28 ( .A1(n218), .A2(B[41]), .ZN(n201) );
  XNOR2_X1 U29 ( .A(n205), .B(B[38]), .ZN(DIFF[38]) );
  NOR2_X1 U30 ( .A1(n222), .A2(B[37]), .ZN(n205) );
  XNOR2_X1 U31 ( .A(n209), .B(B[58]), .ZN(DIFF[58]) );
  NOR2_X1 U32 ( .A1(n200), .A2(B[57]), .ZN(n209) );
  XNOR2_X1 U33 ( .A(n215), .B(B[54]), .ZN(DIFF[54]) );
  NOR2_X1 U34 ( .A1(n204), .A2(B[53]), .ZN(n215) );
  XNOR2_X1 U35 ( .A(B[56]), .B(n203), .ZN(DIFF[56]) );
  NOR2_X1 U36 ( .A1(B[55]), .A2(n202), .ZN(n203) );
  OR3_X1 U37 ( .A1(B[57]), .A2(B[58]), .A3(n200), .ZN(n198) );
  OR3_X1 U38 ( .A1(B[53]), .A2(B[54]), .A3(n204), .ZN(n202) );
  OR3_X1 U39 ( .A1(B[51]), .A2(B[52]), .A3(n206), .ZN(n204) );
  OR3_X1 U40 ( .A1(B[55]), .A2(B[56]), .A3(n202), .ZN(n200) );
  XNOR2_X1 U41 ( .A(B[36]), .B(n225), .ZN(DIFF[36]) );
  NOR2_X1 U42 ( .A1(B[35]), .A2(n224), .ZN(n225) );
  OR3_X1 U43 ( .A1(B[35]), .A2(B[36]), .A3(n224), .ZN(n222) );
  XNOR2_X1 U44 ( .A(n219), .B(B[34]), .ZN(DIFF[34]) );
  NOR2_X1 U45 ( .A1(n226), .A2(B[33]), .ZN(n219) );
  OR3_X1 U46 ( .A1(B[33]), .A2(B[34]), .A3(n226), .ZN(n224) );
  XNOR2_X1 U47 ( .A(B[32]), .B(n229), .ZN(DIFF[32]) );
  NOR2_X1 U48 ( .A1(B[31]), .A2(n228), .ZN(n229) );
  OR3_X1 U49 ( .A1(B[31]), .A2(B[32]), .A3(n228), .ZN(n226) );
  XNOR2_X1 U50 ( .A(n223), .B(B[30]), .ZN(DIFF[30]) );
  NOR2_X1 U51 ( .A1(n230), .A2(B[29]), .ZN(n223) );
  OR3_X1 U52 ( .A1(B[29]), .A2(B[30]), .A3(n230), .ZN(n228) );
  XNOR2_X1 U53 ( .A(B[28]), .B(n234), .ZN(DIFF[28]) );
  NOR2_X1 U54 ( .A1(B[27]), .A2(n233), .ZN(n234) );
  OR3_X1 U55 ( .A1(B[27]), .A2(B[28]), .A3(n233), .ZN(n230) );
  XNOR2_X1 U56 ( .A(n227), .B(B[22]), .ZN(DIFF[22]) );
  NOR2_X1 U57 ( .A1(n239), .A2(B[21]), .ZN(n227) );
  XNOR2_X1 U58 ( .A(n231), .B(B[18]), .ZN(DIFF[18]) );
  NOR2_X1 U59 ( .A1(n243), .A2(B[17]), .ZN(n231) );
  XNOR2_X1 U60 ( .A(n240), .B(B[14]), .ZN(DIFF[14]) );
  NOR2_X1 U61 ( .A1(n247), .A2(B[13]), .ZN(n240) );
  XNOR2_X1 U62 ( .A(n244), .B(B[10]), .ZN(DIFF[10]) );
  NOR2_X1 U63 ( .A1(n190), .A2(B[9]), .ZN(n244) );
  XNOR2_X1 U64 ( .A(n248), .B(B[6]), .ZN(DIFF[6]) );
  NOR2_X1 U65 ( .A1(n194), .A2(B[5]), .ZN(n248) );
  XNOR2_X1 U66 ( .A(B[24]), .B(n238), .ZN(DIFF[24]) );
  NOR2_X1 U67 ( .A1(B[23]), .A2(n237), .ZN(n238) );
  XNOR2_X1 U68 ( .A(B[20]), .B(n242), .ZN(DIFF[20]) );
  NOR2_X1 U69 ( .A1(B[19]), .A2(n241), .ZN(n242) );
  XNOR2_X1 U70 ( .A(B[16]), .B(n246), .ZN(DIFF[16]) );
  NOR2_X1 U71 ( .A1(B[15]), .A2(n245), .ZN(n246) );
  XNOR2_X1 U72 ( .A(B[12]), .B(n250), .ZN(DIFF[12]) );
  NOR2_X1 U73 ( .A1(B[11]), .A2(n249), .ZN(n250) );
  XNOR2_X1 U74 ( .A(B[8]), .B(n191), .ZN(DIFF[8]) );
  NOR2_X1 U75 ( .A1(B[7]), .A2(n192), .ZN(n191) );
  XNOR2_X1 U76 ( .A(B[2]), .B(n232), .ZN(DIFF[2]) );
  NOR2_X1 U77 ( .A1(\B[0] ), .A2(B[1]), .ZN(n232) );
  XNOR2_X1 U78 ( .A(B[4]), .B(n210), .ZN(DIFF[4]) );
  NOR2_X1 U79 ( .A1(B[3]), .A2(n211), .ZN(n210) );
  OR3_X1 U80 ( .A1(B[5]), .A2(B[6]), .A3(n194), .ZN(n192) );
  OR3_X1 U83 ( .A1(B[10]), .A2(B[9]), .A3(n190), .ZN(n249) );
  OR3_X1 U84 ( .A1(B[13]), .A2(B[14]), .A3(n247), .ZN(n245) );
  OR3_X1 U88 ( .A1(B[17]), .A2(B[18]), .A3(n243), .ZN(n241) );
  OR3_X1 U91 ( .A1(B[21]), .A2(B[22]), .A3(n239), .ZN(n237) );
  OR3_X1 U94 ( .A1(B[25]), .A2(B[26]), .A3(n235), .ZN(n233) );
  OR3_X1 U97 ( .A1(B[7]), .A2(B[8]), .A3(n192), .ZN(n190) );
  OR3_X1 U100 ( .A1(B[11]), .A2(B[12]), .A3(n249), .ZN(n247) );
  OR3_X1 U104 ( .A1(B[15]), .A2(B[16]), .A3(n245), .ZN(n243) );
  OR3_X1 U107 ( .A1(B[19]), .A2(B[20]), .A3(n241), .ZN(n239) );
  OR3_X1 U110 ( .A1(B[23]), .A2(B[24]), .A3(n237), .ZN(n235) );
  OR3_X1 U116 ( .A1(B[3]), .A2(B[4]), .A3(n211), .ZN(n194) );
  OR2_X1 U120 ( .A1(n235), .A2(B[25]), .ZN(n236) );
  OR3_X1 U123 ( .A1(B[1]), .A2(B[2]), .A3(\B[0] ), .ZN(n211) );
  INV_X1 U126 ( .A(B[61]), .ZN(n251) );
endmodule


module complementer_N64_5 ( \input , complement2 );
  input [63:0] \input ;
  output [63:0] complement2;


  complementer_N64_5_DW01_sub_0 sub_add_31_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(\input ), .CI(1'b0), .DIFF(complement2) );
endmodule


module ShiftnCompl_N64_3 ( plusA, plus2A_out, minus2A_out, plus4A_out, 
        minus4A_out );
  input [63:0] plusA;
  output [63:0] plus2A_out;
  output [63:0] minus2A_out;
  output [63:0] plus4A_out;
  output [63:0] minus4A_out;
  wire   n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign plus2A_out[0] = 1'b0;
  assign plus4A_out[0] = 1'b0;

  shifter_N64_6 shifter_1 ( .\input (plusA), .shiftLeftOnePos({
        plus2A_out[63:59], n34, n35, n36, plus2A_out[55:1], 
        SYNOPSYS_UNCONNECTED__0}) );
  shifter_N64_5 shifter_2 ( .\input ({plus2A_out[63:1], 1'b0}), 
        .shiftLeftOnePos({plus4A_out[63:57], n37, n38, n39, n40, n41, n42, n43, 
        n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, 
        n58, n59, n60, n61, n62, n63, n64, n65, n66, plus4A_out[26:1], 
        SYNOPSYS_UNCONNECTED__1}) );
  complementer_N64_6 complementer_1 ( .\input ({plus2A_out[63:1], 1'b0}), 
        .complement2(minus2A_out) );
  complementer_N64_5 complementer_2 ( .\input ({plus4A_out[63:1], 1'b0}), 
        .complement2(minus4A_out) );
  BUF_X1 U3 ( .A(n50), .Z(plus4A_out[43]) );
  BUF_X1 U4 ( .A(n54), .Z(plus4A_out[39]) );
  BUF_X1 U5 ( .A(n36), .Z(plus2A_out[56]) );
  BUF_X1 U6 ( .A(n38), .Z(plus4A_out[55]) );
  BUF_X1 U7 ( .A(n42), .Z(plus4A_out[51]) );
  BUF_X1 U8 ( .A(n46), .Z(plus4A_out[47]) );
  BUF_X1 U9 ( .A(n35), .Z(plus2A_out[57]) );
  BUF_X1 U10 ( .A(n34), .Z(plus2A_out[58]) );
  BUF_X1 U11 ( .A(n66), .Z(plus4A_out[27]) );
  BUF_X1 U12 ( .A(n58), .Z(plus4A_out[35]) );
  BUF_X1 U13 ( .A(n62), .Z(plus4A_out[31]) );
  BUF_X1 U14 ( .A(n56), .Z(plus4A_out[37]) );
  BUF_X1 U15 ( .A(n60), .Z(plus4A_out[33]) );
  BUF_X1 U16 ( .A(n64), .Z(plus4A_out[29]) );
  BUF_X1 U17 ( .A(n57), .Z(plus4A_out[36]) );
  BUF_X1 U18 ( .A(n61), .Z(plus4A_out[32]) );
  BUF_X1 U19 ( .A(n65), .Z(plus4A_out[28]) );
  BUF_X1 U20 ( .A(n59), .Z(plus4A_out[34]) );
  BUF_X1 U21 ( .A(n63), .Z(plus4A_out[30]) );
  BUF_X1 U22 ( .A(n48), .Z(plus4A_out[45]) );
  BUF_X1 U23 ( .A(n52), .Z(plus4A_out[41]) );
  BUF_X1 U24 ( .A(n45), .Z(plus4A_out[48]) );
  BUF_X1 U25 ( .A(n49), .Z(plus4A_out[44]) );
  BUF_X1 U26 ( .A(n53), .Z(plus4A_out[40]) );
  BUF_X1 U27 ( .A(n47), .Z(plus4A_out[46]) );
  BUF_X1 U28 ( .A(n51), .Z(plus4A_out[42]) );
  BUF_X1 U29 ( .A(n55), .Z(plus4A_out[38]) );
  BUF_X1 U30 ( .A(n40), .Z(plus4A_out[53]) );
  BUF_X1 U31 ( .A(n44), .Z(plus4A_out[49]) );
  BUF_X1 U32 ( .A(n37), .Z(plus4A_out[56]) );
  BUF_X1 U33 ( .A(n41), .Z(plus4A_out[52]) );
  BUF_X1 U34 ( .A(n39), .Z(plus4A_out[54]) );
  BUF_X1 U35 ( .A(n43), .Z(plus4A_out[50]) );
endmodule


module MUX_GENERIC_N64_RADIX3_3 ( plusA, minusA, plus2A, minus2A, SEL, Y );
  input [63:0] plusA;
  input [63:0] minusA;
  input [63:0] plus2A;
  input [63:0] minus2A;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502;
  tri   [63:0] Y;

  TBUF_X1 \Y_tri[55]  ( .A(n446), .EN(n301), .Z(Y[55]) );
  TBUF_X1 \Y_tri[56]  ( .A(n445), .EN(n301), .Z(Y[56]) );
  TBUF_X1 \Y_tri[57]  ( .A(n444), .EN(n301), .Z(Y[57]) );
  TBUF_X1 \Y_tri[58]  ( .A(n443), .EN(n301), .Z(Y[58]) );
  TBUF_X1 \Y_tri[59]  ( .A(n442), .EN(n301), .Z(Y[59]) );
  TBUF_X1 \Y_tri[60]  ( .A(n441), .EN(n301), .Z(Y[60]) );
  TBUF_X1 \Y_tri[61]  ( .A(n440), .EN(n301), .Z(Y[61]) );
  TBUF_X1 \Y_tri[62]  ( .A(n439), .EN(n301), .Z(Y[62]) );
  TBUF_X1 \Y_tri[63]  ( .A(n438), .EN(n301), .Z(Y[63]) );
  TBUF_X1 \Y_tri[53]  ( .A(n448), .EN(n300), .Z(Y[53]) );
  TBUF_X1 \Y_tri[54]  ( .A(n447), .EN(n300), .Z(Y[54]) );
  TBUF_X1 \Y_tri[22]  ( .A(n479), .EN(n298), .Z(Y[22]) );
  TBUF_X1 \Y_tri[23]  ( .A(n478), .EN(n298), .Z(Y[23]) );
  TBUF_X1 \Y_tri[24]  ( .A(n477), .EN(n298), .Z(Y[24]) );
  TBUF_X1 \Y_tri[25]  ( .A(n476), .EN(n298), .Z(Y[25]) );
  TBUF_X1 \Y_tri[26]  ( .A(n475), .EN(n298), .Z(Y[26]) );
  TBUF_X1 \Y_tri[28]  ( .A(n473), .EN(n298), .Z(Y[28]) );
  TBUF_X1 \Y_tri[29]  ( .A(n472), .EN(n298), .Z(Y[29]) );
  TBUF_X1 \Y_tri[30]  ( .A(n471), .EN(n298), .Z(Y[30]) );
  TBUF_X1 \Y_tri[31]  ( .A(n470), .EN(n298), .Z(Y[31]) );
  TBUF_X1 \Y_tri[32]  ( .A(n469), .EN(n298), .Z(Y[32]) );
  TBUF_X1 \Y_tri[33]  ( .A(n468), .EN(n299), .Z(Y[33]) );
  TBUF_X1 \Y_tri[34]  ( .A(n467), .EN(n299), .Z(Y[34]) );
  TBUF_X1 \Y_tri[35]  ( .A(n466), .EN(n299), .Z(Y[35]) );
  TBUF_X1 \Y_tri[36]  ( .A(n465), .EN(n299), .Z(Y[36]) );
  TBUF_X1 \Y_tri[37]  ( .A(n464), .EN(n299), .Z(Y[37]) );
  TBUF_X1 \Y_tri[38]  ( .A(n463), .EN(n299), .Z(Y[38]) );
  TBUF_X1 \Y_tri[39]  ( .A(n462), .EN(n299), .Z(Y[39]) );
  TBUF_X1 \Y_tri[40]  ( .A(n461), .EN(n299), .Z(Y[40]) );
  TBUF_X1 \Y_tri[41]  ( .A(n460), .EN(n299), .Z(Y[41]) );
  TBUF_X1 \Y_tri[42]  ( .A(n459), .EN(n299), .Z(Y[42]) );
  TBUF_X1 \Y_tri[43]  ( .A(n458), .EN(n299), .Z(Y[43]) );
  TBUF_X1 \Y_tri[44]  ( .A(n457), .EN(n300), .Z(Y[44]) );
  TBUF_X1 \Y_tri[45]  ( .A(n456), .EN(n300), .Z(Y[45]) );
  TBUF_X1 \Y_tri[46]  ( .A(n455), .EN(n300), .Z(Y[46]) );
  TBUF_X1 \Y_tri[47]  ( .A(n454), .EN(n300), .Z(Y[47]) );
  TBUF_X1 \Y_tri[48]  ( .A(n453), .EN(n300), .Z(Y[48]) );
  TBUF_X1 \Y_tri[49]  ( .A(n452), .EN(n300), .Z(Y[49]) );
  TBUF_X1 \Y_tri[50]  ( .A(n451), .EN(n300), .Z(Y[50]) );
  TBUF_X1 \Y_tri[51]  ( .A(n450), .EN(n300), .Z(Y[51]) );
  TBUF_X1 \Y_tri[52]  ( .A(n449), .EN(n300), .Z(Y[52]) );
  TBUF_X1 \Y_tri[12]  ( .A(n489), .EN(n297), .Z(Y[12]) );
  TBUF_X1 \Y_tri[13]  ( .A(n488), .EN(n297), .Z(Y[13]) );
  TBUF_X1 \Y_tri[14]  ( .A(n487), .EN(n297), .Z(Y[14]) );
  TBUF_X1 \Y_tri[15]  ( .A(n486), .EN(n297), .Z(Y[15]) );
  TBUF_X1 \Y_tri[16]  ( .A(n485), .EN(n297), .Z(Y[16]) );
  TBUF_X1 \Y_tri[17]  ( .A(n484), .EN(n297), .Z(Y[17]) );
  TBUF_X1 \Y_tri[18]  ( .A(n483), .EN(n297), .Z(Y[18]) );
  TBUF_X1 \Y_tri[19]  ( .A(n482), .EN(n297), .Z(Y[19]) );
  TBUF_X1 \Y_tri[20]  ( .A(n481), .EN(n297), .Z(Y[20]) );
  TBUF_X1 \Y_tri[21]  ( .A(n480), .EN(n297), .Z(Y[21]) );
  TBUF_X1 \Y_tri[27]  ( .A(n474), .EN(n298), .Z(Y[27]) );
  TBUF_X1 \Y_tri[0]  ( .A(n502), .EN(n296), .Z(Y[0]) );
  TBUF_X1 \Y_tri[1]  ( .A(n501), .EN(n296), .Z(Y[1]) );
  TBUF_X1 \Y_tri[2]  ( .A(n500), .EN(n296), .Z(Y[2]) );
  TBUF_X1 \Y_tri[3]  ( .A(n499), .EN(n296), .Z(Y[3]) );
  TBUF_X1 \Y_tri[5]  ( .A(n497), .EN(n296), .Z(Y[5]) );
  TBUF_X1 \Y_tri[6]  ( .A(n496), .EN(n296), .Z(Y[6]) );
  TBUF_X1 \Y_tri[7]  ( .A(n495), .EN(n296), .Z(Y[7]) );
  TBUF_X1 \Y_tri[8]  ( .A(n494), .EN(n296), .Z(Y[8]) );
  TBUF_X1 \Y_tri[9]  ( .A(n492), .EN(n296), .Z(Y[9]) );
  TBUF_X1 \Y_tri[10]  ( .A(n491), .EN(n296), .Z(Y[10]) );
  TBUF_X1 \Y_tri[11]  ( .A(n490), .EN(n297), .Z(Y[11]) );
  TBUF_X1 \Y_tri[4]  ( .A(n498), .EN(n296), .Z(Y[4]) );
  NAND2_X1 U2 ( .A1(n409), .A2(n408), .ZN(n450) );
  AOI22_X1 U3 ( .A1(plusA[51]), .A2(n282), .B1(plus2A[51]), .B2(n276), .ZN(
        n409) );
  AOI22_X1 U4 ( .A1(minus2A[51]), .A2(n294), .B1(minusA[51]), .B2(n288), .ZN(
        n408) );
  NAND2_X1 U5 ( .A1(n401), .A2(n400), .ZN(n454) );
  AOI22_X1 U6 ( .A1(plusA[47]), .A2(n281), .B1(plus2A[47]), .B2(n275), .ZN(
        n401) );
  AOI22_X1 U7 ( .A1(minus2A[47]), .A2(n293), .B1(minusA[47]), .B2(n287), .ZN(
        n400) );
  NAND2_X1 U8 ( .A1(n393), .A2(n392), .ZN(n458) );
  AOI22_X1 U9 ( .A1(plusA[43]), .A2(n281), .B1(plus2A[43]), .B2(n275), .ZN(
        n393) );
  AOI22_X1 U10 ( .A1(minus2A[43]), .A2(n293), .B1(minusA[43]), .B2(n287), .ZN(
        n392) );
  NAND2_X1 U11 ( .A1(n385), .A2(n384), .ZN(n462) );
  AOI22_X1 U12 ( .A1(plusA[39]), .A2(n281), .B1(plus2A[39]), .B2(n275), .ZN(
        n385) );
  AOI22_X1 U13 ( .A1(minus2A[39]), .A2(n293), .B1(minusA[39]), .B2(n287), .ZN(
        n384) );
  NAND2_X1 U14 ( .A1(n377), .A2(n376), .ZN(n466) );
  AOI22_X1 U15 ( .A1(plusA[35]), .A2(n280), .B1(plus2A[35]), .B2(n274), .ZN(
        n377) );
  AOI22_X1 U16 ( .A1(minus2A[35]), .A2(n292), .B1(minusA[35]), .B2(n286), .ZN(
        n376) );
  NAND2_X1 U17 ( .A1(n369), .A2(n368), .ZN(n470) );
  AOI22_X1 U18 ( .A1(plusA[31]), .A2(n280), .B1(plus2A[31]), .B2(n274), .ZN(
        n369) );
  AOI22_X1 U19 ( .A1(minus2A[31]), .A2(n292), .B1(minusA[31]), .B2(n286), .ZN(
        n368) );
  NAND2_X1 U20 ( .A1(n405), .A2(n404), .ZN(n452) );
  AOI22_X1 U21 ( .A1(plusA[49]), .A2(n282), .B1(plus2A[49]), .B2(n276), .ZN(
        n405) );
  AOI22_X1 U22 ( .A1(minus2A[49]), .A2(n294), .B1(minusA[49]), .B2(n288), .ZN(
        n404) );
  NAND2_X1 U23 ( .A1(n397), .A2(n396), .ZN(n456) );
  AOI22_X1 U24 ( .A1(plusA[45]), .A2(n281), .B1(plus2A[45]), .B2(n275), .ZN(
        n397) );
  AOI22_X1 U25 ( .A1(minus2A[45]), .A2(n293), .B1(minusA[45]), .B2(n287), .ZN(
        n396) );
  NAND2_X1 U26 ( .A1(n389), .A2(n388), .ZN(n460) );
  AOI22_X1 U27 ( .A1(plusA[41]), .A2(n281), .B1(plus2A[41]), .B2(n275), .ZN(
        n389) );
  AOI22_X1 U28 ( .A1(minus2A[41]), .A2(n293), .B1(minusA[41]), .B2(n287), .ZN(
        n388) );
  NAND2_X1 U29 ( .A1(n381), .A2(n380), .ZN(n464) );
  AOI22_X1 U30 ( .A1(plusA[37]), .A2(n281), .B1(plus2A[37]), .B2(n275), .ZN(
        n381) );
  AOI22_X1 U31 ( .A1(minus2A[37]), .A2(n293), .B1(minusA[37]), .B2(n287), .ZN(
        n380) );
  NAND2_X1 U32 ( .A1(n373), .A2(n372), .ZN(n468) );
  AOI22_X1 U33 ( .A1(plusA[33]), .A2(n280), .B1(plus2A[33]), .B2(n274), .ZN(
        n373) );
  AOI22_X1 U34 ( .A1(minus2A[33]), .A2(n292), .B1(minusA[33]), .B2(n286), .ZN(
        n372) );
  NAND2_X1 U35 ( .A1(n411), .A2(n410), .ZN(n449) );
  AOI22_X1 U36 ( .A1(plusA[52]), .A2(n282), .B1(plus2A[52]), .B2(n276), .ZN(
        n411) );
  AOI22_X1 U37 ( .A1(minus2A[52]), .A2(n294), .B1(minusA[52]), .B2(n288), .ZN(
        n410) );
  NAND2_X1 U38 ( .A1(n403), .A2(n402), .ZN(n453) );
  AOI22_X1 U39 ( .A1(plusA[48]), .A2(n282), .B1(plus2A[48]), .B2(n276), .ZN(
        n403) );
  AOI22_X1 U40 ( .A1(minus2A[48]), .A2(n294), .B1(minusA[48]), .B2(n288), .ZN(
        n402) );
  NAND2_X1 U41 ( .A1(n395), .A2(n394), .ZN(n457) );
  AOI22_X1 U42 ( .A1(plusA[44]), .A2(n281), .B1(plus2A[44]), .B2(n275), .ZN(
        n395) );
  AOI22_X1 U43 ( .A1(minus2A[44]), .A2(n293), .B1(minusA[44]), .B2(n287), .ZN(
        n394) );
  NAND2_X1 U44 ( .A1(n387), .A2(n386), .ZN(n461) );
  AOI22_X1 U45 ( .A1(plusA[40]), .A2(n281), .B1(plus2A[40]), .B2(n275), .ZN(
        n387) );
  AOI22_X1 U46 ( .A1(minus2A[40]), .A2(n293), .B1(minusA[40]), .B2(n287), .ZN(
        n386) );
  NAND2_X1 U47 ( .A1(n379), .A2(n378), .ZN(n465) );
  AOI22_X1 U48 ( .A1(plusA[36]), .A2(n281), .B1(plus2A[36]), .B2(n275), .ZN(
        n379) );
  AOI22_X1 U49 ( .A1(minus2A[36]), .A2(n293), .B1(minusA[36]), .B2(n287), .ZN(
        n378) );
  NAND2_X1 U50 ( .A1(n371), .A2(n370), .ZN(n469) );
  AOI22_X1 U51 ( .A1(plusA[32]), .A2(n280), .B1(plus2A[32]), .B2(n274), .ZN(
        n371) );
  AOI22_X1 U52 ( .A1(minus2A[32]), .A2(n292), .B1(minusA[32]), .B2(n286), .ZN(
        n370) );
  NAND2_X1 U53 ( .A1(n407), .A2(n406), .ZN(n451) );
  AOI22_X1 U54 ( .A1(plusA[50]), .A2(n282), .B1(plus2A[50]), .B2(n276), .ZN(
        n407) );
  AOI22_X1 U55 ( .A1(minus2A[50]), .A2(n294), .B1(minusA[50]), .B2(n288), .ZN(
        n406) );
  NAND2_X1 U56 ( .A1(n399), .A2(n398), .ZN(n455) );
  AOI22_X1 U57 ( .A1(plusA[46]), .A2(n281), .B1(plus2A[46]), .B2(n275), .ZN(
        n399) );
  AOI22_X1 U58 ( .A1(minus2A[46]), .A2(n293), .B1(minusA[46]), .B2(n287), .ZN(
        n398) );
  NAND2_X1 U59 ( .A1(n391), .A2(n390), .ZN(n459) );
  AOI22_X1 U60 ( .A1(plusA[42]), .A2(n281), .B1(plus2A[42]), .B2(n275), .ZN(
        n391) );
  AOI22_X1 U61 ( .A1(minus2A[42]), .A2(n293), .B1(minusA[42]), .B2(n287), .ZN(
        n390) );
  NAND2_X1 U62 ( .A1(n383), .A2(n382), .ZN(n463) );
  AOI22_X1 U63 ( .A1(plusA[38]), .A2(n281), .B1(plus2A[38]), .B2(n275), .ZN(
        n383) );
  AOI22_X1 U64 ( .A1(minus2A[38]), .A2(n293), .B1(minusA[38]), .B2(n287), .ZN(
        n382) );
  NAND2_X1 U65 ( .A1(n375), .A2(n374), .ZN(n467) );
  AOI22_X1 U66 ( .A1(plusA[34]), .A2(n280), .B1(plus2A[34]), .B2(n274), .ZN(
        n375) );
  AOI22_X1 U67 ( .A1(minus2A[34]), .A2(n292), .B1(minusA[34]), .B2(n286), .ZN(
        n374) );
  NAND2_X1 U68 ( .A1(n367), .A2(n366), .ZN(n471) );
  AOI22_X1 U69 ( .A1(plusA[30]), .A2(n280), .B1(plus2A[30]), .B2(n274), .ZN(
        n367) );
  AOI22_X1 U70 ( .A1(minus2A[30]), .A2(n292), .B1(minusA[30]), .B2(n286), .ZN(
        n366) );
  NAND2_X1 U71 ( .A1(n425), .A2(n424), .ZN(n442) );
  AOI22_X1 U72 ( .A1(plusA[59]), .A2(n282), .B1(plus2A[59]), .B2(n276), .ZN(
        n425) );
  AOI22_X1 U73 ( .A1(minus2A[59]), .A2(n294), .B1(minusA[59]), .B2(n288), .ZN(
        n424) );
  NAND2_X1 U74 ( .A1(n423), .A2(n422), .ZN(n443) );
  AOI22_X1 U75 ( .A1(plusA[58]), .A2(n282), .B1(plus2A[58]), .B2(n276), .ZN(
        n423) );
  AOI22_X1 U76 ( .A1(minus2A[58]), .A2(n294), .B1(minusA[58]), .B2(n288), .ZN(
        n422) );
  NAND2_X1 U77 ( .A1(n431), .A2(n430), .ZN(n439) );
  AOI22_X1 U78 ( .A1(plusA[62]), .A2(n283), .B1(plus2A[62]), .B2(n277), .ZN(
        n431) );
  AOI22_X1 U79 ( .A1(minus2A[62]), .A2(n295), .B1(minusA[62]), .B2(n289), .ZN(
        n430) );
  NAND2_X1 U80 ( .A1(n427), .A2(n426), .ZN(n441) );
  AOI22_X1 U81 ( .A1(plusA[60]), .A2(n283), .B1(plus2A[60]), .B2(n277), .ZN(
        n427) );
  AOI22_X1 U82 ( .A1(minus2A[60]), .A2(n295), .B1(minusA[60]), .B2(n289), .ZN(
        n426) );
  NAND2_X1 U83 ( .A1(n421), .A2(n420), .ZN(n444) );
  AOI22_X1 U84 ( .A1(plusA[57]), .A2(n282), .B1(plus2A[57]), .B2(n276), .ZN(
        n421) );
  AOI22_X1 U85 ( .A1(minus2A[57]), .A2(n294), .B1(minusA[57]), .B2(n288), .ZN(
        n420) );
  NAND2_X1 U86 ( .A1(n417), .A2(n416), .ZN(n446) );
  AOI22_X1 U87 ( .A1(plusA[55]), .A2(n282), .B1(plus2A[55]), .B2(n276), .ZN(
        n417) );
  AOI22_X1 U88 ( .A1(minus2A[55]), .A2(n294), .B1(minusA[55]), .B2(n288), .ZN(
        n416) );
  NAND2_X1 U89 ( .A1(n413), .A2(n412), .ZN(n448) );
  AOI22_X1 U90 ( .A1(plusA[53]), .A2(n282), .B1(plus2A[53]), .B2(n276), .ZN(
        n413) );
  AOI22_X1 U91 ( .A1(minus2A[53]), .A2(n294), .B1(minusA[53]), .B2(n288), .ZN(
        n412) );
  NAND2_X1 U92 ( .A1(n419), .A2(n418), .ZN(n445) );
  AOI22_X1 U93 ( .A1(plusA[56]), .A2(n282), .B1(plus2A[56]), .B2(n276), .ZN(
        n419) );
  AOI22_X1 U94 ( .A1(minus2A[56]), .A2(n294), .B1(minusA[56]), .B2(n288), .ZN(
        n418) );
  NAND2_X1 U95 ( .A1(n415), .A2(n414), .ZN(n447) );
  AOI22_X1 U96 ( .A1(plusA[54]), .A2(n282), .B1(plus2A[54]), .B2(n276), .ZN(
        n415) );
  AOI22_X1 U97 ( .A1(minus2A[54]), .A2(n294), .B1(minusA[54]), .B2(n288), .ZN(
        n414) );
  NAND2_X1 U98 ( .A1(n437), .A2(n436), .ZN(n438) );
  AOI22_X1 U99 ( .A1(plusA[63]), .A2(n283), .B1(plus2A[63]), .B2(n277), .ZN(
        n437) );
  AOI22_X1 U100 ( .A1(minus2A[63]), .A2(n295), .B1(minusA[63]), .B2(n289), 
        .ZN(n436) );
  NAND2_X1 U101 ( .A1(n429), .A2(n428), .ZN(n440) );
  AOI22_X1 U102 ( .A1(plusA[61]), .A2(n283), .B1(plus2A[61]), .B2(n277), .ZN(
        n429) );
  AOI22_X1 U103 ( .A1(minus2A[61]), .A2(n295), .B1(minusA[61]), .B2(n289), 
        .ZN(n428) );
  BUF_X1 U104 ( .A(n493), .Z(n296) );
  BUF_X1 U105 ( .A(n493), .Z(n297) );
  BUF_X1 U106 ( .A(n433), .Z(n280) );
  BUF_X1 U107 ( .A(n435), .Z(n292) );
  BUF_X1 U108 ( .A(n434), .Z(n286) );
  BUF_X1 U109 ( .A(n432), .Z(n274) );
  BUF_X1 U110 ( .A(n493), .Z(n298) );
  NAND2_X1 U111 ( .A1(n365), .A2(n364), .ZN(n472) );
  AOI22_X1 U112 ( .A1(plusA[29]), .A2(n280), .B1(plus2A[29]), .B2(n274), .ZN(
        n365) );
  AOI22_X1 U113 ( .A1(minus2A[29]), .A2(n292), .B1(minusA[29]), .B2(n286), 
        .ZN(n364) );
  NAND2_X1 U114 ( .A1(n363), .A2(n362), .ZN(n473) );
  AOI22_X1 U115 ( .A1(plusA[28]), .A2(n280), .B1(plus2A[28]), .B2(n274), .ZN(
        n363) );
  AOI22_X1 U116 ( .A1(minus2A[28]), .A2(n292), .B1(minusA[28]), .B2(n286), 
        .ZN(n362) );
  BUF_X1 U117 ( .A(n433), .Z(n281) );
  BUF_X1 U118 ( .A(n435), .Z(n293) );
  BUF_X1 U119 ( .A(n434), .Z(n287) );
  BUF_X1 U120 ( .A(n432), .Z(n275) );
  BUF_X1 U121 ( .A(n493), .Z(n299) );
  BUF_X1 U122 ( .A(n433), .Z(n282) );
  BUF_X1 U123 ( .A(n435), .Z(n294) );
  BUF_X1 U124 ( .A(n434), .Z(n288) );
  BUF_X1 U125 ( .A(n432), .Z(n276) );
  BUF_X1 U126 ( .A(n493), .Z(n300) );
  BUF_X1 U127 ( .A(n493), .Z(n301) );
  BUF_X1 U128 ( .A(n433), .Z(n279) );
  BUF_X1 U129 ( .A(n433), .Z(n278) );
  BUF_X1 U130 ( .A(n435), .Z(n291) );
  BUF_X1 U131 ( .A(n435), .Z(n290) );
  BUF_X1 U132 ( .A(n434), .Z(n285) );
  BUF_X1 U133 ( .A(n432), .Z(n273) );
  BUF_X1 U134 ( .A(n434), .Z(n284) );
  BUF_X1 U135 ( .A(n432), .Z(n272) );
  NOR2_X1 U136 ( .A1(n323), .A2(n304), .ZN(n493) );
  INV_X1 U137 ( .A(SEL[2]), .ZN(n304) );
  NOR2_X1 U138 ( .A1(SEL[1]), .A2(SEL[0]), .ZN(n323) );
  NAND2_X1 U139 ( .A1(n361), .A2(n360), .ZN(n474) );
  AOI22_X1 U140 ( .A1(plusA[27]), .A2(n280), .B1(plus2A[27]), .B2(n274), .ZN(
        n361) );
  AOI22_X1 U141 ( .A1(minus2A[27]), .A2(n292), .B1(minusA[27]), .B2(n286), 
        .ZN(n360) );
  NOR3_X1 U142 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n302), .ZN(n434) );
  NOR3_X1 U143 ( .A1(SEL[1]), .A2(SEL[2]), .A3(n303), .ZN(n433) );
  NOR3_X1 U144 ( .A1(n302), .A2(SEL[2]), .A3(n303), .ZN(n432) );
  AND2_X1 U145 ( .A1(SEL[2]), .A2(n323), .ZN(n435) );
  INV_X1 U146 ( .A(SEL[1]), .ZN(n302) );
  INV_X1 U147 ( .A(SEL[0]), .ZN(n303) );
  NAND2_X1 U148 ( .A1(n359), .A2(n358), .ZN(n475) );
  AOI22_X1 U149 ( .A1(plusA[26]), .A2(n280), .B1(plus2A[26]), .B2(n274), .ZN(
        n359) );
  AOI22_X1 U150 ( .A1(minus2A[26]), .A2(n292), .B1(minusA[26]), .B2(n286), 
        .ZN(n358) );
  NAND2_X1 U151 ( .A1(n357), .A2(n356), .ZN(n476) );
  AOI22_X1 U152 ( .A1(plusA[25]), .A2(n280), .B1(plus2A[25]), .B2(n274), .ZN(
        n357) );
  AOI22_X1 U153 ( .A1(minus2A[25]), .A2(n292), .B1(minusA[25]), .B2(n286), 
        .ZN(n356) );
  NAND2_X1 U154 ( .A1(n353), .A2(n352), .ZN(n478) );
  AOI22_X1 U155 ( .A1(plusA[23]), .A2(n279), .B1(plus2A[23]), .B2(n273), .ZN(
        n353) );
  AOI22_X1 U156 ( .A1(minus2A[23]), .A2(n291), .B1(minusA[23]), .B2(n285), 
        .ZN(n352) );
  NAND2_X1 U157 ( .A1(n351), .A2(n350), .ZN(n479) );
  AOI22_X1 U158 ( .A1(plusA[22]), .A2(n279), .B1(plus2A[22]), .B2(n273), .ZN(
        n351) );
  AOI22_X1 U159 ( .A1(minus2A[22]), .A2(n291), .B1(minusA[22]), .B2(n285), 
        .ZN(n350) );
  NAND2_X1 U160 ( .A1(n349), .A2(n348), .ZN(n480) );
  AOI22_X1 U161 ( .A1(plusA[21]), .A2(n279), .B1(plus2A[21]), .B2(n273), .ZN(
        n349) );
  AOI22_X1 U162 ( .A1(minus2A[21]), .A2(n291), .B1(minusA[21]), .B2(n285), 
        .ZN(n348) );
  NAND2_X1 U163 ( .A1(n345), .A2(n344), .ZN(n482) );
  AOI22_X1 U164 ( .A1(plusA[19]), .A2(n279), .B1(plus2A[19]), .B2(n273), .ZN(
        n345) );
  AOI22_X1 U165 ( .A1(minus2A[19]), .A2(n291), .B1(minusA[19]), .B2(n285), 
        .ZN(n344) );
  NAND2_X1 U166 ( .A1(n343), .A2(n342), .ZN(n483) );
  AOI22_X1 U167 ( .A1(plusA[18]), .A2(n279), .B1(plus2A[18]), .B2(n273), .ZN(
        n343) );
  AOI22_X1 U168 ( .A1(minus2A[18]), .A2(n291), .B1(minusA[18]), .B2(n285), 
        .ZN(n342) );
  NAND2_X1 U169 ( .A1(n341), .A2(n340), .ZN(n484) );
  AOI22_X1 U170 ( .A1(plusA[17]), .A2(n279), .B1(plus2A[17]), .B2(n273), .ZN(
        n341) );
  AOI22_X1 U171 ( .A1(minus2A[17]), .A2(n291), .B1(minusA[17]), .B2(n285), 
        .ZN(n340) );
  NAND2_X1 U172 ( .A1(n337), .A2(n336), .ZN(n486) );
  AOI22_X1 U173 ( .A1(plusA[15]), .A2(n279), .B1(plus2A[15]), .B2(n273), .ZN(
        n337) );
  AOI22_X1 U174 ( .A1(minus2A[15]), .A2(n291), .B1(minusA[15]), .B2(n285), 
        .ZN(n336) );
  NAND2_X1 U175 ( .A1(n335), .A2(n334), .ZN(n487) );
  AOI22_X1 U176 ( .A1(plusA[14]), .A2(n279), .B1(plus2A[14]), .B2(n273), .ZN(
        n335) );
  AOI22_X1 U177 ( .A1(minus2A[14]), .A2(n291), .B1(minusA[14]), .B2(n285), 
        .ZN(n334) );
  NAND2_X1 U178 ( .A1(n333), .A2(n332), .ZN(n488) );
  AOI22_X1 U179 ( .A1(plusA[13]), .A2(n279), .B1(plus2A[13]), .B2(n273), .ZN(
        n333) );
  AOI22_X1 U180 ( .A1(minus2A[13]), .A2(n291), .B1(minusA[13]), .B2(n285), 
        .ZN(n332) );
  NAND2_X1 U181 ( .A1(n329), .A2(n328), .ZN(n490) );
  AOI22_X1 U182 ( .A1(plusA[11]), .A2(n278), .B1(plus2A[11]), .B2(n272), .ZN(
        n329) );
  AOI22_X1 U183 ( .A1(minus2A[11]), .A2(n290), .B1(minusA[11]), .B2(n284), 
        .ZN(n328) );
  NAND2_X1 U184 ( .A1(n327), .A2(n326), .ZN(n491) );
  AOI22_X1 U185 ( .A1(plusA[10]), .A2(n278), .B1(plus2A[10]), .B2(n272), .ZN(
        n327) );
  AOI22_X1 U186 ( .A1(minus2A[10]), .A2(n290), .B1(minusA[10]), .B2(n284), 
        .ZN(n326) );
  NAND2_X1 U187 ( .A1(n325), .A2(n324), .ZN(n492) );
  AOI22_X1 U188 ( .A1(plusA[9]), .A2(n278), .B1(plus2A[9]), .B2(n272), .ZN(
        n325) );
  AOI22_X1 U189 ( .A1(minus2A[9]), .A2(n290), .B1(minusA[9]), .B2(n284), .ZN(
        n324) );
  NAND2_X1 U190 ( .A1(n320), .A2(n319), .ZN(n495) );
  AOI22_X1 U191 ( .A1(plusA[7]), .A2(n278), .B1(plus2A[7]), .B2(n272), .ZN(
        n320) );
  AOI22_X1 U192 ( .A1(minus2A[7]), .A2(n290), .B1(minusA[7]), .B2(n284), .ZN(
        n319) );
  NAND2_X1 U193 ( .A1(n318), .A2(n317), .ZN(n496) );
  AOI22_X1 U194 ( .A1(plusA[6]), .A2(n278), .B1(plus2A[6]), .B2(n272), .ZN(
        n318) );
  AOI22_X1 U195 ( .A1(minus2A[6]), .A2(n290), .B1(minusA[6]), .B2(n284), .ZN(
        n317) );
  NAND2_X1 U196 ( .A1(n316), .A2(n315), .ZN(n497) );
  AOI22_X1 U197 ( .A1(plusA[5]), .A2(n278), .B1(plus2A[5]), .B2(n272), .ZN(
        n316) );
  AOI22_X1 U198 ( .A1(minus2A[5]), .A2(n290), .B1(minusA[5]), .B2(n284), .ZN(
        n315) );
  NAND2_X1 U199 ( .A1(n312), .A2(n311), .ZN(n499) );
  AOI22_X1 U200 ( .A1(plusA[3]), .A2(n278), .B1(plus2A[3]), .B2(n272), .ZN(
        n312) );
  AOI22_X1 U201 ( .A1(minus2A[3]), .A2(n290), .B1(minusA[3]), .B2(n284), .ZN(
        n311) );
  NAND2_X1 U202 ( .A1(n355), .A2(n354), .ZN(n477) );
  AOI22_X1 U203 ( .A1(plusA[24]), .A2(n280), .B1(plus2A[24]), .B2(n274), .ZN(
        n355) );
  AOI22_X1 U204 ( .A1(minus2A[24]), .A2(n292), .B1(minusA[24]), .B2(n286), 
        .ZN(n354) );
  NAND2_X1 U205 ( .A1(n347), .A2(n346), .ZN(n481) );
  AOI22_X1 U206 ( .A1(plusA[20]), .A2(n279), .B1(plus2A[20]), .B2(n273), .ZN(
        n347) );
  AOI22_X1 U207 ( .A1(minus2A[20]), .A2(n291), .B1(minusA[20]), .B2(n285), 
        .ZN(n346) );
  NAND2_X1 U208 ( .A1(n339), .A2(n338), .ZN(n485) );
  AOI22_X1 U209 ( .A1(plusA[16]), .A2(n279), .B1(plus2A[16]), .B2(n273), .ZN(
        n339) );
  AOI22_X1 U210 ( .A1(minus2A[16]), .A2(n291), .B1(minusA[16]), .B2(n285), 
        .ZN(n338) );
  NAND2_X1 U211 ( .A1(n331), .A2(n330), .ZN(n489) );
  AOI22_X1 U212 ( .A1(plusA[12]), .A2(n279), .B1(plus2A[12]), .B2(n273), .ZN(
        n331) );
  AOI22_X1 U213 ( .A1(minus2A[12]), .A2(n291), .B1(minusA[12]), .B2(n285), 
        .ZN(n330) );
  NAND2_X1 U214 ( .A1(n322), .A2(n321), .ZN(n494) );
  AOI22_X1 U215 ( .A1(plusA[8]), .A2(n278), .B1(plus2A[8]), .B2(n272), .ZN(
        n322) );
  AOI22_X1 U216 ( .A1(minus2A[8]), .A2(n290), .B1(minusA[8]), .B2(n284), .ZN(
        n321) );
  NAND2_X1 U217 ( .A1(n314), .A2(n313), .ZN(n498) );
  AOI22_X1 U218 ( .A1(plusA[4]), .A2(n278), .B1(plus2A[4]), .B2(n272), .ZN(
        n314) );
  AOI22_X1 U219 ( .A1(minus2A[4]), .A2(n290), .B1(minusA[4]), .B2(n284), .ZN(
        n313) );
  NAND2_X1 U220 ( .A1(n310), .A2(n309), .ZN(n500) );
  AOI22_X1 U221 ( .A1(plusA[2]), .A2(n278), .B1(plus2A[2]), .B2(n272), .ZN(
        n310) );
  AOI22_X1 U222 ( .A1(minus2A[2]), .A2(n290), .B1(minusA[2]), .B2(n284), .ZN(
        n309) );
  NAND2_X1 U223 ( .A1(n308), .A2(n307), .ZN(n501) );
  AOI22_X1 U224 ( .A1(plusA[1]), .A2(n278), .B1(plus2A[1]), .B2(n272), .ZN(
        n308) );
  AOI22_X1 U225 ( .A1(minus2A[1]), .A2(n290), .B1(minusA[1]), .B2(n284), .ZN(
        n307) );
  NAND2_X1 U226 ( .A1(n306), .A2(n305), .ZN(n502) );
  AOI22_X1 U227 ( .A1(plusA[0]), .A2(n278), .B1(plus2A[0]), .B2(n272), .ZN(
        n306) );
  AOI22_X1 U228 ( .A1(minus2A[0]), .A2(n290), .B1(minusA[0]), .B2(n284), .ZN(
        n305) );
  CLKBUF_X1 U229 ( .A(n432), .Z(n277) );
  CLKBUF_X1 U230 ( .A(n433), .Z(n283) );
  CLKBUF_X1 U231 ( .A(n434), .Z(n289) );
  CLKBUF_X1 U232 ( .A(n435), .Z(n295) );
endmodule


module FA_192 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_191 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_190 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_189 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_188 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  AOI22_X1 U4 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
  INV_X1 U5 ( .A(n7), .ZN(Co) );
endmodule


module FA_187 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_186 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_185 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_184 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_183 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_182 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_181 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_180 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_179 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_178 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_177 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_176 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_175 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_174 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_173 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_172 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_171 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_170 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_169 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_168 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_167 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_166 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_165 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_164 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_163 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_162 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_161 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_160 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_159 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_158 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_157 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_156 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_155 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_154 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_153 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_152 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_151 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_150 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_149 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_148 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_147 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_146 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_145 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_144 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_143 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_142 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_141 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_140 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_139 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_138 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_137 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_136 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_135 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_134 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_133 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_132 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_131 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_130 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_129 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N64_3 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Ci;
  output Co;

  wire   [63:1] CTMP;
  tri   [63:0] A;

  FA_192 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_191 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_190 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_189 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(CTMP[4]) );
  FA_188 FAI_5 ( .A(A[4]), .B(B[4]), .Ci(CTMP[4]), .S(S[4]), .Co(CTMP[5]) );
  FA_187 FAI_6 ( .A(A[5]), .B(B[5]), .Ci(CTMP[5]), .S(S[5]), .Co(CTMP[6]) );
  FA_186 FAI_7 ( .A(A[6]), .B(B[6]), .Ci(CTMP[6]), .S(S[6]), .Co(CTMP[7]) );
  FA_185 FAI_8 ( .A(A[7]), .B(B[7]), .Ci(CTMP[7]), .S(S[7]), .Co(CTMP[8]) );
  FA_184 FAI_9 ( .A(A[8]), .B(B[8]), .Ci(CTMP[8]), .S(S[8]), .Co(CTMP[9]) );
  FA_183 FAI_10 ( .A(A[9]), .B(B[9]), .Ci(CTMP[9]), .S(S[9]), .Co(CTMP[10]) );
  FA_182 FAI_11 ( .A(A[10]), .B(B[10]), .Ci(CTMP[10]), .S(S[10]), .Co(CTMP[11]) );
  FA_181 FAI_12 ( .A(A[11]), .B(B[11]), .Ci(CTMP[11]), .S(S[11]), .Co(CTMP[12]) );
  FA_180 FAI_13 ( .A(A[12]), .B(B[12]), .Ci(CTMP[12]), .S(S[12]), .Co(CTMP[13]) );
  FA_179 FAI_14 ( .A(A[13]), .B(B[13]), .Ci(CTMP[13]), .S(S[13]), .Co(CTMP[14]) );
  FA_178 FAI_15 ( .A(A[14]), .B(B[14]), .Ci(CTMP[14]), .S(S[14]), .Co(CTMP[15]) );
  FA_177 FAI_16 ( .A(A[15]), .B(B[15]), .Ci(CTMP[15]), .S(S[15]), .Co(CTMP[16]) );
  FA_176 FAI_17 ( .A(A[16]), .B(B[16]), .Ci(CTMP[16]), .S(S[16]), .Co(CTMP[17]) );
  FA_175 FAI_18 ( .A(A[17]), .B(B[17]), .Ci(CTMP[17]), .S(S[17]), .Co(CTMP[18]) );
  FA_174 FAI_19 ( .A(A[18]), .B(B[18]), .Ci(CTMP[18]), .S(S[18]), .Co(CTMP[19]) );
  FA_173 FAI_20 ( .A(A[19]), .B(B[19]), .Ci(CTMP[19]), .S(S[19]), .Co(CTMP[20]) );
  FA_172 FAI_21 ( .A(A[20]), .B(B[20]), .Ci(CTMP[20]), .S(S[20]), .Co(CTMP[21]) );
  FA_171 FAI_22 ( .A(A[21]), .B(B[21]), .Ci(CTMP[21]), .S(S[21]), .Co(CTMP[22]) );
  FA_170 FAI_23 ( .A(A[22]), .B(B[22]), .Ci(CTMP[22]), .S(S[22]), .Co(CTMP[23]) );
  FA_169 FAI_24 ( .A(A[23]), .B(B[23]), .Ci(CTMP[23]), .S(S[23]), .Co(CTMP[24]) );
  FA_168 FAI_25 ( .A(A[24]), .B(B[24]), .Ci(CTMP[24]), .S(S[24]), .Co(CTMP[25]) );
  FA_167 FAI_26 ( .A(A[25]), .B(B[25]), .Ci(CTMP[25]), .S(S[25]), .Co(CTMP[26]) );
  FA_166 FAI_27 ( .A(A[26]), .B(B[26]), .Ci(CTMP[26]), .S(S[26]), .Co(CTMP[27]) );
  FA_165 FAI_28 ( .A(A[27]), .B(B[27]), .Ci(CTMP[27]), .S(S[27]), .Co(CTMP[28]) );
  FA_164 FAI_29 ( .A(A[28]), .B(B[28]), .Ci(CTMP[28]), .S(S[28]), .Co(CTMP[29]) );
  FA_163 FAI_30 ( .A(A[29]), .B(B[29]), .Ci(CTMP[29]), .S(S[29]), .Co(CTMP[30]) );
  FA_162 FAI_31 ( .A(A[30]), .B(B[30]), .Ci(CTMP[30]), .S(S[30]), .Co(CTMP[31]) );
  FA_161 FAI_32 ( .A(A[31]), .B(B[31]), .Ci(CTMP[31]), .S(S[31]), .Co(CTMP[32]) );
  FA_160 FAI_33 ( .A(A[32]), .B(B[32]), .Ci(CTMP[32]), .S(S[32]), .Co(CTMP[33]) );
  FA_159 FAI_34 ( .A(A[33]), .B(B[33]), .Ci(CTMP[33]), .S(S[33]), .Co(CTMP[34]) );
  FA_158 FAI_35 ( .A(A[34]), .B(B[34]), .Ci(CTMP[34]), .S(S[34]), .Co(CTMP[35]) );
  FA_157 FAI_36 ( .A(A[35]), .B(B[35]), .Ci(CTMP[35]), .S(S[35]), .Co(CTMP[36]) );
  FA_156 FAI_37 ( .A(A[36]), .B(B[36]), .Ci(CTMP[36]), .S(S[36]), .Co(CTMP[37]) );
  FA_155 FAI_38 ( .A(A[37]), .B(B[37]), .Ci(CTMP[37]), .S(S[37]), .Co(CTMP[38]) );
  FA_154 FAI_39 ( .A(A[38]), .B(B[38]), .Ci(CTMP[38]), .S(S[38]), .Co(CTMP[39]) );
  FA_153 FAI_40 ( .A(A[39]), .B(B[39]), .Ci(CTMP[39]), .S(S[39]), .Co(CTMP[40]) );
  FA_152 FAI_41 ( .A(A[40]), .B(B[40]), .Ci(CTMP[40]), .S(S[40]), .Co(CTMP[41]) );
  FA_151 FAI_42 ( .A(A[41]), .B(B[41]), .Ci(CTMP[41]), .S(S[41]), .Co(CTMP[42]) );
  FA_150 FAI_43 ( .A(A[42]), .B(B[42]), .Ci(CTMP[42]), .S(S[42]), .Co(CTMP[43]) );
  FA_149 FAI_44 ( .A(A[43]), .B(B[43]), .Ci(CTMP[43]), .S(S[43]), .Co(CTMP[44]) );
  FA_148 FAI_45 ( .A(A[44]), .B(B[44]), .Ci(CTMP[44]), .S(S[44]), .Co(CTMP[45]) );
  FA_147 FAI_46 ( .A(A[45]), .B(B[45]), .Ci(CTMP[45]), .S(S[45]), .Co(CTMP[46]) );
  FA_146 FAI_47 ( .A(A[46]), .B(B[46]), .Ci(CTMP[46]), .S(S[46]), .Co(CTMP[47]) );
  FA_145 FAI_48 ( .A(A[47]), .B(B[47]), .Ci(CTMP[47]), .S(S[47]), .Co(CTMP[48]) );
  FA_144 FAI_49 ( .A(A[48]), .B(B[48]), .Ci(CTMP[48]), .S(S[48]), .Co(CTMP[49]) );
  FA_143 FAI_50 ( .A(A[49]), .B(B[49]), .Ci(CTMP[49]), .S(S[49]), .Co(CTMP[50]) );
  FA_142 FAI_51 ( .A(A[50]), .B(B[50]), .Ci(CTMP[50]), .S(S[50]), .Co(CTMP[51]) );
  FA_141 FAI_52 ( .A(A[51]), .B(B[51]), .Ci(CTMP[51]), .S(S[51]), .Co(CTMP[52]) );
  FA_140 FAI_53 ( .A(A[52]), .B(B[52]), .Ci(CTMP[52]), .S(S[52]), .Co(CTMP[53]) );
  FA_139 FAI_54 ( .A(A[53]), .B(B[53]), .Ci(CTMP[53]), .S(S[53]), .Co(CTMP[54]) );
  FA_138 FAI_55 ( .A(A[54]), .B(B[54]), .Ci(CTMP[54]), .S(S[54]), .Co(CTMP[55]) );
  FA_137 FAI_56 ( .A(A[55]), .B(B[55]), .Ci(CTMP[55]), .S(S[55]), .Co(CTMP[56]) );
  FA_136 FAI_57 ( .A(A[56]), .B(B[56]), .Ci(CTMP[56]), .S(S[56]), .Co(CTMP[57]) );
  FA_135 FAI_58 ( .A(A[57]), .B(B[57]), .Ci(CTMP[57]), .S(S[57]), .Co(CTMP[58]) );
  FA_134 FAI_59 ( .A(A[58]), .B(B[58]), .Ci(CTMP[58]), .S(S[58]), .Co(CTMP[59]) );
  FA_133 FAI_60 ( .A(A[59]), .B(B[59]), .Ci(CTMP[59]), .S(S[59]), .Co(CTMP[60]) );
  FA_132 FAI_61 ( .A(A[60]), .B(B[60]), .Ci(CTMP[60]), .S(S[60]), .Co(CTMP[61]) );
  FA_131 FAI_62 ( .A(A[61]), .B(B[61]), .Ci(CTMP[61]), .S(S[61]), .Co(CTMP[62]) );
  FA_130 FAI_63 ( .A(A[62]), .B(B[62]), .Ci(CTMP[62]), .S(S[62]), .Co(CTMP[63]) );
  FA_129 FAI_64 ( .A(A[63]), .B(B[63]), .Ci(CTMP[63]), .S(S[63]), .Co(Co) );
endmodule


module booth_mul_row_N64_RADIX3_3 ( prevA, prevSum, encoderIn, nextA, nextSum
 );
  input [63:0] prevA;
  input [63:0] prevSum;
  input [2:0] encoderIn;
  output [63:0] nextA;
  output [63:0] nextSum;

  wire   [2:0] encoder_to_mux;
  wire   [63:0] plus2A_s;
  wire   [63:0] minus2A_s;
  wire   [63:0] minus4A_s;
  tri   [63:0] mux_to_adder;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign nextA[0] = 1'b0;

  encoder_N64_RADIX3_3 encoder_1 ( .X(encoderIn), .Z(encoder_to_mux) );
  ShiftnCompl_N64_3 ShiftnCompl_1 ( .plusA(prevA), .plus2A_out({plus2A_s[63:1], 
        SYNOPSYS_UNCONNECTED__0}), .minus2A_out(minus2A_s), .plus4A_out({
        nextA[63:1], SYNOPSYS_UNCONNECTED__1}), .minus4A_out(minus4A_s) );
  MUX_GENERIC_N64_RADIX3_3 mux_1 ( .plusA({plus2A_s[63:1], 1'b0}), .minusA(
        minus2A_s), .plus2A({nextA[63:1], 1'b0}), .minus2A(minus4A_s), .SEL(
        encoder_to_mux), .Y(mux_to_adder) );
  RCA_N64_3 rca_1 ( .A(mux_to_adder), .B(prevSum), .Ci(1'b0), .S(nextSum) );
endmodule


module encoder_N64_RADIX3_2 ( X, Z );
  input [2:0] X;
  output [2:0] Z;
  wire   n5, n7, n8;

  OAI22_X1 U1 ( .A1(n8), .A2(n5), .B1(X[2]), .B2(n7), .ZN(Z[1]) );
  INV_X1 U2 ( .A(X[2]), .ZN(n5) );
  AOI21_X1 U3 ( .B1(n8), .B2(n7), .A(X[2]), .ZN(Z[0]) );
  OAI21_X1 U4 ( .B1(X[1]), .B2(X[0]), .A(n7), .ZN(n8) );
  AND3_X1 U5 ( .A1(X[2]), .A2(n7), .A3(n8), .ZN(Z[2]) );
  NAND2_X1 U6 ( .A1(X[1]), .A2(X[0]), .ZN(n7) );
endmodule


module shifter_N64_4 ( \input , shiftLeftOnePos );
  input [63:0] \input ;
  output [63:0] shiftLeftOnePos;
  wire   \input[62] , \input[61] , \input[60] , \input[59] , \input[58] ,
         \input[57] , \input[56] , \input[55] , \input[54] , \input[53] ,
         \input[52] , \input[51] , \input[50] , \input[49] , \input[48] ,
         \input[47] , \input[46] , \input[45] , \input[44] , \input[43] ,
         \input[42] , \input[41] , \input[40] , \input[39] , \input[38] ,
         \input[37] , \input[36] , \input[35] , \input[34] , \input[33] ,
         \input[32] , \input[31] , \input[30] , \input[29] , \input[28] ,
         \input[27] , \input[26] , \input[25] , \input[24] , \input[23] ,
         \input[22] , \input[21] , \input[20] , \input[19] , \input[18] ,
         \input[17] , \input[16] , \input[15] , \input[14] , \input[13] ,
         \input[12] , \input[11] , \input[10] , \input[9] , \input[8] ,
         \input[7] , \input[6] , \input[5] , \input[4] , \input[3] ,
         \input[2] , \input[1] , \input[0] ;
  assign shiftLeftOnePos[0] = 1'b0;
  assign shiftLeftOnePos[63] = \input[62] ;
  assign \input[62]  = \input  [62];
  assign shiftLeftOnePos[62] = \input[61] ;
  assign \input[61]  = \input  [61];
  assign shiftLeftOnePos[61] = \input[60] ;
  assign \input[60]  = \input  [60];
  assign shiftLeftOnePos[60] = \input[59] ;
  assign \input[59]  = \input  [59];
  assign shiftLeftOnePos[59] = \input[58] ;
  assign \input[58]  = \input  [58];
  assign shiftLeftOnePos[58] = \input[57] ;
  assign \input[57]  = \input  [57];
  assign shiftLeftOnePos[57] = \input[56] ;
  assign \input[56]  = \input  [56];
  assign shiftLeftOnePos[56] = \input[55] ;
  assign \input[55]  = \input  [55];
  assign shiftLeftOnePos[55] = \input[54] ;
  assign \input[54]  = \input  [54];
  assign shiftLeftOnePos[54] = \input[53] ;
  assign \input[53]  = \input  [53];
  assign shiftLeftOnePos[53] = \input[52] ;
  assign \input[52]  = \input  [52];
  assign shiftLeftOnePos[52] = \input[51] ;
  assign \input[51]  = \input  [51];
  assign shiftLeftOnePos[51] = \input[50] ;
  assign \input[50]  = \input  [50];
  assign shiftLeftOnePos[50] = \input[49] ;
  assign \input[49]  = \input  [49];
  assign shiftLeftOnePos[49] = \input[48] ;
  assign \input[48]  = \input  [48];
  assign shiftLeftOnePos[48] = \input[47] ;
  assign \input[47]  = \input  [47];
  assign shiftLeftOnePos[47] = \input[46] ;
  assign \input[46]  = \input  [46];
  assign shiftLeftOnePos[46] = \input[45] ;
  assign \input[45]  = \input  [45];
  assign shiftLeftOnePos[45] = \input[44] ;
  assign \input[44]  = \input  [44];
  assign shiftLeftOnePos[44] = \input[43] ;
  assign \input[43]  = \input  [43];
  assign shiftLeftOnePos[43] = \input[42] ;
  assign \input[42]  = \input  [42];
  assign shiftLeftOnePos[42] = \input[41] ;
  assign \input[41]  = \input  [41];
  assign shiftLeftOnePos[41] = \input[40] ;
  assign \input[40]  = \input  [40];
  assign shiftLeftOnePos[40] = \input[39] ;
  assign \input[39]  = \input  [39];
  assign shiftLeftOnePos[39] = \input[38] ;
  assign \input[38]  = \input  [38];
  assign shiftLeftOnePos[38] = \input[37] ;
  assign \input[37]  = \input  [37];
  assign shiftLeftOnePos[37] = \input[36] ;
  assign \input[36]  = \input  [36];
  assign shiftLeftOnePos[36] = \input[35] ;
  assign \input[35]  = \input  [35];
  assign shiftLeftOnePos[35] = \input[34] ;
  assign \input[34]  = \input  [34];
  assign shiftLeftOnePos[34] = \input[33] ;
  assign \input[33]  = \input  [33];
  assign shiftLeftOnePos[33] = \input[32] ;
  assign \input[32]  = \input  [32];
  assign shiftLeftOnePos[32] = \input[31] ;
  assign \input[31]  = \input  [31];
  assign shiftLeftOnePos[31] = \input[30] ;
  assign \input[30]  = \input  [30];
  assign shiftLeftOnePos[30] = \input[29] ;
  assign \input[29]  = \input  [29];
  assign shiftLeftOnePos[29] = \input[28] ;
  assign \input[28]  = \input  [28];
  assign shiftLeftOnePos[28] = \input[27] ;
  assign \input[27]  = \input  [27];
  assign shiftLeftOnePos[27] = \input[26] ;
  assign \input[26]  = \input  [26];
  assign shiftLeftOnePos[26] = \input[25] ;
  assign \input[25]  = \input  [25];
  assign shiftLeftOnePos[25] = \input[24] ;
  assign \input[24]  = \input  [24];
  assign shiftLeftOnePos[24] = \input[23] ;
  assign \input[23]  = \input  [23];
  assign shiftLeftOnePos[23] = \input[22] ;
  assign \input[22]  = \input  [22];
  assign shiftLeftOnePos[22] = \input[21] ;
  assign \input[21]  = \input  [21];
  assign shiftLeftOnePos[21] = \input[20] ;
  assign \input[20]  = \input  [20];
  assign shiftLeftOnePos[20] = \input[19] ;
  assign \input[19]  = \input  [19];
  assign shiftLeftOnePos[19] = \input[18] ;
  assign \input[18]  = \input  [18];
  assign shiftLeftOnePos[18] = \input[17] ;
  assign \input[17]  = \input  [17];
  assign shiftLeftOnePos[17] = \input[16] ;
  assign \input[16]  = \input  [16];
  assign shiftLeftOnePos[16] = \input[15] ;
  assign \input[15]  = \input  [15];
  assign shiftLeftOnePos[15] = \input[14] ;
  assign \input[14]  = \input  [14];
  assign shiftLeftOnePos[14] = \input[13] ;
  assign \input[13]  = \input  [13];
  assign shiftLeftOnePos[13] = \input[12] ;
  assign \input[12]  = \input  [12];
  assign shiftLeftOnePos[12] = \input[11] ;
  assign \input[11]  = \input  [11];
  assign shiftLeftOnePos[11] = \input[10] ;
  assign \input[10]  = \input  [10];
  assign shiftLeftOnePos[10] = \input[9] ;
  assign \input[9]  = \input  [9];
  assign shiftLeftOnePos[9] = \input[8] ;
  assign \input[8]  = \input  [8];
  assign shiftLeftOnePos[8] = \input[7] ;
  assign \input[7]  = \input  [7];
  assign shiftLeftOnePos[7] = \input[6] ;
  assign \input[6]  = \input  [6];
  assign shiftLeftOnePos[6] = \input[5] ;
  assign \input[5]  = \input  [5];
  assign shiftLeftOnePos[5] = \input[4] ;
  assign \input[4]  = \input  [4];
  assign shiftLeftOnePos[4] = \input[3] ;
  assign \input[3]  = \input  [3];
  assign shiftLeftOnePos[3] = \input[2] ;
  assign \input[2]  = \input  [2];
  assign shiftLeftOnePos[2] = \input[1] ;
  assign \input[1]  = \input  [1];
  assign shiftLeftOnePos[1] = \input[0] ;
  assign \input[0]  = \input  [0];

endmodule


module shifter_N64_3 ( \input , shiftLeftOnePos );
  input [63:0] \input ;
  output [63:0] shiftLeftOnePos;
  wire   \input[62] , \input[61] , \input[60] , \input[59] , \input[58] ,
         \input[57] , \input[56] , \input[55] , \input[54] , \input[53] ,
         \input[52] , \input[51] , \input[50] , \input[49] , \input[48] ,
         \input[47] , \input[46] , \input[45] , \input[44] , \input[43] ,
         \input[42] , \input[41] , \input[40] , \input[39] , \input[38] ,
         \input[37] , \input[36] , \input[35] , \input[34] , \input[33] ,
         \input[32] , \input[31] , \input[30] , \input[29] , \input[28] ,
         \input[27] , \input[26] , \input[25] , \input[24] , \input[23] ,
         \input[22] , \input[21] , \input[20] , \input[19] , \input[18] ,
         \input[17] , \input[16] , \input[15] , \input[14] , \input[13] ,
         \input[12] , \input[11] , \input[10] , \input[9] , \input[8] ,
         \input[7] , \input[6] , \input[5] , \input[4] , \input[3] ,
         \input[2] , \input[1] , \input[0] ;
  assign shiftLeftOnePos[0] = 1'b0;
  assign shiftLeftOnePos[63] = \input[62] ;
  assign \input[62]  = \input  [62];
  assign shiftLeftOnePos[62] = \input[61] ;
  assign \input[61]  = \input  [61];
  assign shiftLeftOnePos[61] = \input[60] ;
  assign \input[60]  = \input  [60];
  assign shiftLeftOnePos[60] = \input[59] ;
  assign \input[59]  = \input  [59];
  assign shiftLeftOnePos[59] = \input[58] ;
  assign \input[58]  = \input  [58];
  assign shiftLeftOnePos[58] = \input[57] ;
  assign \input[57]  = \input  [57];
  assign shiftLeftOnePos[57] = \input[56] ;
  assign \input[56]  = \input  [56];
  assign shiftLeftOnePos[56] = \input[55] ;
  assign \input[55]  = \input  [55];
  assign shiftLeftOnePos[55] = \input[54] ;
  assign \input[54]  = \input  [54];
  assign shiftLeftOnePos[54] = \input[53] ;
  assign \input[53]  = \input  [53];
  assign shiftLeftOnePos[53] = \input[52] ;
  assign \input[52]  = \input  [52];
  assign shiftLeftOnePos[52] = \input[51] ;
  assign \input[51]  = \input  [51];
  assign shiftLeftOnePos[51] = \input[50] ;
  assign \input[50]  = \input  [50];
  assign shiftLeftOnePos[50] = \input[49] ;
  assign \input[49]  = \input  [49];
  assign shiftLeftOnePos[49] = \input[48] ;
  assign \input[48]  = \input  [48];
  assign shiftLeftOnePos[48] = \input[47] ;
  assign \input[47]  = \input  [47];
  assign shiftLeftOnePos[47] = \input[46] ;
  assign \input[46]  = \input  [46];
  assign shiftLeftOnePos[46] = \input[45] ;
  assign \input[45]  = \input  [45];
  assign shiftLeftOnePos[45] = \input[44] ;
  assign \input[44]  = \input  [44];
  assign shiftLeftOnePos[44] = \input[43] ;
  assign \input[43]  = \input  [43];
  assign shiftLeftOnePos[43] = \input[42] ;
  assign \input[42]  = \input  [42];
  assign shiftLeftOnePos[42] = \input[41] ;
  assign \input[41]  = \input  [41];
  assign shiftLeftOnePos[41] = \input[40] ;
  assign \input[40]  = \input  [40];
  assign shiftLeftOnePos[40] = \input[39] ;
  assign \input[39]  = \input  [39];
  assign shiftLeftOnePos[39] = \input[38] ;
  assign \input[38]  = \input  [38];
  assign shiftLeftOnePos[38] = \input[37] ;
  assign \input[37]  = \input  [37];
  assign shiftLeftOnePos[37] = \input[36] ;
  assign \input[36]  = \input  [36];
  assign shiftLeftOnePos[36] = \input[35] ;
  assign \input[35]  = \input  [35];
  assign shiftLeftOnePos[35] = \input[34] ;
  assign \input[34]  = \input  [34];
  assign shiftLeftOnePos[34] = \input[33] ;
  assign \input[33]  = \input  [33];
  assign shiftLeftOnePos[33] = \input[32] ;
  assign \input[32]  = \input  [32];
  assign shiftLeftOnePos[32] = \input[31] ;
  assign \input[31]  = \input  [31];
  assign shiftLeftOnePos[31] = \input[30] ;
  assign \input[30]  = \input  [30];
  assign shiftLeftOnePos[30] = \input[29] ;
  assign \input[29]  = \input  [29];
  assign shiftLeftOnePos[29] = \input[28] ;
  assign \input[28]  = \input  [28];
  assign shiftLeftOnePos[28] = \input[27] ;
  assign \input[27]  = \input  [27];
  assign shiftLeftOnePos[27] = \input[26] ;
  assign \input[26]  = \input  [26];
  assign shiftLeftOnePos[26] = \input[25] ;
  assign \input[25]  = \input  [25];
  assign shiftLeftOnePos[25] = \input[24] ;
  assign \input[24]  = \input  [24];
  assign shiftLeftOnePos[24] = \input[23] ;
  assign \input[23]  = \input  [23];
  assign shiftLeftOnePos[23] = \input[22] ;
  assign \input[22]  = \input  [22];
  assign shiftLeftOnePos[22] = \input[21] ;
  assign \input[21]  = \input  [21];
  assign shiftLeftOnePos[21] = \input[20] ;
  assign \input[20]  = \input  [20];
  assign shiftLeftOnePos[20] = \input[19] ;
  assign \input[19]  = \input  [19];
  assign shiftLeftOnePos[19] = \input[18] ;
  assign \input[18]  = \input  [18];
  assign shiftLeftOnePos[18] = \input[17] ;
  assign \input[17]  = \input  [17];
  assign shiftLeftOnePos[17] = \input[16] ;
  assign \input[16]  = \input  [16];
  assign shiftLeftOnePos[16] = \input[15] ;
  assign \input[15]  = \input  [15];
  assign shiftLeftOnePos[15] = \input[14] ;
  assign \input[14]  = \input  [14];
  assign shiftLeftOnePos[14] = \input[13] ;
  assign \input[13]  = \input  [13];
  assign shiftLeftOnePos[13] = \input[12] ;
  assign \input[12]  = \input  [12];
  assign shiftLeftOnePos[12] = \input[11] ;
  assign \input[11]  = \input  [11];
  assign shiftLeftOnePos[11] = \input[10] ;
  assign \input[10]  = \input  [10];
  assign shiftLeftOnePos[10] = \input[9] ;
  assign \input[9]  = \input  [9];
  assign shiftLeftOnePos[9] = \input[8] ;
  assign \input[8]  = \input  [8];
  assign shiftLeftOnePos[8] = \input[7] ;
  assign \input[7]  = \input  [7];
  assign shiftLeftOnePos[7] = \input[6] ;
  assign \input[6]  = \input  [6];
  assign shiftLeftOnePos[6] = \input[5] ;
  assign \input[5]  = \input  [5];
  assign shiftLeftOnePos[5] = \input[4] ;
  assign \input[4]  = \input  [4];
  assign shiftLeftOnePos[4] = \input[3] ;
  assign \input[3]  = \input  [3];
  assign shiftLeftOnePos[3] = \input[2] ;
  assign \input[2]  = \input  [2];
  assign shiftLeftOnePos[2] = \input[1] ;
  assign \input[1]  = \input  [1];
  assign shiftLeftOnePos[1] = \input[0] ;
  assign \input[0]  = \input  [0];

endmodule


module complementer_N64_4_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n190, n191, n192, n193, n194, n196, n197, n198, n199, n200,
         n202, n203, n204, n206, n207, n208, n210, n211, n212, n213, n214,
         n216, n217, n218, n220, n221, n222, n224, n225, n226, n228, n229,
         n230, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n189,
         n195, n201, n205, n209, n215, n219, n223, n227, n231;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U81 ( .A(n190), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U82 ( .A(n192), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U83 ( .A(n193), .B(B[6]), .Z(DIFF[6]) );
  XOR2_X1 U85 ( .A(n196), .B(B[62]), .Z(DIFF[62]) );
  XOR2_X1 U86 ( .A(n194), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U87 ( .A(n198), .B(B[59]), .Z(DIFF[59]) );
  XOR2_X1 U89 ( .A(n200), .B(B[57]), .Z(DIFF[57]) );
  XOR2_X1 U90 ( .A(n202), .B(B[55]), .Z(DIFF[55]) );
  XOR2_X1 U92 ( .A(n204), .B(B[53]), .Z(DIFF[53]) );
  XOR2_X1 U93 ( .A(n206), .B(B[51]), .Z(DIFF[51]) );
  XOR2_X1 U95 ( .A(n208), .B(B[49]), .Z(DIFF[49]) );
  XOR2_X1 U96 ( .A(n212), .B(B[47]), .Z(DIFF[47]) );
  XOR2_X1 U98 ( .A(n214), .B(B[45]), .Z(DIFF[45]) );
  XOR2_X1 U99 ( .A(n216), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U101 ( .A(n218), .B(B[41]), .Z(DIFF[41]) );
  XOR2_X1 U102 ( .A(n211), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U103 ( .A(n220), .B(B[39]), .Z(DIFF[39]) );
  XOR2_X1 U105 ( .A(n222), .B(B[37]), .Z(DIFF[37]) );
  XOR2_X1 U106 ( .A(n224), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U108 ( .A(n226), .B(B[33]), .Z(DIFF[33]) );
  XOR2_X1 U109 ( .A(n228), .B(B[31]), .Z(DIFF[31]) );
  XOR2_X1 U111 ( .A(n230), .B(B[29]), .Z(DIFF[29]) );
  XOR2_X1 U112 ( .A(n233), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U113 ( .A(n236), .B(B[26]), .Z(DIFF[26]) );
  XOR2_X1 U114 ( .A(n235), .B(B[25]), .Z(DIFF[25]) );
  XOR2_X1 U115 ( .A(n237), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U116 ( .A(n240), .B(B[22]), .Z(DIFF[22]) );
  XOR2_X1 U117 ( .A(n239), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U118 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U119 ( .A(n241), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U120 ( .A(n244), .B(B[18]), .Z(DIFF[18]) );
  XOR2_X1 U121 ( .A(n243), .B(B[17]), .Z(DIFF[17]) );
  XOR2_X1 U122 ( .A(n245), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U123 ( .A(n248), .B(B[14]), .Z(DIFF[14]) );
  XOR2_X1 U124 ( .A(n247), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U125 ( .A(n249), .B(B[11]), .Z(DIFF[11]) );
  XOR2_X1 U126 ( .A(n251), .B(B[10]), .Z(DIFF[10]) );
  XOR2_X1 U1 ( .A(n197), .B(n231), .Z(DIFF[61]) );
  NAND2_X1 U2 ( .A1(n197), .A2(n231), .ZN(n196) );
  NOR3_X1 U3 ( .A1(B[59]), .A2(B[60]), .A3(n198), .ZN(n197) );
  XNOR2_X1 U4 ( .A(n189), .B(B[63]), .ZN(DIFF[63]) );
  NOR2_X1 U5 ( .A1(n196), .A2(B[62]), .ZN(n189) );
  XNOR2_X1 U6 ( .A(B[60]), .B(n199), .ZN(DIFF[60]) );
  NOR2_X1 U7 ( .A1(B[59]), .A2(n198), .ZN(n199) );
  XNOR2_X1 U8 ( .A(B[48]), .B(n213), .ZN(DIFF[48]) );
  NOR2_X1 U9 ( .A1(B[47]), .A2(n212), .ZN(n213) );
  XNOR2_X1 U10 ( .A(B[44]), .B(n217), .ZN(DIFF[44]) );
  NOR2_X1 U11 ( .A1(B[43]), .A2(n216), .ZN(n217) );
  XNOR2_X1 U12 ( .A(B[40]), .B(n221), .ZN(DIFF[40]) );
  NOR2_X1 U13 ( .A1(B[39]), .A2(n220), .ZN(n221) );
  OR3_X1 U14 ( .A1(B[41]), .A2(B[42]), .A3(n218), .ZN(n216) );
  OR3_X1 U15 ( .A1(B[45]), .A2(B[46]), .A3(n214), .ZN(n212) );
  OR3_X1 U16 ( .A1(B[39]), .A2(B[40]), .A3(n220), .ZN(n218) );
  OR3_X1 U17 ( .A1(B[43]), .A2(B[44]), .A3(n216), .ZN(n214) );
  XNOR2_X1 U18 ( .A(n195), .B(B[46]), .ZN(DIFF[46]) );
  NOR2_X1 U19 ( .A1(n214), .A2(B[45]), .ZN(n195) );
  XNOR2_X1 U20 ( .A(n201), .B(B[42]), .ZN(DIFF[42]) );
  NOR2_X1 U21 ( .A1(n218), .A2(B[41]), .ZN(n201) );
  XNOR2_X1 U22 ( .A(B[56]), .B(n203), .ZN(DIFF[56]) );
  NOR2_X1 U23 ( .A1(B[55]), .A2(n202), .ZN(n203) );
  XNOR2_X1 U24 ( .A(B[52]), .B(n207), .ZN(DIFF[52]) );
  NOR2_X1 U25 ( .A1(B[51]), .A2(n206), .ZN(n207) );
  OR3_X1 U26 ( .A1(B[57]), .A2(B[58]), .A3(n200), .ZN(n198) );
  OR3_X1 U27 ( .A1(B[49]), .A2(B[50]), .A3(n208), .ZN(n206) );
  OR3_X1 U28 ( .A1(B[53]), .A2(B[54]), .A3(n204), .ZN(n202) );
  OR3_X1 U29 ( .A1(B[47]), .A2(B[48]), .A3(n212), .ZN(n208) );
  OR3_X1 U30 ( .A1(B[51]), .A2(B[52]), .A3(n206), .ZN(n204) );
  OR3_X1 U31 ( .A1(B[55]), .A2(B[56]), .A3(n202), .ZN(n200) );
  XNOR2_X1 U32 ( .A(n205), .B(B[58]), .ZN(DIFF[58]) );
  NOR2_X1 U33 ( .A1(n200), .A2(B[57]), .ZN(n205) );
  XNOR2_X1 U34 ( .A(n209), .B(B[54]), .ZN(DIFF[54]) );
  NOR2_X1 U35 ( .A1(n204), .A2(B[53]), .ZN(n209) );
  XNOR2_X1 U36 ( .A(n215), .B(B[50]), .ZN(DIFF[50]) );
  NOR2_X1 U37 ( .A1(n208), .A2(B[49]), .ZN(n215) );
  OR3_X1 U38 ( .A1(B[37]), .A2(B[38]), .A3(n222), .ZN(n220) );
  XNOR2_X1 U39 ( .A(n219), .B(B[38]), .ZN(DIFF[38]) );
  NOR2_X1 U40 ( .A1(n222), .A2(B[37]), .ZN(n219) );
  XNOR2_X1 U41 ( .A(B[36]), .B(n225), .ZN(DIFF[36]) );
  NOR2_X1 U42 ( .A1(B[35]), .A2(n224), .ZN(n225) );
  OR3_X1 U43 ( .A1(B[35]), .A2(B[36]), .A3(n224), .ZN(n222) );
  OR3_X1 U44 ( .A1(B[33]), .A2(B[34]), .A3(n226), .ZN(n224) );
  XNOR2_X1 U45 ( .A(n223), .B(B[34]), .ZN(DIFF[34]) );
  NOR2_X1 U46 ( .A1(n226), .A2(B[33]), .ZN(n223) );
  XNOR2_X1 U47 ( .A(B[32]), .B(n229), .ZN(DIFF[32]) );
  NOR2_X1 U48 ( .A1(B[31]), .A2(n228), .ZN(n229) );
  OR3_X1 U49 ( .A1(B[31]), .A2(B[32]), .A3(n228), .ZN(n226) );
  OR3_X1 U50 ( .A1(B[29]), .A2(B[30]), .A3(n230), .ZN(n228) );
  XNOR2_X1 U51 ( .A(n227), .B(B[30]), .ZN(DIFF[30]) );
  NOR2_X1 U52 ( .A1(n230), .A2(B[29]), .ZN(n227) );
  OR3_X1 U53 ( .A1(B[27]), .A2(B[28]), .A3(n233), .ZN(n230) );
  XNOR2_X1 U54 ( .A(B[28]), .B(n234), .ZN(DIFF[28]) );
  NOR2_X1 U55 ( .A1(B[27]), .A2(n233), .ZN(n234) );
  NOR2_X1 U56 ( .A1(B[23]), .A2(n237), .ZN(n238) );
  NOR2_X1 U57 ( .A1(B[19]), .A2(n241), .ZN(n242) );
  NOR2_X1 U58 ( .A1(B[15]), .A2(n245), .ZN(n246) );
  NOR2_X1 U59 ( .A1(B[11]), .A2(n249), .ZN(n250) );
  NOR2_X1 U60 ( .A1(B[7]), .A2(n192), .ZN(n191) );
  NOR2_X1 U61 ( .A1(B[3]), .A2(n211), .ZN(n210) );
  OR3_X1 U62 ( .A1(B[25]), .A2(B[26]), .A3(n235), .ZN(n233) );
  OR3_X1 U63 ( .A1(B[21]), .A2(B[22]), .A3(n239), .ZN(n237) );
  OR3_X1 U64 ( .A1(B[17]), .A2(B[18]), .A3(n243), .ZN(n241) );
  OR3_X1 U65 ( .A1(B[13]), .A2(B[14]), .A3(n247), .ZN(n245) );
  OR3_X1 U66 ( .A1(B[10]), .A2(B[9]), .A3(n190), .ZN(n249) );
  OR3_X1 U67 ( .A1(B[5]), .A2(B[6]), .A3(n194), .ZN(n192) );
  OR3_X1 U68 ( .A1(B[23]), .A2(B[24]), .A3(n237), .ZN(n235) );
  OR3_X1 U69 ( .A1(B[19]), .A2(B[20]), .A3(n241), .ZN(n239) );
  OR3_X1 U70 ( .A1(B[15]), .A2(B[16]), .A3(n245), .ZN(n243) );
  OR3_X1 U71 ( .A1(B[11]), .A2(B[12]), .A3(n249), .ZN(n247) );
  OR3_X1 U72 ( .A1(B[7]), .A2(B[8]), .A3(n192), .ZN(n190) );
  OR3_X1 U73 ( .A1(B[3]), .A2(B[4]), .A3(n211), .ZN(n194) );
  XNOR2_X1 U74 ( .A(B[24]), .B(n238), .ZN(DIFF[24]) );
  XNOR2_X1 U75 ( .A(B[20]), .B(n242), .ZN(DIFF[20]) );
  XNOR2_X1 U76 ( .A(B[16]), .B(n246), .ZN(DIFF[16]) );
  XNOR2_X1 U77 ( .A(B[12]), .B(n250), .ZN(DIFF[12]) );
  XNOR2_X1 U78 ( .A(B[8]), .B(n191), .ZN(DIFF[8]) );
  XNOR2_X1 U79 ( .A(B[4]), .B(n210), .ZN(DIFF[4]) );
  XNOR2_X1 U80 ( .A(B[2]), .B(n232), .ZN(DIFF[2]) );
  OR2_X1 U84 ( .A1(n235), .A2(B[25]), .ZN(n236) );
  OR2_X1 U88 ( .A1(n239), .A2(B[21]), .ZN(n240) );
  OR2_X1 U91 ( .A1(n243), .A2(B[17]), .ZN(n244) );
  OR2_X1 U94 ( .A1(n247), .A2(B[13]), .ZN(n248) );
  OR2_X1 U97 ( .A1(n190), .A2(B[9]), .ZN(n251) );
  OR2_X1 U100 ( .A1(n194), .A2(B[5]), .ZN(n193) );
  OR3_X1 U104 ( .A1(B[1]), .A2(B[2]), .A3(\B[0] ), .ZN(n211) );
  NOR2_X1 U107 ( .A1(\B[0] ), .A2(B[1]), .ZN(n232) );
  INV_X1 U110 ( .A(B[61]), .ZN(n231) );
endmodule


module complementer_N64_4 ( \input , complement2 );
  input [63:0] \input ;
  output [63:0] complement2;


  complementer_N64_4_DW01_sub_0 sub_add_31_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(\input ), .CI(1'b0), .DIFF(complement2) );
endmodule


module complementer_N64_3_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n190, n191, n192, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n237, n238, n239, n241, n242, n243, n245, n246, n247,
         n249, n250, n189, n193, n236, n240, n244, n248, n251;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U81 ( .A(n190), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U82 ( .A(n192), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U84 ( .A(n195), .B(B[63]), .Z(DIFF[63]) );
  XOR2_X1 U85 ( .A(n196), .B(B[62]), .Z(DIFF[62]) );
  XOR2_X1 U86 ( .A(n194), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U87 ( .A(n198), .B(B[59]), .Z(DIFF[59]) );
  XOR2_X1 U88 ( .A(n201), .B(B[58]), .Z(DIFF[58]) );
  XOR2_X1 U89 ( .A(n200), .B(B[57]), .Z(DIFF[57]) );
  XOR2_X1 U90 ( .A(n202), .B(B[55]), .Z(DIFF[55]) );
  XOR2_X1 U91 ( .A(n205), .B(B[54]), .Z(DIFF[54]) );
  XOR2_X1 U92 ( .A(n204), .B(B[53]), .Z(DIFF[53]) );
  XOR2_X1 U93 ( .A(n206), .B(B[51]), .Z(DIFF[51]) );
  XOR2_X1 U94 ( .A(n209), .B(B[50]), .Z(DIFF[50]) );
  XOR2_X1 U95 ( .A(n208), .B(B[49]), .Z(DIFF[49]) );
  XOR2_X1 U96 ( .A(n212), .B(B[47]), .Z(DIFF[47]) );
  XOR2_X1 U97 ( .A(n215), .B(B[46]), .Z(DIFF[46]) );
  XOR2_X1 U98 ( .A(n214), .B(B[45]), .Z(DIFF[45]) );
  XOR2_X1 U99 ( .A(n216), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U100 ( .A(n219), .B(B[42]), .Z(DIFF[42]) );
  XOR2_X1 U101 ( .A(n218), .B(B[41]), .Z(DIFF[41]) );
  XOR2_X1 U102 ( .A(n211), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U103 ( .A(n220), .B(B[39]), .Z(DIFF[39]) );
  XOR2_X1 U104 ( .A(n223), .B(B[38]), .Z(DIFF[38]) );
  XOR2_X1 U105 ( .A(n222), .B(B[37]), .Z(DIFF[37]) );
  XOR2_X1 U106 ( .A(n224), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U107 ( .A(n227), .B(B[34]), .Z(DIFF[34]) );
  XOR2_X1 U108 ( .A(n226), .B(B[33]), .Z(DIFF[33]) );
  XOR2_X1 U109 ( .A(n228), .B(B[31]), .Z(DIFF[31]) );
  XOR2_X1 U110 ( .A(n231), .B(B[30]), .Z(DIFF[30]) );
  XOR2_X1 U111 ( .A(n230), .B(B[29]), .Z(DIFF[29]) );
  XOR2_X1 U112 ( .A(n233), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U114 ( .A(n235), .B(B[25]), .Z(DIFF[25]) );
  XOR2_X1 U115 ( .A(n237), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U117 ( .A(n239), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U118 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U119 ( .A(n241), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U121 ( .A(n243), .B(B[17]), .Z(DIFF[17]) );
  XOR2_X1 U122 ( .A(n245), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U124 ( .A(n247), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U125 ( .A(n249), .B(B[11]), .Z(DIFF[11]) );
  OR2_X1 U1 ( .A1(n196), .A2(B[62]), .ZN(n195) );
  NAND2_X1 U2 ( .A1(n197), .A2(n251), .ZN(n196) );
  NOR2_X1 U3 ( .A1(B[43]), .A2(n216), .ZN(n217) );
  NOR2_X1 U4 ( .A1(B[39]), .A2(n220), .ZN(n221) );
  OR3_X1 U5 ( .A1(B[41]), .A2(B[42]), .A3(n218), .ZN(n216) );
  OR3_X1 U6 ( .A1(B[43]), .A2(B[44]), .A3(n216), .ZN(n214) );
  OR3_X1 U7 ( .A1(B[39]), .A2(B[40]), .A3(n220), .ZN(n218) );
  OR2_X1 U8 ( .A1(n218), .A2(B[41]), .ZN(n219) );
  NOR3_X1 U9 ( .A1(B[59]), .A2(B[60]), .A3(n198), .ZN(n197) );
  NOR2_X1 U10 ( .A1(B[59]), .A2(n198), .ZN(n199) );
  NOR2_X1 U11 ( .A1(B[55]), .A2(n202), .ZN(n203) );
  NOR2_X1 U12 ( .A1(B[51]), .A2(n206), .ZN(n207) );
  NOR2_X1 U13 ( .A1(B[47]), .A2(n212), .ZN(n213) );
  OR3_X1 U14 ( .A1(B[57]), .A2(B[58]), .A3(n200), .ZN(n198) );
  OR3_X1 U15 ( .A1(B[53]), .A2(B[54]), .A3(n204), .ZN(n202) );
  OR3_X1 U16 ( .A1(B[49]), .A2(B[50]), .A3(n208), .ZN(n206) );
  OR3_X1 U17 ( .A1(B[45]), .A2(B[46]), .A3(n214), .ZN(n212) );
  OR3_X1 U18 ( .A1(B[55]), .A2(B[56]), .A3(n202), .ZN(n200) );
  OR3_X1 U19 ( .A1(B[51]), .A2(B[52]), .A3(n206), .ZN(n204) );
  OR3_X1 U20 ( .A1(B[47]), .A2(B[48]), .A3(n212), .ZN(n208) );
  OR2_X1 U21 ( .A1(n204), .A2(B[53]), .ZN(n205) );
  OR2_X1 U22 ( .A1(n208), .A2(B[49]), .ZN(n209) );
  OR2_X1 U23 ( .A1(n214), .A2(B[45]), .ZN(n215) );
  OR2_X1 U24 ( .A1(n200), .A2(B[57]), .ZN(n201) );
  OR3_X1 U25 ( .A1(B[37]), .A2(B[38]), .A3(n222), .ZN(n220) );
  OR2_X1 U26 ( .A1(n222), .A2(B[37]), .ZN(n223) );
  NOR2_X1 U27 ( .A1(B[35]), .A2(n224), .ZN(n225) );
  OR3_X1 U28 ( .A1(B[35]), .A2(B[36]), .A3(n224), .ZN(n222) );
  OR3_X1 U29 ( .A1(B[33]), .A2(B[34]), .A3(n226), .ZN(n224) );
  XNOR2_X1 U30 ( .A(B[48]), .B(n213), .ZN(DIFF[48]) );
  XNOR2_X1 U31 ( .A(B[44]), .B(n217), .ZN(DIFF[44]) );
  XNOR2_X1 U32 ( .A(B[40]), .B(n221), .ZN(DIFF[40]) );
  XNOR2_X1 U33 ( .A(B[36]), .B(n225), .ZN(DIFF[36]) );
  XNOR2_X1 U34 ( .A(B[32]), .B(n229), .ZN(DIFF[32]) );
  OR2_X1 U35 ( .A1(n226), .A2(B[33]), .ZN(n227) );
  XNOR2_X1 U36 ( .A(n197), .B(B[61]), .ZN(DIFF[61]) );
  XNOR2_X1 U37 ( .A(B[60]), .B(n199), .ZN(DIFF[60]) );
  XNOR2_X1 U38 ( .A(B[56]), .B(n203), .ZN(DIFF[56]) );
  XNOR2_X1 U39 ( .A(B[52]), .B(n207), .ZN(DIFF[52]) );
  NOR2_X1 U40 ( .A1(B[31]), .A2(n228), .ZN(n229) );
  OR3_X1 U41 ( .A1(B[31]), .A2(B[32]), .A3(n228), .ZN(n226) );
  OR3_X1 U42 ( .A1(B[29]), .A2(B[30]), .A3(n230), .ZN(n228) );
  OR2_X1 U43 ( .A1(n230), .A2(B[29]), .ZN(n231) );
  XNOR2_X1 U44 ( .A(B[28]), .B(n234), .ZN(DIFF[28]) );
  XNOR2_X1 U45 ( .A(n189), .B(B[18]), .ZN(DIFF[18]) );
  NOR2_X1 U46 ( .A1(n243), .A2(B[17]), .ZN(n189) );
  XNOR2_X1 U47 ( .A(n193), .B(B[26]), .ZN(DIFF[26]) );
  NOR2_X1 U48 ( .A1(n235), .A2(B[25]), .ZN(n193) );
  XNOR2_X1 U49 ( .A(n236), .B(B[22]), .ZN(DIFF[22]) );
  NOR2_X1 U50 ( .A1(n239), .A2(B[21]), .ZN(n236) );
  XNOR2_X1 U51 ( .A(n240), .B(B[14]), .ZN(DIFF[14]) );
  NOR2_X1 U52 ( .A1(n247), .A2(B[13]), .ZN(n240) );
  XNOR2_X1 U53 ( .A(n244), .B(B[10]), .ZN(DIFF[10]) );
  NOR2_X1 U54 ( .A1(n190), .A2(B[9]), .ZN(n244) );
  XNOR2_X1 U55 ( .A(n248), .B(B[6]), .ZN(DIFF[6]) );
  NOR2_X1 U56 ( .A1(n194), .A2(B[5]), .ZN(n248) );
  NOR2_X1 U57 ( .A1(B[27]), .A2(n233), .ZN(n234) );
  XNOR2_X1 U58 ( .A(B[24]), .B(n238), .ZN(DIFF[24]) );
  NOR2_X1 U59 ( .A1(B[23]), .A2(n237), .ZN(n238) );
  XNOR2_X1 U60 ( .A(B[20]), .B(n242), .ZN(DIFF[20]) );
  NOR2_X1 U61 ( .A1(B[19]), .A2(n241), .ZN(n242) );
  XNOR2_X1 U62 ( .A(B[16]), .B(n246), .ZN(DIFF[16]) );
  NOR2_X1 U63 ( .A1(B[15]), .A2(n245), .ZN(n246) );
  XNOR2_X1 U64 ( .A(B[12]), .B(n250), .ZN(DIFF[12]) );
  NOR2_X1 U65 ( .A1(B[11]), .A2(n249), .ZN(n250) );
  XNOR2_X1 U66 ( .A(B[8]), .B(n191), .ZN(DIFF[8]) );
  NOR2_X1 U67 ( .A1(B[7]), .A2(n192), .ZN(n191) );
  XNOR2_X1 U68 ( .A(B[2]), .B(n232), .ZN(DIFF[2]) );
  NOR2_X1 U69 ( .A1(\B[0] ), .A2(B[1]), .ZN(n232) );
  XNOR2_X1 U70 ( .A(B[4]), .B(n210), .ZN(DIFF[4]) );
  NOR2_X1 U71 ( .A1(B[3]), .A2(n211), .ZN(n210) );
  OR3_X1 U72 ( .A1(B[5]), .A2(B[6]), .A3(n194), .ZN(n192) );
  OR3_X1 U73 ( .A1(B[10]), .A2(B[9]), .A3(n190), .ZN(n249) );
  OR3_X1 U74 ( .A1(B[13]), .A2(B[14]), .A3(n247), .ZN(n245) );
  OR3_X1 U75 ( .A1(B[17]), .A2(B[18]), .A3(n243), .ZN(n241) );
  OR3_X1 U76 ( .A1(B[21]), .A2(B[22]), .A3(n239), .ZN(n237) );
  OR3_X1 U77 ( .A1(B[25]), .A2(B[26]), .A3(n235), .ZN(n233) );
  OR3_X1 U78 ( .A1(B[7]), .A2(B[8]), .A3(n192), .ZN(n190) );
  OR3_X1 U79 ( .A1(B[11]), .A2(B[12]), .A3(n249), .ZN(n247) );
  OR3_X1 U80 ( .A1(B[15]), .A2(B[16]), .A3(n245), .ZN(n243) );
  OR3_X1 U83 ( .A1(B[19]), .A2(B[20]), .A3(n241), .ZN(n239) );
  OR3_X1 U113 ( .A1(B[23]), .A2(B[24]), .A3(n237), .ZN(n235) );
  OR3_X1 U116 ( .A1(B[27]), .A2(B[28]), .A3(n233), .ZN(n230) );
  OR3_X1 U120 ( .A1(B[3]), .A2(B[4]), .A3(n211), .ZN(n194) );
  OR3_X1 U123 ( .A1(B[1]), .A2(B[2]), .A3(\B[0] ), .ZN(n211) );
  INV_X1 U126 ( .A(B[61]), .ZN(n251) );
endmodule


module complementer_N64_3 ( \input , complement2 );
  input [63:0] \input ;
  output [63:0] complement2;


  complementer_N64_3_DW01_sub_0 sub_add_31_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(\input ), .CI(1'b0), .DIFF(complement2) );
endmodule


module ShiftnCompl_N64_2 ( plusA, plus2A_out, minus2A_out, plus4A_out, 
        minus4A_out );
  input [63:0] plusA;
  output [63:0] plus2A_out;
  output [63:0] minus2A_out;
  output [63:0] plus4A_out;
  output [63:0] minus4A_out;

  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign plus2A_out[0] = 1'b0;
  assign plus4A_out[0] = 1'b0;

  shifter_N64_4 shifter_1 ( .\input (plusA), .shiftLeftOnePos({
        plus2A_out[63:1], SYNOPSYS_UNCONNECTED__0}) );
  shifter_N64_3 shifter_2 ( .\input ({plus2A_out[63:1], 1'b0}), 
        .shiftLeftOnePos({plus4A_out[63:1], SYNOPSYS_UNCONNECTED__1}) );
  complementer_N64_4 complementer_1 ( .\input ({plus2A_out[63:1], 1'b0}), 
        .complement2(minus2A_out) );
  complementer_N64_3 complementer_2 ( .\input ({plus4A_out[63:1], 1'b0}), 
        .complement2(minus4A_out) );
endmodule


module MUX_GENERIC_N64_RADIX3_2 ( plusA, minusA, plus2A, minus2A, SEL, Y );
  input [63:0] plusA;
  input [63:0] minusA;
  input [63:0] plus2A;
  input [63:0] minus2A;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502;
  tri   [63:0] Y;

  TBUF_X1 \Y_tri[55]  ( .A(n446), .EN(n301), .Z(Y[55]) );
  TBUF_X1 \Y_tri[56]  ( .A(n445), .EN(n301), .Z(Y[56]) );
  TBUF_X1 \Y_tri[57]  ( .A(n444), .EN(n301), .Z(Y[57]) );
  TBUF_X1 \Y_tri[58]  ( .A(n443), .EN(n301), .Z(Y[58]) );
  TBUF_X1 \Y_tri[59]  ( .A(n442), .EN(n301), .Z(Y[59]) );
  TBUF_X1 \Y_tri[60]  ( .A(n441), .EN(n301), .Z(Y[60]) );
  TBUF_X1 \Y_tri[61]  ( .A(n440), .EN(n301), .Z(Y[61]) );
  TBUF_X1 \Y_tri[62]  ( .A(n439), .EN(n301), .Z(Y[62]) );
  TBUF_X1 \Y_tri[63]  ( .A(n438), .EN(n301), .Z(Y[63]) );
  TBUF_X1 \Y_tri[49]  ( .A(n452), .EN(n300), .Z(Y[49]) );
  TBUF_X1 \Y_tri[50]  ( .A(n451), .EN(n300), .Z(Y[50]) );
  TBUF_X1 \Y_tri[51]  ( .A(n450), .EN(n300), .Z(Y[51]) );
  TBUF_X1 \Y_tri[52]  ( .A(n449), .EN(n300), .Z(Y[52]) );
  TBUF_X1 \Y_tri[53]  ( .A(n448), .EN(n300), .Z(Y[53]) );
  TBUF_X1 \Y_tri[54]  ( .A(n447), .EN(n300), .Z(Y[54]) );
  TBUF_X1 \Y_tri[20]  ( .A(n481), .EN(n297), .Z(Y[20]) );
  TBUF_X1 \Y_tri[21]  ( .A(n480), .EN(n297), .Z(Y[21]) );
  TBUF_X1 \Y_tri[22]  ( .A(n479), .EN(n298), .Z(Y[22]) );
  TBUF_X1 \Y_tri[23]  ( .A(n478), .EN(n298), .Z(Y[23]) );
  TBUF_X1 \Y_tri[24]  ( .A(n477), .EN(n298), .Z(Y[24]) );
  TBUF_X1 \Y_tri[25]  ( .A(n476), .EN(n298), .Z(Y[25]) );
  TBUF_X1 \Y_tri[26]  ( .A(n475), .EN(n298), .Z(Y[26]) );
  TBUF_X1 \Y_tri[27]  ( .A(n474), .EN(n298), .Z(Y[27]) );
  TBUF_X1 \Y_tri[28]  ( .A(n473), .EN(n298), .Z(Y[28]) );
  TBUF_X1 \Y_tri[29]  ( .A(n472), .EN(n298), .Z(Y[29]) );
  TBUF_X1 \Y_tri[30]  ( .A(n471), .EN(n298), .Z(Y[30]) );
  TBUF_X1 \Y_tri[31]  ( .A(n470), .EN(n298), .Z(Y[31]) );
  TBUF_X1 \Y_tri[32]  ( .A(n469), .EN(n298), .Z(Y[32]) );
  TBUF_X1 \Y_tri[33]  ( .A(n468), .EN(n299), .Z(Y[33]) );
  TBUF_X1 \Y_tri[34]  ( .A(n467), .EN(n299), .Z(Y[34]) );
  TBUF_X1 \Y_tri[35]  ( .A(n466), .EN(n299), .Z(Y[35]) );
  TBUF_X1 \Y_tri[36]  ( .A(n465), .EN(n299), .Z(Y[36]) );
  TBUF_X1 \Y_tri[37]  ( .A(n464), .EN(n299), .Z(Y[37]) );
  TBUF_X1 \Y_tri[38]  ( .A(n463), .EN(n299), .Z(Y[38]) );
  TBUF_X1 \Y_tri[39]  ( .A(n462), .EN(n299), .Z(Y[39]) );
  TBUF_X1 \Y_tri[40]  ( .A(n461), .EN(n299), .Z(Y[40]) );
  TBUF_X1 \Y_tri[41]  ( .A(n460), .EN(n299), .Z(Y[41]) );
  TBUF_X1 \Y_tri[42]  ( .A(n459), .EN(n299), .Z(Y[42]) );
  TBUF_X1 \Y_tri[43]  ( .A(n458), .EN(n299), .Z(Y[43]) );
  TBUF_X1 \Y_tri[44]  ( .A(n457), .EN(n300), .Z(Y[44]) );
  TBUF_X1 \Y_tri[45]  ( .A(n456), .EN(n300), .Z(Y[45]) );
  TBUF_X1 \Y_tri[46]  ( .A(n455), .EN(n300), .Z(Y[46]) );
  TBUF_X1 \Y_tri[47]  ( .A(n454), .EN(n300), .Z(Y[47]) );
  TBUF_X1 \Y_tri[48]  ( .A(n453), .EN(n300), .Z(Y[48]) );
  TBUF_X1 \Y_tri[10]  ( .A(n491), .EN(n296), .Z(Y[10]) );
  TBUF_X1 \Y_tri[11]  ( .A(n490), .EN(n297), .Z(Y[11]) );
  TBUF_X1 \Y_tri[12]  ( .A(n489), .EN(n297), .Z(Y[12]) );
  TBUF_X1 \Y_tri[13]  ( .A(n488), .EN(n297), .Z(Y[13]) );
  TBUF_X1 \Y_tri[14]  ( .A(n487), .EN(n297), .Z(Y[14]) );
  TBUF_X1 \Y_tri[15]  ( .A(n486), .EN(n297), .Z(Y[15]) );
  TBUF_X1 \Y_tri[16]  ( .A(n485), .EN(n297), .Z(Y[16]) );
  TBUF_X1 \Y_tri[17]  ( .A(n484), .EN(n297), .Z(Y[17]) );
  TBUF_X1 \Y_tri[18]  ( .A(n483), .EN(n297), .Z(Y[18]) );
  TBUF_X1 \Y_tri[19]  ( .A(n482), .EN(n297), .Z(Y[19]) );
  TBUF_X1 \Y_tri[0]  ( .A(n502), .EN(n296), .Z(Y[0]) );
  TBUF_X1 \Y_tri[1]  ( .A(n501), .EN(n296), .Z(Y[1]) );
  TBUF_X1 \Y_tri[3]  ( .A(n499), .EN(n296), .Z(Y[3]) );
  TBUF_X1 \Y_tri[4]  ( .A(n498), .EN(n296), .Z(Y[4]) );
  TBUF_X1 \Y_tri[5]  ( .A(n497), .EN(n296), .Z(Y[5]) );
  TBUF_X1 \Y_tri[6]  ( .A(n496), .EN(n296), .Z(Y[6]) );
  TBUF_X1 \Y_tri[7]  ( .A(n495), .EN(n296), .Z(Y[7]) );
  TBUF_X1 \Y_tri[8]  ( .A(n494), .EN(n296), .Z(Y[8]) );
  TBUF_X1 \Y_tri[9]  ( .A(n492), .EN(n296), .Z(Y[9]) );
  TBUF_X1 \Y_tri[2]  ( .A(n500), .EN(n296), .Z(Y[2]) );
  NAND2_X1 U2 ( .A1(n397), .A2(n396), .ZN(n456) );
  AOI22_X1 U3 ( .A1(plusA[45]), .A2(n281), .B1(plus2A[45]), .B2(n275), .ZN(
        n397) );
  AOI22_X1 U4 ( .A1(minus2A[45]), .A2(n293), .B1(minusA[45]), .B2(n287), .ZN(
        n396) );
  NAND2_X1 U5 ( .A1(n389), .A2(n388), .ZN(n460) );
  AOI22_X1 U6 ( .A1(plusA[41]), .A2(n281), .B1(plus2A[41]), .B2(n275), .ZN(
        n389) );
  AOI22_X1 U7 ( .A1(minus2A[41]), .A2(n293), .B1(minusA[41]), .B2(n287), .ZN(
        n388) );
  NAND2_X1 U8 ( .A1(n381), .A2(n380), .ZN(n464) );
  AOI22_X1 U9 ( .A1(plusA[37]), .A2(n281), .B1(plus2A[37]), .B2(n275), .ZN(
        n381) );
  AOI22_X1 U10 ( .A1(minus2A[37]), .A2(n293), .B1(minusA[37]), .B2(n287), .ZN(
        n380) );
  NAND2_X1 U11 ( .A1(n373), .A2(n372), .ZN(n468) );
  AOI22_X1 U12 ( .A1(plusA[33]), .A2(n280), .B1(plus2A[33]), .B2(n274), .ZN(
        n373) );
  AOI22_X1 U13 ( .A1(minus2A[33]), .A2(n292), .B1(minusA[33]), .B2(n286), .ZN(
        n372) );
  NAND2_X1 U14 ( .A1(n401), .A2(n400), .ZN(n454) );
  AOI22_X1 U15 ( .A1(plusA[47]), .A2(n281), .B1(plus2A[47]), .B2(n275), .ZN(
        n401) );
  AOI22_X1 U16 ( .A1(minus2A[47]), .A2(n293), .B1(minusA[47]), .B2(n287), .ZN(
        n400) );
  NAND2_X1 U17 ( .A1(n393), .A2(n392), .ZN(n458) );
  AOI22_X1 U18 ( .A1(plusA[43]), .A2(n281), .B1(plus2A[43]), .B2(n275), .ZN(
        n393) );
  AOI22_X1 U19 ( .A1(minus2A[43]), .A2(n293), .B1(minusA[43]), .B2(n287), .ZN(
        n392) );
  NAND2_X1 U20 ( .A1(n385), .A2(n384), .ZN(n462) );
  AOI22_X1 U21 ( .A1(plusA[39]), .A2(n281), .B1(plus2A[39]), .B2(n275), .ZN(
        n385) );
  AOI22_X1 U22 ( .A1(minus2A[39]), .A2(n293), .B1(minusA[39]), .B2(n287), .ZN(
        n384) );
  NAND2_X1 U23 ( .A1(n377), .A2(n376), .ZN(n466) );
  AOI22_X1 U24 ( .A1(plusA[35]), .A2(n280), .B1(plus2A[35]), .B2(n274), .ZN(
        n377) );
  AOI22_X1 U25 ( .A1(minus2A[35]), .A2(n292), .B1(minusA[35]), .B2(n286), .ZN(
        n376) );
  NAND2_X1 U26 ( .A1(n399), .A2(n398), .ZN(n455) );
  AOI22_X1 U27 ( .A1(plusA[46]), .A2(n281), .B1(plus2A[46]), .B2(n275), .ZN(
        n399) );
  AOI22_X1 U28 ( .A1(minus2A[46]), .A2(n293), .B1(minusA[46]), .B2(n287), .ZN(
        n398) );
  NAND2_X1 U29 ( .A1(n391), .A2(n390), .ZN(n459) );
  AOI22_X1 U30 ( .A1(plusA[42]), .A2(n281), .B1(plus2A[42]), .B2(n275), .ZN(
        n391) );
  AOI22_X1 U31 ( .A1(minus2A[42]), .A2(n293), .B1(minusA[42]), .B2(n287), .ZN(
        n390) );
  NAND2_X1 U32 ( .A1(n383), .A2(n382), .ZN(n463) );
  AOI22_X1 U33 ( .A1(plusA[38]), .A2(n281), .B1(plus2A[38]), .B2(n275), .ZN(
        n383) );
  AOI22_X1 U34 ( .A1(minus2A[38]), .A2(n293), .B1(minusA[38]), .B2(n287), .ZN(
        n382) );
  NAND2_X1 U35 ( .A1(n375), .A2(n374), .ZN(n467) );
  AOI22_X1 U36 ( .A1(plusA[34]), .A2(n280), .B1(plus2A[34]), .B2(n274), .ZN(
        n375) );
  AOI22_X1 U37 ( .A1(minus2A[34]), .A2(n292), .B1(minusA[34]), .B2(n286), .ZN(
        n374) );
  NAND2_X1 U38 ( .A1(n403), .A2(n402), .ZN(n453) );
  AOI22_X1 U39 ( .A1(plusA[48]), .A2(n282), .B1(plus2A[48]), .B2(n276), .ZN(
        n403) );
  AOI22_X1 U40 ( .A1(minus2A[48]), .A2(n294), .B1(minusA[48]), .B2(n288), .ZN(
        n402) );
  NAND2_X1 U41 ( .A1(n395), .A2(n394), .ZN(n457) );
  AOI22_X1 U42 ( .A1(plusA[44]), .A2(n281), .B1(plus2A[44]), .B2(n275), .ZN(
        n395) );
  AOI22_X1 U43 ( .A1(minus2A[44]), .A2(n293), .B1(minusA[44]), .B2(n287), .ZN(
        n394) );
  NAND2_X1 U44 ( .A1(n387), .A2(n386), .ZN(n461) );
  AOI22_X1 U45 ( .A1(plusA[40]), .A2(n281), .B1(plus2A[40]), .B2(n275), .ZN(
        n387) );
  AOI22_X1 U46 ( .A1(minus2A[40]), .A2(n293), .B1(minusA[40]), .B2(n287), .ZN(
        n386) );
  NAND2_X1 U47 ( .A1(n379), .A2(n378), .ZN(n465) );
  AOI22_X1 U48 ( .A1(plusA[36]), .A2(n281), .B1(plus2A[36]), .B2(n275), .ZN(
        n379) );
  AOI22_X1 U49 ( .A1(minus2A[36]), .A2(n293), .B1(minusA[36]), .B2(n287), .ZN(
        n378) );
  NAND2_X1 U50 ( .A1(n371), .A2(n370), .ZN(n469) );
  AOI22_X1 U51 ( .A1(plusA[32]), .A2(n280), .B1(plus2A[32]), .B2(n274), .ZN(
        n371) );
  AOI22_X1 U52 ( .A1(minus2A[32]), .A2(n292), .B1(minusA[32]), .B2(n286), .ZN(
        n370) );
  NAND2_X1 U53 ( .A1(n423), .A2(n422), .ZN(n443) );
  AOI22_X1 U54 ( .A1(plusA[58]), .A2(n282), .B1(plus2A[58]), .B2(n276), .ZN(
        n423) );
  AOI22_X1 U55 ( .A1(minus2A[58]), .A2(n294), .B1(minusA[58]), .B2(n288), .ZN(
        n422) );
  NAND2_X1 U56 ( .A1(n437), .A2(n436), .ZN(n438) );
  AOI22_X1 U57 ( .A1(plusA[63]), .A2(n283), .B1(plus2A[63]), .B2(n277), .ZN(
        n437) );
  AOI22_X1 U58 ( .A1(minus2A[63]), .A2(n295), .B1(minusA[63]), .B2(n289), .ZN(
        n436) );
  NAND2_X1 U59 ( .A1(n429), .A2(n428), .ZN(n440) );
  AOI22_X1 U60 ( .A1(plusA[61]), .A2(n283), .B1(plus2A[61]), .B2(n277), .ZN(
        n429) );
  AOI22_X1 U61 ( .A1(minus2A[61]), .A2(n295), .B1(minusA[61]), .B2(n289), .ZN(
        n428) );
  NAND2_X1 U62 ( .A1(n427), .A2(n426), .ZN(n441) );
  AOI22_X1 U63 ( .A1(plusA[60]), .A2(n283), .B1(plus2A[60]), .B2(n277), .ZN(
        n427) );
  AOI22_X1 U64 ( .A1(minus2A[60]), .A2(n295), .B1(minusA[60]), .B2(n289), .ZN(
        n426) );
  NAND2_X1 U65 ( .A1(n425), .A2(n424), .ZN(n442) );
  AOI22_X1 U66 ( .A1(plusA[59]), .A2(n282), .B1(plus2A[59]), .B2(n276), .ZN(
        n425) );
  AOI22_X1 U67 ( .A1(minus2A[59]), .A2(n294), .B1(minusA[59]), .B2(n288), .ZN(
        n424) );
  NAND2_X1 U68 ( .A1(n413), .A2(n412), .ZN(n448) );
  AOI22_X1 U69 ( .A1(plusA[53]), .A2(n282), .B1(plus2A[53]), .B2(n276), .ZN(
        n413) );
  AOI22_X1 U70 ( .A1(minus2A[53]), .A2(n294), .B1(minusA[53]), .B2(n288), .ZN(
        n412) );
  NAND2_X1 U71 ( .A1(n405), .A2(n404), .ZN(n452) );
  AOI22_X1 U72 ( .A1(plusA[49]), .A2(n282), .B1(plus2A[49]), .B2(n276), .ZN(
        n405) );
  AOI22_X1 U73 ( .A1(minus2A[49]), .A2(n294), .B1(minusA[49]), .B2(n288), .ZN(
        n404) );
  NAND2_X1 U74 ( .A1(n421), .A2(n420), .ZN(n444) );
  AOI22_X1 U75 ( .A1(plusA[57]), .A2(n282), .B1(plus2A[57]), .B2(n276), .ZN(
        n421) );
  AOI22_X1 U76 ( .A1(minus2A[57]), .A2(n294), .B1(minusA[57]), .B2(n288), .ZN(
        n420) );
  NAND2_X1 U77 ( .A1(n417), .A2(n416), .ZN(n446) );
  AOI22_X1 U78 ( .A1(plusA[55]), .A2(n282), .B1(plus2A[55]), .B2(n276), .ZN(
        n417) );
  AOI22_X1 U79 ( .A1(minus2A[55]), .A2(n294), .B1(minusA[55]), .B2(n288), .ZN(
        n416) );
  NAND2_X1 U80 ( .A1(n409), .A2(n408), .ZN(n450) );
  AOI22_X1 U81 ( .A1(plusA[51]), .A2(n282), .B1(plus2A[51]), .B2(n276), .ZN(
        n409) );
  AOI22_X1 U82 ( .A1(minus2A[51]), .A2(n294), .B1(minusA[51]), .B2(n288), .ZN(
        n408) );
  NAND2_X1 U83 ( .A1(n415), .A2(n414), .ZN(n447) );
  AOI22_X1 U84 ( .A1(plusA[54]), .A2(n282), .B1(plus2A[54]), .B2(n276), .ZN(
        n415) );
  AOI22_X1 U85 ( .A1(minus2A[54]), .A2(n294), .B1(minusA[54]), .B2(n288), .ZN(
        n414) );
  NAND2_X1 U86 ( .A1(n407), .A2(n406), .ZN(n451) );
  AOI22_X1 U87 ( .A1(plusA[50]), .A2(n282), .B1(plus2A[50]), .B2(n276), .ZN(
        n407) );
  AOI22_X1 U88 ( .A1(minus2A[50]), .A2(n294), .B1(minusA[50]), .B2(n288), .ZN(
        n406) );
  NAND2_X1 U89 ( .A1(n419), .A2(n418), .ZN(n445) );
  AOI22_X1 U90 ( .A1(plusA[56]), .A2(n282), .B1(plus2A[56]), .B2(n276), .ZN(
        n419) );
  AOI22_X1 U91 ( .A1(minus2A[56]), .A2(n294), .B1(minusA[56]), .B2(n288), .ZN(
        n418) );
  NAND2_X1 U92 ( .A1(n411), .A2(n410), .ZN(n449) );
  AOI22_X1 U93 ( .A1(plusA[52]), .A2(n282), .B1(plus2A[52]), .B2(n276), .ZN(
        n411) );
  AOI22_X1 U94 ( .A1(minus2A[52]), .A2(n294), .B1(minusA[52]), .B2(n288), .ZN(
        n410) );
  NAND2_X1 U95 ( .A1(n431), .A2(n430), .ZN(n439) );
  AOI22_X1 U96 ( .A1(plusA[62]), .A2(n283), .B1(plus2A[62]), .B2(n277), .ZN(
        n431) );
  AOI22_X1 U97 ( .A1(minus2A[62]), .A2(n295), .B1(minusA[62]), .B2(n289), .ZN(
        n430) );
  BUF_X1 U98 ( .A(n493), .Z(n296) );
  BUF_X1 U99 ( .A(n493), .Z(n297) );
  BUF_X1 U100 ( .A(n433), .Z(n280) );
  BUF_X1 U101 ( .A(n435), .Z(n292) );
  BUF_X1 U102 ( .A(n434), .Z(n286) );
  BUF_X1 U103 ( .A(n432), .Z(n274) );
  BUF_X1 U104 ( .A(n493), .Z(n298) );
  NAND2_X1 U105 ( .A1(n369), .A2(n368), .ZN(n470) );
  AOI22_X1 U106 ( .A1(plusA[31]), .A2(n280), .B1(plus2A[31]), .B2(n274), .ZN(
        n369) );
  AOI22_X1 U107 ( .A1(minus2A[31]), .A2(n292), .B1(minusA[31]), .B2(n286), 
        .ZN(n368) );
  NAND2_X1 U108 ( .A1(n367), .A2(n366), .ZN(n471) );
  AOI22_X1 U109 ( .A1(plusA[30]), .A2(n280), .B1(plus2A[30]), .B2(n274), .ZN(
        n367) );
  AOI22_X1 U110 ( .A1(minus2A[30]), .A2(n292), .B1(minusA[30]), .B2(n286), 
        .ZN(n366) );
  BUF_X1 U111 ( .A(n433), .Z(n281) );
  BUF_X1 U112 ( .A(n435), .Z(n293) );
  BUF_X1 U113 ( .A(n434), .Z(n287) );
  BUF_X1 U114 ( .A(n432), .Z(n275) );
  BUF_X1 U115 ( .A(n493), .Z(n299) );
  BUF_X1 U116 ( .A(n433), .Z(n282) );
  BUF_X1 U117 ( .A(n435), .Z(n294) );
  BUF_X1 U118 ( .A(n434), .Z(n288) );
  BUF_X1 U119 ( .A(n432), .Z(n276) );
  BUF_X1 U120 ( .A(n493), .Z(n300) );
  BUF_X1 U121 ( .A(n493), .Z(n301) );
  BUF_X1 U122 ( .A(n433), .Z(n279) );
  BUF_X1 U123 ( .A(n433), .Z(n278) );
  BUF_X1 U124 ( .A(n435), .Z(n291) );
  BUF_X1 U125 ( .A(n435), .Z(n290) );
  BUF_X1 U126 ( .A(n434), .Z(n285) );
  BUF_X1 U127 ( .A(n432), .Z(n273) );
  BUF_X1 U128 ( .A(n434), .Z(n284) );
  BUF_X1 U129 ( .A(n432), .Z(n272) );
  NOR2_X1 U130 ( .A1(n323), .A2(n304), .ZN(n493) );
  INV_X1 U131 ( .A(SEL[2]), .ZN(n304) );
  NOR2_X1 U132 ( .A1(SEL[1]), .A2(SEL[0]), .ZN(n323) );
  NOR3_X1 U133 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n302), .ZN(n434) );
  NOR3_X1 U134 ( .A1(SEL[1]), .A2(SEL[2]), .A3(n303), .ZN(n433) );
  NOR3_X1 U135 ( .A1(n302), .A2(SEL[2]), .A3(n303), .ZN(n432) );
  AND2_X1 U136 ( .A1(SEL[2]), .A2(n323), .ZN(n435) );
  INV_X1 U137 ( .A(SEL[1]), .ZN(n302) );
  INV_X1 U138 ( .A(SEL[0]), .ZN(n303) );
  NAND2_X1 U139 ( .A1(n365), .A2(n364), .ZN(n472) );
  AOI22_X1 U140 ( .A1(plusA[29]), .A2(n280), .B1(plus2A[29]), .B2(n274), .ZN(
        n365) );
  AOI22_X1 U141 ( .A1(minus2A[29]), .A2(n292), .B1(minusA[29]), .B2(n286), 
        .ZN(n364) );
  NAND2_X1 U142 ( .A1(n363), .A2(n362), .ZN(n473) );
  AOI22_X1 U143 ( .A1(plusA[28]), .A2(n280), .B1(plus2A[28]), .B2(n274), .ZN(
        n363) );
  AOI22_X1 U144 ( .A1(minus2A[28]), .A2(n292), .B1(minusA[28]), .B2(n286), 
        .ZN(n362) );
  NAND2_X1 U145 ( .A1(n361), .A2(n360), .ZN(n474) );
  AOI22_X1 U146 ( .A1(plusA[27]), .A2(n280), .B1(plus2A[27]), .B2(n274), .ZN(
        n361) );
  AOI22_X1 U147 ( .A1(minus2A[27]), .A2(n292), .B1(minusA[27]), .B2(n286), 
        .ZN(n360) );
  NAND2_X1 U148 ( .A1(n359), .A2(n358), .ZN(n475) );
  AOI22_X1 U149 ( .A1(plusA[26]), .A2(n280), .B1(plus2A[26]), .B2(n274), .ZN(
        n359) );
  AOI22_X1 U150 ( .A1(minus2A[26]), .A2(n292), .B1(minusA[26]), .B2(n286), 
        .ZN(n358) );
  NAND2_X1 U151 ( .A1(n357), .A2(n356), .ZN(n476) );
  AOI22_X1 U152 ( .A1(plusA[25]), .A2(n280), .B1(plus2A[25]), .B2(n274), .ZN(
        n357) );
  AOI22_X1 U153 ( .A1(minus2A[25]), .A2(n292), .B1(minusA[25]), .B2(n286), 
        .ZN(n356) );
  NAND2_X1 U154 ( .A1(n353), .A2(n352), .ZN(n478) );
  AOI22_X1 U155 ( .A1(plusA[23]), .A2(n279), .B1(plus2A[23]), .B2(n273), .ZN(
        n353) );
  AOI22_X1 U156 ( .A1(minus2A[23]), .A2(n291), .B1(minusA[23]), .B2(n285), 
        .ZN(n352) );
  NAND2_X1 U157 ( .A1(n351), .A2(n350), .ZN(n479) );
  AOI22_X1 U158 ( .A1(plusA[22]), .A2(n279), .B1(plus2A[22]), .B2(n273), .ZN(
        n351) );
  AOI22_X1 U159 ( .A1(minus2A[22]), .A2(n291), .B1(minusA[22]), .B2(n285), 
        .ZN(n350) );
  NAND2_X1 U160 ( .A1(n349), .A2(n348), .ZN(n480) );
  AOI22_X1 U161 ( .A1(plusA[21]), .A2(n279), .B1(plus2A[21]), .B2(n273), .ZN(
        n349) );
  AOI22_X1 U162 ( .A1(minus2A[21]), .A2(n291), .B1(minusA[21]), .B2(n285), 
        .ZN(n348) );
  NAND2_X1 U163 ( .A1(n345), .A2(n344), .ZN(n482) );
  AOI22_X1 U164 ( .A1(plusA[19]), .A2(n279), .B1(plus2A[19]), .B2(n273), .ZN(
        n345) );
  AOI22_X1 U165 ( .A1(minus2A[19]), .A2(n291), .B1(minusA[19]), .B2(n285), 
        .ZN(n344) );
  NAND2_X1 U166 ( .A1(n343), .A2(n342), .ZN(n483) );
  AOI22_X1 U167 ( .A1(plusA[18]), .A2(n279), .B1(plus2A[18]), .B2(n273), .ZN(
        n343) );
  AOI22_X1 U168 ( .A1(minus2A[18]), .A2(n291), .B1(minusA[18]), .B2(n285), 
        .ZN(n342) );
  NAND2_X1 U169 ( .A1(n341), .A2(n340), .ZN(n484) );
  AOI22_X1 U170 ( .A1(plusA[17]), .A2(n279), .B1(plus2A[17]), .B2(n273), .ZN(
        n341) );
  AOI22_X1 U171 ( .A1(minus2A[17]), .A2(n291), .B1(minusA[17]), .B2(n285), 
        .ZN(n340) );
  NAND2_X1 U172 ( .A1(n337), .A2(n336), .ZN(n486) );
  AOI22_X1 U173 ( .A1(plusA[15]), .A2(n279), .B1(plus2A[15]), .B2(n273), .ZN(
        n337) );
  AOI22_X1 U174 ( .A1(minus2A[15]), .A2(n291), .B1(minusA[15]), .B2(n285), 
        .ZN(n336) );
  NAND2_X1 U175 ( .A1(n335), .A2(n334), .ZN(n487) );
  AOI22_X1 U176 ( .A1(plusA[14]), .A2(n279), .B1(plus2A[14]), .B2(n273), .ZN(
        n335) );
  AOI22_X1 U177 ( .A1(minus2A[14]), .A2(n291), .B1(minusA[14]), .B2(n285), 
        .ZN(n334) );
  NAND2_X1 U178 ( .A1(n333), .A2(n332), .ZN(n488) );
  AOI22_X1 U179 ( .A1(plusA[13]), .A2(n279), .B1(plus2A[13]), .B2(n273), .ZN(
        n333) );
  AOI22_X1 U180 ( .A1(minus2A[13]), .A2(n291), .B1(minusA[13]), .B2(n285), 
        .ZN(n332) );
  NAND2_X1 U181 ( .A1(n329), .A2(n328), .ZN(n490) );
  AOI22_X1 U182 ( .A1(plusA[11]), .A2(n278), .B1(plus2A[11]), .B2(n272), .ZN(
        n329) );
  AOI22_X1 U183 ( .A1(minus2A[11]), .A2(n290), .B1(minusA[11]), .B2(n284), 
        .ZN(n328) );
  NAND2_X1 U184 ( .A1(n327), .A2(n326), .ZN(n491) );
  AOI22_X1 U185 ( .A1(plusA[10]), .A2(n278), .B1(plus2A[10]), .B2(n272), .ZN(
        n327) );
  AOI22_X1 U186 ( .A1(minus2A[10]), .A2(n290), .B1(minusA[10]), .B2(n284), 
        .ZN(n326) );
  NAND2_X1 U187 ( .A1(n325), .A2(n324), .ZN(n492) );
  AOI22_X1 U188 ( .A1(plusA[9]), .A2(n278), .B1(plus2A[9]), .B2(n272), .ZN(
        n325) );
  AOI22_X1 U189 ( .A1(minus2A[9]), .A2(n290), .B1(minusA[9]), .B2(n284), .ZN(
        n324) );
  NAND2_X1 U190 ( .A1(n320), .A2(n319), .ZN(n495) );
  AOI22_X1 U191 ( .A1(plusA[7]), .A2(n278), .B1(plus2A[7]), .B2(n272), .ZN(
        n320) );
  AOI22_X1 U192 ( .A1(minus2A[7]), .A2(n290), .B1(minusA[7]), .B2(n284), .ZN(
        n319) );
  NAND2_X1 U193 ( .A1(n318), .A2(n317), .ZN(n496) );
  AOI22_X1 U194 ( .A1(plusA[6]), .A2(n278), .B1(plus2A[6]), .B2(n272), .ZN(
        n318) );
  AOI22_X1 U195 ( .A1(minus2A[6]), .A2(n290), .B1(minusA[6]), .B2(n284), .ZN(
        n317) );
  NAND2_X1 U196 ( .A1(n316), .A2(n315), .ZN(n497) );
  AOI22_X1 U197 ( .A1(plusA[5]), .A2(n278), .B1(plus2A[5]), .B2(n272), .ZN(
        n316) );
  AOI22_X1 U198 ( .A1(minus2A[5]), .A2(n290), .B1(minusA[5]), .B2(n284), .ZN(
        n315) );
  NAND2_X1 U199 ( .A1(n312), .A2(n311), .ZN(n499) );
  AOI22_X1 U200 ( .A1(plusA[3]), .A2(n278), .B1(plus2A[3]), .B2(n272), .ZN(
        n312) );
  AOI22_X1 U201 ( .A1(minus2A[3]), .A2(n290), .B1(minusA[3]), .B2(n284), .ZN(
        n311) );
  NAND2_X1 U202 ( .A1(n355), .A2(n354), .ZN(n477) );
  AOI22_X1 U203 ( .A1(plusA[24]), .A2(n280), .B1(plus2A[24]), .B2(n274), .ZN(
        n355) );
  AOI22_X1 U204 ( .A1(minus2A[24]), .A2(n292), .B1(minusA[24]), .B2(n286), 
        .ZN(n354) );
  NAND2_X1 U205 ( .A1(n347), .A2(n346), .ZN(n481) );
  AOI22_X1 U206 ( .A1(plusA[20]), .A2(n279), .B1(plus2A[20]), .B2(n273), .ZN(
        n347) );
  AOI22_X1 U207 ( .A1(minus2A[20]), .A2(n291), .B1(minusA[20]), .B2(n285), 
        .ZN(n346) );
  NAND2_X1 U208 ( .A1(n339), .A2(n338), .ZN(n485) );
  AOI22_X1 U209 ( .A1(plusA[16]), .A2(n279), .B1(plus2A[16]), .B2(n273), .ZN(
        n339) );
  AOI22_X1 U210 ( .A1(minus2A[16]), .A2(n291), .B1(minusA[16]), .B2(n285), 
        .ZN(n338) );
  NAND2_X1 U211 ( .A1(n331), .A2(n330), .ZN(n489) );
  AOI22_X1 U212 ( .A1(plusA[12]), .A2(n279), .B1(plus2A[12]), .B2(n273), .ZN(
        n331) );
  AOI22_X1 U213 ( .A1(minus2A[12]), .A2(n291), .B1(minusA[12]), .B2(n285), 
        .ZN(n330) );
  NAND2_X1 U214 ( .A1(n322), .A2(n321), .ZN(n494) );
  AOI22_X1 U215 ( .A1(plusA[8]), .A2(n278), .B1(plus2A[8]), .B2(n272), .ZN(
        n322) );
  AOI22_X1 U216 ( .A1(minus2A[8]), .A2(n290), .B1(minusA[8]), .B2(n284), .ZN(
        n321) );
  NAND2_X1 U217 ( .A1(n314), .A2(n313), .ZN(n498) );
  AOI22_X1 U218 ( .A1(plusA[4]), .A2(n278), .B1(plus2A[4]), .B2(n272), .ZN(
        n314) );
  AOI22_X1 U219 ( .A1(minus2A[4]), .A2(n290), .B1(minusA[4]), .B2(n284), .ZN(
        n313) );
  NAND2_X1 U220 ( .A1(n310), .A2(n309), .ZN(n500) );
  AOI22_X1 U221 ( .A1(plusA[2]), .A2(n278), .B1(plus2A[2]), .B2(n272), .ZN(
        n310) );
  AOI22_X1 U222 ( .A1(minus2A[2]), .A2(n290), .B1(minusA[2]), .B2(n284), .ZN(
        n309) );
  NAND2_X1 U223 ( .A1(n308), .A2(n307), .ZN(n501) );
  AOI22_X1 U224 ( .A1(plusA[1]), .A2(n278), .B1(plus2A[1]), .B2(n272), .ZN(
        n308) );
  AOI22_X1 U225 ( .A1(minus2A[1]), .A2(n290), .B1(minusA[1]), .B2(n284), .ZN(
        n307) );
  NAND2_X1 U226 ( .A1(n306), .A2(n305), .ZN(n502) );
  AOI22_X1 U227 ( .A1(plusA[0]), .A2(n278), .B1(plus2A[0]), .B2(n272), .ZN(
        n306) );
  AOI22_X1 U228 ( .A1(minus2A[0]), .A2(n290), .B1(minusA[0]), .B2(n284), .ZN(
        n305) );
  CLKBUF_X1 U229 ( .A(n432), .Z(n277) );
  CLKBUF_X1 U230 ( .A(n433), .Z(n283) );
  CLKBUF_X1 U231 ( .A(n434), .Z(n289) );
  CLKBUF_X1 U232 ( .A(n435), .Z(n295) );
endmodule


module FA_128 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_127 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_126 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_125 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_124 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_123 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_122 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_121 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_120 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_119 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_118 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_117 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_116 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_115 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_114 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_113 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_112 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_111 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_110 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_109 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_108 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_107 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_106 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_105 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_104 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_103 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_102 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_101 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_100 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_99 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_98 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_97 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_96 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_95 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_94 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_93 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_92 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_91 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_90 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_89 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_88 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_87 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_86 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_85 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_84 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_83 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_82 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_81 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_80 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_79 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_78 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_77 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_76 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_75 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_74 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_73 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_72 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_71 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_70 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_69 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_68 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_67 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_66 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_65 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N64_2 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Ci;
  output Co;

  wire   [63:1] CTMP;
  tri   [63:0] A;

  FA_128 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_127 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_126 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_125 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(CTMP[4]) );
  FA_124 FAI_5 ( .A(A[4]), .B(B[4]), .Ci(CTMP[4]), .S(S[4]), .Co(CTMP[5]) );
  FA_123 FAI_6 ( .A(A[5]), .B(B[5]), .Ci(CTMP[5]), .S(S[5]), .Co(CTMP[6]) );
  FA_122 FAI_7 ( .A(A[6]), .B(B[6]), .Ci(CTMP[6]), .S(S[6]), .Co(CTMP[7]) );
  FA_121 FAI_8 ( .A(A[7]), .B(B[7]), .Ci(CTMP[7]), .S(S[7]), .Co(CTMP[8]) );
  FA_120 FAI_9 ( .A(A[8]), .B(B[8]), .Ci(CTMP[8]), .S(S[8]), .Co(CTMP[9]) );
  FA_119 FAI_10 ( .A(A[9]), .B(B[9]), .Ci(CTMP[9]), .S(S[9]), .Co(CTMP[10]) );
  FA_118 FAI_11 ( .A(A[10]), .B(B[10]), .Ci(CTMP[10]), .S(S[10]), .Co(CTMP[11]) );
  FA_117 FAI_12 ( .A(A[11]), .B(B[11]), .Ci(CTMP[11]), .S(S[11]), .Co(CTMP[12]) );
  FA_116 FAI_13 ( .A(A[12]), .B(B[12]), .Ci(CTMP[12]), .S(S[12]), .Co(CTMP[13]) );
  FA_115 FAI_14 ( .A(A[13]), .B(B[13]), .Ci(CTMP[13]), .S(S[13]), .Co(CTMP[14]) );
  FA_114 FAI_15 ( .A(A[14]), .B(B[14]), .Ci(CTMP[14]), .S(S[14]), .Co(CTMP[15]) );
  FA_113 FAI_16 ( .A(A[15]), .B(B[15]), .Ci(CTMP[15]), .S(S[15]), .Co(CTMP[16]) );
  FA_112 FAI_17 ( .A(A[16]), .B(B[16]), .Ci(CTMP[16]), .S(S[16]), .Co(CTMP[17]) );
  FA_111 FAI_18 ( .A(A[17]), .B(B[17]), .Ci(CTMP[17]), .S(S[17]), .Co(CTMP[18]) );
  FA_110 FAI_19 ( .A(A[18]), .B(B[18]), .Ci(CTMP[18]), .S(S[18]), .Co(CTMP[19]) );
  FA_109 FAI_20 ( .A(A[19]), .B(B[19]), .Ci(CTMP[19]), .S(S[19]), .Co(CTMP[20]) );
  FA_108 FAI_21 ( .A(A[20]), .B(B[20]), .Ci(CTMP[20]), .S(S[20]), .Co(CTMP[21]) );
  FA_107 FAI_22 ( .A(A[21]), .B(B[21]), .Ci(CTMP[21]), .S(S[21]), .Co(CTMP[22]) );
  FA_106 FAI_23 ( .A(A[22]), .B(B[22]), .Ci(CTMP[22]), .S(S[22]), .Co(CTMP[23]) );
  FA_105 FAI_24 ( .A(A[23]), .B(B[23]), .Ci(CTMP[23]), .S(S[23]), .Co(CTMP[24]) );
  FA_104 FAI_25 ( .A(A[24]), .B(B[24]), .Ci(CTMP[24]), .S(S[24]), .Co(CTMP[25]) );
  FA_103 FAI_26 ( .A(A[25]), .B(B[25]), .Ci(CTMP[25]), .S(S[25]), .Co(CTMP[26]) );
  FA_102 FAI_27 ( .A(A[26]), .B(B[26]), .Ci(CTMP[26]), .S(S[26]), .Co(CTMP[27]) );
  FA_101 FAI_28 ( .A(A[27]), .B(B[27]), .Ci(CTMP[27]), .S(S[27]), .Co(CTMP[28]) );
  FA_100 FAI_29 ( .A(A[28]), .B(B[28]), .Ci(CTMP[28]), .S(S[28]), .Co(CTMP[29]) );
  FA_99 FAI_30 ( .A(A[29]), .B(B[29]), .Ci(CTMP[29]), .S(S[29]), .Co(CTMP[30])
         );
  FA_98 FAI_31 ( .A(A[30]), .B(B[30]), .Ci(CTMP[30]), .S(S[30]), .Co(CTMP[31])
         );
  FA_97 FAI_32 ( .A(A[31]), .B(B[31]), .Ci(CTMP[31]), .S(S[31]), .Co(CTMP[32])
         );
  FA_96 FAI_33 ( .A(A[32]), .B(B[32]), .Ci(CTMP[32]), .S(S[32]), .Co(CTMP[33])
         );
  FA_95 FAI_34 ( .A(A[33]), .B(B[33]), .Ci(CTMP[33]), .S(S[33]), .Co(CTMP[34])
         );
  FA_94 FAI_35 ( .A(A[34]), .B(B[34]), .Ci(CTMP[34]), .S(S[34]), .Co(CTMP[35])
         );
  FA_93 FAI_36 ( .A(A[35]), .B(B[35]), .Ci(CTMP[35]), .S(S[35]), .Co(CTMP[36])
         );
  FA_92 FAI_37 ( .A(A[36]), .B(B[36]), .Ci(CTMP[36]), .S(S[36]), .Co(CTMP[37])
         );
  FA_91 FAI_38 ( .A(A[37]), .B(B[37]), .Ci(CTMP[37]), .S(S[37]), .Co(CTMP[38])
         );
  FA_90 FAI_39 ( .A(A[38]), .B(B[38]), .Ci(CTMP[38]), .S(S[38]), .Co(CTMP[39])
         );
  FA_89 FAI_40 ( .A(A[39]), .B(B[39]), .Ci(CTMP[39]), .S(S[39]), .Co(CTMP[40])
         );
  FA_88 FAI_41 ( .A(A[40]), .B(B[40]), .Ci(CTMP[40]), .S(S[40]), .Co(CTMP[41])
         );
  FA_87 FAI_42 ( .A(A[41]), .B(B[41]), .Ci(CTMP[41]), .S(S[41]), .Co(CTMP[42])
         );
  FA_86 FAI_43 ( .A(A[42]), .B(B[42]), .Ci(CTMP[42]), .S(S[42]), .Co(CTMP[43])
         );
  FA_85 FAI_44 ( .A(A[43]), .B(B[43]), .Ci(CTMP[43]), .S(S[43]), .Co(CTMP[44])
         );
  FA_84 FAI_45 ( .A(A[44]), .B(B[44]), .Ci(CTMP[44]), .S(S[44]), .Co(CTMP[45])
         );
  FA_83 FAI_46 ( .A(A[45]), .B(B[45]), .Ci(CTMP[45]), .S(S[45]), .Co(CTMP[46])
         );
  FA_82 FAI_47 ( .A(A[46]), .B(B[46]), .Ci(CTMP[46]), .S(S[46]), .Co(CTMP[47])
         );
  FA_81 FAI_48 ( .A(A[47]), .B(B[47]), .Ci(CTMP[47]), .S(S[47]), .Co(CTMP[48])
         );
  FA_80 FAI_49 ( .A(A[48]), .B(B[48]), .Ci(CTMP[48]), .S(S[48]), .Co(CTMP[49])
         );
  FA_79 FAI_50 ( .A(A[49]), .B(B[49]), .Ci(CTMP[49]), .S(S[49]), .Co(CTMP[50])
         );
  FA_78 FAI_51 ( .A(A[50]), .B(B[50]), .Ci(CTMP[50]), .S(S[50]), .Co(CTMP[51])
         );
  FA_77 FAI_52 ( .A(A[51]), .B(B[51]), .Ci(CTMP[51]), .S(S[51]), .Co(CTMP[52])
         );
  FA_76 FAI_53 ( .A(A[52]), .B(B[52]), .Ci(CTMP[52]), .S(S[52]), .Co(CTMP[53])
         );
  FA_75 FAI_54 ( .A(A[53]), .B(B[53]), .Ci(CTMP[53]), .S(S[53]), .Co(CTMP[54])
         );
  FA_74 FAI_55 ( .A(A[54]), .B(B[54]), .Ci(CTMP[54]), .S(S[54]), .Co(CTMP[55])
         );
  FA_73 FAI_56 ( .A(A[55]), .B(B[55]), .Ci(CTMP[55]), .S(S[55]), .Co(CTMP[56])
         );
  FA_72 FAI_57 ( .A(A[56]), .B(B[56]), .Ci(CTMP[56]), .S(S[56]), .Co(CTMP[57])
         );
  FA_71 FAI_58 ( .A(A[57]), .B(B[57]), .Ci(CTMP[57]), .S(S[57]), .Co(CTMP[58])
         );
  FA_70 FAI_59 ( .A(A[58]), .B(B[58]), .Ci(CTMP[58]), .S(S[58]), .Co(CTMP[59])
         );
  FA_69 FAI_60 ( .A(A[59]), .B(B[59]), .Ci(CTMP[59]), .S(S[59]), .Co(CTMP[60])
         );
  FA_68 FAI_61 ( .A(A[60]), .B(B[60]), .Ci(CTMP[60]), .S(S[60]), .Co(CTMP[61])
         );
  FA_67 FAI_62 ( .A(A[61]), .B(B[61]), .Ci(CTMP[61]), .S(S[61]), .Co(CTMP[62])
         );
  FA_66 FAI_63 ( .A(A[62]), .B(B[62]), .Ci(CTMP[62]), .S(S[62]), .Co(CTMP[63])
         );
  FA_65 FAI_64 ( .A(A[63]), .B(B[63]), .Ci(CTMP[63]), .S(S[63]), .Co(Co) );
endmodule


module booth_mul_row_N64_RADIX3_2 ( prevA, prevSum, encoderIn, nextA, nextSum
 );
  input [63:0] prevA;
  input [63:0] prevSum;
  input [2:0] encoderIn;
  output [63:0] nextA;
  output [63:0] nextSum;

  wire   [2:0] encoder_to_mux;
  wire   [63:0] plus2A_s;
  wire   [63:0] minus2A_s;
  wire   [63:0] minus4A_s;
  tri   [63:0] mux_to_adder;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign nextA[0] = 1'b0;

  encoder_N64_RADIX3_2 encoder_1 ( .X(encoderIn), .Z(encoder_to_mux) );
  ShiftnCompl_N64_2 ShiftnCompl_1 ( .plusA(prevA), .plus2A_out({plus2A_s[63:1], 
        SYNOPSYS_UNCONNECTED__0}), .minus2A_out(minus2A_s), .plus4A_out({
        nextA[63:1], SYNOPSYS_UNCONNECTED__1}), .minus4A_out(minus4A_s) );
  MUX_GENERIC_N64_RADIX3_2 mux_1 ( .plusA({plus2A_s[63:1], 1'b0}), .minusA(
        minus2A_s), .plus2A({nextA[63:1], 1'b0}), .minus2A(minus4A_s), .SEL(
        encoder_to_mux), .Y(mux_to_adder) );
  RCA_N64_2 rca_1 ( .A(mux_to_adder), .B(prevSum), .Ci(1'b0), .S(nextSum) );
endmodule


module encoder_N64_RADIX3_1 ( X, Z );
  input [2:0] X;
  output [2:0] Z;
  wire   n5, n7, n8;

  OAI22_X1 U1 ( .A1(n8), .A2(n5), .B1(X[2]), .B2(n7), .ZN(Z[1]) );
  INV_X1 U2 ( .A(X[2]), .ZN(n5) );
  AOI21_X1 U3 ( .B1(n8), .B2(n7), .A(X[2]), .ZN(Z[0]) );
  OAI21_X1 U4 ( .B1(X[1]), .B2(X[0]), .A(n7), .ZN(n8) );
  AND3_X1 U5 ( .A1(X[2]), .A2(n7), .A3(n8), .ZN(Z[2]) );
  NAND2_X1 U6 ( .A1(X[1]), .A2(X[0]), .ZN(n7) );
endmodule


module shifter_N64_2 ( \input , shiftLeftOnePos );
  input [63:0] \input ;
  output [63:0] shiftLeftOnePos;
  wire   \input[62] , \input[61] , \input[60] , \input[59] , \input[58] ,
         \input[57] , \input[56] , \input[55] , \input[54] , \input[53] ,
         \input[52] , \input[51] , \input[50] , \input[49] , \input[48] ,
         \input[47] , \input[46] , \input[45] , \input[44] , \input[43] ,
         \input[42] , \input[41] , \input[40] , \input[39] , \input[38] ,
         \input[37] , \input[36] , \input[35] , \input[34] , \input[33] ,
         \input[32] , \input[31] , \input[30] , \input[29] , \input[28] ,
         \input[27] , \input[26] , \input[25] , \input[24] , \input[23] ,
         \input[22] , \input[21] , \input[20] , \input[19] , \input[18] ,
         \input[17] , \input[16] , \input[15] , \input[14] , \input[13] ,
         \input[12] , \input[11] , \input[10] , \input[9] , \input[8] ,
         \input[7] , \input[6] , \input[5] , \input[4] , \input[3] ,
         \input[2] , \input[1] , \input[0] ;
  assign shiftLeftOnePos[0] = 1'b0;
  assign shiftLeftOnePos[63] = \input[62] ;
  assign \input[62]  = \input  [62];
  assign shiftLeftOnePos[62] = \input[61] ;
  assign \input[61]  = \input  [61];
  assign shiftLeftOnePos[61] = \input[60] ;
  assign \input[60]  = \input  [60];
  assign shiftLeftOnePos[60] = \input[59] ;
  assign \input[59]  = \input  [59];
  assign shiftLeftOnePos[59] = \input[58] ;
  assign \input[58]  = \input  [58];
  assign shiftLeftOnePos[58] = \input[57] ;
  assign \input[57]  = \input  [57];
  assign shiftLeftOnePos[57] = \input[56] ;
  assign \input[56]  = \input  [56];
  assign shiftLeftOnePos[56] = \input[55] ;
  assign \input[55]  = \input  [55];
  assign shiftLeftOnePos[55] = \input[54] ;
  assign \input[54]  = \input  [54];
  assign shiftLeftOnePos[54] = \input[53] ;
  assign \input[53]  = \input  [53];
  assign shiftLeftOnePos[53] = \input[52] ;
  assign \input[52]  = \input  [52];
  assign shiftLeftOnePos[52] = \input[51] ;
  assign \input[51]  = \input  [51];
  assign shiftLeftOnePos[51] = \input[50] ;
  assign \input[50]  = \input  [50];
  assign shiftLeftOnePos[50] = \input[49] ;
  assign \input[49]  = \input  [49];
  assign shiftLeftOnePos[49] = \input[48] ;
  assign \input[48]  = \input  [48];
  assign shiftLeftOnePos[48] = \input[47] ;
  assign \input[47]  = \input  [47];
  assign shiftLeftOnePos[47] = \input[46] ;
  assign \input[46]  = \input  [46];
  assign shiftLeftOnePos[46] = \input[45] ;
  assign \input[45]  = \input  [45];
  assign shiftLeftOnePos[45] = \input[44] ;
  assign \input[44]  = \input  [44];
  assign shiftLeftOnePos[44] = \input[43] ;
  assign \input[43]  = \input  [43];
  assign shiftLeftOnePos[43] = \input[42] ;
  assign \input[42]  = \input  [42];
  assign shiftLeftOnePos[42] = \input[41] ;
  assign \input[41]  = \input  [41];
  assign shiftLeftOnePos[41] = \input[40] ;
  assign \input[40]  = \input  [40];
  assign shiftLeftOnePos[40] = \input[39] ;
  assign \input[39]  = \input  [39];
  assign shiftLeftOnePos[39] = \input[38] ;
  assign \input[38]  = \input  [38];
  assign shiftLeftOnePos[38] = \input[37] ;
  assign \input[37]  = \input  [37];
  assign shiftLeftOnePos[37] = \input[36] ;
  assign \input[36]  = \input  [36];
  assign shiftLeftOnePos[36] = \input[35] ;
  assign \input[35]  = \input  [35];
  assign shiftLeftOnePos[35] = \input[34] ;
  assign \input[34]  = \input  [34];
  assign shiftLeftOnePos[34] = \input[33] ;
  assign \input[33]  = \input  [33];
  assign shiftLeftOnePos[33] = \input[32] ;
  assign \input[32]  = \input  [32];
  assign shiftLeftOnePos[32] = \input[31] ;
  assign \input[31]  = \input  [31];
  assign shiftLeftOnePos[31] = \input[30] ;
  assign \input[30]  = \input  [30];
  assign shiftLeftOnePos[30] = \input[29] ;
  assign \input[29]  = \input  [29];
  assign shiftLeftOnePos[29] = \input[28] ;
  assign \input[28]  = \input  [28];
  assign shiftLeftOnePos[28] = \input[27] ;
  assign \input[27]  = \input  [27];
  assign shiftLeftOnePos[27] = \input[26] ;
  assign \input[26]  = \input  [26];
  assign shiftLeftOnePos[26] = \input[25] ;
  assign \input[25]  = \input  [25];
  assign shiftLeftOnePos[25] = \input[24] ;
  assign \input[24]  = \input  [24];
  assign shiftLeftOnePos[24] = \input[23] ;
  assign \input[23]  = \input  [23];
  assign shiftLeftOnePos[23] = \input[22] ;
  assign \input[22]  = \input  [22];
  assign shiftLeftOnePos[22] = \input[21] ;
  assign \input[21]  = \input  [21];
  assign shiftLeftOnePos[21] = \input[20] ;
  assign \input[20]  = \input  [20];
  assign shiftLeftOnePos[20] = \input[19] ;
  assign \input[19]  = \input  [19];
  assign shiftLeftOnePos[19] = \input[18] ;
  assign \input[18]  = \input  [18];
  assign shiftLeftOnePos[18] = \input[17] ;
  assign \input[17]  = \input  [17];
  assign shiftLeftOnePos[17] = \input[16] ;
  assign \input[16]  = \input  [16];
  assign shiftLeftOnePos[16] = \input[15] ;
  assign \input[15]  = \input  [15];
  assign shiftLeftOnePos[15] = \input[14] ;
  assign \input[14]  = \input  [14];
  assign shiftLeftOnePos[14] = \input[13] ;
  assign \input[13]  = \input  [13];
  assign shiftLeftOnePos[13] = \input[12] ;
  assign \input[12]  = \input  [12];
  assign shiftLeftOnePos[12] = \input[11] ;
  assign \input[11]  = \input  [11];
  assign shiftLeftOnePos[11] = \input[10] ;
  assign \input[10]  = \input  [10];
  assign shiftLeftOnePos[10] = \input[9] ;
  assign \input[9]  = \input  [9];
  assign shiftLeftOnePos[9] = \input[8] ;
  assign \input[8]  = \input  [8];
  assign shiftLeftOnePos[8] = \input[7] ;
  assign \input[7]  = \input  [7];
  assign shiftLeftOnePos[7] = \input[6] ;
  assign \input[6]  = \input  [6];
  assign shiftLeftOnePos[6] = \input[5] ;
  assign \input[5]  = \input  [5];
  assign shiftLeftOnePos[5] = \input[4] ;
  assign \input[4]  = \input  [4];
  assign shiftLeftOnePos[4] = \input[3] ;
  assign \input[3]  = \input  [3];
  assign shiftLeftOnePos[3] = \input[2] ;
  assign \input[2]  = \input  [2];
  assign shiftLeftOnePos[2] = \input[1] ;
  assign \input[1]  = \input  [1];
  assign shiftLeftOnePos[1] = \input[0] ;
  assign \input[0]  = \input  [0];

endmodule


module shifter_N64_1 ( \input , shiftLeftOnePos );
  input [63:0] \input ;
  output [63:0] shiftLeftOnePos;
  wire   \input[62] , \input[61] , \input[60] , \input[59] , \input[58] ,
         \input[57] , \input[56] , \input[55] , \input[54] , \input[53] ,
         \input[52] , \input[51] , \input[50] , \input[49] , \input[48] ,
         \input[47] , \input[46] , \input[45] , \input[44] , \input[43] ,
         \input[42] , \input[41] , \input[40] , \input[39] , \input[38] ,
         \input[37] , \input[36] , \input[35] , \input[34] , \input[33] ,
         \input[32] , \input[31] , \input[30] , \input[29] , \input[28] ,
         \input[27] , \input[26] , \input[25] , \input[24] , \input[23] ,
         \input[22] , \input[21] , \input[20] , \input[19] , \input[18] ,
         \input[17] , \input[16] , \input[15] , \input[14] , \input[13] ,
         \input[12] , \input[11] , \input[10] , \input[9] , \input[8] ,
         \input[7] , \input[6] , \input[5] , \input[4] , \input[3] ,
         \input[2] , \input[1] , \input[0] ;
  assign shiftLeftOnePos[0] = 1'b0;
  assign shiftLeftOnePos[63] = \input[62] ;
  assign \input[62]  = \input  [62];
  assign shiftLeftOnePos[62] = \input[61] ;
  assign \input[61]  = \input  [61];
  assign shiftLeftOnePos[61] = \input[60] ;
  assign \input[60]  = \input  [60];
  assign shiftLeftOnePos[60] = \input[59] ;
  assign \input[59]  = \input  [59];
  assign shiftLeftOnePos[59] = \input[58] ;
  assign \input[58]  = \input  [58];
  assign shiftLeftOnePos[58] = \input[57] ;
  assign \input[57]  = \input  [57];
  assign shiftLeftOnePos[57] = \input[56] ;
  assign \input[56]  = \input  [56];
  assign shiftLeftOnePos[56] = \input[55] ;
  assign \input[55]  = \input  [55];
  assign shiftLeftOnePos[55] = \input[54] ;
  assign \input[54]  = \input  [54];
  assign shiftLeftOnePos[54] = \input[53] ;
  assign \input[53]  = \input  [53];
  assign shiftLeftOnePos[53] = \input[52] ;
  assign \input[52]  = \input  [52];
  assign shiftLeftOnePos[52] = \input[51] ;
  assign \input[51]  = \input  [51];
  assign shiftLeftOnePos[51] = \input[50] ;
  assign \input[50]  = \input  [50];
  assign shiftLeftOnePos[50] = \input[49] ;
  assign \input[49]  = \input  [49];
  assign shiftLeftOnePos[49] = \input[48] ;
  assign \input[48]  = \input  [48];
  assign shiftLeftOnePos[48] = \input[47] ;
  assign \input[47]  = \input  [47];
  assign shiftLeftOnePos[47] = \input[46] ;
  assign \input[46]  = \input  [46];
  assign shiftLeftOnePos[46] = \input[45] ;
  assign \input[45]  = \input  [45];
  assign shiftLeftOnePos[45] = \input[44] ;
  assign \input[44]  = \input  [44];
  assign shiftLeftOnePos[44] = \input[43] ;
  assign \input[43]  = \input  [43];
  assign shiftLeftOnePos[43] = \input[42] ;
  assign \input[42]  = \input  [42];
  assign shiftLeftOnePos[42] = \input[41] ;
  assign \input[41]  = \input  [41];
  assign shiftLeftOnePos[41] = \input[40] ;
  assign \input[40]  = \input  [40];
  assign shiftLeftOnePos[40] = \input[39] ;
  assign \input[39]  = \input  [39];
  assign shiftLeftOnePos[39] = \input[38] ;
  assign \input[38]  = \input  [38];
  assign shiftLeftOnePos[38] = \input[37] ;
  assign \input[37]  = \input  [37];
  assign shiftLeftOnePos[37] = \input[36] ;
  assign \input[36]  = \input  [36];
  assign shiftLeftOnePos[36] = \input[35] ;
  assign \input[35]  = \input  [35];
  assign shiftLeftOnePos[35] = \input[34] ;
  assign \input[34]  = \input  [34];
  assign shiftLeftOnePos[34] = \input[33] ;
  assign \input[33]  = \input  [33];
  assign shiftLeftOnePos[33] = \input[32] ;
  assign \input[32]  = \input  [32];
  assign shiftLeftOnePos[32] = \input[31] ;
  assign \input[31]  = \input  [31];
  assign shiftLeftOnePos[31] = \input[30] ;
  assign \input[30]  = \input  [30];
  assign shiftLeftOnePos[30] = \input[29] ;
  assign \input[29]  = \input  [29];
  assign shiftLeftOnePos[29] = \input[28] ;
  assign \input[28]  = \input  [28];
  assign shiftLeftOnePos[28] = \input[27] ;
  assign \input[27]  = \input  [27];
  assign shiftLeftOnePos[27] = \input[26] ;
  assign \input[26]  = \input  [26];
  assign shiftLeftOnePos[26] = \input[25] ;
  assign \input[25]  = \input  [25];
  assign shiftLeftOnePos[25] = \input[24] ;
  assign \input[24]  = \input  [24];
  assign shiftLeftOnePos[24] = \input[23] ;
  assign \input[23]  = \input  [23];
  assign shiftLeftOnePos[23] = \input[22] ;
  assign \input[22]  = \input  [22];
  assign shiftLeftOnePos[22] = \input[21] ;
  assign \input[21]  = \input  [21];
  assign shiftLeftOnePos[21] = \input[20] ;
  assign \input[20]  = \input  [20];
  assign shiftLeftOnePos[20] = \input[19] ;
  assign \input[19]  = \input  [19];
  assign shiftLeftOnePos[19] = \input[18] ;
  assign \input[18]  = \input  [18];
  assign shiftLeftOnePos[18] = \input[17] ;
  assign \input[17]  = \input  [17];
  assign shiftLeftOnePos[17] = \input[16] ;
  assign \input[16]  = \input  [16];
  assign shiftLeftOnePos[16] = \input[15] ;
  assign \input[15]  = \input  [15];
  assign shiftLeftOnePos[15] = \input[14] ;
  assign \input[14]  = \input  [14];
  assign shiftLeftOnePos[14] = \input[13] ;
  assign \input[13]  = \input  [13];
  assign shiftLeftOnePos[13] = \input[12] ;
  assign \input[12]  = \input  [12];
  assign shiftLeftOnePos[12] = \input[11] ;
  assign \input[11]  = \input  [11];
  assign shiftLeftOnePos[11] = \input[10] ;
  assign \input[10]  = \input  [10];
  assign shiftLeftOnePos[10] = \input[9] ;
  assign \input[9]  = \input  [9];
  assign shiftLeftOnePos[9] = \input[8] ;
  assign \input[8]  = \input  [8];
  assign shiftLeftOnePos[8] = \input[7] ;
  assign \input[7]  = \input  [7];
  assign shiftLeftOnePos[7] = \input[6] ;
  assign \input[6]  = \input  [6];
  assign shiftLeftOnePos[6] = \input[5] ;
  assign \input[5]  = \input  [5];
  assign shiftLeftOnePos[5] = \input[4] ;
  assign \input[4]  = \input  [4];
  assign shiftLeftOnePos[4] = \input[3] ;
  assign \input[3]  = \input  [3];
  assign shiftLeftOnePos[3] = \input[2] ;
  assign \input[2]  = \input  [2];
  assign shiftLeftOnePos[2] = \input[1] ;
  assign \input[1]  = \input  [1];
  assign shiftLeftOnePos[1] = \input[0] ;
  assign \input[0]  = \input  [0];

endmodule


module complementer_N64_2_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n190, n191, n192, n193, n194, n196, n197, n198, n199, n200,
         n202, n203, n204, n206, n207, n208, n210, n211, n212, n213, n214,
         n216, n217, n218, n220, n221, n222, n224, n225, n226, n228, n229,
         n230, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n189,
         n195, n201, n205, n209, n215, n219, n223, n227, n231;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U81 ( .A(n190), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U82 ( .A(n192), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U83 ( .A(n193), .B(B[6]), .Z(DIFF[6]) );
  XOR2_X1 U85 ( .A(n196), .B(B[62]), .Z(DIFF[62]) );
  XOR2_X1 U86 ( .A(n194), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U87 ( .A(n198), .B(B[59]), .Z(DIFF[59]) );
  XOR2_X1 U89 ( .A(n200), .B(B[57]), .Z(DIFF[57]) );
  XOR2_X1 U90 ( .A(n202), .B(B[55]), .Z(DIFF[55]) );
  XOR2_X1 U92 ( .A(n204), .B(B[53]), .Z(DIFF[53]) );
  XOR2_X1 U93 ( .A(n206), .B(B[51]), .Z(DIFF[51]) );
  XOR2_X1 U95 ( .A(n208), .B(B[49]), .Z(DIFF[49]) );
  XOR2_X1 U96 ( .A(n212), .B(B[47]), .Z(DIFF[47]) );
  XOR2_X1 U98 ( .A(n214), .B(B[45]), .Z(DIFF[45]) );
  XOR2_X1 U99 ( .A(n216), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U101 ( .A(n218), .B(B[41]), .Z(DIFF[41]) );
  XOR2_X1 U102 ( .A(n211), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U103 ( .A(n220), .B(B[39]), .Z(DIFF[39]) );
  XOR2_X1 U105 ( .A(n222), .B(B[37]), .Z(DIFF[37]) );
  XOR2_X1 U106 ( .A(n224), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U108 ( .A(n226), .B(B[33]), .Z(DIFF[33]) );
  XOR2_X1 U109 ( .A(n228), .B(B[31]), .Z(DIFF[31]) );
  XOR2_X1 U111 ( .A(n230), .B(B[29]), .Z(DIFF[29]) );
  XOR2_X1 U112 ( .A(n233), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U113 ( .A(n236), .B(B[26]), .Z(DIFF[26]) );
  XOR2_X1 U114 ( .A(n235), .B(B[25]), .Z(DIFF[25]) );
  XOR2_X1 U115 ( .A(n237), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U116 ( .A(n240), .B(B[22]), .Z(DIFF[22]) );
  XOR2_X1 U117 ( .A(n239), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U118 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U119 ( .A(n241), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U120 ( .A(n244), .B(B[18]), .Z(DIFF[18]) );
  XOR2_X1 U121 ( .A(n243), .B(B[17]), .Z(DIFF[17]) );
  XOR2_X1 U122 ( .A(n245), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U123 ( .A(n248), .B(B[14]), .Z(DIFF[14]) );
  XOR2_X1 U124 ( .A(n247), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U125 ( .A(n249), .B(B[11]), .Z(DIFF[11]) );
  XOR2_X1 U126 ( .A(n251), .B(B[10]), .Z(DIFF[10]) );
  XNOR2_X1 U1 ( .A(n189), .B(B[63]), .ZN(DIFF[63]) );
  NOR2_X1 U2 ( .A1(n196), .A2(B[62]), .ZN(n189) );
  XOR2_X1 U3 ( .A(n197), .B(n231), .Z(DIFF[61]) );
  NAND2_X1 U4 ( .A1(n197), .A2(n231), .ZN(n196) );
  NOR3_X1 U5 ( .A1(B[59]), .A2(B[60]), .A3(n198), .ZN(n197) );
  XNOR2_X1 U6 ( .A(n195), .B(B[54]), .ZN(DIFF[54]) );
  NOR2_X1 U7 ( .A1(n204), .A2(B[53]), .ZN(n195) );
  XNOR2_X1 U8 ( .A(n201), .B(B[50]), .ZN(DIFF[50]) );
  NOR2_X1 U9 ( .A1(n208), .A2(B[49]), .ZN(n201) );
  XNOR2_X1 U10 ( .A(n205), .B(B[42]), .ZN(DIFF[42]) );
  NOR2_X1 U11 ( .A1(n218), .A2(B[41]), .ZN(n205) );
  XNOR2_X1 U12 ( .A(n209), .B(B[58]), .ZN(DIFF[58]) );
  NOR2_X1 U13 ( .A1(n200), .A2(B[57]), .ZN(n209) );
  XNOR2_X1 U14 ( .A(B[60]), .B(n199), .ZN(DIFF[60]) );
  NOR2_X1 U15 ( .A1(B[59]), .A2(n198), .ZN(n199) );
  XNOR2_X1 U16 ( .A(B[56]), .B(n203), .ZN(DIFF[56]) );
  NOR2_X1 U17 ( .A1(B[55]), .A2(n202), .ZN(n203) );
  XNOR2_X1 U18 ( .A(B[52]), .B(n207), .ZN(DIFF[52]) );
  NOR2_X1 U19 ( .A1(B[51]), .A2(n206), .ZN(n207) );
  XNOR2_X1 U20 ( .A(B[48]), .B(n213), .ZN(DIFF[48]) );
  NOR2_X1 U21 ( .A1(B[47]), .A2(n212), .ZN(n213) );
  XNOR2_X1 U22 ( .A(B[44]), .B(n217), .ZN(DIFF[44]) );
  NOR2_X1 U23 ( .A1(B[43]), .A2(n216), .ZN(n217) );
  OR3_X1 U24 ( .A1(B[57]), .A2(B[58]), .A3(n200), .ZN(n198) );
  OR3_X1 U25 ( .A1(B[41]), .A2(B[42]), .A3(n218), .ZN(n216) );
  OR3_X1 U26 ( .A1(B[45]), .A2(B[46]), .A3(n214), .ZN(n212) );
  OR3_X1 U27 ( .A1(B[49]), .A2(B[50]), .A3(n208), .ZN(n206) );
  OR3_X1 U28 ( .A1(B[53]), .A2(B[54]), .A3(n204), .ZN(n202) );
  OR3_X1 U29 ( .A1(B[43]), .A2(B[44]), .A3(n216), .ZN(n214) );
  OR3_X1 U30 ( .A1(B[47]), .A2(B[48]), .A3(n212), .ZN(n208) );
  OR3_X1 U31 ( .A1(B[51]), .A2(B[52]), .A3(n206), .ZN(n204) );
  OR3_X1 U32 ( .A1(B[55]), .A2(B[56]), .A3(n202), .ZN(n200) );
  XNOR2_X1 U33 ( .A(n215), .B(B[46]), .ZN(DIFF[46]) );
  NOR2_X1 U34 ( .A1(n214), .A2(B[45]), .ZN(n215) );
  XNOR2_X1 U35 ( .A(B[40]), .B(n221), .ZN(DIFF[40]) );
  NOR2_X1 U36 ( .A1(B[39]), .A2(n220), .ZN(n221) );
  OR3_X1 U37 ( .A1(B[39]), .A2(B[40]), .A3(n220), .ZN(n218) );
  XNOR2_X1 U38 ( .A(n219), .B(B[38]), .ZN(DIFF[38]) );
  NOR2_X1 U39 ( .A1(n222), .A2(B[37]), .ZN(n219) );
  OR3_X1 U40 ( .A1(B[37]), .A2(B[38]), .A3(n222), .ZN(n220) );
  XNOR2_X1 U41 ( .A(B[36]), .B(n225), .ZN(DIFF[36]) );
  NOR2_X1 U42 ( .A1(B[35]), .A2(n224), .ZN(n225) );
  OR3_X1 U43 ( .A1(B[35]), .A2(B[36]), .A3(n224), .ZN(n222) );
  XNOR2_X1 U44 ( .A(n223), .B(B[34]), .ZN(DIFF[34]) );
  NOR2_X1 U45 ( .A1(n226), .A2(B[33]), .ZN(n223) );
  OR3_X1 U46 ( .A1(B[33]), .A2(B[34]), .A3(n226), .ZN(n224) );
  XNOR2_X1 U47 ( .A(B[32]), .B(n229), .ZN(DIFF[32]) );
  NOR2_X1 U48 ( .A1(B[31]), .A2(n228), .ZN(n229) );
  OR3_X1 U49 ( .A1(B[31]), .A2(B[32]), .A3(n228), .ZN(n226) );
  XNOR2_X1 U50 ( .A(n227), .B(B[30]), .ZN(DIFF[30]) );
  NOR2_X1 U51 ( .A1(n230), .A2(B[29]), .ZN(n227) );
  OR3_X1 U52 ( .A1(B[29]), .A2(B[30]), .A3(n230), .ZN(n228) );
  NOR2_X1 U53 ( .A1(B[27]), .A2(n233), .ZN(n234) );
  NOR2_X1 U54 ( .A1(B[23]), .A2(n237), .ZN(n238) );
  NOR2_X1 U55 ( .A1(B[19]), .A2(n241), .ZN(n242) );
  NOR2_X1 U56 ( .A1(B[15]), .A2(n245), .ZN(n246) );
  NOR2_X1 U57 ( .A1(B[11]), .A2(n249), .ZN(n250) );
  NOR2_X1 U58 ( .A1(B[7]), .A2(n192), .ZN(n191) );
  NOR2_X1 U59 ( .A1(B[3]), .A2(n211), .ZN(n210) );
  OR3_X1 U60 ( .A1(B[25]), .A2(B[26]), .A3(n235), .ZN(n233) );
  OR3_X1 U61 ( .A1(B[21]), .A2(B[22]), .A3(n239), .ZN(n237) );
  OR3_X1 U62 ( .A1(B[17]), .A2(B[18]), .A3(n243), .ZN(n241) );
  OR3_X1 U63 ( .A1(B[13]), .A2(B[14]), .A3(n247), .ZN(n245) );
  OR3_X1 U64 ( .A1(B[10]), .A2(B[9]), .A3(n190), .ZN(n249) );
  OR3_X1 U65 ( .A1(B[5]), .A2(B[6]), .A3(n194), .ZN(n192) );
  OR3_X1 U66 ( .A1(B[27]), .A2(B[28]), .A3(n233), .ZN(n230) );
  OR3_X1 U67 ( .A1(B[23]), .A2(B[24]), .A3(n237), .ZN(n235) );
  OR3_X1 U68 ( .A1(B[19]), .A2(B[20]), .A3(n241), .ZN(n239) );
  OR3_X1 U69 ( .A1(B[15]), .A2(B[16]), .A3(n245), .ZN(n243) );
  OR3_X1 U70 ( .A1(B[11]), .A2(B[12]), .A3(n249), .ZN(n247) );
  OR3_X1 U71 ( .A1(B[7]), .A2(B[8]), .A3(n192), .ZN(n190) );
  OR3_X1 U72 ( .A1(B[3]), .A2(B[4]), .A3(n211), .ZN(n194) );
  XNOR2_X1 U73 ( .A(B[28]), .B(n234), .ZN(DIFF[28]) );
  XNOR2_X1 U74 ( .A(B[24]), .B(n238), .ZN(DIFF[24]) );
  XNOR2_X1 U75 ( .A(B[20]), .B(n242), .ZN(DIFF[20]) );
  XNOR2_X1 U76 ( .A(B[16]), .B(n246), .ZN(DIFF[16]) );
  XNOR2_X1 U77 ( .A(B[12]), .B(n250), .ZN(DIFF[12]) );
  XNOR2_X1 U78 ( .A(B[8]), .B(n191), .ZN(DIFF[8]) );
  XNOR2_X1 U79 ( .A(B[4]), .B(n210), .ZN(DIFF[4]) );
  XNOR2_X1 U80 ( .A(B[2]), .B(n232), .ZN(DIFF[2]) );
  OR2_X1 U84 ( .A1(n235), .A2(B[25]), .ZN(n236) );
  OR2_X1 U88 ( .A1(n239), .A2(B[21]), .ZN(n240) );
  OR2_X1 U91 ( .A1(n243), .A2(B[17]), .ZN(n244) );
  OR2_X1 U94 ( .A1(n247), .A2(B[13]), .ZN(n248) );
  OR2_X1 U97 ( .A1(n190), .A2(B[9]), .ZN(n251) );
  OR2_X1 U100 ( .A1(n194), .A2(B[5]), .ZN(n193) );
  OR3_X1 U104 ( .A1(B[1]), .A2(B[2]), .A3(\B[0] ), .ZN(n211) );
  NOR2_X1 U107 ( .A1(\B[0] ), .A2(B[1]), .ZN(n232) );
  INV_X1 U110 ( .A(B[61]), .ZN(n231) );
endmodule


module complementer_N64_2 ( \input , complement2 );
  input [63:0] \input ;
  output [63:0] complement2;


  complementer_N64_2_DW01_sub_0 sub_add_31_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(\input ), .CI(1'b0), .DIFF(complement2) );
endmodule


module complementer_N64_1_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n190, n191, n192, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n237, n238, n239, n241, n242, n243, n245, n246, n247,
         n249, n250, n189, n193, n236, n240, n244, n248, n251;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U81 ( .A(n190), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U82 ( .A(n192), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U84 ( .A(n195), .B(B[63]), .Z(DIFF[63]) );
  XOR2_X1 U85 ( .A(n196), .B(B[62]), .Z(DIFF[62]) );
  XOR2_X1 U86 ( .A(n194), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U87 ( .A(n198), .B(B[59]), .Z(DIFF[59]) );
  XOR2_X1 U88 ( .A(n201), .B(B[58]), .Z(DIFF[58]) );
  XOR2_X1 U89 ( .A(n200), .B(B[57]), .Z(DIFF[57]) );
  XOR2_X1 U90 ( .A(n202), .B(B[55]), .Z(DIFF[55]) );
  XOR2_X1 U91 ( .A(n205), .B(B[54]), .Z(DIFF[54]) );
  XOR2_X1 U92 ( .A(n204), .B(B[53]), .Z(DIFF[53]) );
  XOR2_X1 U93 ( .A(n206), .B(B[51]), .Z(DIFF[51]) );
  XOR2_X1 U94 ( .A(n209), .B(B[50]), .Z(DIFF[50]) );
  XOR2_X1 U95 ( .A(n208), .B(B[49]), .Z(DIFF[49]) );
  XOR2_X1 U96 ( .A(n212), .B(B[47]), .Z(DIFF[47]) );
  XOR2_X1 U97 ( .A(n215), .B(B[46]), .Z(DIFF[46]) );
  XOR2_X1 U98 ( .A(n214), .B(B[45]), .Z(DIFF[45]) );
  XOR2_X1 U99 ( .A(n216), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U100 ( .A(n219), .B(B[42]), .Z(DIFF[42]) );
  XOR2_X1 U101 ( .A(n218), .B(B[41]), .Z(DIFF[41]) );
  XOR2_X1 U102 ( .A(n211), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U103 ( .A(n220), .B(B[39]), .Z(DIFF[39]) );
  XOR2_X1 U104 ( .A(n223), .B(B[38]), .Z(DIFF[38]) );
  XOR2_X1 U105 ( .A(n222), .B(B[37]), .Z(DIFF[37]) );
  XOR2_X1 U106 ( .A(n224), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U107 ( .A(n227), .B(B[34]), .Z(DIFF[34]) );
  XOR2_X1 U108 ( .A(n226), .B(B[33]), .Z(DIFF[33]) );
  XOR2_X1 U109 ( .A(n228), .B(B[31]), .Z(DIFF[31]) );
  XOR2_X1 U110 ( .A(n231), .B(B[30]), .Z(DIFF[30]) );
  XOR2_X1 U111 ( .A(n230), .B(B[29]), .Z(DIFF[29]) );
  XOR2_X1 U112 ( .A(n233), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U114 ( .A(n235), .B(B[25]), .Z(DIFF[25]) );
  XOR2_X1 U115 ( .A(n237), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U117 ( .A(n239), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U118 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U119 ( .A(n241), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U121 ( .A(n243), .B(B[17]), .Z(DIFF[17]) );
  XOR2_X1 U122 ( .A(n245), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U124 ( .A(n247), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U125 ( .A(n249), .B(B[11]), .Z(DIFF[11]) );
  OR2_X1 U1 ( .A1(n196), .A2(B[62]), .ZN(n195) );
  NAND2_X1 U2 ( .A1(n197), .A2(n251), .ZN(n196) );
  NOR3_X1 U3 ( .A1(B[59]), .A2(B[60]), .A3(n198), .ZN(n197) );
  NOR2_X1 U4 ( .A1(B[55]), .A2(n202), .ZN(n203) );
  NOR2_X1 U5 ( .A1(B[51]), .A2(n206), .ZN(n207) );
  NOR2_X1 U6 ( .A1(B[47]), .A2(n212), .ZN(n213) );
  NOR2_X1 U7 ( .A1(B[43]), .A2(n216), .ZN(n217) );
  NOR2_X1 U8 ( .A1(B[59]), .A2(n198), .ZN(n199) );
  OR3_X1 U9 ( .A1(B[57]), .A2(B[58]), .A3(n200), .ZN(n198) );
  OR3_X1 U10 ( .A1(B[53]), .A2(B[54]), .A3(n204), .ZN(n202) );
  OR3_X1 U11 ( .A1(B[49]), .A2(B[50]), .A3(n208), .ZN(n206) );
  OR3_X1 U12 ( .A1(B[45]), .A2(B[46]), .A3(n214), .ZN(n212) );
  OR3_X1 U13 ( .A1(B[41]), .A2(B[42]), .A3(n218), .ZN(n216) );
  OR3_X1 U14 ( .A1(B[55]), .A2(B[56]), .A3(n202), .ZN(n200) );
  OR3_X1 U15 ( .A1(B[51]), .A2(B[52]), .A3(n206), .ZN(n204) );
  OR3_X1 U16 ( .A1(B[47]), .A2(B[48]), .A3(n212), .ZN(n208) );
  OR3_X1 U17 ( .A1(B[43]), .A2(B[44]), .A3(n216), .ZN(n214) );
  OR2_X1 U18 ( .A1(n200), .A2(B[57]), .ZN(n201) );
  OR2_X1 U19 ( .A1(n204), .A2(B[53]), .ZN(n205) );
  OR2_X1 U20 ( .A1(n208), .A2(B[49]), .ZN(n209) );
  OR2_X1 U21 ( .A1(n214), .A2(B[45]), .ZN(n215) );
  OR2_X1 U22 ( .A1(n218), .A2(B[41]), .ZN(n219) );
  NOR2_X1 U23 ( .A1(B[39]), .A2(n220), .ZN(n221) );
  OR3_X1 U24 ( .A1(B[39]), .A2(B[40]), .A3(n220), .ZN(n218) );
  OR2_X1 U25 ( .A1(n222), .A2(B[37]), .ZN(n223) );
  OR3_X1 U26 ( .A1(B[37]), .A2(B[38]), .A3(n222), .ZN(n220) );
  NOR2_X1 U27 ( .A1(B[35]), .A2(n224), .ZN(n225) );
  OR3_X1 U28 ( .A1(B[35]), .A2(B[36]), .A3(n224), .ZN(n222) );
  XNOR2_X1 U29 ( .A(B[40]), .B(n221), .ZN(DIFF[40]) );
  XNOR2_X1 U30 ( .A(B[36]), .B(n225), .ZN(DIFF[36]) );
  XNOR2_X1 U31 ( .A(n197), .B(B[61]), .ZN(DIFF[61]) );
  XNOR2_X1 U32 ( .A(B[60]), .B(n199), .ZN(DIFF[60]) );
  XNOR2_X1 U33 ( .A(B[56]), .B(n203), .ZN(DIFF[56]) );
  XNOR2_X1 U34 ( .A(B[52]), .B(n207), .ZN(DIFF[52]) );
  XNOR2_X1 U35 ( .A(B[48]), .B(n213), .ZN(DIFF[48]) );
  XNOR2_X1 U36 ( .A(B[44]), .B(n217), .ZN(DIFF[44]) );
  OR3_X1 U37 ( .A1(B[33]), .A2(B[34]), .A3(n226), .ZN(n224) );
  XNOR2_X1 U38 ( .A(B[32]), .B(n229), .ZN(DIFF[32]) );
  OR2_X1 U39 ( .A1(n226), .A2(B[33]), .ZN(n227) );
  NOR2_X1 U40 ( .A1(B[31]), .A2(n228), .ZN(n229) );
  OR3_X1 U41 ( .A1(B[31]), .A2(B[32]), .A3(n228), .ZN(n226) );
  XNOR2_X1 U42 ( .A(n189), .B(B[22]), .ZN(DIFF[22]) );
  NOR2_X1 U43 ( .A1(n239), .A2(B[21]), .ZN(n189) );
  XNOR2_X1 U44 ( .A(n193), .B(B[26]), .ZN(DIFF[26]) );
  NOR2_X1 U45 ( .A1(n235), .A2(B[25]), .ZN(n193) );
  XNOR2_X1 U46 ( .A(n236), .B(B[18]), .ZN(DIFF[18]) );
  NOR2_X1 U47 ( .A1(n243), .A2(B[17]), .ZN(n236) );
  XNOR2_X1 U48 ( .A(n240), .B(B[14]), .ZN(DIFF[14]) );
  NOR2_X1 U49 ( .A1(n247), .A2(B[13]), .ZN(n240) );
  XNOR2_X1 U50 ( .A(n244), .B(B[10]), .ZN(DIFF[10]) );
  NOR2_X1 U51 ( .A1(n190), .A2(B[9]), .ZN(n244) );
  XNOR2_X1 U52 ( .A(n248), .B(B[6]), .ZN(DIFF[6]) );
  NOR2_X1 U53 ( .A1(n194), .A2(B[5]), .ZN(n248) );
  XNOR2_X1 U54 ( .A(B[28]), .B(n234), .ZN(DIFF[28]) );
  NOR2_X1 U55 ( .A1(B[27]), .A2(n233), .ZN(n234) );
  XNOR2_X1 U56 ( .A(B[24]), .B(n238), .ZN(DIFF[24]) );
  NOR2_X1 U57 ( .A1(B[23]), .A2(n237), .ZN(n238) );
  XNOR2_X1 U58 ( .A(B[20]), .B(n242), .ZN(DIFF[20]) );
  NOR2_X1 U59 ( .A1(B[19]), .A2(n241), .ZN(n242) );
  XNOR2_X1 U60 ( .A(B[16]), .B(n246), .ZN(DIFF[16]) );
  NOR2_X1 U61 ( .A1(B[15]), .A2(n245), .ZN(n246) );
  XNOR2_X1 U62 ( .A(B[12]), .B(n250), .ZN(DIFF[12]) );
  NOR2_X1 U63 ( .A1(B[11]), .A2(n249), .ZN(n250) );
  XNOR2_X1 U64 ( .A(B[8]), .B(n191), .ZN(DIFF[8]) );
  NOR2_X1 U65 ( .A1(B[7]), .A2(n192), .ZN(n191) );
  XNOR2_X1 U66 ( .A(B[2]), .B(n232), .ZN(DIFF[2]) );
  NOR2_X1 U67 ( .A1(\B[0] ), .A2(B[1]), .ZN(n232) );
  XNOR2_X1 U68 ( .A(B[4]), .B(n210), .ZN(DIFF[4]) );
  NOR2_X1 U69 ( .A1(B[3]), .A2(n211), .ZN(n210) );
  OR3_X1 U70 ( .A1(B[5]), .A2(B[6]), .A3(n194), .ZN(n192) );
  OR3_X1 U71 ( .A1(B[10]), .A2(B[9]), .A3(n190), .ZN(n249) );
  OR3_X1 U72 ( .A1(B[13]), .A2(B[14]), .A3(n247), .ZN(n245) );
  OR3_X1 U73 ( .A1(B[17]), .A2(B[18]), .A3(n243), .ZN(n241) );
  OR3_X1 U74 ( .A1(B[21]), .A2(B[22]), .A3(n239), .ZN(n237) );
  OR3_X1 U75 ( .A1(B[25]), .A2(B[26]), .A3(n235), .ZN(n233) );
  OR3_X1 U76 ( .A1(B[29]), .A2(B[30]), .A3(n230), .ZN(n228) );
  OR3_X1 U77 ( .A1(B[7]), .A2(B[8]), .A3(n192), .ZN(n190) );
  OR3_X1 U78 ( .A1(B[11]), .A2(B[12]), .A3(n249), .ZN(n247) );
  OR3_X1 U79 ( .A1(B[15]), .A2(B[16]), .A3(n245), .ZN(n243) );
  OR3_X1 U80 ( .A1(B[19]), .A2(B[20]), .A3(n241), .ZN(n239) );
  OR3_X1 U83 ( .A1(B[23]), .A2(B[24]), .A3(n237), .ZN(n235) );
  OR3_X1 U113 ( .A1(B[27]), .A2(B[28]), .A3(n233), .ZN(n230) );
  OR3_X1 U116 ( .A1(B[3]), .A2(B[4]), .A3(n211), .ZN(n194) );
  OR2_X1 U120 ( .A1(n230), .A2(B[29]), .ZN(n231) );
  OR3_X1 U123 ( .A1(B[1]), .A2(B[2]), .A3(\B[0] ), .ZN(n211) );
  INV_X1 U126 ( .A(B[61]), .ZN(n251) );
endmodule


module complementer_N64_1 ( \input , complement2 );
  input [63:0] \input ;
  output [63:0] complement2;


  complementer_N64_1_DW01_sub_0 sub_add_31_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(\input ), .CI(1'b0), .DIFF(complement2) );
endmodule


module ShiftnCompl_N64_1 ( plusA, plus2A_out, minus2A_out, plus4A_out, 
        minus4A_out );
  input [63:0] plusA;
  output [63:0] plus2A_out;
  output [63:0] minus2A_out;
  output [63:0] plus4A_out;
  output [63:0] minus4A_out;

  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign plus2A_out[0] = 1'b0;
  assign plus4A_out[0] = 1'b0;

  shifter_N64_2 shifter_1 ( .\input (plusA), .shiftLeftOnePos({
        plus2A_out[63:1], SYNOPSYS_UNCONNECTED__0}) );
  shifter_N64_1 shifter_2 ( .\input ({plus2A_out[63:1], 1'b0}), 
        .shiftLeftOnePos({plus4A_out[63:1], SYNOPSYS_UNCONNECTED__1}) );
  complementer_N64_2 complementer_1 ( .\input ({plus2A_out[63:1], 1'b0}), 
        .complement2(minus2A_out) );
  complementer_N64_1 complementer_2 ( .\input ({plus4A_out[63:1], 1'b0}), 
        .complement2(minus4A_out) );
endmodule


module MUX_GENERIC_N64_RADIX3_1 ( plusA, minusA, plus2A, minus2A, SEL, Y );
  input [63:0] plusA;
  input [63:0] minusA;
  input [63:0] plus2A;
  input [63:0] minus2A;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502;
  tri   [63:0] Y;

  TBUF_X1 \Y_tri[55]  ( .A(n446), .EN(n301), .Z(Y[55]) );
  TBUF_X1 \Y_tri[56]  ( .A(n445), .EN(n301), .Z(Y[56]) );
  TBUF_X1 \Y_tri[57]  ( .A(n444), .EN(n301), .Z(Y[57]) );
  TBUF_X1 \Y_tri[58]  ( .A(n443), .EN(n301), .Z(Y[58]) );
  TBUF_X1 \Y_tri[59]  ( .A(n442), .EN(n301), .Z(Y[59]) );
  TBUF_X1 \Y_tri[60]  ( .A(n441), .EN(n301), .Z(Y[60]) );
  TBUF_X1 \Y_tri[61]  ( .A(n440), .EN(n301), .Z(Y[61]) );
  TBUF_X1 \Y_tri[62]  ( .A(n439), .EN(n301), .Z(Y[62]) );
  TBUF_X1 \Y_tri[63]  ( .A(n438), .EN(n301), .Z(Y[63]) );
  TBUF_X1 \Y_tri[29]  ( .A(n472), .EN(n298), .Z(Y[29]) );
  TBUF_X1 \Y_tri[42]  ( .A(n459), .EN(n299), .Z(Y[42]) );
  TBUF_X1 \Y_tri[43]  ( .A(n458), .EN(n299), .Z(Y[43]) );
  TBUF_X1 \Y_tri[44]  ( .A(n457), .EN(n300), .Z(Y[44]) );
  TBUF_X1 \Y_tri[45]  ( .A(n456), .EN(n300), .Z(Y[45]) );
  TBUF_X1 \Y_tri[46]  ( .A(n455), .EN(n300), .Z(Y[46]) );
  TBUF_X1 \Y_tri[47]  ( .A(n454), .EN(n300), .Z(Y[47]) );
  TBUF_X1 \Y_tri[48]  ( .A(n453), .EN(n300), .Z(Y[48]) );
  TBUF_X1 \Y_tri[49]  ( .A(n452), .EN(n300), .Z(Y[49]) );
  TBUF_X1 \Y_tri[50]  ( .A(n451), .EN(n300), .Z(Y[50]) );
  TBUF_X1 \Y_tri[51]  ( .A(n450), .EN(n300), .Z(Y[51]) );
  TBUF_X1 \Y_tri[52]  ( .A(n449), .EN(n300), .Z(Y[52]) );
  TBUF_X1 \Y_tri[53]  ( .A(n448), .EN(n300), .Z(Y[53]) );
  TBUF_X1 \Y_tri[54]  ( .A(n447), .EN(n300), .Z(Y[54]) );
  TBUF_X1 \Y_tri[18]  ( .A(n483), .EN(n297), .Z(Y[18]) );
  TBUF_X1 \Y_tri[19]  ( .A(n482), .EN(n297), .Z(Y[19]) );
  TBUF_X1 \Y_tri[20]  ( .A(n481), .EN(n297), .Z(Y[20]) );
  TBUF_X1 \Y_tri[21]  ( .A(n480), .EN(n297), .Z(Y[21]) );
  TBUF_X1 \Y_tri[22]  ( .A(n479), .EN(n298), .Z(Y[22]) );
  TBUF_X1 \Y_tri[23]  ( .A(n478), .EN(n298), .Z(Y[23]) );
  TBUF_X1 \Y_tri[24]  ( .A(n477), .EN(n298), .Z(Y[24]) );
  TBUF_X1 \Y_tri[25]  ( .A(n476), .EN(n298), .Z(Y[25]) );
  TBUF_X1 \Y_tri[26]  ( .A(n475), .EN(n298), .Z(Y[26]) );
  TBUF_X1 \Y_tri[27]  ( .A(n474), .EN(n298), .Z(Y[27]) );
  TBUF_X1 \Y_tri[28]  ( .A(n473), .EN(n298), .Z(Y[28]) );
  TBUF_X1 \Y_tri[30]  ( .A(n471), .EN(n298), .Z(Y[30]) );
  TBUF_X1 \Y_tri[31]  ( .A(n470), .EN(n298), .Z(Y[31]) );
  TBUF_X1 \Y_tri[32]  ( .A(n469), .EN(n298), .Z(Y[32]) );
  TBUF_X1 \Y_tri[33]  ( .A(n468), .EN(n299), .Z(Y[33]) );
  TBUF_X1 \Y_tri[34]  ( .A(n467), .EN(n299), .Z(Y[34]) );
  TBUF_X1 \Y_tri[35]  ( .A(n466), .EN(n299), .Z(Y[35]) );
  TBUF_X1 \Y_tri[36]  ( .A(n465), .EN(n299), .Z(Y[36]) );
  TBUF_X1 \Y_tri[37]  ( .A(n464), .EN(n299), .Z(Y[37]) );
  TBUF_X1 \Y_tri[38]  ( .A(n463), .EN(n299), .Z(Y[38]) );
  TBUF_X1 \Y_tri[39]  ( .A(n462), .EN(n299), .Z(Y[39]) );
  TBUF_X1 \Y_tri[40]  ( .A(n461), .EN(n299), .Z(Y[40]) );
  TBUF_X1 \Y_tri[41]  ( .A(n460), .EN(n299), .Z(Y[41]) );
  TBUF_X1 \Y_tri[8]  ( .A(n494), .EN(n296), .Z(Y[8]) );
  TBUF_X1 \Y_tri[9]  ( .A(n492), .EN(n296), .Z(Y[9]) );
  TBUF_X1 \Y_tri[10]  ( .A(n491), .EN(n296), .Z(Y[10]) );
  TBUF_X1 \Y_tri[11]  ( .A(n490), .EN(n297), .Z(Y[11]) );
  TBUF_X1 \Y_tri[12]  ( .A(n489), .EN(n297), .Z(Y[12]) );
  TBUF_X1 \Y_tri[13]  ( .A(n488), .EN(n297), .Z(Y[13]) );
  TBUF_X1 \Y_tri[14]  ( .A(n487), .EN(n297), .Z(Y[14]) );
  TBUF_X1 \Y_tri[15]  ( .A(n486), .EN(n297), .Z(Y[15]) );
  TBUF_X1 \Y_tri[16]  ( .A(n485), .EN(n297), .Z(Y[16]) );
  TBUF_X1 \Y_tri[17]  ( .A(n484), .EN(n297), .Z(Y[17]) );
  TBUF_X1 \Y_tri[1]  ( .A(n501), .EN(n296), .Z(Y[1]) );
  TBUF_X1 \Y_tri[2]  ( .A(n500), .EN(n296), .Z(Y[2]) );
  TBUF_X1 \Y_tri[3]  ( .A(n499), .EN(n296), .Z(Y[3]) );
  TBUF_X1 \Y_tri[4]  ( .A(n498), .EN(n296), .Z(Y[4]) );
  TBUF_X1 \Y_tri[5]  ( .A(n497), .EN(n296), .Z(Y[5]) );
  TBUF_X1 \Y_tri[6]  ( .A(n496), .EN(n296), .Z(Y[6]) );
  TBUF_X1 \Y_tri[7]  ( .A(n495), .EN(n296), .Z(Y[7]) );
  TBUF_X1 \Y_tri[0]  ( .A(n502), .EN(n296), .Z(Y[0]) );
  NAND2_X1 U2 ( .A1(n385), .A2(n384), .ZN(n462) );
  AOI22_X1 U3 ( .A1(plusA[39]), .A2(n281), .B1(plus2A[39]), .B2(n275), .ZN(
        n385) );
  AOI22_X1 U4 ( .A1(minus2A[39]), .A2(n293), .B1(minusA[39]), .B2(n287), .ZN(
        n384) );
  NAND2_X1 U5 ( .A1(n377), .A2(n376), .ZN(n466) );
  AOI22_X1 U6 ( .A1(plusA[35]), .A2(n280), .B1(plus2A[35]), .B2(n274), .ZN(
        n377) );
  AOI22_X1 U7 ( .A1(minus2A[35]), .A2(n292), .B1(minusA[35]), .B2(n286), .ZN(
        n376) );
  NAND2_X1 U8 ( .A1(n389), .A2(n388), .ZN(n460) );
  AOI22_X1 U9 ( .A1(plusA[41]), .A2(n281), .B1(plus2A[41]), .B2(n275), .ZN(
        n389) );
  AOI22_X1 U10 ( .A1(minus2A[41]), .A2(n293), .B1(minusA[41]), .B2(n287), .ZN(
        n388) );
  NAND2_X1 U11 ( .A1(n381), .A2(n380), .ZN(n464) );
  AOI22_X1 U12 ( .A1(plusA[37]), .A2(n281), .B1(plus2A[37]), .B2(n275), .ZN(
        n381) );
  AOI22_X1 U13 ( .A1(minus2A[37]), .A2(n293), .B1(minusA[37]), .B2(n287), .ZN(
        n380) );
  NAND2_X1 U14 ( .A1(n387), .A2(n386), .ZN(n461) );
  AOI22_X1 U15 ( .A1(plusA[40]), .A2(n281), .B1(plus2A[40]), .B2(n275), .ZN(
        n387) );
  AOI22_X1 U16 ( .A1(minus2A[40]), .A2(n293), .B1(minusA[40]), .B2(n287), .ZN(
        n386) );
  NAND2_X1 U17 ( .A1(n379), .A2(n378), .ZN(n465) );
  AOI22_X1 U18 ( .A1(plusA[36]), .A2(n281), .B1(plus2A[36]), .B2(n275), .ZN(
        n379) );
  AOI22_X1 U19 ( .A1(minus2A[36]), .A2(n293), .B1(minusA[36]), .B2(n287), .ZN(
        n378) );
  NAND2_X1 U20 ( .A1(n383), .A2(n382), .ZN(n463) );
  AOI22_X1 U21 ( .A1(plusA[38]), .A2(n281), .B1(plus2A[38]), .B2(n275), .ZN(
        n383) );
  AOI22_X1 U22 ( .A1(minus2A[38]), .A2(n293), .B1(minusA[38]), .B2(n287), .ZN(
        n382) );
  NAND2_X1 U23 ( .A1(n375), .A2(n374), .ZN(n467) );
  AOI22_X1 U24 ( .A1(plusA[34]), .A2(n280), .B1(plus2A[34]), .B2(n274), .ZN(
        n375) );
  AOI22_X1 U25 ( .A1(minus2A[34]), .A2(n292), .B1(minusA[34]), .B2(n286), .ZN(
        n374) );
  NAND2_X1 U26 ( .A1(n417), .A2(n416), .ZN(n446) );
  AOI22_X1 U27 ( .A1(plusA[55]), .A2(n282), .B1(plus2A[55]), .B2(n276), .ZN(
        n417) );
  AOI22_X1 U28 ( .A1(minus2A[55]), .A2(n294), .B1(minusA[55]), .B2(n288), .ZN(
        n416) );
  NAND2_X1 U29 ( .A1(n437), .A2(n436), .ZN(n438) );
  AOI22_X1 U30 ( .A1(plusA[63]), .A2(n283), .B1(plus2A[63]), .B2(n277), .ZN(
        n437) );
  AOI22_X1 U31 ( .A1(minus2A[63]), .A2(n295), .B1(minusA[63]), .B2(n289), .ZN(
        n436) );
  NAND2_X1 U32 ( .A1(n431), .A2(n430), .ZN(n439) );
  AOI22_X1 U33 ( .A1(plusA[62]), .A2(n283), .B1(plus2A[62]), .B2(n277), .ZN(
        n431) );
  AOI22_X1 U34 ( .A1(minus2A[62]), .A2(n295), .B1(minusA[62]), .B2(n289), .ZN(
        n430) );
  NAND2_X1 U35 ( .A1(n429), .A2(n428), .ZN(n440) );
  AOI22_X1 U36 ( .A1(plusA[61]), .A2(n283), .B1(plus2A[61]), .B2(n277), .ZN(
        n429) );
  AOI22_X1 U37 ( .A1(minus2A[61]), .A2(n295), .B1(minusA[61]), .B2(n289), .ZN(
        n428) );
  NAND2_X1 U38 ( .A1(n409), .A2(n408), .ZN(n450) );
  AOI22_X1 U39 ( .A1(plusA[51]), .A2(n282), .B1(plus2A[51]), .B2(n276), .ZN(
        n409) );
  AOI22_X1 U40 ( .A1(minus2A[51]), .A2(n294), .B1(minusA[51]), .B2(n288), .ZN(
        n408) );
  NAND2_X1 U41 ( .A1(n401), .A2(n400), .ZN(n454) );
  AOI22_X1 U42 ( .A1(plusA[47]), .A2(n281), .B1(plus2A[47]), .B2(n275), .ZN(
        n401) );
  AOI22_X1 U43 ( .A1(minus2A[47]), .A2(n293), .B1(minusA[47]), .B2(n287), .ZN(
        n400) );
  NAND2_X1 U44 ( .A1(n393), .A2(n392), .ZN(n458) );
  AOI22_X1 U45 ( .A1(plusA[43]), .A2(n281), .B1(plus2A[43]), .B2(n275), .ZN(
        n393) );
  AOI22_X1 U46 ( .A1(minus2A[43]), .A2(n293), .B1(minusA[43]), .B2(n287), .ZN(
        n392) );
  NAND2_X1 U47 ( .A1(n425), .A2(n424), .ZN(n442) );
  AOI22_X1 U48 ( .A1(plusA[59]), .A2(n282), .B1(plus2A[59]), .B2(n276), .ZN(
        n425) );
  AOI22_X1 U49 ( .A1(minus2A[59]), .A2(n294), .B1(minusA[59]), .B2(n288), .ZN(
        n424) );
  NAND2_X1 U50 ( .A1(n421), .A2(n420), .ZN(n444) );
  AOI22_X1 U51 ( .A1(plusA[57]), .A2(n282), .B1(plus2A[57]), .B2(n276), .ZN(
        n421) );
  AOI22_X1 U52 ( .A1(minus2A[57]), .A2(n294), .B1(minusA[57]), .B2(n288), .ZN(
        n420) );
  NAND2_X1 U53 ( .A1(n413), .A2(n412), .ZN(n448) );
  AOI22_X1 U54 ( .A1(plusA[53]), .A2(n282), .B1(plus2A[53]), .B2(n276), .ZN(
        n413) );
  AOI22_X1 U55 ( .A1(minus2A[53]), .A2(n294), .B1(minusA[53]), .B2(n288), .ZN(
        n412) );
  NAND2_X1 U56 ( .A1(n405), .A2(n404), .ZN(n452) );
  AOI22_X1 U57 ( .A1(plusA[49]), .A2(n282), .B1(plus2A[49]), .B2(n276), .ZN(
        n405) );
  AOI22_X1 U58 ( .A1(minus2A[49]), .A2(n294), .B1(minusA[49]), .B2(n288), .ZN(
        n404) );
  NAND2_X1 U59 ( .A1(n397), .A2(n396), .ZN(n456) );
  AOI22_X1 U60 ( .A1(plusA[45]), .A2(n281), .B1(plus2A[45]), .B2(n275), .ZN(
        n397) );
  AOI22_X1 U61 ( .A1(minus2A[45]), .A2(n293), .B1(minusA[45]), .B2(n287), .ZN(
        n396) );
  NAND2_X1 U62 ( .A1(n427), .A2(n426), .ZN(n441) );
  AOI22_X1 U63 ( .A1(plusA[60]), .A2(n283), .B1(plus2A[60]), .B2(n277), .ZN(
        n427) );
  AOI22_X1 U64 ( .A1(minus2A[60]), .A2(n295), .B1(minusA[60]), .B2(n289), .ZN(
        n426) );
  NAND2_X1 U65 ( .A1(n419), .A2(n418), .ZN(n445) );
  AOI22_X1 U66 ( .A1(plusA[56]), .A2(n282), .B1(plus2A[56]), .B2(n276), .ZN(
        n419) );
  AOI22_X1 U67 ( .A1(minus2A[56]), .A2(n294), .B1(minusA[56]), .B2(n288), .ZN(
        n418) );
  NAND2_X1 U68 ( .A1(n411), .A2(n410), .ZN(n449) );
  AOI22_X1 U69 ( .A1(plusA[52]), .A2(n282), .B1(plus2A[52]), .B2(n276), .ZN(
        n411) );
  AOI22_X1 U70 ( .A1(minus2A[52]), .A2(n294), .B1(minusA[52]), .B2(n288), .ZN(
        n410) );
  NAND2_X1 U71 ( .A1(n403), .A2(n402), .ZN(n453) );
  AOI22_X1 U72 ( .A1(plusA[48]), .A2(n282), .B1(plus2A[48]), .B2(n276), .ZN(
        n403) );
  AOI22_X1 U73 ( .A1(minus2A[48]), .A2(n294), .B1(minusA[48]), .B2(n288), .ZN(
        n402) );
  NAND2_X1 U74 ( .A1(n395), .A2(n394), .ZN(n457) );
  AOI22_X1 U75 ( .A1(plusA[44]), .A2(n281), .B1(plus2A[44]), .B2(n275), .ZN(
        n395) );
  AOI22_X1 U76 ( .A1(minus2A[44]), .A2(n293), .B1(minusA[44]), .B2(n287), .ZN(
        n394) );
  NAND2_X1 U77 ( .A1(n423), .A2(n422), .ZN(n443) );
  AOI22_X1 U78 ( .A1(plusA[58]), .A2(n282), .B1(plus2A[58]), .B2(n276), .ZN(
        n423) );
  AOI22_X1 U79 ( .A1(minus2A[58]), .A2(n294), .B1(minusA[58]), .B2(n288), .ZN(
        n422) );
  NAND2_X1 U80 ( .A1(n415), .A2(n414), .ZN(n447) );
  AOI22_X1 U81 ( .A1(plusA[54]), .A2(n282), .B1(plus2A[54]), .B2(n276), .ZN(
        n415) );
  AOI22_X1 U82 ( .A1(minus2A[54]), .A2(n294), .B1(minusA[54]), .B2(n288), .ZN(
        n414) );
  NAND2_X1 U83 ( .A1(n407), .A2(n406), .ZN(n451) );
  AOI22_X1 U84 ( .A1(plusA[50]), .A2(n282), .B1(plus2A[50]), .B2(n276), .ZN(
        n407) );
  AOI22_X1 U85 ( .A1(minus2A[50]), .A2(n294), .B1(minusA[50]), .B2(n288), .ZN(
        n406) );
  NAND2_X1 U86 ( .A1(n399), .A2(n398), .ZN(n455) );
  AOI22_X1 U87 ( .A1(plusA[46]), .A2(n281), .B1(plus2A[46]), .B2(n275), .ZN(
        n399) );
  AOI22_X1 U88 ( .A1(minus2A[46]), .A2(n293), .B1(minusA[46]), .B2(n287), .ZN(
        n398) );
  NAND2_X1 U89 ( .A1(n391), .A2(n390), .ZN(n459) );
  AOI22_X1 U90 ( .A1(plusA[42]), .A2(n281), .B1(plus2A[42]), .B2(n275), .ZN(
        n391) );
  AOI22_X1 U91 ( .A1(minus2A[42]), .A2(n293), .B1(minusA[42]), .B2(n287), .ZN(
        n390) );
  BUF_X1 U92 ( .A(n493), .Z(n296) );
  BUF_X1 U93 ( .A(n493), .Z(n297) );
  BUF_X1 U94 ( .A(n493), .Z(n298) );
  NAND2_X1 U95 ( .A1(n373), .A2(n372), .ZN(n468) );
  AOI22_X1 U96 ( .A1(plusA[33]), .A2(n280), .B1(plus2A[33]), .B2(n274), .ZN(
        n373) );
  AOI22_X1 U97 ( .A1(minus2A[33]), .A2(n292), .B1(minusA[33]), .B2(n286), .ZN(
        n372) );
  NAND2_X1 U98 ( .A1(n371), .A2(n370), .ZN(n469) );
  AOI22_X1 U99 ( .A1(plusA[32]), .A2(n280), .B1(plus2A[32]), .B2(n274), .ZN(
        n371) );
  AOI22_X1 U100 ( .A1(minus2A[32]), .A2(n292), .B1(minusA[32]), .B2(n286), 
        .ZN(n370) );
  BUF_X1 U101 ( .A(n433), .Z(n281) );
  BUF_X1 U102 ( .A(n433), .Z(n280) );
  BUF_X1 U103 ( .A(n435), .Z(n293) );
  BUF_X1 U104 ( .A(n435), .Z(n292) );
  BUF_X1 U105 ( .A(n434), .Z(n287) );
  BUF_X1 U106 ( .A(n432), .Z(n275) );
  BUF_X1 U107 ( .A(n434), .Z(n286) );
  BUF_X1 U108 ( .A(n432), .Z(n274) );
  BUF_X1 U109 ( .A(n493), .Z(n299) );
  BUF_X1 U110 ( .A(n433), .Z(n282) );
  BUF_X1 U111 ( .A(n435), .Z(n294) );
  BUF_X1 U112 ( .A(n434), .Z(n288) );
  BUF_X1 U113 ( .A(n432), .Z(n276) );
  BUF_X1 U114 ( .A(n493), .Z(n300) );
  BUF_X1 U115 ( .A(n493), .Z(n301) );
  BUF_X1 U116 ( .A(n433), .Z(n279) );
  BUF_X1 U117 ( .A(n433), .Z(n278) );
  BUF_X1 U118 ( .A(n435), .Z(n291) );
  BUF_X1 U119 ( .A(n435), .Z(n290) );
  BUF_X1 U120 ( .A(n434), .Z(n285) );
  BUF_X1 U121 ( .A(n432), .Z(n273) );
  BUF_X1 U122 ( .A(n434), .Z(n284) );
  BUF_X1 U123 ( .A(n432), .Z(n272) );
  NOR2_X1 U124 ( .A1(n323), .A2(n304), .ZN(n493) );
  INV_X1 U125 ( .A(SEL[2]), .ZN(n304) );
  NOR2_X1 U126 ( .A1(SEL[1]), .A2(SEL[0]), .ZN(n323) );
  NAND2_X1 U127 ( .A1(n369), .A2(n368), .ZN(n470) );
  AOI22_X1 U128 ( .A1(plusA[31]), .A2(n280), .B1(plus2A[31]), .B2(n274), .ZN(
        n369) );
  AOI22_X1 U129 ( .A1(minus2A[31]), .A2(n292), .B1(minusA[31]), .B2(n286), 
        .ZN(n368) );
  NOR3_X1 U130 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n302), .ZN(n434) );
  NOR3_X1 U131 ( .A1(SEL[1]), .A2(SEL[2]), .A3(n303), .ZN(n433) );
  NOR3_X1 U132 ( .A1(n302), .A2(SEL[2]), .A3(n303), .ZN(n432) );
  AND2_X1 U133 ( .A1(SEL[2]), .A2(n323), .ZN(n435) );
  INV_X1 U134 ( .A(SEL[1]), .ZN(n302) );
  INV_X1 U135 ( .A(SEL[0]), .ZN(n303) );
  NAND2_X1 U136 ( .A1(n367), .A2(n366), .ZN(n471) );
  AOI22_X1 U137 ( .A1(plusA[30]), .A2(n280), .B1(plus2A[30]), .B2(n274), .ZN(
        n367) );
  AOI22_X1 U138 ( .A1(minus2A[30]), .A2(n292), .B1(minusA[30]), .B2(n286), 
        .ZN(n366) );
  NAND2_X1 U139 ( .A1(n365), .A2(n364), .ZN(n472) );
  AOI22_X1 U140 ( .A1(plusA[29]), .A2(n280), .B1(plus2A[29]), .B2(n274), .ZN(
        n365) );
  AOI22_X1 U141 ( .A1(minus2A[29]), .A2(n292), .B1(minusA[29]), .B2(n286), 
        .ZN(n364) );
  NAND2_X1 U142 ( .A1(n361), .A2(n360), .ZN(n474) );
  AOI22_X1 U143 ( .A1(plusA[27]), .A2(n280), .B1(plus2A[27]), .B2(n274), .ZN(
        n361) );
  AOI22_X1 U144 ( .A1(minus2A[27]), .A2(n292), .B1(minusA[27]), .B2(n286), 
        .ZN(n360) );
  NAND2_X1 U145 ( .A1(n359), .A2(n358), .ZN(n475) );
  AOI22_X1 U146 ( .A1(plusA[26]), .A2(n280), .B1(plus2A[26]), .B2(n274), .ZN(
        n359) );
  AOI22_X1 U147 ( .A1(minus2A[26]), .A2(n292), .B1(minusA[26]), .B2(n286), 
        .ZN(n358) );
  NAND2_X1 U148 ( .A1(n357), .A2(n356), .ZN(n476) );
  AOI22_X1 U149 ( .A1(plusA[25]), .A2(n280), .B1(plus2A[25]), .B2(n274), .ZN(
        n357) );
  AOI22_X1 U150 ( .A1(minus2A[25]), .A2(n292), .B1(minusA[25]), .B2(n286), 
        .ZN(n356) );
  NAND2_X1 U151 ( .A1(n353), .A2(n352), .ZN(n478) );
  AOI22_X1 U152 ( .A1(plusA[23]), .A2(n279), .B1(plus2A[23]), .B2(n273), .ZN(
        n353) );
  AOI22_X1 U153 ( .A1(minus2A[23]), .A2(n291), .B1(minusA[23]), .B2(n285), 
        .ZN(n352) );
  NAND2_X1 U154 ( .A1(n351), .A2(n350), .ZN(n479) );
  AOI22_X1 U155 ( .A1(plusA[22]), .A2(n279), .B1(plus2A[22]), .B2(n273), .ZN(
        n351) );
  AOI22_X1 U156 ( .A1(minus2A[22]), .A2(n291), .B1(minusA[22]), .B2(n285), 
        .ZN(n350) );
  NAND2_X1 U157 ( .A1(n349), .A2(n348), .ZN(n480) );
  AOI22_X1 U158 ( .A1(plusA[21]), .A2(n279), .B1(plus2A[21]), .B2(n273), .ZN(
        n349) );
  AOI22_X1 U159 ( .A1(minus2A[21]), .A2(n291), .B1(minusA[21]), .B2(n285), 
        .ZN(n348) );
  NAND2_X1 U160 ( .A1(n345), .A2(n344), .ZN(n482) );
  AOI22_X1 U161 ( .A1(plusA[19]), .A2(n279), .B1(plus2A[19]), .B2(n273), .ZN(
        n345) );
  AOI22_X1 U162 ( .A1(minus2A[19]), .A2(n291), .B1(minusA[19]), .B2(n285), 
        .ZN(n344) );
  NAND2_X1 U163 ( .A1(n343), .A2(n342), .ZN(n483) );
  AOI22_X1 U164 ( .A1(plusA[18]), .A2(n279), .B1(plus2A[18]), .B2(n273), .ZN(
        n343) );
  AOI22_X1 U165 ( .A1(minus2A[18]), .A2(n291), .B1(minusA[18]), .B2(n285), 
        .ZN(n342) );
  NAND2_X1 U166 ( .A1(n341), .A2(n340), .ZN(n484) );
  AOI22_X1 U167 ( .A1(plusA[17]), .A2(n279), .B1(plus2A[17]), .B2(n273), .ZN(
        n341) );
  AOI22_X1 U168 ( .A1(minus2A[17]), .A2(n291), .B1(minusA[17]), .B2(n285), 
        .ZN(n340) );
  NAND2_X1 U169 ( .A1(n337), .A2(n336), .ZN(n486) );
  AOI22_X1 U170 ( .A1(plusA[15]), .A2(n279), .B1(plus2A[15]), .B2(n273), .ZN(
        n337) );
  AOI22_X1 U171 ( .A1(minus2A[15]), .A2(n291), .B1(minusA[15]), .B2(n285), 
        .ZN(n336) );
  NAND2_X1 U172 ( .A1(n335), .A2(n334), .ZN(n487) );
  AOI22_X1 U173 ( .A1(plusA[14]), .A2(n279), .B1(plus2A[14]), .B2(n273), .ZN(
        n335) );
  AOI22_X1 U174 ( .A1(minus2A[14]), .A2(n291), .B1(minusA[14]), .B2(n285), 
        .ZN(n334) );
  NAND2_X1 U175 ( .A1(n333), .A2(n332), .ZN(n488) );
  AOI22_X1 U176 ( .A1(plusA[13]), .A2(n279), .B1(plus2A[13]), .B2(n273), .ZN(
        n333) );
  AOI22_X1 U177 ( .A1(minus2A[13]), .A2(n291), .B1(minusA[13]), .B2(n285), 
        .ZN(n332) );
  NAND2_X1 U178 ( .A1(n329), .A2(n328), .ZN(n490) );
  AOI22_X1 U179 ( .A1(plusA[11]), .A2(n278), .B1(plus2A[11]), .B2(n272), .ZN(
        n329) );
  AOI22_X1 U180 ( .A1(minus2A[11]), .A2(n290), .B1(minusA[11]), .B2(n284), 
        .ZN(n328) );
  NAND2_X1 U181 ( .A1(n327), .A2(n326), .ZN(n491) );
  AOI22_X1 U182 ( .A1(plusA[10]), .A2(n278), .B1(plus2A[10]), .B2(n272), .ZN(
        n327) );
  AOI22_X1 U183 ( .A1(minus2A[10]), .A2(n290), .B1(minusA[10]), .B2(n284), 
        .ZN(n326) );
  NAND2_X1 U184 ( .A1(n325), .A2(n324), .ZN(n492) );
  AOI22_X1 U185 ( .A1(plusA[9]), .A2(n278), .B1(plus2A[9]), .B2(n272), .ZN(
        n325) );
  AOI22_X1 U186 ( .A1(minus2A[9]), .A2(n290), .B1(minusA[9]), .B2(n284), .ZN(
        n324) );
  NAND2_X1 U187 ( .A1(n320), .A2(n319), .ZN(n495) );
  AOI22_X1 U188 ( .A1(plusA[7]), .A2(n278), .B1(plus2A[7]), .B2(n272), .ZN(
        n320) );
  AOI22_X1 U189 ( .A1(minus2A[7]), .A2(n290), .B1(minusA[7]), .B2(n284), .ZN(
        n319) );
  NAND2_X1 U190 ( .A1(n318), .A2(n317), .ZN(n496) );
  AOI22_X1 U191 ( .A1(plusA[6]), .A2(n278), .B1(plus2A[6]), .B2(n272), .ZN(
        n318) );
  AOI22_X1 U192 ( .A1(minus2A[6]), .A2(n290), .B1(minusA[6]), .B2(n284), .ZN(
        n317) );
  NAND2_X1 U193 ( .A1(n316), .A2(n315), .ZN(n497) );
  AOI22_X1 U194 ( .A1(plusA[5]), .A2(n278), .B1(plus2A[5]), .B2(n272), .ZN(
        n316) );
  AOI22_X1 U195 ( .A1(minus2A[5]), .A2(n290), .B1(minusA[5]), .B2(n284), .ZN(
        n315) );
  NAND2_X1 U196 ( .A1(n312), .A2(n311), .ZN(n499) );
  AOI22_X1 U197 ( .A1(plusA[3]), .A2(n278), .B1(plus2A[3]), .B2(n272), .ZN(
        n312) );
  AOI22_X1 U198 ( .A1(minus2A[3]), .A2(n290), .B1(minusA[3]), .B2(n284), .ZN(
        n311) );
  NAND2_X1 U199 ( .A1(n363), .A2(n362), .ZN(n473) );
  AOI22_X1 U200 ( .A1(plusA[28]), .A2(n280), .B1(plus2A[28]), .B2(n274), .ZN(
        n363) );
  AOI22_X1 U201 ( .A1(minus2A[28]), .A2(n292), .B1(minusA[28]), .B2(n286), 
        .ZN(n362) );
  NAND2_X1 U202 ( .A1(n355), .A2(n354), .ZN(n477) );
  AOI22_X1 U203 ( .A1(plusA[24]), .A2(n280), .B1(plus2A[24]), .B2(n274), .ZN(
        n355) );
  AOI22_X1 U204 ( .A1(minus2A[24]), .A2(n292), .B1(minusA[24]), .B2(n286), 
        .ZN(n354) );
  NAND2_X1 U205 ( .A1(n347), .A2(n346), .ZN(n481) );
  AOI22_X1 U206 ( .A1(plusA[20]), .A2(n279), .B1(plus2A[20]), .B2(n273), .ZN(
        n347) );
  AOI22_X1 U207 ( .A1(minus2A[20]), .A2(n291), .B1(minusA[20]), .B2(n285), 
        .ZN(n346) );
  NAND2_X1 U208 ( .A1(n339), .A2(n338), .ZN(n485) );
  AOI22_X1 U209 ( .A1(plusA[16]), .A2(n279), .B1(plus2A[16]), .B2(n273), .ZN(
        n339) );
  AOI22_X1 U210 ( .A1(minus2A[16]), .A2(n291), .B1(minusA[16]), .B2(n285), 
        .ZN(n338) );
  NAND2_X1 U211 ( .A1(n331), .A2(n330), .ZN(n489) );
  AOI22_X1 U212 ( .A1(plusA[12]), .A2(n279), .B1(plus2A[12]), .B2(n273), .ZN(
        n331) );
  AOI22_X1 U213 ( .A1(minus2A[12]), .A2(n291), .B1(minusA[12]), .B2(n285), 
        .ZN(n330) );
  NAND2_X1 U214 ( .A1(n322), .A2(n321), .ZN(n494) );
  AOI22_X1 U215 ( .A1(plusA[8]), .A2(n278), .B1(plus2A[8]), .B2(n272), .ZN(
        n322) );
  AOI22_X1 U216 ( .A1(minus2A[8]), .A2(n290), .B1(minusA[8]), .B2(n284), .ZN(
        n321) );
  NAND2_X1 U217 ( .A1(n314), .A2(n313), .ZN(n498) );
  AOI22_X1 U218 ( .A1(plusA[4]), .A2(n278), .B1(plus2A[4]), .B2(n272), .ZN(
        n314) );
  AOI22_X1 U219 ( .A1(minus2A[4]), .A2(n290), .B1(minusA[4]), .B2(n284), .ZN(
        n313) );
  NAND2_X1 U220 ( .A1(n310), .A2(n309), .ZN(n500) );
  AOI22_X1 U221 ( .A1(plusA[2]), .A2(n278), .B1(plus2A[2]), .B2(n272), .ZN(
        n310) );
  AOI22_X1 U222 ( .A1(minus2A[2]), .A2(n290), .B1(minusA[2]), .B2(n284), .ZN(
        n309) );
  NAND2_X1 U223 ( .A1(n308), .A2(n307), .ZN(n501) );
  AOI22_X1 U224 ( .A1(plusA[1]), .A2(n278), .B1(plus2A[1]), .B2(n272), .ZN(
        n308) );
  AOI22_X1 U225 ( .A1(minus2A[1]), .A2(n290), .B1(minusA[1]), .B2(n284), .ZN(
        n307) );
  NAND2_X1 U226 ( .A1(n306), .A2(n305), .ZN(n502) );
  AOI22_X1 U227 ( .A1(plusA[0]), .A2(n278), .B1(plus2A[0]), .B2(n272), .ZN(
        n306) );
  AOI22_X1 U228 ( .A1(minus2A[0]), .A2(n290), .B1(minusA[0]), .B2(n284), .ZN(
        n305) );
  CLKBUF_X1 U229 ( .A(n432), .Z(n277) );
  CLKBUF_X1 U230 ( .A(n433), .Z(n283) );
  CLKBUF_X1 U231 ( .A(n434), .Z(n289) );
  CLKBUF_X1 U232 ( .A(n435), .Z(n295) );
endmodule


module FA_64 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_63 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_62 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_61 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_60 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_59 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_58 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_57 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_56 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_55 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_54 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_53 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n6, n7;
  tri   A;

  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  XNOR2_X1 U1 ( .A(Ci), .B(n4), .ZN(S) );
  INV_X1 U2 ( .A(n6), .ZN(n4) );
  INV_X1 U3 ( .A(n7), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n7) );
endmodule


module FA_52 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_51 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_50 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_49 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_48 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_47 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_46 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_45 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_44 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_43 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_42 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_41 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_40 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_39 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_38 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_37 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_36 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_35 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_34 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_33 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_32 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_31 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_30 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_29 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_28 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_27 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_26 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_25 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_24 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_23 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_22 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_21 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_20 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_19 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_18 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_17 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_16 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_15 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_14 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_13 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_12 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_11 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_10 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_9 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_8 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_7 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_6 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_5 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_4 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
  INV_X1 U2 ( .A(n6), .ZN(Co) );
endmodule


module FA_3 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n5), .ZN(n6) );
endmodule


module FA_2 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module FA_1 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5, n6;
  tri   A;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n6), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n6) );
endmodule


module RCA_N64_1 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Ci;
  output Co;

  wire   [63:1] CTMP;
  tri   [63:0] A;

  FA_64 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_63 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_62 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_61 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(CTMP[4]) );
  FA_60 FAI_5 ( .A(A[4]), .B(B[4]), .Ci(CTMP[4]), .S(S[4]), .Co(CTMP[5]) );
  FA_59 FAI_6 ( .A(A[5]), .B(B[5]), .Ci(CTMP[5]), .S(S[5]), .Co(CTMP[6]) );
  FA_58 FAI_7 ( .A(A[6]), .B(B[6]), .Ci(CTMP[6]), .S(S[6]), .Co(CTMP[7]) );
  FA_57 FAI_8 ( .A(A[7]), .B(B[7]), .Ci(CTMP[7]), .S(S[7]), .Co(CTMP[8]) );
  FA_56 FAI_9 ( .A(A[8]), .B(B[8]), .Ci(CTMP[8]), .S(S[8]), .Co(CTMP[9]) );
  FA_55 FAI_10 ( .A(A[9]), .B(B[9]), .Ci(CTMP[9]), .S(S[9]), .Co(CTMP[10]) );
  FA_54 FAI_11 ( .A(A[10]), .B(B[10]), .Ci(CTMP[10]), .S(S[10]), .Co(CTMP[11])
         );
  FA_53 FAI_12 ( .A(A[11]), .B(B[11]), .Ci(CTMP[11]), .S(S[11]), .Co(CTMP[12])
         );
  FA_52 FAI_13 ( .A(A[12]), .B(B[12]), .Ci(CTMP[12]), .S(S[12]), .Co(CTMP[13])
         );
  FA_51 FAI_14 ( .A(A[13]), .B(B[13]), .Ci(CTMP[13]), .S(S[13]), .Co(CTMP[14])
         );
  FA_50 FAI_15 ( .A(A[14]), .B(B[14]), .Ci(CTMP[14]), .S(S[14]), .Co(CTMP[15])
         );
  FA_49 FAI_16 ( .A(A[15]), .B(B[15]), .Ci(CTMP[15]), .S(S[15]), .Co(CTMP[16])
         );
  FA_48 FAI_17 ( .A(A[16]), .B(B[16]), .Ci(CTMP[16]), .S(S[16]), .Co(CTMP[17])
         );
  FA_47 FAI_18 ( .A(A[17]), .B(B[17]), .Ci(CTMP[17]), .S(S[17]), .Co(CTMP[18])
         );
  FA_46 FAI_19 ( .A(A[18]), .B(B[18]), .Ci(CTMP[18]), .S(S[18]), .Co(CTMP[19])
         );
  FA_45 FAI_20 ( .A(A[19]), .B(B[19]), .Ci(CTMP[19]), .S(S[19]), .Co(CTMP[20])
         );
  FA_44 FAI_21 ( .A(A[20]), .B(B[20]), .Ci(CTMP[20]), .S(S[20]), .Co(CTMP[21])
         );
  FA_43 FAI_22 ( .A(A[21]), .B(B[21]), .Ci(CTMP[21]), .S(S[21]), .Co(CTMP[22])
         );
  FA_42 FAI_23 ( .A(A[22]), .B(B[22]), .Ci(CTMP[22]), .S(S[22]), .Co(CTMP[23])
         );
  FA_41 FAI_24 ( .A(A[23]), .B(B[23]), .Ci(CTMP[23]), .S(S[23]), .Co(CTMP[24])
         );
  FA_40 FAI_25 ( .A(A[24]), .B(B[24]), .Ci(CTMP[24]), .S(S[24]), .Co(CTMP[25])
         );
  FA_39 FAI_26 ( .A(A[25]), .B(B[25]), .Ci(CTMP[25]), .S(S[25]), .Co(CTMP[26])
         );
  FA_38 FAI_27 ( .A(A[26]), .B(B[26]), .Ci(CTMP[26]), .S(S[26]), .Co(CTMP[27])
         );
  FA_37 FAI_28 ( .A(A[27]), .B(B[27]), .Ci(CTMP[27]), .S(S[27]), .Co(CTMP[28])
         );
  FA_36 FAI_29 ( .A(A[28]), .B(B[28]), .Ci(CTMP[28]), .S(S[28]), .Co(CTMP[29])
         );
  FA_35 FAI_30 ( .A(A[29]), .B(B[29]), .Ci(CTMP[29]), .S(S[29]), .Co(CTMP[30])
         );
  FA_34 FAI_31 ( .A(A[30]), .B(B[30]), .Ci(CTMP[30]), .S(S[30]), .Co(CTMP[31])
         );
  FA_33 FAI_32 ( .A(A[31]), .B(B[31]), .Ci(CTMP[31]), .S(S[31]), .Co(CTMP[32])
         );
  FA_32 FAI_33 ( .A(A[32]), .B(B[32]), .Ci(CTMP[32]), .S(S[32]), .Co(CTMP[33])
         );
  FA_31 FAI_34 ( .A(A[33]), .B(B[33]), .Ci(CTMP[33]), .S(S[33]), .Co(CTMP[34])
         );
  FA_30 FAI_35 ( .A(A[34]), .B(B[34]), .Ci(CTMP[34]), .S(S[34]), .Co(CTMP[35])
         );
  FA_29 FAI_36 ( .A(A[35]), .B(B[35]), .Ci(CTMP[35]), .S(S[35]), .Co(CTMP[36])
         );
  FA_28 FAI_37 ( .A(A[36]), .B(B[36]), .Ci(CTMP[36]), .S(S[36]), .Co(CTMP[37])
         );
  FA_27 FAI_38 ( .A(A[37]), .B(B[37]), .Ci(CTMP[37]), .S(S[37]), .Co(CTMP[38])
         );
  FA_26 FAI_39 ( .A(A[38]), .B(B[38]), .Ci(CTMP[38]), .S(S[38]), .Co(CTMP[39])
         );
  FA_25 FAI_40 ( .A(A[39]), .B(B[39]), .Ci(CTMP[39]), .S(S[39]), .Co(CTMP[40])
         );
  FA_24 FAI_41 ( .A(A[40]), .B(B[40]), .Ci(CTMP[40]), .S(S[40]), .Co(CTMP[41])
         );
  FA_23 FAI_42 ( .A(A[41]), .B(B[41]), .Ci(CTMP[41]), .S(S[41]), .Co(CTMP[42])
         );
  FA_22 FAI_43 ( .A(A[42]), .B(B[42]), .Ci(CTMP[42]), .S(S[42]), .Co(CTMP[43])
         );
  FA_21 FAI_44 ( .A(A[43]), .B(B[43]), .Ci(CTMP[43]), .S(S[43]), .Co(CTMP[44])
         );
  FA_20 FAI_45 ( .A(A[44]), .B(B[44]), .Ci(CTMP[44]), .S(S[44]), .Co(CTMP[45])
         );
  FA_19 FAI_46 ( .A(A[45]), .B(B[45]), .Ci(CTMP[45]), .S(S[45]), .Co(CTMP[46])
         );
  FA_18 FAI_47 ( .A(A[46]), .B(B[46]), .Ci(CTMP[46]), .S(S[46]), .Co(CTMP[47])
         );
  FA_17 FAI_48 ( .A(A[47]), .B(B[47]), .Ci(CTMP[47]), .S(S[47]), .Co(CTMP[48])
         );
  FA_16 FAI_49 ( .A(A[48]), .B(B[48]), .Ci(CTMP[48]), .S(S[48]), .Co(CTMP[49])
         );
  FA_15 FAI_50 ( .A(A[49]), .B(B[49]), .Ci(CTMP[49]), .S(S[49]), .Co(CTMP[50])
         );
  FA_14 FAI_51 ( .A(A[50]), .B(B[50]), .Ci(CTMP[50]), .S(S[50]), .Co(CTMP[51])
         );
  FA_13 FAI_52 ( .A(A[51]), .B(B[51]), .Ci(CTMP[51]), .S(S[51]), .Co(CTMP[52])
         );
  FA_12 FAI_53 ( .A(A[52]), .B(B[52]), .Ci(CTMP[52]), .S(S[52]), .Co(CTMP[53])
         );
  FA_11 FAI_54 ( .A(A[53]), .B(B[53]), .Ci(CTMP[53]), .S(S[53]), .Co(CTMP[54])
         );
  FA_10 FAI_55 ( .A(A[54]), .B(B[54]), .Ci(CTMP[54]), .S(S[54]), .Co(CTMP[55])
         );
  FA_9 FAI_56 ( .A(A[55]), .B(B[55]), .Ci(CTMP[55]), .S(S[55]), .Co(CTMP[56])
         );
  FA_8 FAI_57 ( .A(A[56]), .B(B[56]), .Ci(CTMP[56]), .S(S[56]), .Co(CTMP[57])
         );
  FA_7 FAI_58 ( .A(A[57]), .B(B[57]), .Ci(CTMP[57]), .S(S[57]), .Co(CTMP[58])
         );
  FA_6 FAI_59 ( .A(A[58]), .B(B[58]), .Ci(CTMP[58]), .S(S[58]), .Co(CTMP[59])
         );
  FA_5 FAI_60 ( .A(A[59]), .B(B[59]), .Ci(CTMP[59]), .S(S[59]), .Co(CTMP[60])
         );
  FA_4 FAI_61 ( .A(A[60]), .B(B[60]), .Ci(CTMP[60]), .S(S[60]), .Co(CTMP[61])
         );
  FA_3 FAI_62 ( .A(A[61]), .B(B[61]), .Ci(CTMP[61]), .S(S[61]), .Co(CTMP[62])
         );
  FA_2 FAI_63 ( .A(A[62]), .B(B[62]), .Ci(CTMP[62]), .S(S[62]), .Co(CTMP[63])
         );
  FA_1 FAI_64 ( .A(A[63]), .B(B[63]), .Ci(CTMP[63]), .S(S[63]), .Co(Co) );
endmodule


module booth_mul_row_N64_RADIX3_1 ( prevA, prevSum, encoderIn, nextA, nextSum
 );
  input [63:0] prevA;
  input [63:0] prevSum;
  input [2:0] encoderIn;
  output [63:0] nextA;
  output [63:0] nextSum;

  wire   [2:0] encoder_to_mux;
  wire   [63:0] plus2A_s;
  wire   [63:0] minus2A_s;
  wire   [63:0] minus4A_s;
  tri   [63:0] mux_to_adder;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign nextA[0] = 1'b0;

  encoder_N64_RADIX3_1 encoder_1 ( .X(encoderIn), .Z(encoder_to_mux) );
  ShiftnCompl_N64_1 ShiftnCompl_1 ( .plusA(prevA), .plus2A_out({plus2A_s[63:1], 
        SYNOPSYS_UNCONNECTED__0}), .minus2A_out(minus2A_s), .plus4A_out({
        nextA[63:1], SYNOPSYS_UNCONNECTED__1}), .minus4A_out(minus4A_s) );
  MUX_GENERIC_N64_RADIX3_1 mux_1 ( .plusA({plus2A_s[63:1], 1'b0}), .minusA(
        minus2A_s), .plus2A({nextA[63:1], 1'b0}), .minus2A(minus4A_s), .SEL(
        encoder_to_mux), .Y(mux_to_adder) );
  RCA_N64_1 rca_1 ( .A(mux_to_adder), .B(prevSum), .Ci(1'b0), .S(nextSum) );
endmodule


module registers_N32_1 ( Clk, Rst, A, B, A_out, B_out );
  input [31:0] A;
  input [31:0] B;
  output [31:0] A_out;
  output [31:0] B_out;
  input Clk, Rst;
  wire   n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203;

  DFF_X1 \B_out_reg[1]  ( .D(n193), .CK(Clk), .Q(B_out[1]) );
  DFF_X1 \B_out_reg[0]  ( .D(n192), .CK(Clk), .Q(B_out[0]) );
  DFF_X1 \B_out_reg[2]  ( .D(n191), .CK(Clk), .Q(B_out[2]) );
  DFF_X1 \B_out_reg[3]  ( .D(n190), .CK(Clk), .Q(B_out[3]) );
  DFF_X1 \B_out_reg[4]  ( .D(n189), .CK(Clk), .Q(B_out[4]) );
  DFF_X1 \B_out_reg[5]  ( .D(n188), .CK(Clk), .Q(B_out[5]) );
  DFF_X1 \B_out_reg[6]  ( .D(n187), .CK(Clk), .Q(B_out[6]) );
  DFF_X1 \B_out_reg[7]  ( .D(n186), .CK(Clk), .Q(B_out[7]) );
  DFF_X1 \B_out_reg[8]  ( .D(n185), .CK(Clk), .Q(B_out[8]) );
  DFF_X1 \B_out_reg[9]  ( .D(n184), .CK(Clk), .Q(B_out[9]) );
  DFF_X1 \B_out_reg[10]  ( .D(n183), .CK(Clk), .Q(B_out[10]) );
  DFF_X1 \B_out_reg[11]  ( .D(n182), .CK(Clk), .Q(B_out[11]) );
  DFF_X1 \B_out_reg[12]  ( .D(n181), .CK(Clk), .Q(B_out[12]) );
  DFF_X1 \B_out_reg[13]  ( .D(n180), .CK(Clk), .Q(B_out[13]) );
  DFF_X1 \B_out_reg[14]  ( .D(n179), .CK(Clk), .Q(B_out[14]) );
  DFF_X1 \B_out_reg[15]  ( .D(n178), .CK(Clk), .Q(B_out[15]) );
  DFF_X1 \B_out_reg[16]  ( .D(n177), .CK(Clk), .Q(B_out[16]) );
  DFF_X1 \B_out_reg[17]  ( .D(n176), .CK(Clk), .Q(B_out[17]) );
  DFF_X1 \B_out_reg[18]  ( .D(n175), .CK(Clk), .Q(B_out[18]) );
  DFF_X1 \B_out_reg[19]  ( .D(n174), .CK(Clk), .Q(B_out[19]) );
  DFF_X1 \B_out_reg[20]  ( .D(n173), .CK(Clk), .Q(B_out[20]) );
  DFF_X1 \B_out_reg[21]  ( .D(n172), .CK(Clk), .Q(B_out[21]) );
  DFF_X1 \B_out_reg[22]  ( .D(n171), .CK(Clk), .Q(B_out[22]) );
  DFF_X1 \B_out_reg[23]  ( .D(n170), .CK(Clk), .Q(B_out[23]) );
  DFF_X1 \B_out_reg[24]  ( .D(n169), .CK(Clk), .Q(B_out[24]) );
  DFF_X1 \B_out_reg[25]  ( .D(n168), .CK(Clk), .Q(B_out[25]) );
  DFF_X1 \B_out_reg[26]  ( .D(n167), .CK(Clk), .Q(B_out[26]) );
  DFF_X1 \B_out_reg[27]  ( .D(n166), .CK(Clk), .Q(B_out[27]) );
  DFF_X1 \B_out_reg[28]  ( .D(n165), .CK(Clk), .Q(B_out[28]) );
  DFF_X1 \B_out_reg[29]  ( .D(n164), .CK(Clk), .Q(B_out[29]) );
  DFF_X1 \B_out_reg[30]  ( .D(n163), .CK(Clk), .Q(B_out[30]) );
  DFF_X1 \B_out_reg[31]  ( .D(n162), .CK(Clk), .Q(B_out[31]) );
  DFF_X1 \A_out_reg[0]  ( .D(n161), .CK(Clk), .Q(A_out[0]) );
  DFF_X1 \A_out_reg[1]  ( .D(n160), .CK(Clk), .Q(A_out[1]) );
  DFF_X1 \A_out_reg[2]  ( .D(n159), .CK(Clk), .Q(A_out[2]) );
  DFF_X1 \A_out_reg[3]  ( .D(n158), .CK(Clk), .Q(A_out[3]) );
  DFF_X1 \A_out_reg[4]  ( .D(n157), .CK(Clk), .Q(A_out[4]) );
  DFF_X1 \A_out_reg[5]  ( .D(n156), .CK(Clk), .Q(A_out[5]) );
  DFF_X1 \A_out_reg[6]  ( .D(n155), .CK(Clk), .Q(A_out[6]) );
  DFF_X1 \A_out_reg[7]  ( .D(n154), .CK(Clk), .Q(A_out[7]) );
  DFF_X1 \A_out_reg[8]  ( .D(n153), .CK(Clk), .Q(A_out[8]) );
  DFF_X1 \A_out_reg[9]  ( .D(n152), .CK(Clk), .Q(A_out[9]) );
  DFF_X1 \A_out_reg[10]  ( .D(n151), .CK(Clk), .Q(A_out[10]) );
  DFF_X1 \A_out_reg[11]  ( .D(n150), .CK(Clk), .Q(A_out[11]) );
  DFF_X1 \A_out_reg[12]  ( .D(n149), .CK(Clk), .Q(A_out[12]) );
  DFF_X1 \A_out_reg[13]  ( .D(n148), .CK(Clk), .Q(A_out[13]) );
  DFF_X1 \A_out_reg[14]  ( .D(n147), .CK(Clk), .Q(A_out[14]) );
  DFF_X1 \A_out_reg[15]  ( .D(n146), .CK(Clk), .Q(A_out[15]) );
  DFF_X1 \A_out_reg[16]  ( .D(n145), .CK(Clk), .Q(A_out[16]) );
  DFF_X1 \A_out_reg[17]  ( .D(n144), .CK(Clk), .Q(A_out[17]) );
  DFF_X1 \A_out_reg[18]  ( .D(n143), .CK(Clk), .Q(A_out[18]) );
  DFF_X1 \A_out_reg[19]  ( .D(n142), .CK(Clk), .Q(A_out[19]) );
  DFF_X1 \A_out_reg[20]  ( .D(n141), .CK(Clk), .Q(A_out[20]) );
  DFF_X1 \A_out_reg[21]  ( .D(n140), .CK(Clk), .Q(A_out[21]) );
  DFF_X1 \A_out_reg[22]  ( .D(n139), .CK(Clk), .Q(A_out[22]) );
  DFF_X1 \A_out_reg[23]  ( .D(n138), .CK(Clk), .Q(A_out[23]) );
  DFF_X1 \A_out_reg[24]  ( .D(n137), .CK(Clk), .Q(A_out[24]) );
  DFF_X1 \A_out_reg[25]  ( .D(n136), .CK(Clk), .Q(A_out[25]) );
  DFF_X1 \A_out_reg[26]  ( .D(n135), .CK(Clk), .Q(A_out[26]) );
  DFF_X1 \A_out_reg[27]  ( .D(n134), .CK(Clk), .Q(A_out[27]) );
  DFF_X1 \A_out_reg[28]  ( .D(n133), .CK(Clk), .Q(A_out[28]) );
  DFF_X1 \A_out_reg[29]  ( .D(n132), .CK(Clk), .Q(A_out[29]) );
  DFF_X1 \A_out_reg[30]  ( .D(n131), .CK(Clk), .Q(A_out[30]) );
  DFF_X1 \A_out_reg[31]  ( .D(n130), .CK(Clk), .Q(A_out[31]) );
  AND2_X1 U3 ( .A1(A[31]), .A2(n195), .ZN(n130) );
  AND2_X1 U4 ( .A1(A[30]), .A2(n195), .ZN(n131) );
  AND2_X1 U5 ( .A1(A[29]), .A2(n195), .ZN(n132) );
  AND2_X1 U6 ( .A1(A[28]), .A2(n195), .ZN(n133) );
  AND2_X1 U7 ( .A1(A[27]), .A2(n195), .ZN(n134) );
  AND2_X1 U8 ( .A1(A[26]), .A2(n195), .ZN(n135) );
  AND2_X1 U9 ( .A1(A[25]), .A2(n195), .ZN(n136) );
  AND2_X1 U10 ( .A1(A[24]), .A2(n195), .ZN(n137) );
  AND2_X1 U11 ( .A1(A[23]), .A2(n195), .ZN(n138) );
  AND2_X1 U12 ( .A1(A[22]), .A2(n195), .ZN(n139) );
  AND2_X1 U13 ( .A1(A[21]), .A2(n196), .ZN(n140) );
  AND2_X1 U14 ( .A1(A[20]), .A2(n196), .ZN(n141) );
  AND2_X1 U15 ( .A1(A[19]), .A2(n196), .ZN(n142) );
  AND2_X1 U16 ( .A1(A[18]), .A2(n196), .ZN(n143) );
  AND2_X1 U17 ( .A1(A[17]), .A2(n196), .ZN(n144) );
  AND2_X1 U18 ( .A1(A[16]), .A2(n196), .ZN(n145) );
  AND2_X1 U19 ( .A1(A[15]), .A2(n196), .ZN(n146) );
  AND2_X1 U20 ( .A1(A[14]), .A2(n196), .ZN(n147) );
  AND2_X1 U21 ( .A1(A[13]), .A2(n196), .ZN(n148) );
  AND2_X1 U22 ( .A1(A[12]), .A2(n196), .ZN(n149) );
  AND2_X1 U23 ( .A1(A[11]), .A2(n197), .ZN(n150) );
  AND2_X1 U24 ( .A1(A[10]), .A2(n197), .ZN(n151) );
  AND2_X1 U25 ( .A1(A[9]), .A2(n197), .ZN(n152) );
  AND2_X1 U26 ( .A1(A[8]), .A2(n197), .ZN(n153) );
  AND2_X1 U27 ( .A1(A[7]), .A2(n197), .ZN(n154) );
  AND2_X1 U28 ( .A1(A[6]), .A2(n197), .ZN(n155) );
  AND2_X1 U29 ( .A1(A[5]), .A2(n197), .ZN(n156) );
  AND2_X1 U30 ( .A1(A[4]), .A2(n197), .ZN(n157) );
  AND2_X1 U31 ( .A1(A[3]), .A2(n197), .ZN(n158) );
  AND2_X1 U32 ( .A1(A[2]), .A2(n197), .ZN(n159) );
  AND2_X1 U33 ( .A1(A[1]), .A2(n198), .ZN(n160) );
  AND2_X1 U34 ( .A1(A[0]), .A2(n198), .ZN(n161) );
  AND2_X1 U35 ( .A1(B[31]), .A2(n198), .ZN(n162) );
  AND2_X1 U36 ( .A1(B[30]), .A2(n198), .ZN(n163) );
  AND2_X1 U37 ( .A1(B[29]), .A2(n198), .ZN(n164) );
  AND2_X1 U38 ( .A1(B[28]), .A2(n198), .ZN(n165) );
  AND2_X1 U39 ( .A1(B[27]), .A2(n198), .ZN(n166) );
  AND2_X1 U40 ( .A1(B[26]), .A2(n198), .ZN(n167) );
  AND2_X1 U41 ( .A1(B[25]), .A2(n198), .ZN(n168) );
  AND2_X1 U42 ( .A1(B[24]), .A2(n198), .ZN(n169) );
  AND2_X1 U43 ( .A1(B[23]), .A2(n199), .ZN(n170) );
  AND2_X1 U44 ( .A1(B[22]), .A2(n199), .ZN(n171) );
  AND2_X1 U45 ( .A1(B[21]), .A2(n199), .ZN(n172) );
  AND2_X1 U46 ( .A1(B[20]), .A2(n199), .ZN(n173) );
  AND2_X1 U47 ( .A1(B[19]), .A2(n199), .ZN(n174) );
  AND2_X1 U48 ( .A1(B[18]), .A2(n199), .ZN(n175) );
  AND2_X1 U49 ( .A1(B[17]), .A2(n199), .ZN(n176) );
  AND2_X1 U50 ( .A1(B[16]), .A2(n199), .ZN(n177) );
  AND2_X1 U51 ( .A1(B[15]), .A2(n199), .ZN(n178) );
  AND2_X1 U52 ( .A1(B[14]), .A2(n199), .ZN(n179) );
  AND2_X1 U53 ( .A1(B[13]), .A2(n200), .ZN(n180) );
  AND2_X1 U54 ( .A1(B[12]), .A2(n200), .ZN(n181) );
  AND2_X1 U55 ( .A1(B[11]), .A2(n200), .ZN(n182) );
  AND2_X1 U56 ( .A1(B[10]), .A2(n200), .ZN(n183) );
  AND2_X1 U57 ( .A1(B[9]), .A2(n194), .ZN(n184) );
  AND2_X1 U58 ( .A1(B[8]), .A2(n194), .ZN(n185) );
  AND2_X1 U59 ( .A1(B[7]), .A2(n194), .ZN(n186) );
  AND2_X1 U60 ( .A1(B[6]), .A2(n194), .ZN(n187) );
  AND2_X1 U61 ( .A1(B[5]), .A2(n194), .ZN(n188) );
  AND2_X1 U62 ( .A1(B[4]), .A2(n194), .ZN(n189) );
  AND2_X1 U63 ( .A1(B[3]), .A2(n194), .ZN(n190) );
  AND2_X1 U64 ( .A1(B[2]), .A2(n194), .ZN(n191) );
  AND2_X1 U65 ( .A1(B[0]), .A2(n194), .ZN(n192) );
  AND2_X1 U66 ( .A1(B[1]), .A2(n194), .ZN(n193) );
  BUF_X1 U67 ( .A(n201), .Z(n197) );
  BUF_X1 U68 ( .A(n201), .Z(n199) );
  BUF_X1 U69 ( .A(n201), .Z(n198) );
  BUF_X1 U70 ( .A(n202), .Z(n196) );
  BUF_X1 U71 ( .A(n202), .Z(n195) );
  BUF_X1 U72 ( .A(n202), .Z(n194) );
  BUF_X1 U73 ( .A(n203), .Z(n201) );
  BUF_X1 U74 ( .A(n203), .Z(n202) );
  INV_X1 U75 ( .A(Rst), .ZN(n203) );
  CLKBUF_X1 U76 ( .A(n201), .Z(n200) );
endmodule


module Booth ( Clk, Rst, A, B, P );
  input [31:0] A;
  input [31:0] B;
  output [63:0] P;
  input Clk, Rst;
  wire   \sigMatrix[0][127] , \sigMatrix[0][126] , \sigMatrix[0][125] ,
         \sigMatrix[0][124] , \sigMatrix[0][123] , \sigMatrix[0][122] ,
         \sigMatrix[0][121] , \sigMatrix[0][120] , \sigMatrix[0][119] ,
         \sigMatrix[0][118] , \sigMatrix[0][117] , \sigMatrix[0][116] ,
         \sigMatrix[0][115] , \sigMatrix[0][114] , \sigMatrix[0][113] ,
         \sigMatrix[0][112] , \sigMatrix[0][111] , \sigMatrix[0][110] ,
         \sigMatrix[0][109] , \sigMatrix[0][108] , \sigMatrix[0][107] ,
         \sigMatrix[0][106] , \sigMatrix[0][105] , \sigMatrix[0][104] ,
         \sigMatrix[0][103] , \sigMatrix[0][102] , \sigMatrix[0][101] ,
         \sigMatrix[0][100] , \sigMatrix[0][99] , \sigMatrix[0][98] ,
         \sigMatrix[0][97] , \sigMatrix[0][96] , \sigMatrix[0][95] ,
         \sigMatrix[0][94] , \sigMatrix[0][93] , \sigMatrix[0][92] ,
         \sigMatrix[0][91] , \sigMatrix[0][90] , \sigMatrix[0][89] ,
         \sigMatrix[0][88] , \sigMatrix[0][87] , \sigMatrix[0][86] ,
         \sigMatrix[0][85] , \sigMatrix[0][84] , \sigMatrix[0][83] ,
         \sigMatrix[0][82] , \sigMatrix[0][81] , \sigMatrix[0][80] ,
         \sigMatrix[0][79] , \sigMatrix[0][78] , \sigMatrix[0][77] ,
         \sigMatrix[0][76] , \sigMatrix[0][75] , \sigMatrix[0][74] ,
         \sigMatrix[0][73] , \sigMatrix[0][72] , \sigMatrix[0][71] ,
         \sigMatrix[0][70] , \sigMatrix[0][69] , \sigMatrix[0][68] ,
         \sigMatrix[0][67] , \sigMatrix[0][66] , \sigMatrix[0][65] ,
         \sigMatrix[1][127] , \sigMatrix[1][126] , \sigMatrix[1][125] ,
         \sigMatrix[1][124] , \sigMatrix[1][123] , \sigMatrix[1][122] ,
         \sigMatrix[1][121] , \sigMatrix[1][120] , \sigMatrix[1][119] ,
         \sigMatrix[1][118] , \sigMatrix[1][117] , \sigMatrix[1][116] ,
         \sigMatrix[1][115] , \sigMatrix[1][114] , \sigMatrix[1][113] ,
         \sigMatrix[1][112] , \sigMatrix[1][111] , \sigMatrix[1][110] ,
         \sigMatrix[1][109] , \sigMatrix[1][108] , \sigMatrix[1][107] ,
         \sigMatrix[1][106] , \sigMatrix[1][105] , \sigMatrix[1][104] ,
         \sigMatrix[1][103] , \sigMatrix[1][102] , \sigMatrix[1][101] ,
         \sigMatrix[1][100] , \sigMatrix[1][99] , \sigMatrix[1][98] ,
         \sigMatrix[1][97] , \sigMatrix[1][96] , \sigMatrix[1][95] ,
         \sigMatrix[1][94] , \sigMatrix[1][93] , \sigMatrix[1][92] ,
         \sigMatrix[1][91] , \sigMatrix[1][90] , \sigMatrix[1][89] ,
         \sigMatrix[1][88] , \sigMatrix[1][87] , \sigMatrix[1][86] ,
         \sigMatrix[1][85] , \sigMatrix[1][84] , \sigMatrix[1][83] ,
         \sigMatrix[1][82] , \sigMatrix[1][81] , \sigMatrix[1][80] ,
         \sigMatrix[1][79] , \sigMatrix[1][78] , \sigMatrix[1][77] ,
         \sigMatrix[1][76] , \sigMatrix[1][75] , \sigMatrix[1][74] ,
         \sigMatrix[1][73] , \sigMatrix[1][72] , \sigMatrix[1][71] ,
         \sigMatrix[1][70] , \sigMatrix[1][69] , \sigMatrix[1][68] ,
         \sigMatrix[1][67] , \sigMatrix[1][66] , \sigMatrix[1][65] ,
         \sigMatrix[1][63] , \sigMatrix[1][62] , \sigMatrix[1][61] ,
         \sigMatrix[1][60] , \sigMatrix[1][59] , \sigMatrix[1][58] ,
         \sigMatrix[1][57] , \sigMatrix[1][56] , \sigMatrix[1][55] ,
         \sigMatrix[1][54] , \sigMatrix[1][53] , \sigMatrix[1][52] ,
         \sigMatrix[1][51] , \sigMatrix[1][50] , \sigMatrix[1][49] ,
         \sigMatrix[1][48] , \sigMatrix[1][47] , \sigMatrix[1][46] ,
         \sigMatrix[1][45] , \sigMatrix[1][44] , \sigMatrix[1][43] ,
         \sigMatrix[1][42] , \sigMatrix[1][41] , \sigMatrix[1][40] ,
         \sigMatrix[1][39] , \sigMatrix[1][38] , \sigMatrix[1][37] ,
         \sigMatrix[1][36] , \sigMatrix[1][35] , \sigMatrix[1][34] ,
         \sigMatrix[1][33] , \sigMatrix[1][32] , \sigMatrix[1][31] ,
         \sigMatrix[1][30] , \sigMatrix[1][29] , \sigMatrix[1][28] ,
         \sigMatrix[1][27] , \sigMatrix[1][26] , \sigMatrix[1][25] ,
         \sigMatrix[1][24] , \sigMatrix[1][23] , \sigMatrix[1][22] ,
         \sigMatrix[1][21] , \sigMatrix[1][20] , \sigMatrix[1][19] ,
         \sigMatrix[1][18] , \sigMatrix[1][17] , \sigMatrix[1][16] ,
         \sigMatrix[1][15] , \sigMatrix[1][14] , \sigMatrix[1][13] ,
         \sigMatrix[1][12] , \sigMatrix[1][11] , \sigMatrix[1][10] ,
         \sigMatrix[1][9] , \sigMatrix[1][8] , \sigMatrix[1][7] ,
         \sigMatrix[1][6] , \sigMatrix[1][5] , \sigMatrix[1][4] ,
         \sigMatrix[1][3] , \sigMatrix[1][2] , \sigMatrix[1][1] ,
         \sigMatrix[1][0] , \sigMatrix[2][127] , \sigMatrix[2][126] ,
         \sigMatrix[2][125] , \sigMatrix[2][124] , \sigMatrix[2][123] ,
         \sigMatrix[2][122] , \sigMatrix[2][121] , \sigMatrix[2][120] ,
         \sigMatrix[2][119] , \sigMatrix[2][118] , \sigMatrix[2][117] ,
         \sigMatrix[2][116] , \sigMatrix[2][115] , \sigMatrix[2][114] ,
         \sigMatrix[2][113] , \sigMatrix[2][112] , \sigMatrix[2][111] ,
         \sigMatrix[2][110] , \sigMatrix[2][109] , \sigMatrix[2][108] ,
         \sigMatrix[2][107] , \sigMatrix[2][106] , \sigMatrix[2][105] ,
         \sigMatrix[2][104] , \sigMatrix[2][103] , \sigMatrix[2][102] ,
         \sigMatrix[2][101] , \sigMatrix[2][100] , \sigMatrix[2][99] ,
         \sigMatrix[2][98] , \sigMatrix[2][97] , \sigMatrix[2][96] ,
         \sigMatrix[2][95] , \sigMatrix[2][94] , \sigMatrix[2][93] ,
         \sigMatrix[2][92] , \sigMatrix[2][91] , \sigMatrix[2][90] ,
         \sigMatrix[2][89] , \sigMatrix[2][88] , \sigMatrix[2][87] ,
         \sigMatrix[2][86] , \sigMatrix[2][85] , \sigMatrix[2][84] ,
         \sigMatrix[2][83] , \sigMatrix[2][82] , \sigMatrix[2][81] ,
         \sigMatrix[2][80] , \sigMatrix[2][79] , \sigMatrix[2][78] ,
         \sigMatrix[2][77] , \sigMatrix[2][76] , \sigMatrix[2][75] ,
         \sigMatrix[2][74] , \sigMatrix[2][73] , \sigMatrix[2][72] ,
         \sigMatrix[2][71] , \sigMatrix[2][70] , \sigMatrix[2][69] ,
         \sigMatrix[2][68] , \sigMatrix[2][67] , \sigMatrix[2][66] ,
         \sigMatrix[2][65] , \sigMatrix[2][63] , \sigMatrix[2][62] ,
         \sigMatrix[2][61] , \sigMatrix[2][60] , \sigMatrix[2][59] ,
         \sigMatrix[2][58] , \sigMatrix[2][57] , \sigMatrix[2][56] ,
         \sigMatrix[2][55] , \sigMatrix[2][54] , \sigMatrix[2][53] ,
         \sigMatrix[2][52] , \sigMatrix[2][51] , \sigMatrix[2][50] ,
         \sigMatrix[2][49] , \sigMatrix[2][48] , \sigMatrix[2][47] ,
         \sigMatrix[2][46] , \sigMatrix[2][45] , \sigMatrix[2][44] ,
         \sigMatrix[2][43] , \sigMatrix[2][42] , \sigMatrix[2][41] ,
         \sigMatrix[2][40] , \sigMatrix[2][39] , \sigMatrix[2][38] ,
         \sigMatrix[2][37] , \sigMatrix[2][36] , \sigMatrix[2][35] ,
         \sigMatrix[2][34] , \sigMatrix[2][33] , \sigMatrix[2][32] ,
         \sigMatrix[2][31] , \sigMatrix[2][30] , \sigMatrix[2][29] ,
         \sigMatrix[2][28] , \sigMatrix[2][27] , \sigMatrix[2][26] ,
         \sigMatrix[2][25] , \sigMatrix[2][24] , \sigMatrix[2][23] ,
         \sigMatrix[2][22] , \sigMatrix[2][21] , \sigMatrix[2][20] ,
         \sigMatrix[2][19] , \sigMatrix[2][18] , \sigMatrix[2][17] ,
         \sigMatrix[2][16] , \sigMatrix[2][15] , \sigMatrix[2][14] ,
         \sigMatrix[2][13] , \sigMatrix[2][12] , \sigMatrix[2][11] ,
         \sigMatrix[2][10] , \sigMatrix[2][9] , \sigMatrix[2][8] ,
         \sigMatrix[2][7] , \sigMatrix[2][6] , \sigMatrix[2][5] ,
         \sigMatrix[2][4] , \sigMatrix[2][3] , \sigMatrix[2][2] ,
         \sigMatrix[2][1] , \sigMatrix[2][0] , \sigMatrix[3][127] ,
         \sigMatrix[3][126] , \sigMatrix[3][125] , \sigMatrix[3][124] ,
         \sigMatrix[3][123] , \sigMatrix[3][122] , \sigMatrix[3][121] ,
         \sigMatrix[3][120] , \sigMatrix[3][119] , \sigMatrix[3][118] ,
         \sigMatrix[3][117] , \sigMatrix[3][116] , \sigMatrix[3][115] ,
         \sigMatrix[3][114] , \sigMatrix[3][113] , \sigMatrix[3][112] ,
         \sigMatrix[3][111] , \sigMatrix[3][110] , \sigMatrix[3][109] ,
         \sigMatrix[3][108] , \sigMatrix[3][107] , \sigMatrix[3][106] ,
         \sigMatrix[3][105] , \sigMatrix[3][104] , \sigMatrix[3][103] ,
         \sigMatrix[3][102] , \sigMatrix[3][101] , \sigMatrix[3][100] ,
         \sigMatrix[3][99] , \sigMatrix[3][98] , \sigMatrix[3][97] ,
         \sigMatrix[3][96] , \sigMatrix[3][95] , \sigMatrix[3][94] ,
         \sigMatrix[3][93] , \sigMatrix[3][92] , \sigMatrix[3][91] ,
         \sigMatrix[3][90] , \sigMatrix[3][89] , \sigMatrix[3][88] ,
         \sigMatrix[3][87] , \sigMatrix[3][86] , \sigMatrix[3][85] ,
         \sigMatrix[3][84] , \sigMatrix[3][83] , \sigMatrix[3][82] ,
         \sigMatrix[3][81] , \sigMatrix[3][80] , \sigMatrix[3][79] ,
         \sigMatrix[3][78] , \sigMatrix[3][77] , \sigMatrix[3][76] ,
         \sigMatrix[3][75] , \sigMatrix[3][74] , \sigMatrix[3][73] ,
         \sigMatrix[3][72] , \sigMatrix[3][71] , \sigMatrix[3][70] ,
         \sigMatrix[3][69] , \sigMatrix[3][68] , \sigMatrix[3][67] ,
         \sigMatrix[3][66] , \sigMatrix[3][65] , \sigMatrix[3][63] ,
         \sigMatrix[3][62] , \sigMatrix[3][61] , \sigMatrix[3][60] ,
         \sigMatrix[3][59] , \sigMatrix[3][58] , \sigMatrix[3][57] ,
         \sigMatrix[3][56] , \sigMatrix[3][55] , \sigMatrix[3][54] ,
         \sigMatrix[3][53] , \sigMatrix[3][52] , \sigMatrix[3][51] ,
         \sigMatrix[3][50] , \sigMatrix[3][49] , \sigMatrix[3][48] ,
         \sigMatrix[3][47] , \sigMatrix[3][46] , \sigMatrix[3][45] ,
         \sigMatrix[3][44] , \sigMatrix[3][43] , \sigMatrix[3][42] ,
         \sigMatrix[3][41] , \sigMatrix[3][40] , \sigMatrix[3][39] ,
         \sigMatrix[3][38] , \sigMatrix[3][37] , \sigMatrix[3][36] ,
         \sigMatrix[3][35] , \sigMatrix[3][34] , \sigMatrix[3][33] ,
         \sigMatrix[3][32] , \sigMatrix[3][31] , \sigMatrix[3][30] ,
         \sigMatrix[3][29] , \sigMatrix[3][28] , \sigMatrix[3][27] ,
         \sigMatrix[3][26] , \sigMatrix[3][25] , \sigMatrix[3][24] ,
         \sigMatrix[3][23] , \sigMatrix[3][22] , \sigMatrix[3][21] ,
         \sigMatrix[3][20] , \sigMatrix[3][19] , \sigMatrix[3][18] ,
         \sigMatrix[3][17] , \sigMatrix[3][16] , \sigMatrix[3][15] ,
         \sigMatrix[3][14] , \sigMatrix[3][13] , \sigMatrix[3][12] ,
         \sigMatrix[3][11] , \sigMatrix[3][10] , \sigMatrix[3][9] ,
         \sigMatrix[3][8] , \sigMatrix[3][7] , \sigMatrix[3][6] ,
         \sigMatrix[3][5] , \sigMatrix[3][4] , \sigMatrix[3][3] ,
         \sigMatrix[3][2] , \sigMatrix[3][1] , \sigMatrix[3][0] ,
         \sigMatrix[4][127] , \sigMatrix[4][126] , \sigMatrix[4][125] ,
         \sigMatrix[4][124] , \sigMatrix[4][123] , \sigMatrix[4][122] ,
         \sigMatrix[4][121] , \sigMatrix[4][120] , \sigMatrix[4][119] ,
         \sigMatrix[4][118] , \sigMatrix[4][117] , \sigMatrix[4][116] ,
         \sigMatrix[4][115] , \sigMatrix[4][114] , \sigMatrix[4][113] ,
         \sigMatrix[4][112] , \sigMatrix[4][111] , \sigMatrix[4][110] ,
         \sigMatrix[4][109] , \sigMatrix[4][108] , \sigMatrix[4][107] ,
         \sigMatrix[4][106] , \sigMatrix[4][105] , \sigMatrix[4][104] ,
         \sigMatrix[4][103] , \sigMatrix[4][102] , \sigMatrix[4][101] ,
         \sigMatrix[4][100] , \sigMatrix[4][99] , \sigMatrix[4][98] ,
         \sigMatrix[4][97] , \sigMatrix[4][96] , \sigMatrix[4][95] ,
         \sigMatrix[4][94] , \sigMatrix[4][93] , \sigMatrix[4][92] ,
         \sigMatrix[4][91] , \sigMatrix[4][90] , \sigMatrix[4][89] ,
         \sigMatrix[4][88] , \sigMatrix[4][87] , \sigMatrix[4][86] ,
         \sigMatrix[4][85] , \sigMatrix[4][84] , \sigMatrix[4][83] ,
         \sigMatrix[4][82] , \sigMatrix[4][81] , \sigMatrix[4][80] ,
         \sigMatrix[4][79] , \sigMatrix[4][78] , \sigMatrix[4][77] ,
         \sigMatrix[4][76] , \sigMatrix[4][75] , \sigMatrix[4][74] ,
         \sigMatrix[4][73] , \sigMatrix[4][72] , \sigMatrix[4][71] ,
         \sigMatrix[4][70] , \sigMatrix[4][69] , \sigMatrix[4][68] ,
         \sigMatrix[4][67] , \sigMatrix[4][66] , \sigMatrix[4][65] ,
         \sigMatrix[4][63] , \sigMatrix[4][62] , \sigMatrix[4][61] ,
         \sigMatrix[4][60] , \sigMatrix[4][59] , \sigMatrix[4][58] ,
         \sigMatrix[4][57] , \sigMatrix[4][56] , \sigMatrix[4][55] ,
         \sigMatrix[4][54] , \sigMatrix[4][53] , \sigMatrix[4][52] ,
         \sigMatrix[4][51] , \sigMatrix[4][50] , \sigMatrix[4][49] ,
         \sigMatrix[4][48] , \sigMatrix[4][47] , \sigMatrix[4][46] ,
         \sigMatrix[4][45] , \sigMatrix[4][44] , \sigMatrix[4][43] ,
         \sigMatrix[4][42] , \sigMatrix[4][41] , \sigMatrix[4][40] ,
         \sigMatrix[4][39] , \sigMatrix[4][38] , \sigMatrix[4][37] ,
         \sigMatrix[4][36] , \sigMatrix[4][35] , \sigMatrix[4][34] ,
         \sigMatrix[4][33] , \sigMatrix[4][32] , \sigMatrix[4][31] ,
         \sigMatrix[4][30] , \sigMatrix[4][29] , \sigMatrix[4][28] ,
         \sigMatrix[4][27] , \sigMatrix[4][26] , \sigMatrix[4][25] ,
         \sigMatrix[4][24] , \sigMatrix[4][23] , \sigMatrix[4][22] ,
         \sigMatrix[4][21] , \sigMatrix[4][20] , \sigMatrix[4][19] ,
         \sigMatrix[4][18] , \sigMatrix[4][17] , \sigMatrix[4][16] ,
         \sigMatrix[4][15] , \sigMatrix[4][14] , \sigMatrix[4][13] ,
         \sigMatrix[4][12] , \sigMatrix[4][11] , \sigMatrix[4][10] ,
         \sigMatrix[4][9] , \sigMatrix[4][8] , \sigMatrix[4][7] ,
         \sigMatrix[4][6] , \sigMatrix[4][5] , \sigMatrix[4][4] ,
         \sigMatrix[4][3] , \sigMatrix[4][2] , \sigMatrix[4][1] ,
         \sigMatrix[4][0] , \sigMatrix[5][127] , \sigMatrix[5][126] ,
         \sigMatrix[5][125] , \sigMatrix[5][124] , \sigMatrix[5][123] ,
         \sigMatrix[5][122] , \sigMatrix[5][121] , \sigMatrix[5][120] ,
         \sigMatrix[5][119] , \sigMatrix[5][118] , \sigMatrix[5][117] ,
         \sigMatrix[5][116] , \sigMatrix[5][115] , \sigMatrix[5][114] ,
         \sigMatrix[5][113] , \sigMatrix[5][112] , \sigMatrix[5][111] ,
         \sigMatrix[5][110] , \sigMatrix[5][109] , \sigMatrix[5][108] ,
         \sigMatrix[5][107] , \sigMatrix[5][106] , \sigMatrix[5][105] ,
         \sigMatrix[5][104] , \sigMatrix[5][103] , \sigMatrix[5][102] ,
         \sigMatrix[5][101] , \sigMatrix[5][100] , \sigMatrix[5][99] ,
         \sigMatrix[5][98] , \sigMatrix[5][97] , \sigMatrix[5][96] ,
         \sigMatrix[5][95] , \sigMatrix[5][94] , \sigMatrix[5][93] ,
         \sigMatrix[5][92] , \sigMatrix[5][91] , \sigMatrix[5][90] ,
         \sigMatrix[5][89] , \sigMatrix[5][88] , \sigMatrix[5][87] ,
         \sigMatrix[5][86] , \sigMatrix[5][85] , \sigMatrix[5][84] ,
         \sigMatrix[5][83] , \sigMatrix[5][82] , \sigMatrix[5][81] ,
         \sigMatrix[5][80] , \sigMatrix[5][79] , \sigMatrix[5][78] ,
         \sigMatrix[5][77] , \sigMatrix[5][76] , \sigMatrix[5][75] ,
         \sigMatrix[5][74] , \sigMatrix[5][73] , \sigMatrix[5][72] ,
         \sigMatrix[5][71] , \sigMatrix[5][70] , \sigMatrix[5][69] ,
         \sigMatrix[5][68] , \sigMatrix[5][67] , \sigMatrix[5][66] ,
         \sigMatrix[5][65] , \sigMatrix[5][63] , \sigMatrix[5][62] ,
         \sigMatrix[5][61] , \sigMatrix[5][60] , \sigMatrix[5][59] ,
         \sigMatrix[5][58] , \sigMatrix[5][57] , \sigMatrix[5][56] ,
         \sigMatrix[5][55] , \sigMatrix[5][54] , \sigMatrix[5][53] ,
         \sigMatrix[5][52] , \sigMatrix[5][51] , \sigMatrix[5][50] ,
         \sigMatrix[5][49] , \sigMatrix[5][48] , \sigMatrix[5][47] ,
         \sigMatrix[5][46] , \sigMatrix[5][45] , \sigMatrix[5][44] ,
         \sigMatrix[5][43] , \sigMatrix[5][42] , \sigMatrix[5][41] ,
         \sigMatrix[5][40] , \sigMatrix[5][39] , \sigMatrix[5][38] ,
         \sigMatrix[5][37] , \sigMatrix[5][36] , \sigMatrix[5][35] ,
         \sigMatrix[5][34] , \sigMatrix[5][33] , \sigMatrix[5][32] ,
         \sigMatrix[5][31] , \sigMatrix[5][30] , \sigMatrix[5][29] ,
         \sigMatrix[5][28] , \sigMatrix[5][27] , \sigMatrix[5][26] ,
         \sigMatrix[5][25] , \sigMatrix[5][24] , \sigMatrix[5][23] ,
         \sigMatrix[5][22] , \sigMatrix[5][21] , \sigMatrix[5][20] ,
         \sigMatrix[5][19] , \sigMatrix[5][18] , \sigMatrix[5][17] ,
         \sigMatrix[5][16] , \sigMatrix[5][15] , \sigMatrix[5][14] ,
         \sigMatrix[5][13] , \sigMatrix[5][12] , \sigMatrix[5][11] ,
         \sigMatrix[5][10] , \sigMatrix[5][9] , \sigMatrix[5][8] ,
         \sigMatrix[5][7] , \sigMatrix[5][6] , \sigMatrix[5][5] ,
         \sigMatrix[5][4] , \sigMatrix[5][3] , \sigMatrix[5][2] ,
         \sigMatrix[5][1] , \sigMatrix[5][0] , \sigMatrix[6][127] ,
         \sigMatrix[6][126] , \sigMatrix[6][125] , \sigMatrix[6][124] ,
         \sigMatrix[6][123] , \sigMatrix[6][122] , \sigMatrix[6][121] ,
         \sigMatrix[6][120] , \sigMatrix[6][119] , \sigMatrix[6][118] ,
         \sigMatrix[6][117] , \sigMatrix[6][116] , \sigMatrix[6][115] ,
         \sigMatrix[6][114] , \sigMatrix[6][113] , \sigMatrix[6][112] ,
         \sigMatrix[6][111] , \sigMatrix[6][110] , \sigMatrix[6][109] ,
         \sigMatrix[6][108] , \sigMatrix[6][107] , \sigMatrix[6][106] ,
         \sigMatrix[6][105] , \sigMatrix[6][104] , \sigMatrix[6][103] ,
         \sigMatrix[6][102] , \sigMatrix[6][101] , \sigMatrix[6][100] ,
         \sigMatrix[6][99] , \sigMatrix[6][98] , \sigMatrix[6][97] ,
         \sigMatrix[6][96] , \sigMatrix[6][95] , \sigMatrix[6][94] ,
         \sigMatrix[6][93] , \sigMatrix[6][92] , \sigMatrix[6][91] ,
         \sigMatrix[6][90] , \sigMatrix[6][89] , \sigMatrix[6][88] ,
         \sigMatrix[6][87] , \sigMatrix[6][86] , \sigMatrix[6][85] ,
         \sigMatrix[6][84] , \sigMatrix[6][83] , \sigMatrix[6][82] ,
         \sigMatrix[6][81] , \sigMatrix[6][80] , \sigMatrix[6][79] ,
         \sigMatrix[6][78] , \sigMatrix[6][77] , \sigMatrix[6][76] ,
         \sigMatrix[6][75] , \sigMatrix[6][74] , \sigMatrix[6][73] ,
         \sigMatrix[6][72] , \sigMatrix[6][71] , \sigMatrix[6][70] ,
         \sigMatrix[6][69] , \sigMatrix[6][68] , \sigMatrix[6][67] ,
         \sigMatrix[6][66] , \sigMatrix[6][65] , \sigMatrix[6][63] ,
         \sigMatrix[6][62] , \sigMatrix[6][61] , \sigMatrix[6][60] ,
         \sigMatrix[6][59] , \sigMatrix[6][58] , \sigMatrix[6][57] ,
         \sigMatrix[6][56] , \sigMatrix[6][55] , \sigMatrix[6][54] ,
         \sigMatrix[6][53] , \sigMatrix[6][52] , \sigMatrix[6][51] ,
         \sigMatrix[6][50] , \sigMatrix[6][49] , \sigMatrix[6][48] ,
         \sigMatrix[6][47] , \sigMatrix[6][46] , \sigMatrix[6][45] ,
         \sigMatrix[6][44] , \sigMatrix[6][43] , \sigMatrix[6][42] ,
         \sigMatrix[6][41] , \sigMatrix[6][40] , \sigMatrix[6][39] ,
         \sigMatrix[6][38] , \sigMatrix[6][37] , \sigMatrix[6][36] ,
         \sigMatrix[6][35] , \sigMatrix[6][34] , \sigMatrix[6][33] ,
         \sigMatrix[6][32] , \sigMatrix[6][31] , \sigMatrix[6][30] ,
         \sigMatrix[6][29] , \sigMatrix[6][28] , \sigMatrix[6][27] ,
         \sigMatrix[6][26] , \sigMatrix[6][25] , \sigMatrix[6][24] ,
         \sigMatrix[6][23] , \sigMatrix[6][22] , \sigMatrix[6][21] ,
         \sigMatrix[6][20] , \sigMatrix[6][19] , \sigMatrix[6][18] ,
         \sigMatrix[6][17] , \sigMatrix[6][16] , \sigMatrix[6][15] ,
         \sigMatrix[6][14] , \sigMatrix[6][13] , \sigMatrix[6][12] ,
         \sigMatrix[6][11] , \sigMatrix[6][10] , \sigMatrix[6][9] ,
         \sigMatrix[6][8] , \sigMatrix[6][7] , \sigMatrix[6][6] ,
         \sigMatrix[6][5] , \sigMatrix[6][4] , \sigMatrix[6][3] ,
         \sigMatrix[6][2] , \sigMatrix[6][1] , \sigMatrix[6][0] ,
         \sigMatrix[7][127] , \sigMatrix[7][126] , \sigMatrix[7][125] ,
         \sigMatrix[7][124] , \sigMatrix[7][123] , \sigMatrix[7][122] ,
         \sigMatrix[7][121] , \sigMatrix[7][120] , \sigMatrix[7][119] ,
         \sigMatrix[7][118] , \sigMatrix[7][117] , \sigMatrix[7][116] ,
         \sigMatrix[7][115] , \sigMatrix[7][114] , \sigMatrix[7][113] ,
         \sigMatrix[7][112] , \sigMatrix[7][111] , \sigMatrix[7][110] ,
         \sigMatrix[7][109] , \sigMatrix[7][108] , \sigMatrix[7][107] ,
         \sigMatrix[7][106] , \sigMatrix[7][105] , \sigMatrix[7][104] ,
         \sigMatrix[7][103] , \sigMatrix[7][102] , \sigMatrix[7][101] ,
         \sigMatrix[7][100] , \sigMatrix[7][99] , \sigMatrix[7][98] ,
         \sigMatrix[7][97] , \sigMatrix[7][96] , \sigMatrix[7][95] ,
         \sigMatrix[7][94] , \sigMatrix[7][93] , \sigMatrix[7][92] ,
         \sigMatrix[7][91] , \sigMatrix[7][90] , \sigMatrix[7][89] ,
         \sigMatrix[7][88] , \sigMatrix[7][87] , \sigMatrix[7][86] ,
         \sigMatrix[7][85] , \sigMatrix[7][84] , \sigMatrix[7][83] ,
         \sigMatrix[7][82] , \sigMatrix[7][81] , \sigMatrix[7][80] ,
         \sigMatrix[7][79] , \sigMatrix[7][78] , \sigMatrix[7][77] ,
         \sigMatrix[7][76] , \sigMatrix[7][75] , \sigMatrix[7][74] ,
         \sigMatrix[7][73] , \sigMatrix[7][72] , \sigMatrix[7][71] ,
         \sigMatrix[7][70] , \sigMatrix[7][69] , \sigMatrix[7][68] ,
         \sigMatrix[7][67] , \sigMatrix[7][66] , \sigMatrix[7][65] ,
         \sigMatrix[7][63] , \sigMatrix[7][62] , \sigMatrix[7][61] ,
         \sigMatrix[7][60] , \sigMatrix[7][59] , \sigMatrix[7][58] ,
         \sigMatrix[7][57] , \sigMatrix[7][56] , \sigMatrix[7][55] ,
         \sigMatrix[7][54] , \sigMatrix[7][53] , \sigMatrix[7][52] ,
         \sigMatrix[7][51] , \sigMatrix[7][50] , \sigMatrix[7][49] ,
         \sigMatrix[7][48] , \sigMatrix[7][47] , \sigMatrix[7][46] ,
         \sigMatrix[7][45] , \sigMatrix[7][44] , \sigMatrix[7][43] ,
         \sigMatrix[7][42] , \sigMatrix[7][41] , \sigMatrix[7][40] ,
         \sigMatrix[7][39] , \sigMatrix[7][38] , \sigMatrix[7][37] ,
         \sigMatrix[7][36] , \sigMatrix[7][35] , \sigMatrix[7][34] ,
         \sigMatrix[7][33] , \sigMatrix[7][32] , \sigMatrix[7][31] ,
         \sigMatrix[7][30] , \sigMatrix[7][29] , \sigMatrix[7][28] ,
         \sigMatrix[7][27] , \sigMatrix[7][26] , \sigMatrix[7][25] ,
         \sigMatrix[7][24] , \sigMatrix[7][23] , \sigMatrix[7][22] ,
         \sigMatrix[7][21] , \sigMatrix[7][20] , \sigMatrix[7][19] ,
         \sigMatrix[7][18] , \sigMatrix[7][17] , \sigMatrix[7][16] ,
         \sigMatrix[7][15] , \sigMatrix[7][14] , \sigMatrix[7][13] ,
         \sigMatrix[7][12] , \sigMatrix[7][11] , \sigMatrix[7][10] ,
         \sigMatrix[7][9] , \sigMatrix[7][8] , \sigMatrix[7][7] ,
         \sigMatrix[7][6] , \sigMatrix[7][5] , \sigMatrix[7][4] ,
         \sigMatrix[7][3] , \sigMatrix[7][2] , \sigMatrix[7][1] ,
         \sigMatrix[7][0] , \sigMatrix[8][127] , \sigMatrix[8][126] ,
         \sigMatrix[8][125] , \sigMatrix[8][124] , \sigMatrix[8][123] ,
         \sigMatrix[8][122] , \sigMatrix[8][121] , \sigMatrix[8][120] ,
         \sigMatrix[8][119] , \sigMatrix[8][118] , \sigMatrix[8][117] ,
         \sigMatrix[8][116] , \sigMatrix[8][115] , \sigMatrix[8][114] ,
         \sigMatrix[8][113] , \sigMatrix[8][112] , \sigMatrix[8][111] ,
         \sigMatrix[8][110] , \sigMatrix[8][109] , \sigMatrix[8][108] ,
         \sigMatrix[8][107] , \sigMatrix[8][106] , \sigMatrix[8][105] ,
         \sigMatrix[8][104] , \sigMatrix[8][103] , \sigMatrix[8][102] ,
         \sigMatrix[8][101] , \sigMatrix[8][100] , \sigMatrix[8][99] ,
         \sigMatrix[8][98] , \sigMatrix[8][97] , \sigMatrix[8][96] ,
         \sigMatrix[8][95] , \sigMatrix[8][94] , \sigMatrix[8][93] ,
         \sigMatrix[8][92] , \sigMatrix[8][91] , \sigMatrix[8][90] ,
         \sigMatrix[8][89] , \sigMatrix[8][88] , \sigMatrix[8][87] ,
         \sigMatrix[8][86] , \sigMatrix[8][85] , \sigMatrix[8][84] ,
         \sigMatrix[8][83] , \sigMatrix[8][82] , \sigMatrix[8][81] ,
         \sigMatrix[8][80] , \sigMatrix[8][79] , \sigMatrix[8][78] ,
         \sigMatrix[8][77] , \sigMatrix[8][76] , \sigMatrix[8][75] ,
         \sigMatrix[8][74] , \sigMatrix[8][73] , \sigMatrix[8][72] ,
         \sigMatrix[8][71] , \sigMatrix[8][70] , \sigMatrix[8][69] ,
         \sigMatrix[8][68] , \sigMatrix[8][67] , \sigMatrix[8][66] ,
         \sigMatrix[8][65] , \sigMatrix[8][63] , \sigMatrix[8][62] ,
         \sigMatrix[8][61] , \sigMatrix[8][60] , \sigMatrix[8][59] ,
         \sigMatrix[8][58] , \sigMatrix[8][57] , \sigMatrix[8][56] ,
         \sigMatrix[8][55] , \sigMatrix[8][54] , \sigMatrix[8][53] ,
         \sigMatrix[8][52] , \sigMatrix[8][51] , \sigMatrix[8][50] ,
         \sigMatrix[8][49] , \sigMatrix[8][48] , \sigMatrix[8][47] ,
         \sigMatrix[8][46] , \sigMatrix[8][45] , \sigMatrix[8][44] ,
         \sigMatrix[8][43] , \sigMatrix[8][42] , \sigMatrix[8][41] ,
         \sigMatrix[8][40] , \sigMatrix[8][39] , \sigMatrix[8][38] ,
         \sigMatrix[8][37] , \sigMatrix[8][36] , \sigMatrix[8][35] ,
         \sigMatrix[8][34] , \sigMatrix[8][33] , \sigMatrix[8][32] ,
         \sigMatrix[8][31] , \sigMatrix[8][30] , \sigMatrix[8][29] ,
         \sigMatrix[8][28] , \sigMatrix[8][27] , \sigMatrix[8][26] ,
         \sigMatrix[8][25] , \sigMatrix[8][24] , \sigMatrix[8][23] ,
         \sigMatrix[8][22] , \sigMatrix[8][21] , \sigMatrix[8][20] ,
         \sigMatrix[8][19] , \sigMatrix[8][18] , \sigMatrix[8][17] ,
         \sigMatrix[8][16] , \sigMatrix[8][15] , \sigMatrix[8][14] ,
         \sigMatrix[8][13] , \sigMatrix[8][12] , \sigMatrix[8][11] ,
         \sigMatrix[8][10] , \sigMatrix[8][9] , \sigMatrix[8][8] ,
         \sigMatrix[8][7] , \sigMatrix[8][6] , \sigMatrix[8][5] ,
         \sigMatrix[8][4] , \sigMatrix[8][3] , \sigMatrix[8][2] ,
         \sigMatrix[8][1] , \sigMatrix[8][0] , \sigMatrix[9][127] ,
         \sigMatrix[9][126] , \sigMatrix[9][125] , \sigMatrix[9][124] ,
         \sigMatrix[9][123] , \sigMatrix[9][122] , \sigMatrix[9][121] ,
         \sigMatrix[9][120] , \sigMatrix[9][119] , \sigMatrix[9][118] ,
         \sigMatrix[9][117] , \sigMatrix[9][116] , \sigMatrix[9][115] ,
         \sigMatrix[9][114] , \sigMatrix[9][113] , \sigMatrix[9][112] ,
         \sigMatrix[9][111] , \sigMatrix[9][110] , \sigMatrix[9][109] ,
         \sigMatrix[9][108] , \sigMatrix[9][107] , \sigMatrix[9][106] ,
         \sigMatrix[9][105] , \sigMatrix[9][104] , \sigMatrix[9][103] ,
         \sigMatrix[9][102] , \sigMatrix[9][101] , \sigMatrix[9][100] ,
         \sigMatrix[9][99] , \sigMatrix[9][98] , \sigMatrix[9][97] ,
         \sigMatrix[9][96] , \sigMatrix[9][95] , \sigMatrix[9][94] ,
         \sigMatrix[9][93] , \sigMatrix[9][92] , \sigMatrix[9][91] ,
         \sigMatrix[9][90] , \sigMatrix[9][89] , \sigMatrix[9][88] ,
         \sigMatrix[9][87] , \sigMatrix[9][86] , \sigMatrix[9][85] ,
         \sigMatrix[9][84] , \sigMatrix[9][83] , \sigMatrix[9][82] ,
         \sigMatrix[9][81] , \sigMatrix[9][80] , \sigMatrix[9][79] ,
         \sigMatrix[9][78] , \sigMatrix[9][77] , \sigMatrix[9][76] ,
         \sigMatrix[9][75] , \sigMatrix[9][74] , \sigMatrix[9][73] ,
         \sigMatrix[9][72] , \sigMatrix[9][71] , \sigMatrix[9][70] ,
         \sigMatrix[9][69] , \sigMatrix[9][68] , \sigMatrix[9][67] ,
         \sigMatrix[9][66] , \sigMatrix[9][65] , \sigMatrix[9][63] ,
         \sigMatrix[9][62] , \sigMatrix[9][61] , \sigMatrix[9][60] ,
         \sigMatrix[9][59] , \sigMatrix[9][58] , \sigMatrix[9][57] ,
         \sigMatrix[9][56] , \sigMatrix[9][55] , \sigMatrix[9][54] ,
         \sigMatrix[9][53] , \sigMatrix[9][52] , \sigMatrix[9][51] ,
         \sigMatrix[9][50] , \sigMatrix[9][49] , \sigMatrix[9][48] ,
         \sigMatrix[9][47] , \sigMatrix[9][46] , \sigMatrix[9][45] ,
         \sigMatrix[9][44] , \sigMatrix[9][43] , \sigMatrix[9][42] ,
         \sigMatrix[9][41] , \sigMatrix[9][40] , \sigMatrix[9][39] ,
         \sigMatrix[9][38] , \sigMatrix[9][37] , \sigMatrix[9][36] ,
         \sigMatrix[9][35] , \sigMatrix[9][34] , \sigMatrix[9][33] ,
         \sigMatrix[9][32] , \sigMatrix[9][31] , \sigMatrix[9][30] ,
         \sigMatrix[9][29] , \sigMatrix[9][28] , \sigMatrix[9][27] ,
         \sigMatrix[9][26] , \sigMatrix[9][25] , \sigMatrix[9][24] ,
         \sigMatrix[9][23] , \sigMatrix[9][22] , \sigMatrix[9][21] ,
         \sigMatrix[9][20] , \sigMatrix[9][19] , \sigMatrix[9][18] ,
         \sigMatrix[9][17] , \sigMatrix[9][16] , \sigMatrix[9][15] ,
         \sigMatrix[9][14] , \sigMatrix[9][13] , \sigMatrix[9][12] ,
         \sigMatrix[9][11] , \sigMatrix[9][10] , \sigMatrix[9][9] ,
         \sigMatrix[9][8] , \sigMatrix[9][7] , \sigMatrix[9][6] ,
         \sigMatrix[9][5] , \sigMatrix[9][4] , \sigMatrix[9][3] ,
         \sigMatrix[9][2] , \sigMatrix[9][1] , \sigMatrix[9][0] ,
         \sigMatrix[10][127] , \sigMatrix[10][126] , \sigMatrix[10][125] ,
         \sigMatrix[10][124] , \sigMatrix[10][123] , \sigMatrix[10][122] ,
         \sigMatrix[10][121] , \sigMatrix[10][120] , \sigMatrix[10][119] ,
         \sigMatrix[10][118] , \sigMatrix[10][117] , \sigMatrix[10][116] ,
         \sigMatrix[10][115] , \sigMatrix[10][114] , \sigMatrix[10][113] ,
         \sigMatrix[10][112] , \sigMatrix[10][111] , \sigMatrix[10][110] ,
         \sigMatrix[10][109] , \sigMatrix[10][108] , \sigMatrix[10][107] ,
         \sigMatrix[10][106] , \sigMatrix[10][105] , \sigMatrix[10][104] ,
         \sigMatrix[10][103] , \sigMatrix[10][102] , \sigMatrix[10][101] ,
         \sigMatrix[10][100] , \sigMatrix[10][99] , \sigMatrix[10][98] ,
         \sigMatrix[10][97] , \sigMatrix[10][96] , \sigMatrix[10][95] ,
         \sigMatrix[10][94] , \sigMatrix[10][93] , \sigMatrix[10][92] ,
         \sigMatrix[10][91] , \sigMatrix[10][90] , \sigMatrix[10][89] ,
         \sigMatrix[10][88] , \sigMatrix[10][87] , \sigMatrix[10][86] ,
         \sigMatrix[10][85] , \sigMatrix[10][84] , \sigMatrix[10][83] ,
         \sigMatrix[10][82] , \sigMatrix[10][81] , \sigMatrix[10][80] ,
         \sigMatrix[10][79] , \sigMatrix[10][78] , \sigMatrix[10][77] ,
         \sigMatrix[10][76] , \sigMatrix[10][75] , \sigMatrix[10][74] ,
         \sigMatrix[10][73] , \sigMatrix[10][72] , \sigMatrix[10][71] ,
         \sigMatrix[10][70] , \sigMatrix[10][69] , \sigMatrix[10][68] ,
         \sigMatrix[10][67] , \sigMatrix[10][66] , \sigMatrix[10][65] ,
         \sigMatrix[10][63] , \sigMatrix[10][62] , \sigMatrix[10][61] ,
         \sigMatrix[10][60] , \sigMatrix[10][59] , \sigMatrix[10][58] ,
         \sigMatrix[10][57] , \sigMatrix[10][56] , \sigMatrix[10][55] ,
         \sigMatrix[10][54] , \sigMatrix[10][53] , \sigMatrix[10][52] ,
         \sigMatrix[10][51] , \sigMatrix[10][50] , \sigMatrix[10][49] ,
         \sigMatrix[10][48] , \sigMatrix[10][47] , \sigMatrix[10][46] ,
         \sigMatrix[10][45] , \sigMatrix[10][44] , \sigMatrix[10][43] ,
         \sigMatrix[10][42] , \sigMatrix[10][41] , \sigMatrix[10][40] ,
         \sigMatrix[10][39] , \sigMatrix[10][38] , \sigMatrix[10][37] ,
         \sigMatrix[10][36] , \sigMatrix[10][35] , \sigMatrix[10][34] ,
         \sigMatrix[10][33] , \sigMatrix[10][32] , \sigMatrix[10][31] ,
         \sigMatrix[10][30] , \sigMatrix[10][29] , \sigMatrix[10][28] ,
         \sigMatrix[10][27] , \sigMatrix[10][26] , \sigMatrix[10][25] ,
         \sigMatrix[10][24] , \sigMatrix[10][23] , \sigMatrix[10][22] ,
         \sigMatrix[10][21] , \sigMatrix[10][20] , \sigMatrix[10][19] ,
         \sigMatrix[10][18] , \sigMatrix[10][17] , \sigMatrix[10][16] ,
         \sigMatrix[10][15] , \sigMatrix[10][14] , \sigMatrix[10][13] ,
         \sigMatrix[10][12] , \sigMatrix[10][11] , \sigMatrix[10][10] ,
         \sigMatrix[10][9] , \sigMatrix[10][8] , \sigMatrix[10][7] ,
         \sigMatrix[10][6] , \sigMatrix[10][5] , \sigMatrix[10][4] ,
         \sigMatrix[10][3] , \sigMatrix[10][2] , \sigMatrix[10][1] ,
         \sigMatrix[10][0] , \sigMatrix[11][127] , \sigMatrix[11][126] ,
         \sigMatrix[11][125] , \sigMatrix[11][124] , \sigMatrix[11][123] ,
         \sigMatrix[11][122] , \sigMatrix[11][121] , \sigMatrix[11][120] ,
         \sigMatrix[11][119] , \sigMatrix[11][118] , \sigMatrix[11][117] ,
         \sigMatrix[11][116] , \sigMatrix[11][115] , \sigMatrix[11][114] ,
         \sigMatrix[11][113] , \sigMatrix[11][112] , \sigMatrix[11][111] ,
         \sigMatrix[11][110] , \sigMatrix[11][109] , \sigMatrix[11][108] ,
         \sigMatrix[11][107] , \sigMatrix[11][106] , \sigMatrix[11][105] ,
         \sigMatrix[11][104] , \sigMatrix[11][103] , \sigMatrix[11][102] ,
         \sigMatrix[11][101] , \sigMatrix[11][100] , \sigMatrix[11][99] ,
         \sigMatrix[11][98] , \sigMatrix[11][97] , \sigMatrix[11][96] ,
         \sigMatrix[11][95] , \sigMatrix[11][94] , \sigMatrix[11][93] ,
         \sigMatrix[11][92] , \sigMatrix[11][91] , \sigMatrix[11][90] ,
         \sigMatrix[11][89] , \sigMatrix[11][88] , \sigMatrix[11][87] ,
         \sigMatrix[11][86] , \sigMatrix[11][85] , \sigMatrix[11][84] ,
         \sigMatrix[11][83] , \sigMatrix[11][82] , \sigMatrix[11][81] ,
         \sigMatrix[11][80] , \sigMatrix[11][79] , \sigMatrix[11][78] ,
         \sigMatrix[11][77] , \sigMatrix[11][76] , \sigMatrix[11][75] ,
         \sigMatrix[11][74] , \sigMatrix[11][73] , \sigMatrix[11][72] ,
         \sigMatrix[11][71] , \sigMatrix[11][70] , \sigMatrix[11][69] ,
         \sigMatrix[11][68] , \sigMatrix[11][67] , \sigMatrix[11][66] ,
         \sigMatrix[11][65] , \sigMatrix[11][63] , \sigMatrix[11][62] ,
         \sigMatrix[11][61] , \sigMatrix[11][60] , \sigMatrix[11][59] ,
         \sigMatrix[11][58] , \sigMatrix[11][57] , \sigMatrix[11][56] ,
         \sigMatrix[11][55] , \sigMatrix[11][54] , \sigMatrix[11][53] ,
         \sigMatrix[11][52] , \sigMatrix[11][51] , \sigMatrix[11][50] ,
         \sigMatrix[11][49] , \sigMatrix[11][48] , \sigMatrix[11][47] ,
         \sigMatrix[11][46] , \sigMatrix[11][45] , \sigMatrix[11][44] ,
         \sigMatrix[11][43] , \sigMatrix[11][42] , \sigMatrix[11][41] ,
         \sigMatrix[11][40] , \sigMatrix[11][39] , \sigMatrix[11][38] ,
         \sigMatrix[11][37] , \sigMatrix[11][36] , \sigMatrix[11][35] ,
         \sigMatrix[11][34] , \sigMatrix[11][33] , \sigMatrix[11][32] ,
         \sigMatrix[11][31] , \sigMatrix[11][30] , \sigMatrix[11][29] ,
         \sigMatrix[11][28] , \sigMatrix[11][27] , \sigMatrix[11][26] ,
         \sigMatrix[11][25] , \sigMatrix[11][24] , \sigMatrix[11][23] ,
         \sigMatrix[11][22] , \sigMatrix[11][21] , \sigMatrix[11][20] ,
         \sigMatrix[11][19] , \sigMatrix[11][18] , \sigMatrix[11][17] ,
         \sigMatrix[11][16] , \sigMatrix[11][15] , \sigMatrix[11][14] ,
         \sigMatrix[11][13] , \sigMatrix[11][12] , \sigMatrix[11][11] ,
         \sigMatrix[11][10] , \sigMatrix[11][9] , \sigMatrix[11][8] ,
         \sigMatrix[11][7] , \sigMatrix[11][6] , \sigMatrix[11][5] ,
         \sigMatrix[11][4] , \sigMatrix[11][3] , \sigMatrix[11][2] ,
         \sigMatrix[11][1] , \sigMatrix[11][0] , \sigMatrix[12][127] ,
         \sigMatrix[12][126] , \sigMatrix[12][125] , \sigMatrix[12][124] ,
         \sigMatrix[12][123] , \sigMatrix[12][122] , \sigMatrix[12][121] ,
         \sigMatrix[12][120] , \sigMatrix[12][119] , \sigMatrix[12][118] ,
         \sigMatrix[12][117] , \sigMatrix[12][116] , \sigMatrix[12][115] ,
         \sigMatrix[12][114] , \sigMatrix[12][113] , \sigMatrix[12][112] ,
         \sigMatrix[12][111] , \sigMatrix[12][110] , \sigMatrix[12][109] ,
         \sigMatrix[12][108] , \sigMatrix[12][107] , \sigMatrix[12][106] ,
         \sigMatrix[12][105] , \sigMatrix[12][104] , \sigMatrix[12][103] ,
         \sigMatrix[12][102] , \sigMatrix[12][101] , \sigMatrix[12][100] ,
         \sigMatrix[12][99] , \sigMatrix[12][98] , \sigMatrix[12][97] ,
         \sigMatrix[12][96] , \sigMatrix[12][95] , \sigMatrix[12][94] ,
         \sigMatrix[12][93] , \sigMatrix[12][92] , \sigMatrix[12][91] ,
         \sigMatrix[12][90] , \sigMatrix[12][89] , \sigMatrix[12][88] ,
         \sigMatrix[12][87] , \sigMatrix[12][86] , \sigMatrix[12][85] ,
         \sigMatrix[12][84] , \sigMatrix[12][83] , \sigMatrix[12][82] ,
         \sigMatrix[12][81] , \sigMatrix[12][80] , \sigMatrix[12][79] ,
         \sigMatrix[12][78] , \sigMatrix[12][77] , \sigMatrix[12][76] ,
         \sigMatrix[12][75] , \sigMatrix[12][74] , \sigMatrix[12][73] ,
         \sigMatrix[12][72] , \sigMatrix[12][71] , \sigMatrix[12][70] ,
         \sigMatrix[12][69] , \sigMatrix[12][68] , \sigMatrix[12][67] ,
         \sigMatrix[12][66] , \sigMatrix[12][65] , \sigMatrix[12][63] ,
         \sigMatrix[12][62] , \sigMatrix[12][61] , \sigMatrix[12][60] ,
         \sigMatrix[12][59] , \sigMatrix[12][58] , \sigMatrix[12][57] ,
         \sigMatrix[12][56] , \sigMatrix[12][55] , \sigMatrix[12][54] ,
         \sigMatrix[12][53] , \sigMatrix[12][52] , \sigMatrix[12][51] ,
         \sigMatrix[12][50] , \sigMatrix[12][49] , \sigMatrix[12][48] ,
         \sigMatrix[12][47] , \sigMatrix[12][46] , \sigMatrix[12][45] ,
         \sigMatrix[12][44] , \sigMatrix[12][43] , \sigMatrix[12][42] ,
         \sigMatrix[12][41] , \sigMatrix[12][40] , \sigMatrix[12][39] ,
         \sigMatrix[12][38] , \sigMatrix[12][37] , \sigMatrix[12][36] ,
         \sigMatrix[12][35] , \sigMatrix[12][34] , \sigMatrix[12][33] ,
         \sigMatrix[12][32] , \sigMatrix[12][31] , \sigMatrix[12][30] ,
         \sigMatrix[12][29] , \sigMatrix[12][28] , \sigMatrix[12][27] ,
         \sigMatrix[12][26] , \sigMatrix[12][25] , \sigMatrix[12][24] ,
         \sigMatrix[12][23] , \sigMatrix[12][22] , \sigMatrix[12][21] ,
         \sigMatrix[12][20] , \sigMatrix[12][19] , \sigMatrix[12][18] ,
         \sigMatrix[12][17] , \sigMatrix[12][16] , \sigMatrix[12][15] ,
         \sigMatrix[12][14] , \sigMatrix[12][13] , \sigMatrix[12][12] ,
         \sigMatrix[12][11] , \sigMatrix[12][10] , \sigMatrix[12][9] ,
         \sigMatrix[12][8] , \sigMatrix[12][7] , \sigMatrix[12][6] ,
         \sigMatrix[12][5] , \sigMatrix[12][4] , \sigMatrix[12][3] ,
         \sigMatrix[12][2] , \sigMatrix[12][1] , \sigMatrix[12][0] ,
         \sigMatrix[13][127] , \sigMatrix[13][126] , \sigMatrix[13][125] ,
         \sigMatrix[13][124] , \sigMatrix[13][123] , \sigMatrix[13][122] ,
         \sigMatrix[13][121] , \sigMatrix[13][120] , \sigMatrix[13][119] ,
         \sigMatrix[13][118] , \sigMatrix[13][117] , \sigMatrix[13][116] ,
         \sigMatrix[13][115] , \sigMatrix[13][114] , \sigMatrix[13][113] ,
         \sigMatrix[13][112] , \sigMatrix[13][111] , \sigMatrix[13][110] ,
         \sigMatrix[13][109] , \sigMatrix[13][108] , \sigMatrix[13][107] ,
         \sigMatrix[13][106] , \sigMatrix[13][105] , \sigMatrix[13][104] ,
         \sigMatrix[13][103] , \sigMatrix[13][102] , \sigMatrix[13][101] ,
         \sigMatrix[13][100] , \sigMatrix[13][99] , \sigMatrix[13][98] ,
         \sigMatrix[13][97] , \sigMatrix[13][96] , \sigMatrix[13][95] ,
         \sigMatrix[13][94] , \sigMatrix[13][93] , \sigMatrix[13][92] ,
         \sigMatrix[13][91] , \sigMatrix[13][90] , \sigMatrix[13][89] ,
         \sigMatrix[13][88] , \sigMatrix[13][87] , \sigMatrix[13][86] ,
         \sigMatrix[13][85] , \sigMatrix[13][84] , \sigMatrix[13][83] ,
         \sigMatrix[13][82] , \sigMatrix[13][81] , \sigMatrix[13][80] ,
         \sigMatrix[13][79] , \sigMatrix[13][78] , \sigMatrix[13][77] ,
         \sigMatrix[13][76] , \sigMatrix[13][75] , \sigMatrix[13][74] ,
         \sigMatrix[13][73] , \sigMatrix[13][72] , \sigMatrix[13][71] ,
         \sigMatrix[13][70] , \sigMatrix[13][69] , \sigMatrix[13][68] ,
         \sigMatrix[13][67] , \sigMatrix[13][66] , \sigMatrix[13][65] ,
         \sigMatrix[13][63] , \sigMatrix[13][62] , \sigMatrix[13][61] ,
         \sigMatrix[13][60] , \sigMatrix[13][59] , \sigMatrix[13][58] ,
         \sigMatrix[13][57] , \sigMatrix[13][56] , \sigMatrix[13][55] ,
         \sigMatrix[13][54] , \sigMatrix[13][53] , \sigMatrix[13][52] ,
         \sigMatrix[13][51] , \sigMatrix[13][50] , \sigMatrix[13][49] ,
         \sigMatrix[13][48] , \sigMatrix[13][47] , \sigMatrix[13][46] ,
         \sigMatrix[13][45] , \sigMatrix[13][44] , \sigMatrix[13][43] ,
         \sigMatrix[13][42] , \sigMatrix[13][41] , \sigMatrix[13][40] ,
         \sigMatrix[13][39] , \sigMatrix[13][38] , \sigMatrix[13][37] ,
         \sigMatrix[13][36] , \sigMatrix[13][35] , \sigMatrix[13][34] ,
         \sigMatrix[13][33] , \sigMatrix[13][32] , \sigMatrix[13][31] ,
         \sigMatrix[13][30] , \sigMatrix[13][29] , \sigMatrix[13][28] ,
         \sigMatrix[13][27] , \sigMatrix[13][26] , \sigMatrix[13][25] ,
         \sigMatrix[13][24] , \sigMatrix[13][23] , \sigMatrix[13][22] ,
         \sigMatrix[13][21] , \sigMatrix[13][20] , \sigMatrix[13][19] ,
         \sigMatrix[13][18] , \sigMatrix[13][17] , \sigMatrix[13][16] ,
         \sigMatrix[13][15] , \sigMatrix[13][14] , \sigMatrix[13][13] ,
         \sigMatrix[13][12] , \sigMatrix[13][11] , \sigMatrix[13][10] ,
         \sigMatrix[13][9] , \sigMatrix[13][8] , \sigMatrix[13][7] ,
         \sigMatrix[13][6] , \sigMatrix[13][5] , \sigMatrix[13][4] ,
         \sigMatrix[13][3] , \sigMatrix[13][2] , \sigMatrix[13][1] ,
         \sigMatrix[13][0] , \sigMatrix[14][127] , \sigMatrix[14][126] ,
         \sigMatrix[14][125] , \sigMatrix[14][124] , \sigMatrix[14][123] ,
         \sigMatrix[14][122] , \sigMatrix[14][121] , \sigMatrix[14][120] ,
         \sigMatrix[14][119] , \sigMatrix[14][118] , \sigMatrix[14][117] ,
         \sigMatrix[14][116] , \sigMatrix[14][115] , \sigMatrix[14][114] ,
         \sigMatrix[14][113] , \sigMatrix[14][112] , \sigMatrix[14][111] ,
         \sigMatrix[14][110] , \sigMatrix[14][109] , \sigMatrix[14][108] ,
         \sigMatrix[14][107] , \sigMatrix[14][106] , \sigMatrix[14][105] ,
         \sigMatrix[14][104] , \sigMatrix[14][103] , \sigMatrix[14][102] ,
         \sigMatrix[14][101] , \sigMatrix[14][100] , \sigMatrix[14][99] ,
         \sigMatrix[14][98] , \sigMatrix[14][97] , \sigMatrix[14][96] ,
         \sigMatrix[14][95] , \sigMatrix[14][94] , \sigMatrix[14][93] ,
         \sigMatrix[14][92] , \sigMatrix[14][91] , \sigMatrix[14][90] ,
         \sigMatrix[14][89] , \sigMatrix[14][88] , \sigMatrix[14][87] ,
         \sigMatrix[14][86] , \sigMatrix[14][85] , \sigMatrix[14][84] ,
         \sigMatrix[14][83] , \sigMatrix[14][82] , \sigMatrix[14][81] ,
         \sigMatrix[14][80] , \sigMatrix[14][79] , \sigMatrix[14][78] ,
         \sigMatrix[14][77] , \sigMatrix[14][76] , \sigMatrix[14][75] ,
         \sigMatrix[14][74] , \sigMatrix[14][73] , \sigMatrix[14][72] ,
         \sigMatrix[14][71] , \sigMatrix[14][70] , \sigMatrix[14][69] ,
         \sigMatrix[14][68] , \sigMatrix[14][67] , \sigMatrix[14][66] ,
         \sigMatrix[14][65] , \sigMatrix[14][63] , \sigMatrix[14][62] ,
         \sigMatrix[14][61] , \sigMatrix[14][60] , \sigMatrix[14][59] ,
         \sigMatrix[14][58] , \sigMatrix[14][57] , \sigMatrix[14][56] ,
         \sigMatrix[14][55] , \sigMatrix[14][54] , \sigMatrix[14][53] ,
         \sigMatrix[14][52] , \sigMatrix[14][51] , \sigMatrix[14][50] ,
         \sigMatrix[14][49] , \sigMatrix[14][48] , \sigMatrix[14][47] ,
         \sigMatrix[14][46] , \sigMatrix[14][45] , \sigMatrix[14][44] ,
         \sigMatrix[14][43] , \sigMatrix[14][42] , \sigMatrix[14][41] ,
         \sigMatrix[14][40] , \sigMatrix[14][39] , \sigMatrix[14][38] ,
         \sigMatrix[14][37] , \sigMatrix[14][36] , \sigMatrix[14][35] ,
         \sigMatrix[14][34] , \sigMatrix[14][33] , \sigMatrix[14][32] ,
         \sigMatrix[14][31] , \sigMatrix[14][30] , \sigMatrix[14][29] ,
         \sigMatrix[14][28] , \sigMatrix[14][27] , \sigMatrix[14][26] ,
         \sigMatrix[14][25] , \sigMatrix[14][24] , \sigMatrix[14][23] ,
         \sigMatrix[14][22] , \sigMatrix[14][21] , \sigMatrix[14][20] ,
         \sigMatrix[14][19] , \sigMatrix[14][18] , \sigMatrix[14][17] ,
         \sigMatrix[14][16] , \sigMatrix[14][15] , \sigMatrix[14][14] ,
         \sigMatrix[14][13] , \sigMatrix[14][12] , \sigMatrix[14][11] ,
         \sigMatrix[14][10] , \sigMatrix[14][9] , \sigMatrix[14][8] ,
         \sigMatrix[14][7] , \sigMatrix[14][6] , \sigMatrix[14][5] ,
         \sigMatrix[14][4] , \sigMatrix[14][3] , \sigMatrix[14][2] ,
         \sigMatrix[14][1] , \sigMatrix[14][0] , n8, n9, n10, n11, n12, n13,
         n14, n15;
  wire   [31:0] A_out_s;
  wire   [31:0] B_out_s;
  wire   [63:0] P_s;
  tri   \sigMatrix[0][63] ;
  tri   \sigMatrix[0][62] ;
  tri   \sigMatrix[0][61] ;
  tri   \sigMatrix[0][60] ;
  tri   \sigMatrix[0][59] ;
  tri   \sigMatrix[0][58] ;
  tri   \sigMatrix[0][57] ;
  tri   \sigMatrix[0][56] ;
  tri   \sigMatrix[0][55] ;
  tri   \sigMatrix[0][54] ;
  tri   \sigMatrix[0][53] ;
  tri   \sigMatrix[0][52] ;
  tri   \sigMatrix[0][51] ;
  tri   \sigMatrix[0][50] ;
  tri   \sigMatrix[0][49] ;
  tri   \sigMatrix[0][48] ;
  tri   \sigMatrix[0][47] ;
  tri   \sigMatrix[0][46] ;
  tri   \sigMatrix[0][45] ;
  tri   \sigMatrix[0][44] ;
  tri   \sigMatrix[0][43] ;
  tri   \sigMatrix[0][42] ;
  tri   \sigMatrix[0][41] ;
  tri   \sigMatrix[0][40] ;
  tri   \sigMatrix[0][39] ;
  tri   \sigMatrix[0][38] ;
  tri   \sigMatrix[0][37] ;
  tri   \sigMatrix[0][36] ;
  tri   \sigMatrix[0][35] ;
  tri   \sigMatrix[0][34] ;
  tri   \sigMatrix[0][33] ;
  tri   \sigMatrix[0][32] ;
  tri   \sigMatrix[0][31] ;
  tri   \sigMatrix[0][30] ;
  tri   \sigMatrix[0][29] ;
  tri   \sigMatrix[0][28] ;
  tri   \sigMatrix[0][27] ;
  tri   \sigMatrix[0][26] ;
  tri   \sigMatrix[0][25] ;
  tri   \sigMatrix[0][24] ;
  tri   \sigMatrix[0][23] ;
  tri   \sigMatrix[0][22] ;
  tri   \sigMatrix[0][21] ;
  tri   \sigMatrix[0][20] ;
  tri   \sigMatrix[0][19] ;
  tri   \sigMatrix[0][18] ;
  tri   \sigMatrix[0][17] ;
  tri   \sigMatrix[0][16] ;
  tri   \sigMatrix[0][15] ;
  tri   \sigMatrix[0][14] ;
  tri   \sigMatrix[0][13] ;
  tri   \sigMatrix[0][12] ;
  tri   \sigMatrix[0][11] ;
  tri   \sigMatrix[0][10] ;
  tri   \sigMatrix[0][9] ;
  tri   \sigMatrix[0][8] ;
  tri   \sigMatrix[0][7] ;
  tri   \sigMatrix[0][6] ;
  tri   \sigMatrix[0][5] ;
  tri   \sigMatrix[0][4] ;
  tri   \sigMatrix[0][3] ;
  tri   \sigMatrix[0][2] ;
  tri   \sigMatrix[0][1] ;
  tri   \sigMatrix[0][0] ;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14;

  registers_N32_0 regs ( .Clk(Clk), .Rst(Rst), .A(A), .B(B), .A_out(A_out_s), 
        .B_out(B_out_s) );
  booth_mul_row_special_N64_RADIX3 booth_mul_row_special_1_0 ( .A({n11, n14, 
        n12, n13, n10, n15, n15, n14, n11, n10, n14, n15, n13, n13, n12, n15, 
        n13, n14, n12, n11, n10, n15, n14, n13, n11, n15, n14, n14, n12, n10, 
        n11, n15, n14, A_out_s[30:0]}), .encoderIn({B_out_s[1:0], 1'b0}), 
        .nextA({\sigMatrix[0][127] , \sigMatrix[0][126] , \sigMatrix[0][125] , 
        \sigMatrix[0][124] , \sigMatrix[0][123] , \sigMatrix[0][122] , 
        \sigMatrix[0][121] , \sigMatrix[0][120] , \sigMatrix[0][119] , 
        \sigMatrix[0][118] , \sigMatrix[0][117] , \sigMatrix[0][116] , 
        \sigMatrix[0][115] , \sigMatrix[0][114] , \sigMatrix[0][113] , 
        \sigMatrix[0][112] , \sigMatrix[0][111] , \sigMatrix[0][110] , 
        \sigMatrix[0][109] , \sigMatrix[0][108] , \sigMatrix[0][107] , 
        \sigMatrix[0][106] , \sigMatrix[0][105] , \sigMatrix[0][104] , 
        \sigMatrix[0][103] , \sigMatrix[0][102] , \sigMatrix[0][101] , 
        \sigMatrix[0][100] , \sigMatrix[0][99] , \sigMatrix[0][98] , 
        \sigMatrix[0][97] , \sigMatrix[0][96] , \sigMatrix[0][95] , 
        \sigMatrix[0][94] , \sigMatrix[0][93] , \sigMatrix[0][92] , 
        \sigMatrix[0][91] , \sigMatrix[0][90] , \sigMatrix[0][89] , 
        \sigMatrix[0][88] , \sigMatrix[0][87] , \sigMatrix[0][86] , 
        \sigMatrix[0][85] , \sigMatrix[0][84] , \sigMatrix[0][83] , 
        \sigMatrix[0][82] , \sigMatrix[0][81] , \sigMatrix[0][80] , 
        \sigMatrix[0][79] , \sigMatrix[0][78] , \sigMatrix[0][77] , 
        \sigMatrix[0][76] , \sigMatrix[0][75] , \sigMatrix[0][74] , 
        \sigMatrix[0][73] , \sigMatrix[0][72] , \sigMatrix[0][71] , 
        \sigMatrix[0][70] , \sigMatrix[0][69] , \sigMatrix[0][68] , 
        \sigMatrix[0][67] , \sigMatrix[0][66] , \sigMatrix[0][65] , 
        SYNOPSYS_UNCONNECTED__0}), .nextSum({\sigMatrix[0][63] , 
        \sigMatrix[0][62] , \sigMatrix[0][61] , \sigMatrix[0][60] , 
        \sigMatrix[0][59] , \sigMatrix[0][58] , \sigMatrix[0][57] , 
        \sigMatrix[0][56] , \sigMatrix[0][55] , \sigMatrix[0][54] , 
        \sigMatrix[0][53] , \sigMatrix[0][52] , \sigMatrix[0][51] , 
        \sigMatrix[0][50] , \sigMatrix[0][49] , \sigMatrix[0][48] , 
        \sigMatrix[0][47] , \sigMatrix[0][46] , \sigMatrix[0][45] , 
        \sigMatrix[0][44] , \sigMatrix[0][43] , \sigMatrix[0][42] , 
        \sigMatrix[0][41] , \sigMatrix[0][40] , \sigMatrix[0][39] , 
        \sigMatrix[0][38] , \sigMatrix[0][37] , \sigMatrix[0][36] , 
        \sigMatrix[0][35] , \sigMatrix[0][34] , \sigMatrix[0][33] , 
        \sigMatrix[0][32] , \sigMatrix[0][31] , \sigMatrix[0][30] , 
        \sigMatrix[0][29] , \sigMatrix[0][28] , \sigMatrix[0][27] , 
        \sigMatrix[0][26] , \sigMatrix[0][25] , \sigMatrix[0][24] , 
        \sigMatrix[0][23] , \sigMatrix[0][22] , \sigMatrix[0][21] , 
        \sigMatrix[0][20] , \sigMatrix[0][19] , \sigMatrix[0][18] , 
        \sigMatrix[0][17] , \sigMatrix[0][16] , \sigMatrix[0][15] , 
        \sigMatrix[0][14] , \sigMatrix[0][13] , \sigMatrix[0][12] , 
        \sigMatrix[0][11] , \sigMatrix[0][10] , \sigMatrix[0][9] , 
        \sigMatrix[0][8] , \sigMatrix[0][7] , \sigMatrix[0][6] , 
        \sigMatrix[0][5] , \sigMatrix[0][4] , \sigMatrix[0][3] , 
        \sigMatrix[0][2] , \sigMatrix[0][1] , \sigMatrix[0][0] }) );
  booth_mul_row_N64_RADIX3_0 booth_mul_row_1_1 ( .prevA({\sigMatrix[0][127] , 
        \sigMatrix[0][126] , \sigMatrix[0][125] , \sigMatrix[0][124] , 
        \sigMatrix[0][123] , \sigMatrix[0][122] , \sigMatrix[0][121] , 
        \sigMatrix[0][120] , \sigMatrix[0][119] , \sigMatrix[0][118] , 
        \sigMatrix[0][117] , \sigMatrix[0][116] , \sigMatrix[0][115] , 
        \sigMatrix[0][114] , \sigMatrix[0][113] , \sigMatrix[0][112] , 
        \sigMatrix[0][111] , \sigMatrix[0][110] , \sigMatrix[0][109] , 
        \sigMatrix[0][108] , \sigMatrix[0][107] , \sigMatrix[0][106] , 
        \sigMatrix[0][105] , \sigMatrix[0][104] , \sigMatrix[0][103] , 
        \sigMatrix[0][102] , \sigMatrix[0][101] , \sigMatrix[0][100] , 
        \sigMatrix[0][99] , \sigMatrix[0][98] , \sigMatrix[0][97] , 
        \sigMatrix[0][96] , \sigMatrix[0][95] , \sigMatrix[0][94] , 
        \sigMatrix[0][93] , \sigMatrix[0][92] , \sigMatrix[0][91] , 
        \sigMatrix[0][90] , \sigMatrix[0][89] , \sigMatrix[0][88] , 
        \sigMatrix[0][87] , \sigMatrix[0][86] , \sigMatrix[0][85] , 
        \sigMatrix[0][84] , \sigMatrix[0][83] , \sigMatrix[0][82] , 
        \sigMatrix[0][81] , \sigMatrix[0][80] , \sigMatrix[0][79] , 
        \sigMatrix[0][78] , \sigMatrix[0][77] , \sigMatrix[0][76] , 
        \sigMatrix[0][75] , \sigMatrix[0][74] , \sigMatrix[0][73] , 
        \sigMatrix[0][72] , \sigMatrix[0][71] , \sigMatrix[0][70] , 
        \sigMatrix[0][69] , \sigMatrix[0][68] , \sigMatrix[0][67] , 
        \sigMatrix[0][66] , \sigMatrix[0][65] , 1'b0}), .prevSum({
        \sigMatrix[0][63] , \sigMatrix[0][62] , \sigMatrix[0][61] , 
        \sigMatrix[0][60] , \sigMatrix[0][59] , \sigMatrix[0][58] , 
        \sigMatrix[0][57] , \sigMatrix[0][56] , \sigMatrix[0][55] , 
        \sigMatrix[0][54] , \sigMatrix[0][53] , \sigMatrix[0][52] , 
        \sigMatrix[0][51] , \sigMatrix[0][50] , \sigMatrix[0][49] , 
        \sigMatrix[0][48] , \sigMatrix[0][47] , \sigMatrix[0][46] , 
        \sigMatrix[0][45] , \sigMatrix[0][44] , \sigMatrix[0][43] , 
        \sigMatrix[0][42] , \sigMatrix[0][41] , \sigMatrix[0][40] , 
        \sigMatrix[0][39] , \sigMatrix[0][38] , \sigMatrix[0][37] , 
        \sigMatrix[0][36] , \sigMatrix[0][35] , \sigMatrix[0][34] , 
        \sigMatrix[0][33] , \sigMatrix[0][32] , \sigMatrix[0][31] , 
        \sigMatrix[0][30] , \sigMatrix[0][29] , \sigMatrix[0][28] , 
        \sigMatrix[0][27] , \sigMatrix[0][26] , \sigMatrix[0][25] , 
        \sigMatrix[0][24] , \sigMatrix[0][23] , \sigMatrix[0][22] , 
        \sigMatrix[0][21] , \sigMatrix[0][20] , \sigMatrix[0][19] , 
        \sigMatrix[0][18] , \sigMatrix[0][17] , \sigMatrix[0][16] , 
        \sigMatrix[0][15] , \sigMatrix[0][14] , \sigMatrix[0][13] , 
        \sigMatrix[0][12] , \sigMatrix[0][11] , \sigMatrix[0][10] , 
        \sigMatrix[0][9] , \sigMatrix[0][8] , \sigMatrix[0][7] , 
        \sigMatrix[0][6] , \sigMatrix[0][5] , \sigMatrix[0][4] , 
        \sigMatrix[0][3] , \sigMatrix[0][2] , \sigMatrix[0][1] , 
        \sigMatrix[0][0] }), .encoderIn(B_out_s[3:1]), .nextA({
        \sigMatrix[1][127] , \sigMatrix[1][126] , \sigMatrix[1][125] , 
        \sigMatrix[1][124] , \sigMatrix[1][123] , \sigMatrix[1][122] , 
        \sigMatrix[1][121] , \sigMatrix[1][120] , \sigMatrix[1][119] , 
        \sigMatrix[1][118] , \sigMatrix[1][117] , \sigMatrix[1][116] , 
        \sigMatrix[1][115] , \sigMatrix[1][114] , \sigMatrix[1][113] , 
        \sigMatrix[1][112] , \sigMatrix[1][111] , \sigMatrix[1][110] , 
        \sigMatrix[1][109] , \sigMatrix[1][108] , \sigMatrix[1][107] , 
        \sigMatrix[1][106] , \sigMatrix[1][105] , \sigMatrix[1][104] , 
        \sigMatrix[1][103] , \sigMatrix[1][102] , \sigMatrix[1][101] , 
        \sigMatrix[1][100] , \sigMatrix[1][99] , \sigMatrix[1][98] , 
        \sigMatrix[1][97] , \sigMatrix[1][96] , \sigMatrix[1][95] , 
        \sigMatrix[1][94] , \sigMatrix[1][93] , \sigMatrix[1][92] , 
        \sigMatrix[1][91] , \sigMatrix[1][90] , \sigMatrix[1][89] , 
        \sigMatrix[1][88] , \sigMatrix[1][87] , \sigMatrix[1][86] , 
        \sigMatrix[1][85] , \sigMatrix[1][84] , \sigMatrix[1][83] , 
        \sigMatrix[1][82] , \sigMatrix[1][81] , \sigMatrix[1][80] , 
        \sigMatrix[1][79] , \sigMatrix[1][78] , \sigMatrix[1][77] , 
        \sigMatrix[1][76] , \sigMatrix[1][75] , \sigMatrix[1][74] , 
        \sigMatrix[1][73] , \sigMatrix[1][72] , \sigMatrix[1][71] , 
        \sigMatrix[1][70] , \sigMatrix[1][69] , \sigMatrix[1][68] , 
        \sigMatrix[1][67] , \sigMatrix[1][66] , \sigMatrix[1][65] , 
        SYNOPSYS_UNCONNECTED__1}), .nextSum({\sigMatrix[1][63] , 
        \sigMatrix[1][62] , \sigMatrix[1][61] , \sigMatrix[1][60] , 
        \sigMatrix[1][59] , \sigMatrix[1][58] , \sigMatrix[1][57] , 
        \sigMatrix[1][56] , \sigMatrix[1][55] , \sigMatrix[1][54] , 
        \sigMatrix[1][53] , \sigMatrix[1][52] , \sigMatrix[1][51] , 
        \sigMatrix[1][50] , \sigMatrix[1][49] , \sigMatrix[1][48] , 
        \sigMatrix[1][47] , \sigMatrix[1][46] , \sigMatrix[1][45] , 
        \sigMatrix[1][44] , \sigMatrix[1][43] , \sigMatrix[1][42] , 
        \sigMatrix[1][41] , \sigMatrix[1][40] , \sigMatrix[1][39] , 
        \sigMatrix[1][38] , \sigMatrix[1][37] , \sigMatrix[1][36] , 
        \sigMatrix[1][35] , \sigMatrix[1][34] , \sigMatrix[1][33] , 
        \sigMatrix[1][32] , \sigMatrix[1][31] , \sigMatrix[1][30] , 
        \sigMatrix[1][29] , \sigMatrix[1][28] , \sigMatrix[1][27] , 
        \sigMatrix[1][26] , \sigMatrix[1][25] , \sigMatrix[1][24] , 
        \sigMatrix[1][23] , \sigMatrix[1][22] , \sigMatrix[1][21] , 
        \sigMatrix[1][20] , \sigMatrix[1][19] , \sigMatrix[1][18] , 
        \sigMatrix[1][17] , \sigMatrix[1][16] , \sigMatrix[1][15] , 
        \sigMatrix[1][14] , \sigMatrix[1][13] , \sigMatrix[1][12] , 
        \sigMatrix[1][11] , \sigMatrix[1][10] , \sigMatrix[1][9] , 
        \sigMatrix[1][8] , \sigMatrix[1][7] , \sigMatrix[1][6] , 
        \sigMatrix[1][5] , \sigMatrix[1][4] , \sigMatrix[1][3] , 
        \sigMatrix[1][2] , \sigMatrix[1][1] , \sigMatrix[1][0] }) );
  booth_mul_row_N64_RADIX3_14 booth_mul_row_1_2 ( .prevA({\sigMatrix[1][127] , 
        \sigMatrix[1][126] , \sigMatrix[1][125] , \sigMatrix[1][124] , 
        \sigMatrix[1][123] , \sigMatrix[1][122] , \sigMatrix[1][121] , 
        \sigMatrix[1][120] , \sigMatrix[1][119] , \sigMatrix[1][118] , 
        \sigMatrix[1][117] , \sigMatrix[1][116] , \sigMatrix[1][115] , 
        \sigMatrix[1][114] , \sigMatrix[1][113] , \sigMatrix[1][112] , 
        \sigMatrix[1][111] , \sigMatrix[1][110] , \sigMatrix[1][109] , 
        \sigMatrix[1][108] , \sigMatrix[1][107] , \sigMatrix[1][106] , 
        \sigMatrix[1][105] , \sigMatrix[1][104] , \sigMatrix[1][103] , 
        \sigMatrix[1][102] , \sigMatrix[1][101] , \sigMatrix[1][100] , 
        \sigMatrix[1][99] , \sigMatrix[1][98] , \sigMatrix[1][97] , 
        \sigMatrix[1][96] , \sigMatrix[1][95] , \sigMatrix[1][94] , 
        \sigMatrix[1][93] , \sigMatrix[1][92] , \sigMatrix[1][91] , 
        \sigMatrix[1][90] , \sigMatrix[1][89] , \sigMatrix[1][88] , 
        \sigMatrix[1][87] , \sigMatrix[1][86] , \sigMatrix[1][85] , 
        \sigMatrix[1][84] , \sigMatrix[1][83] , \sigMatrix[1][82] , 
        \sigMatrix[1][81] , \sigMatrix[1][80] , \sigMatrix[1][79] , 
        \sigMatrix[1][78] , \sigMatrix[1][77] , \sigMatrix[1][76] , 
        \sigMatrix[1][75] , \sigMatrix[1][74] , \sigMatrix[1][73] , 
        \sigMatrix[1][72] , \sigMatrix[1][71] , \sigMatrix[1][70] , 
        \sigMatrix[1][69] , \sigMatrix[1][68] , \sigMatrix[1][67] , 
        \sigMatrix[1][66] , \sigMatrix[1][65] , 1'b0}), .prevSum({
        \sigMatrix[1][63] , \sigMatrix[1][62] , \sigMatrix[1][61] , 
        \sigMatrix[1][60] , \sigMatrix[1][59] , \sigMatrix[1][58] , 
        \sigMatrix[1][57] , \sigMatrix[1][56] , \sigMatrix[1][55] , 
        \sigMatrix[1][54] , \sigMatrix[1][53] , \sigMatrix[1][52] , 
        \sigMatrix[1][51] , \sigMatrix[1][50] , \sigMatrix[1][49] , 
        \sigMatrix[1][48] , \sigMatrix[1][47] , \sigMatrix[1][46] , 
        \sigMatrix[1][45] , \sigMatrix[1][44] , \sigMatrix[1][43] , 
        \sigMatrix[1][42] , \sigMatrix[1][41] , \sigMatrix[1][40] , 
        \sigMatrix[1][39] , \sigMatrix[1][38] , \sigMatrix[1][37] , 
        \sigMatrix[1][36] , \sigMatrix[1][35] , \sigMatrix[1][34] , 
        \sigMatrix[1][33] , \sigMatrix[1][32] , \sigMatrix[1][31] , 
        \sigMatrix[1][30] , \sigMatrix[1][29] , \sigMatrix[1][28] , 
        \sigMatrix[1][27] , \sigMatrix[1][26] , \sigMatrix[1][25] , 
        \sigMatrix[1][24] , \sigMatrix[1][23] , \sigMatrix[1][22] , 
        \sigMatrix[1][21] , \sigMatrix[1][20] , \sigMatrix[1][19] , 
        \sigMatrix[1][18] , \sigMatrix[1][17] , \sigMatrix[1][16] , 
        \sigMatrix[1][15] , \sigMatrix[1][14] , \sigMatrix[1][13] , 
        \sigMatrix[1][12] , \sigMatrix[1][11] , \sigMatrix[1][10] , 
        \sigMatrix[1][9] , \sigMatrix[1][8] , \sigMatrix[1][7] , 
        \sigMatrix[1][6] , \sigMatrix[1][5] , \sigMatrix[1][4] , 
        \sigMatrix[1][3] , \sigMatrix[1][2] , \sigMatrix[1][1] , 
        \sigMatrix[1][0] }), .encoderIn(B_out_s[5:3]), .nextA({
        \sigMatrix[2][127] , \sigMatrix[2][126] , \sigMatrix[2][125] , 
        \sigMatrix[2][124] , \sigMatrix[2][123] , \sigMatrix[2][122] , 
        \sigMatrix[2][121] , \sigMatrix[2][120] , \sigMatrix[2][119] , 
        \sigMatrix[2][118] , \sigMatrix[2][117] , \sigMatrix[2][116] , 
        \sigMatrix[2][115] , \sigMatrix[2][114] , \sigMatrix[2][113] , 
        \sigMatrix[2][112] , \sigMatrix[2][111] , \sigMatrix[2][110] , 
        \sigMatrix[2][109] , \sigMatrix[2][108] , \sigMatrix[2][107] , 
        \sigMatrix[2][106] , \sigMatrix[2][105] , \sigMatrix[2][104] , 
        \sigMatrix[2][103] , \sigMatrix[2][102] , \sigMatrix[2][101] , 
        \sigMatrix[2][100] , \sigMatrix[2][99] , \sigMatrix[2][98] , 
        \sigMatrix[2][97] , \sigMatrix[2][96] , \sigMatrix[2][95] , 
        \sigMatrix[2][94] , \sigMatrix[2][93] , \sigMatrix[2][92] , 
        \sigMatrix[2][91] , \sigMatrix[2][90] , \sigMatrix[2][89] , 
        \sigMatrix[2][88] , \sigMatrix[2][87] , \sigMatrix[2][86] , 
        \sigMatrix[2][85] , \sigMatrix[2][84] , \sigMatrix[2][83] , 
        \sigMatrix[2][82] , \sigMatrix[2][81] , \sigMatrix[2][80] , 
        \sigMatrix[2][79] , \sigMatrix[2][78] , \sigMatrix[2][77] , 
        \sigMatrix[2][76] , \sigMatrix[2][75] , \sigMatrix[2][74] , 
        \sigMatrix[2][73] , \sigMatrix[2][72] , \sigMatrix[2][71] , 
        \sigMatrix[2][70] , \sigMatrix[2][69] , \sigMatrix[2][68] , 
        \sigMatrix[2][67] , \sigMatrix[2][66] , \sigMatrix[2][65] , 
        SYNOPSYS_UNCONNECTED__2}), .nextSum({\sigMatrix[2][63] , 
        \sigMatrix[2][62] , \sigMatrix[2][61] , \sigMatrix[2][60] , 
        \sigMatrix[2][59] , \sigMatrix[2][58] , \sigMatrix[2][57] , 
        \sigMatrix[2][56] , \sigMatrix[2][55] , \sigMatrix[2][54] , 
        \sigMatrix[2][53] , \sigMatrix[2][52] , \sigMatrix[2][51] , 
        \sigMatrix[2][50] , \sigMatrix[2][49] , \sigMatrix[2][48] , 
        \sigMatrix[2][47] , \sigMatrix[2][46] , \sigMatrix[2][45] , 
        \sigMatrix[2][44] , \sigMatrix[2][43] , \sigMatrix[2][42] , 
        \sigMatrix[2][41] , \sigMatrix[2][40] , \sigMatrix[2][39] , 
        \sigMatrix[2][38] , \sigMatrix[2][37] , \sigMatrix[2][36] , 
        \sigMatrix[2][35] , \sigMatrix[2][34] , \sigMatrix[2][33] , 
        \sigMatrix[2][32] , \sigMatrix[2][31] , \sigMatrix[2][30] , 
        \sigMatrix[2][29] , \sigMatrix[2][28] , \sigMatrix[2][27] , 
        \sigMatrix[2][26] , \sigMatrix[2][25] , \sigMatrix[2][24] , 
        \sigMatrix[2][23] , \sigMatrix[2][22] , \sigMatrix[2][21] , 
        \sigMatrix[2][20] , \sigMatrix[2][19] , \sigMatrix[2][18] , 
        \sigMatrix[2][17] , \sigMatrix[2][16] , \sigMatrix[2][15] , 
        \sigMatrix[2][14] , \sigMatrix[2][13] , \sigMatrix[2][12] , 
        \sigMatrix[2][11] , \sigMatrix[2][10] , \sigMatrix[2][9] , 
        \sigMatrix[2][8] , \sigMatrix[2][7] , \sigMatrix[2][6] , 
        \sigMatrix[2][5] , \sigMatrix[2][4] , \sigMatrix[2][3] , 
        \sigMatrix[2][2] , \sigMatrix[2][1] , \sigMatrix[2][0] }) );
  booth_mul_row_N64_RADIX3_13 booth_mul_row_1_3 ( .prevA({\sigMatrix[2][127] , 
        \sigMatrix[2][126] , \sigMatrix[2][125] , \sigMatrix[2][124] , 
        \sigMatrix[2][123] , \sigMatrix[2][122] , \sigMatrix[2][121] , 
        \sigMatrix[2][120] , \sigMatrix[2][119] , \sigMatrix[2][118] , 
        \sigMatrix[2][117] , \sigMatrix[2][116] , \sigMatrix[2][115] , 
        \sigMatrix[2][114] , \sigMatrix[2][113] , \sigMatrix[2][112] , 
        \sigMatrix[2][111] , \sigMatrix[2][110] , \sigMatrix[2][109] , 
        \sigMatrix[2][108] , \sigMatrix[2][107] , \sigMatrix[2][106] , 
        \sigMatrix[2][105] , \sigMatrix[2][104] , \sigMatrix[2][103] , 
        \sigMatrix[2][102] , \sigMatrix[2][101] , \sigMatrix[2][100] , 
        \sigMatrix[2][99] , \sigMatrix[2][98] , \sigMatrix[2][97] , 
        \sigMatrix[2][96] , \sigMatrix[2][95] , \sigMatrix[2][94] , 
        \sigMatrix[2][93] , \sigMatrix[2][92] , \sigMatrix[2][91] , 
        \sigMatrix[2][90] , \sigMatrix[2][89] , \sigMatrix[2][88] , 
        \sigMatrix[2][87] , \sigMatrix[2][86] , \sigMatrix[2][85] , 
        \sigMatrix[2][84] , \sigMatrix[2][83] , \sigMatrix[2][82] , 
        \sigMatrix[2][81] , \sigMatrix[2][80] , \sigMatrix[2][79] , 
        \sigMatrix[2][78] , \sigMatrix[2][77] , \sigMatrix[2][76] , 
        \sigMatrix[2][75] , \sigMatrix[2][74] , \sigMatrix[2][73] , 
        \sigMatrix[2][72] , \sigMatrix[2][71] , \sigMatrix[2][70] , 
        \sigMatrix[2][69] , \sigMatrix[2][68] , \sigMatrix[2][67] , 
        \sigMatrix[2][66] , \sigMatrix[2][65] , 1'b0}), .prevSum({
        \sigMatrix[2][63] , \sigMatrix[2][62] , \sigMatrix[2][61] , 
        \sigMatrix[2][60] , \sigMatrix[2][59] , \sigMatrix[2][58] , 
        \sigMatrix[2][57] , \sigMatrix[2][56] , \sigMatrix[2][55] , 
        \sigMatrix[2][54] , \sigMatrix[2][53] , \sigMatrix[2][52] , 
        \sigMatrix[2][51] , \sigMatrix[2][50] , \sigMatrix[2][49] , 
        \sigMatrix[2][48] , \sigMatrix[2][47] , \sigMatrix[2][46] , 
        \sigMatrix[2][45] , \sigMatrix[2][44] , \sigMatrix[2][43] , 
        \sigMatrix[2][42] , \sigMatrix[2][41] , \sigMatrix[2][40] , 
        \sigMatrix[2][39] , \sigMatrix[2][38] , \sigMatrix[2][37] , 
        \sigMatrix[2][36] , \sigMatrix[2][35] , \sigMatrix[2][34] , 
        \sigMatrix[2][33] , \sigMatrix[2][32] , \sigMatrix[2][31] , 
        \sigMatrix[2][30] , \sigMatrix[2][29] , \sigMatrix[2][28] , 
        \sigMatrix[2][27] , \sigMatrix[2][26] , \sigMatrix[2][25] , 
        \sigMatrix[2][24] , \sigMatrix[2][23] , \sigMatrix[2][22] , 
        \sigMatrix[2][21] , \sigMatrix[2][20] , \sigMatrix[2][19] , 
        \sigMatrix[2][18] , \sigMatrix[2][17] , \sigMatrix[2][16] , 
        \sigMatrix[2][15] , \sigMatrix[2][14] , \sigMatrix[2][13] , 
        \sigMatrix[2][12] , \sigMatrix[2][11] , \sigMatrix[2][10] , 
        \sigMatrix[2][9] , \sigMatrix[2][8] , \sigMatrix[2][7] , 
        \sigMatrix[2][6] , \sigMatrix[2][5] , \sigMatrix[2][4] , 
        \sigMatrix[2][3] , \sigMatrix[2][2] , \sigMatrix[2][1] , 
        \sigMatrix[2][0] }), .encoderIn(B_out_s[7:5]), .nextA({
        \sigMatrix[3][127] , \sigMatrix[3][126] , \sigMatrix[3][125] , 
        \sigMatrix[3][124] , \sigMatrix[3][123] , \sigMatrix[3][122] , 
        \sigMatrix[3][121] , \sigMatrix[3][120] , \sigMatrix[3][119] , 
        \sigMatrix[3][118] , \sigMatrix[3][117] , \sigMatrix[3][116] , 
        \sigMatrix[3][115] , \sigMatrix[3][114] , \sigMatrix[3][113] , 
        \sigMatrix[3][112] , \sigMatrix[3][111] , \sigMatrix[3][110] , 
        \sigMatrix[3][109] , \sigMatrix[3][108] , \sigMatrix[3][107] , 
        \sigMatrix[3][106] , \sigMatrix[3][105] , \sigMatrix[3][104] , 
        \sigMatrix[3][103] , \sigMatrix[3][102] , \sigMatrix[3][101] , 
        \sigMatrix[3][100] , \sigMatrix[3][99] , \sigMatrix[3][98] , 
        \sigMatrix[3][97] , \sigMatrix[3][96] , \sigMatrix[3][95] , 
        \sigMatrix[3][94] , \sigMatrix[3][93] , \sigMatrix[3][92] , 
        \sigMatrix[3][91] , \sigMatrix[3][90] , \sigMatrix[3][89] , 
        \sigMatrix[3][88] , \sigMatrix[3][87] , \sigMatrix[3][86] , 
        \sigMatrix[3][85] , \sigMatrix[3][84] , \sigMatrix[3][83] , 
        \sigMatrix[3][82] , \sigMatrix[3][81] , \sigMatrix[3][80] , 
        \sigMatrix[3][79] , \sigMatrix[3][78] , \sigMatrix[3][77] , 
        \sigMatrix[3][76] , \sigMatrix[3][75] , \sigMatrix[3][74] , 
        \sigMatrix[3][73] , \sigMatrix[3][72] , \sigMatrix[3][71] , 
        \sigMatrix[3][70] , \sigMatrix[3][69] , \sigMatrix[3][68] , 
        \sigMatrix[3][67] , \sigMatrix[3][66] , \sigMatrix[3][65] , 
        SYNOPSYS_UNCONNECTED__3}), .nextSum({\sigMatrix[3][63] , 
        \sigMatrix[3][62] , \sigMatrix[3][61] , \sigMatrix[3][60] , 
        \sigMatrix[3][59] , \sigMatrix[3][58] , \sigMatrix[3][57] , 
        \sigMatrix[3][56] , \sigMatrix[3][55] , \sigMatrix[3][54] , 
        \sigMatrix[3][53] , \sigMatrix[3][52] , \sigMatrix[3][51] , 
        \sigMatrix[3][50] , \sigMatrix[3][49] , \sigMatrix[3][48] , 
        \sigMatrix[3][47] , \sigMatrix[3][46] , \sigMatrix[3][45] , 
        \sigMatrix[3][44] , \sigMatrix[3][43] , \sigMatrix[3][42] , 
        \sigMatrix[3][41] , \sigMatrix[3][40] , \sigMatrix[3][39] , 
        \sigMatrix[3][38] , \sigMatrix[3][37] , \sigMatrix[3][36] , 
        \sigMatrix[3][35] , \sigMatrix[3][34] , \sigMatrix[3][33] , 
        \sigMatrix[3][32] , \sigMatrix[3][31] , \sigMatrix[3][30] , 
        \sigMatrix[3][29] , \sigMatrix[3][28] , \sigMatrix[3][27] , 
        \sigMatrix[3][26] , \sigMatrix[3][25] , \sigMatrix[3][24] , 
        \sigMatrix[3][23] , \sigMatrix[3][22] , \sigMatrix[3][21] , 
        \sigMatrix[3][20] , \sigMatrix[3][19] , \sigMatrix[3][18] , 
        \sigMatrix[3][17] , \sigMatrix[3][16] , \sigMatrix[3][15] , 
        \sigMatrix[3][14] , \sigMatrix[3][13] , \sigMatrix[3][12] , 
        \sigMatrix[3][11] , \sigMatrix[3][10] , \sigMatrix[3][9] , 
        \sigMatrix[3][8] , \sigMatrix[3][7] , \sigMatrix[3][6] , 
        \sigMatrix[3][5] , \sigMatrix[3][4] , \sigMatrix[3][3] , 
        \sigMatrix[3][2] , \sigMatrix[3][1] , \sigMatrix[3][0] }) );
  booth_mul_row_N64_RADIX3_12 booth_mul_row_1_4 ( .prevA({\sigMatrix[3][127] , 
        \sigMatrix[3][126] , \sigMatrix[3][125] , \sigMatrix[3][124] , 
        \sigMatrix[3][123] , \sigMatrix[3][122] , \sigMatrix[3][121] , 
        \sigMatrix[3][120] , \sigMatrix[3][119] , \sigMatrix[3][118] , 
        \sigMatrix[3][117] , \sigMatrix[3][116] , \sigMatrix[3][115] , 
        \sigMatrix[3][114] , \sigMatrix[3][113] , \sigMatrix[3][112] , 
        \sigMatrix[3][111] , \sigMatrix[3][110] , \sigMatrix[3][109] , 
        \sigMatrix[3][108] , \sigMatrix[3][107] , \sigMatrix[3][106] , 
        \sigMatrix[3][105] , \sigMatrix[3][104] , \sigMatrix[3][103] , 
        \sigMatrix[3][102] , \sigMatrix[3][101] , \sigMatrix[3][100] , 
        \sigMatrix[3][99] , \sigMatrix[3][98] , \sigMatrix[3][97] , 
        \sigMatrix[3][96] , \sigMatrix[3][95] , \sigMatrix[3][94] , 
        \sigMatrix[3][93] , \sigMatrix[3][92] , \sigMatrix[3][91] , 
        \sigMatrix[3][90] , \sigMatrix[3][89] , \sigMatrix[3][88] , 
        \sigMatrix[3][87] , \sigMatrix[3][86] , \sigMatrix[3][85] , 
        \sigMatrix[3][84] , \sigMatrix[3][83] , \sigMatrix[3][82] , 
        \sigMatrix[3][81] , \sigMatrix[3][80] , \sigMatrix[3][79] , 
        \sigMatrix[3][78] , \sigMatrix[3][77] , \sigMatrix[3][76] , 
        \sigMatrix[3][75] , \sigMatrix[3][74] , \sigMatrix[3][73] , 
        \sigMatrix[3][72] , \sigMatrix[3][71] , \sigMatrix[3][70] , 
        \sigMatrix[3][69] , \sigMatrix[3][68] , \sigMatrix[3][67] , 
        \sigMatrix[3][66] , \sigMatrix[3][65] , 1'b0}), .prevSum({
        \sigMatrix[3][63] , \sigMatrix[3][62] , \sigMatrix[3][61] , 
        \sigMatrix[3][60] , \sigMatrix[3][59] , \sigMatrix[3][58] , 
        \sigMatrix[3][57] , \sigMatrix[3][56] , \sigMatrix[3][55] , 
        \sigMatrix[3][54] , \sigMatrix[3][53] , \sigMatrix[3][52] , 
        \sigMatrix[3][51] , \sigMatrix[3][50] , \sigMatrix[3][49] , 
        \sigMatrix[3][48] , \sigMatrix[3][47] , \sigMatrix[3][46] , 
        \sigMatrix[3][45] , \sigMatrix[3][44] , \sigMatrix[3][43] , 
        \sigMatrix[3][42] , \sigMatrix[3][41] , \sigMatrix[3][40] , 
        \sigMatrix[3][39] , \sigMatrix[3][38] , \sigMatrix[3][37] , 
        \sigMatrix[3][36] , \sigMatrix[3][35] , \sigMatrix[3][34] , 
        \sigMatrix[3][33] , \sigMatrix[3][32] , \sigMatrix[3][31] , 
        \sigMatrix[3][30] , \sigMatrix[3][29] , \sigMatrix[3][28] , 
        \sigMatrix[3][27] , \sigMatrix[3][26] , \sigMatrix[3][25] , 
        \sigMatrix[3][24] , \sigMatrix[3][23] , \sigMatrix[3][22] , 
        \sigMatrix[3][21] , \sigMatrix[3][20] , \sigMatrix[3][19] , 
        \sigMatrix[3][18] , \sigMatrix[3][17] , \sigMatrix[3][16] , 
        \sigMatrix[3][15] , \sigMatrix[3][14] , \sigMatrix[3][13] , 
        \sigMatrix[3][12] , \sigMatrix[3][11] , \sigMatrix[3][10] , 
        \sigMatrix[3][9] , \sigMatrix[3][8] , \sigMatrix[3][7] , 
        \sigMatrix[3][6] , \sigMatrix[3][5] , \sigMatrix[3][4] , 
        \sigMatrix[3][3] , \sigMatrix[3][2] , \sigMatrix[3][1] , 
        \sigMatrix[3][0] }), .encoderIn(B_out_s[9:7]), .nextA({
        \sigMatrix[4][127] , \sigMatrix[4][126] , \sigMatrix[4][125] , 
        \sigMatrix[4][124] , \sigMatrix[4][123] , \sigMatrix[4][122] , 
        \sigMatrix[4][121] , \sigMatrix[4][120] , \sigMatrix[4][119] , 
        \sigMatrix[4][118] , \sigMatrix[4][117] , \sigMatrix[4][116] , 
        \sigMatrix[4][115] , \sigMatrix[4][114] , \sigMatrix[4][113] , 
        \sigMatrix[4][112] , \sigMatrix[4][111] , \sigMatrix[4][110] , 
        \sigMatrix[4][109] , \sigMatrix[4][108] , \sigMatrix[4][107] , 
        \sigMatrix[4][106] , \sigMatrix[4][105] , \sigMatrix[4][104] , 
        \sigMatrix[4][103] , \sigMatrix[4][102] , \sigMatrix[4][101] , 
        \sigMatrix[4][100] , \sigMatrix[4][99] , \sigMatrix[4][98] , 
        \sigMatrix[4][97] , \sigMatrix[4][96] , \sigMatrix[4][95] , 
        \sigMatrix[4][94] , \sigMatrix[4][93] , \sigMatrix[4][92] , 
        \sigMatrix[4][91] , \sigMatrix[4][90] , \sigMatrix[4][89] , 
        \sigMatrix[4][88] , \sigMatrix[4][87] , \sigMatrix[4][86] , 
        \sigMatrix[4][85] , \sigMatrix[4][84] , \sigMatrix[4][83] , 
        \sigMatrix[4][82] , \sigMatrix[4][81] , \sigMatrix[4][80] , 
        \sigMatrix[4][79] , \sigMatrix[4][78] , \sigMatrix[4][77] , 
        \sigMatrix[4][76] , \sigMatrix[4][75] , \sigMatrix[4][74] , 
        \sigMatrix[4][73] , \sigMatrix[4][72] , \sigMatrix[4][71] , 
        \sigMatrix[4][70] , \sigMatrix[4][69] , \sigMatrix[4][68] , 
        \sigMatrix[4][67] , \sigMatrix[4][66] , \sigMatrix[4][65] , 
        SYNOPSYS_UNCONNECTED__4}), .nextSum({\sigMatrix[4][63] , 
        \sigMatrix[4][62] , \sigMatrix[4][61] , \sigMatrix[4][60] , 
        \sigMatrix[4][59] , \sigMatrix[4][58] , \sigMatrix[4][57] , 
        \sigMatrix[4][56] , \sigMatrix[4][55] , \sigMatrix[4][54] , 
        \sigMatrix[4][53] , \sigMatrix[4][52] , \sigMatrix[4][51] , 
        \sigMatrix[4][50] , \sigMatrix[4][49] , \sigMatrix[4][48] , 
        \sigMatrix[4][47] , \sigMatrix[4][46] , \sigMatrix[4][45] , 
        \sigMatrix[4][44] , \sigMatrix[4][43] , \sigMatrix[4][42] , 
        \sigMatrix[4][41] , \sigMatrix[4][40] , \sigMatrix[4][39] , 
        \sigMatrix[4][38] , \sigMatrix[4][37] , \sigMatrix[4][36] , 
        \sigMatrix[4][35] , \sigMatrix[4][34] , \sigMatrix[4][33] , 
        \sigMatrix[4][32] , \sigMatrix[4][31] , \sigMatrix[4][30] , 
        \sigMatrix[4][29] , \sigMatrix[4][28] , \sigMatrix[4][27] , 
        \sigMatrix[4][26] , \sigMatrix[4][25] , \sigMatrix[4][24] , 
        \sigMatrix[4][23] , \sigMatrix[4][22] , \sigMatrix[4][21] , 
        \sigMatrix[4][20] , \sigMatrix[4][19] , \sigMatrix[4][18] , 
        \sigMatrix[4][17] , \sigMatrix[4][16] , \sigMatrix[4][15] , 
        \sigMatrix[4][14] , \sigMatrix[4][13] , \sigMatrix[4][12] , 
        \sigMatrix[4][11] , \sigMatrix[4][10] , \sigMatrix[4][9] , 
        \sigMatrix[4][8] , \sigMatrix[4][7] , \sigMatrix[4][6] , 
        \sigMatrix[4][5] , \sigMatrix[4][4] , \sigMatrix[4][3] , 
        \sigMatrix[4][2] , \sigMatrix[4][1] , \sigMatrix[4][0] }) );
  booth_mul_row_N64_RADIX3_11 booth_mul_row_1_5 ( .prevA({\sigMatrix[4][127] , 
        \sigMatrix[4][126] , \sigMatrix[4][125] , \sigMatrix[4][124] , 
        \sigMatrix[4][123] , \sigMatrix[4][122] , \sigMatrix[4][121] , 
        \sigMatrix[4][120] , \sigMatrix[4][119] , \sigMatrix[4][118] , 
        \sigMatrix[4][117] , \sigMatrix[4][116] , \sigMatrix[4][115] , 
        \sigMatrix[4][114] , \sigMatrix[4][113] , \sigMatrix[4][112] , 
        \sigMatrix[4][111] , \sigMatrix[4][110] , \sigMatrix[4][109] , 
        \sigMatrix[4][108] , \sigMatrix[4][107] , \sigMatrix[4][106] , 
        \sigMatrix[4][105] , \sigMatrix[4][104] , \sigMatrix[4][103] , 
        \sigMatrix[4][102] , \sigMatrix[4][101] , \sigMatrix[4][100] , 
        \sigMatrix[4][99] , \sigMatrix[4][98] , \sigMatrix[4][97] , 
        \sigMatrix[4][96] , \sigMatrix[4][95] , \sigMatrix[4][94] , 
        \sigMatrix[4][93] , \sigMatrix[4][92] , \sigMatrix[4][91] , 
        \sigMatrix[4][90] , \sigMatrix[4][89] , \sigMatrix[4][88] , 
        \sigMatrix[4][87] , \sigMatrix[4][86] , \sigMatrix[4][85] , 
        \sigMatrix[4][84] , \sigMatrix[4][83] , \sigMatrix[4][82] , 
        \sigMatrix[4][81] , \sigMatrix[4][80] , \sigMatrix[4][79] , 
        \sigMatrix[4][78] , \sigMatrix[4][77] , \sigMatrix[4][76] , 
        \sigMatrix[4][75] , \sigMatrix[4][74] , \sigMatrix[4][73] , 
        \sigMatrix[4][72] , \sigMatrix[4][71] , \sigMatrix[4][70] , 
        \sigMatrix[4][69] , \sigMatrix[4][68] , \sigMatrix[4][67] , 
        \sigMatrix[4][66] , \sigMatrix[4][65] , 1'b0}), .prevSum({
        \sigMatrix[4][63] , \sigMatrix[4][62] , \sigMatrix[4][61] , 
        \sigMatrix[4][60] , \sigMatrix[4][59] , \sigMatrix[4][58] , 
        \sigMatrix[4][57] , \sigMatrix[4][56] , \sigMatrix[4][55] , 
        \sigMatrix[4][54] , \sigMatrix[4][53] , \sigMatrix[4][52] , 
        \sigMatrix[4][51] , \sigMatrix[4][50] , \sigMatrix[4][49] , 
        \sigMatrix[4][48] , \sigMatrix[4][47] , \sigMatrix[4][46] , 
        \sigMatrix[4][45] , \sigMatrix[4][44] , \sigMatrix[4][43] , 
        \sigMatrix[4][42] , \sigMatrix[4][41] , \sigMatrix[4][40] , 
        \sigMatrix[4][39] , \sigMatrix[4][38] , \sigMatrix[4][37] , 
        \sigMatrix[4][36] , \sigMatrix[4][35] , \sigMatrix[4][34] , 
        \sigMatrix[4][33] , \sigMatrix[4][32] , \sigMatrix[4][31] , 
        \sigMatrix[4][30] , \sigMatrix[4][29] , \sigMatrix[4][28] , 
        \sigMatrix[4][27] , \sigMatrix[4][26] , \sigMatrix[4][25] , 
        \sigMatrix[4][24] , \sigMatrix[4][23] , \sigMatrix[4][22] , 
        \sigMatrix[4][21] , \sigMatrix[4][20] , \sigMatrix[4][19] , 
        \sigMatrix[4][18] , \sigMatrix[4][17] , \sigMatrix[4][16] , 
        \sigMatrix[4][15] , \sigMatrix[4][14] , \sigMatrix[4][13] , 
        \sigMatrix[4][12] , \sigMatrix[4][11] , \sigMatrix[4][10] , 
        \sigMatrix[4][9] , \sigMatrix[4][8] , \sigMatrix[4][7] , 
        \sigMatrix[4][6] , \sigMatrix[4][5] , \sigMatrix[4][4] , 
        \sigMatrix[4][3] , \sigMatrix[4][2] , \sigMatrix[4][1] , 
        \sigMatrix[4][0] }), .encoderIn(B_out_s[11:9]), .nextA({
        \sigMatrix[5][127] , \sigMatrix[5][126] , \sigMatrix[5][125] , 
        \sigMatrix[5][124] , \sigMatrix[5][123] , \sigMatrix[5][122] , 
        \sigMatrix[5][121] , \sigMatrix[5][120] , \sigMatrix[5][119] , 
        \sigMatrix[5][118] , \sigMatrix[5][117] , \sigMatrix[5][116] , 
        \sigMatrix[5][115] , \sigMatrix[5][114] , \sigMatrix[5][113] , 
        \sigMatrix[5][112] , \sigMatrix[5][111] , \sigMatrix[5][110] , 
        \sigMatrix[5][109] , \sigMatrix[5][108] , \sigMatrix[5][107] , 
        \sigMatrix[5][106] , \sigMatrix[5][105] , \sigMatrix[5][104] , 
        \sigMatrix[5][103] , \sigMatrix[5][102] , \sigMatrix[5][101] , 
        \sigMatrix[5][100] , \sigMatrix[5][99] , \sigMatrix[5][98] , 
        \sigMatrix[5][97] , \sigMatrix[5][96] , \sigMatrix[5][95] , 
        \sigMatrix[5][94] , \sigMatrix[5][93] , \sigMatrix[5][92] , 
        \sigMatrix[5][91] , \sigMatrix[5][90] , \sigMatrix[5][89] , 
        \sigMatrix[5][88] , \sigMatrix[5][87] , \sigMatrix[5][86] , 
        \sigMatrix[5][85] , \sigMatrix[5][84] , \sigMatrix[5][83] , 
        \sigMatrix[5][82] , \sigMatrix[5][81] , \sigMatrix[5][80] , 
        \sigMatrix[5][79] , \sigMatrix[5][78] , \sigMatrix[5][77] , 
        \sigMatrix[5][76] , \sigMatrix[5][75] , \sigMatrix[5][74] , 
        \sigMatrix[5][73] , \sigMatrix[5][72] , \sigMatrix[5][71] , 
        \sigMatrix[5][70] , \sigMatrix[5][69] , \sigMatrix[5][68] , 
        \sigMatrix[5][67] , \sigMatrix[5][66] , \sigMatrix[5][65] , 
        SYNOPSYS_UNCONNECTED__5}), .nextSum({\sigMatrix[5][63] , 
        \sigMatrix[5][62] , \sigMatrix[5][61] , \sigMatrix[5][60] , 
        \sigMatrix[5][59] , \sigMatrix[5][58] , \sigMatrix[5][57] , 
        \sigMatrix[5][56] , \sigMatrix[5][55] , \sigMatrix[5][54] , 
        \sigMatrix[5][53] , \sigMatrix[5][52] , \sigMatrix[5][51] , 
        \sigMatrix[5][50] , \sigMatrix[5][49] , \sigMatrix[5][48] , 
        \sigMatrix[5][47] , \sigMatrix[5][46] , \sigMatrix[5][45] , 
        \sigMatrix[5][44] , \sigMatrix[5][43] , \sigMatrix[5][42] , 
        \sigMatrix[5][41] , \sigMatrix[5][40] , \sigMatrix[5][39] , 
        \sigMatrix[5][38] , \sigMatrix[5][37] , \sigMatrix[5][36] , 
        \sigMatrix[5][35] , \sigMatrix[5][34] , \sigMatrix[5][33] , 
        \sigMatrix[5][32] , \sigMatrix[5][31] , \sigMatrix[5][30] , 
        \sigMatrix[5][29] , \sigMatrix[5][28] , \sigMatrix[5][27] , 
        \sigMatrix[5][26] , \sigMatrix[5][25] , \sigMatrix[5][24] , 
        \sigMatrix[5][23] , \sigMatrix[5][22] , \sigMatrix[5][21] , 
        \sigMatrix[5][20] , \sigMatrix[5][19] , \sigMatrix[5][18] , 
        \sigMatrix[5][17] , \sigMatrix[5][16] , \sigMatrix[5][15] , 
        \sigMatrix[5][14] , \sigMatrix[5][13] , \sigMatrix[5][12] , 
        \sigMatrix[5][11] , \sigMatrix[5][10] , \sigMatrix[5][9] , 
        \sigMatrix[5][8] , \sigMatrix[5][7] , \sigMatrix[5][6] , 
        \sigMatrix[5][5] , \sigMatrix[5][4] , \sigMatrix[5][3] , 
        \sigMatrix[5][2] , \sigMatrix[5][1] , \sigMatrix[5][0] }) );
  booth_mul_row_N64_RADIX3_10 booth_mul_row_1_6 ( .prevA({\sigMatrix[5][127] , 
        \sigMatrix[5][126] , \sigMatrix[5][125] , \sigMatrix[5][124] , 
        \sigMatrix[5][123] , \sigMatrix[5][122] , \sigMatrix[5][121] , 
        \sigMatrix[5][120] , \sigMatrix[5][119] , \sigMatrix[5][118] , 
        \sigMatrix[5][117] , \sigMatrix[5][116] , \sigMatrix[5][115] , 
        \sigMatrix[5][114] , \sigMatrix[5][113] , \sigMatrix[5][112] , 
        \sigMatrix[5][111] , \sigMatrix[5][110] , \sigMatrix[5][109] , 
        \sigMatrix[5][108] , \sigMatrix[5][107] , \sigMatrix[5][106] , 
        \sigMatrix[5][105] , \sigMatrix[5][104] , \sigMatrix[5][103] , 
        \sigMatrix[5][102] , \sigMatrix[5][101] , \sigMatrix[5][100] , 
        \sigMatrix[5][99] , \sigMatrix[5][98] , \sigMatrix[5][97] , 
        \sigMatrix[5][96] , \sigMatrix[5][95] , \sigMatrix[5][94] , 
        \sigMatrix[5][93] , \sigMatrix[5][92] , \sigMatrix[5][91] , 
        \sigMatrix[5][90] , \sigMatrix[5][89] , \sigMatrix[5][88] , 
        \sigMatrix[5][87] , \sigMatrix[5][86] , \sigMatrix[5][85] , 
        \sigMatrix[5][84] , \sigMatrix[5][83] , \sigMatrix[5][82] , 
        \sigMatrix[5][81] , \sigMatrix[5][80] , \sigMatrix[5][79] , 
        \sigMatrix[5][78] , \sigMatrix[5][77] , \sigMatrix[5][76] , 
        \sigMatrix[5][75] , \sigMatrix[5][74] , \sigMatrix[5][73] , 
        \sigMatrix[5][72] , \sigMatrix[5][71] , \sigMatrix[5][70] , 
        \sigMatrix[5][69] , \sigMatrix[5][68] , \sigMatrix[5][67] , 
        \sigMatrix[5][66] , \sigMatrix[5][65] , 1'b0}), .prevSum({
        \sigMatrix[5][63] , \sigMatrix[5][62] , \sigMatrix[5][61] , 
        \sigMatrix[5][60] , \sigMatrix[5][59] , \sigMatrix[5][58] , 
        \sigMatrix[5][57] , \sigMatrix[5][56] , \sigMatrix[5][55] , 
        \sigMatrix[5][54] , \sigMatrix[5][53] , \sigMatrix[5][52] , 
        \sigMatrix[5][51] , \sigMatrix[5][50] , \sigMatrix[5][49] , 
        \sigMatrix[5][48] , \sigMatrix[5][47] , \sigMatrix[5][46] , 
        \sigMatrix[5][45] , \sigMatrix[5][44] , \sigMatrix[5][43] , 
        \sigMatrix[5][42] , \sigMatrix[5][41] , \sigMatrix[5][40] , 
        \sigMatrix[5][39] , \sigMatrix[5][38] , \sigMatrix[5][37] , 
        \sigMatrix[5][36] , \sigMatrix[5][35] , \sigMatrix[5][34] , 
        \sigMatrix[5][33] , \sigMatrix[5][32] , \sigMatrix[5][31] , 
        \sigMatrix[5][30] , \sigMatrix[5][29] , \sigMatrix[5][28] , 
        \sigMatrix[5][27] , \sigMatrix[5][26] , \sigMatrix[5][25] , 
        \sigMatrix[5][24] , \sigMatrix[5][23] , \sigMatrix[5][22] , 
        \sigMatrix[5][21] , \sigMatrix[5][20] , \sigMatrix[5][19] , 
        \sigMatrix[5][18] , \sigMatrix[5][17] , \sigMatrix[5][16] , 
        \sigMatrix[5][15] , \sigMatrix[5][14] , \sigMatrix[5][13] , 
        \sigMatrix[5][12] , \sigMatrix[5][11] , \sigMatrix[5][10] , 
        \sigMatrix[5][9] , \sigMatrix[5][8] , \sigMatrix[5][7] , 
        \sigMatrix[5][6] , \sigMatrix[5][5] , \sigMatrix[5][4] , 
        \sigMatrix[5][3] , \sigMatrix[5][2] , \sigMatrix[5][1] , 
        \sigMatrix[5][0] }), .encoderIn(B_out_s[13:11]), .nextA({
        \sigMatrix[6][127] , \sigMatrix[6][126] , \sigMatrix[6][125] , 
        \sigMatrix[6][124] , \sigMatrix[6][123] , \sigMatrix[6][122] , 
        \sigMatrix[6][121] , \sigMatrix[6][120] , \sigMatrix[6][119] , 
        \sigMatrix[6][118] , \sigMatrix[6][117] , \sigMatrix[6][116] , 
        \sigMatrix[6][115] , \sigMatrix[6][114] , \sigMatrix[6][113] , 
        \sigMatrix[6][112] , \sigMatrix[6][111] , \sigMatrix[6][110] , 
        \sigMatrix[6][109] , \sigMatrix[6][108] , \sigMatrix[6][107] , 
        \sigMatrix[6][106] , \sigMatrix[6][105] , \sigMatrix[6][104] , 
        \sigMatrix[6][103] , \sigMatrix[6][102] , \sigMatrix[6][101] , 
        \sigMatrix[6][100] , \sigMatrix[6][99] , \sigMatrix[6][98] , 
        \sigMatrix[6][97] , \sigMatrix[6][96] , \sigMatrix[6][95] , 
        \sigMatrix[6][94] , \sigMatrix[6][93] , \sigMatrix[6][92] , 
        \sigMatrix[6][91] , \sigMatrix[6][90] , \sigMatrix[6][89] , 
        \sigMatrix[6][88] , \sigMatrix[6][87] , \sigMatrix[6][86] , 
        \sigMatrix[6][85] , \sigMatrix[6][84] , \sigMatrix[6][83] , 
        \sigMatrix[6][82] , \sigMatrix[6][81] , \sigMatrix[6][80] , 
        \sigMatrix[6][79] , \sigMatrix[6][78] , \sigMatrix[6][77] , 
        \sigMatrix[6][76] , \sigMatrix[6][75] , \sigMatrix[6][74] , 
        \sigMatrix[6][73] , \sigMatrix[6][72] , \sigMatrix[6][71] , 
        \sigMatrix[6][70] , \sigMatrix[6][69] , \sigMatrix[6][68] , 
        \sigMatrix[6][67] , \sigMatrix[6][66] , \sigMatrix[6][65] , 
        SYNOPSYS_UNCONNECTED__6}), .nextSum({\sigMatrix[6][63] , 
        \sigMatrix[6][62] , \sigMatrix[6][61] , \sigMatrix[6][60] , 
        \sigMatrix[6][59] , \sigMatrix[6][58] , \sigMatrix[6][57] , 
        \sigMatrix[6][56] , \sigMatrix[6][55] , \sigMatrix[6][54] , 
        \sigMatrix[6][53] , \sigMatrix[6][52] , \sigMatrix[6][51] , 
        \sigMatrix[6][50] , \sigMatrix[6][49] , \sigMatrix[6][48] , 
        \sigMatrix[6][47] , \sigMatrix[6][46] , \sigMatrix[6][45] , 
        \sigMatrix[6][44] , \sigMatrix[6][43] , \sigMatrix[6][42] , 
        \sigMatrix[6][41] , \sigMatrix[6][40] , \sigMatrix[6][39] , 
        \sigMatrix[6][38] , \sigMatrix[6][37] , \sigMatrix[6][36] , 
        \sigMatrix[6][35] , \sigMatrix[6][34] , \sigMatrix[6][33] , 
        \sigMatrix[6][32] , \sigMatrix[6][31] , \sigMatrix[6][30] , 
        \sigMatrix[6][29] , \sigMatrix[6][28] , \sigMatrix[6][27] , 
        \sigMatrix[6][26] , \sigMatrix[6][25] , \sigMatrix[6][24] , 
        \sigMatrix[6][23] , \sigMatrix[6][22] , \sigMatrix[6][21] , 
        \sigMatrix[6][20] , \sigMatrix[6][19] , \sigMatrix[6][18] , 
        \sigMatrix[6][17] , \sigMatrix[6][16] , \sigMatrix[6][15] , 
        \sigMatrix[6][14] , \sigMatrix[6][13] , \sigMatrix[6][12] , 
        \sigMatrix[6][11] , \sigMatrix[6][10] , \sigMatrix[6][9] , 
        \sigMatrix[6][8] , \sigMatrix[6][7] , \sigMatrix[6][6] , 
        \sigMatrix[6][5] , \sigMatrix[6][4] , \sigMatrix[6][3] , 
        \sigMatrix[6][2] , \sigMatrix[6][1] , \sigMatrix[6][0] }) );
  booth_mul_row_N64_RADIX3_9 booth_mul_row_1_7 ( .prevA({\sigMatrix[6][127] , 
        \sigMatrix[6][126] , \sigMatrix[6][125] , \sigMatrix[6][124] , 
        \sigMatrix[6][123] , \sigMatrix[6][122] , \sigMatrix[6][121] , 
        \sigMatrix[6][120] , \sigMatrix[6][119] , \sigMatrix[6][118] , 
        \sigMatrix[6][117] , \sigMatrix[6][116] , \sigMatrix[6][115] , 
        \sigMatrix[6][114] , \sigMatrix[6][113] , \sigMatrix[6][112] , 
        \sigMatrix[6][111] , \sigMatrix[6][110] , \sigMatrix[6][109] , 
        \sigMatrix[6][108] , \sigMatrix[6][107] , \sigMatrix[6][106] , 
        \sigMatrix[6][105] , \sigMatrix[6][104] , \sigMatrix[6][103] , 
        \sigMatrix[6][102] , \sigMatrix[6][101] , \sigMatrix[6][100] , 
        \sigMatrix[6][99] , \sigMatrix[6][98] , \sigMatrix[6][97] , 
        \sigMatrix[6][96] , \sigMatrix[6][95] , \sigMatrix[6][94] , 
        \sigMatrix[6][93] , \sigMatrix[6][92] , \sigMatrix[6][91] , 
        \sigMatrix[6][90] , \sigMatrix[6][89] , \sigMatrix[6][88] , 
        \sigMatrix[6][87] , \sigMatrix[6][86] , \sigMatrix[6][85] , 
        \sigMatrix[6][84] , \sigMatrix[6][83] , \sigMatrix[6][82] , 
        \sigMatrix[6][81] , \sigMatrix[6][80] , \sigMatrix[6][79] , 
        \sigMatrix[6][78] , \sigMatrix[6][77] , \sigMatrix[6][76] , 
        \sigMatrix[6][75] , \sigMatrix[6][74] , \sigMatrix[6][73] , 
        \sigMatrix[6][72] , \sigMatrix[6][71] , \sigMatrix[6][70] , 
        \sigMatrix[6][69] , \sigMatrix[6][68] , \sigMatrix[6][67] , 
        \sigMatrix[6][66] , \sigMatrix[6][65] , 1'b0}), .prevSum({
        \sigMatrix[6][63] , \sigMatrix[6][62] , \sigMatrix[6][61] , 
        \sigMatrix[6][60] , \sigMatrix[6][59] , \sigMatrix[6][58] , 
        \sigMatrix[6][57] , \sigMatrix[6][56] , \sigMatrix[6][55] , 
        \sigMatrix[6][54] , \sigMatrix[6][53] , \sigMatrix[6][52] , 
        \sigMatrix[6][51] , \sigMatrix[6][50] , \sigMatrix[6][49] , 
        \sigMatrix[6][48] , \sigMatrix[6][47] , \sigMatrix[6][46] , 
        \sigMatrix[6][45] , \sigMatrix[6][44] , \sigMatrix[6][43] , 
        \sigMatrix[6][42] , \sigMatrix[6][41] , \sigMatrix[6][40] , 
        \sigMatrix[6][39] , \sigMatrix[6][38] , \sigMatrix[6][37] , 
        \sigMatrix[6][36] , \sigMatrix[6][35] , \sigMatrix[6][34] , 
        \sigMatrix[6][33] , \sigMatrix[6][32] , \sigMatrix[6][31] , 
        \sigMatrix[6][30] , \sigMatrix[6][29] , \sigMatrix[6][28] , 
        \sigMatrix[6][27] , \sigMatrix[6][26] , \sigMatrix[6][25] , 
        \sigMatrix[6][24] , \sigMatrix[6][23] , \sigMatrix[6][22] , 
        \sigMatrix[6][21] , \sigMatrix[6][20] , \sigMatrix[6][19] , 
        \sigMatrix[6][18] , \sigMatrix[6][17] , \sigMatrix[6][16] , 
        \sigMatrix[6][15] , \sigMatrix[6][14] , \sigMatrix[6][13] , 
        \sigMatrix[6][12] , \sigMatrix[6][11] , \sigMatrix[6][10] , 
        \sigMatrix[6][9] , \sigMatrix[6][8] , \sigMatrix[6][7] , 
        \sigMatrix[6][6] , \sigMatrix[6][5] , \sigMatrix[6][4] , 
        \sigMatrix[6][3] , \sigMatrix[6][2] , \sigMatrix[6][1] , 
        \sigMatrix[6][0] }), .encoderIn(B_out_s[15:13]), .nextA({
        \sigMatrix[7][127] , \sigMatrix[7][126] , \sigMatrix[7][125] , 
        \sigMatrix[7][124] , \sigMatrix[7][123] , \sigMatrix[7][122] , 
        \sigMatrix[7][121] , \sigMatrix[7][120] , \sigMatrix[7][119] , 
        \sigMatrix[7][118] , \sigMatrix[7][117] , \sigMatrix[7][116] , 
        \sigMatrix[7][115] , \sigMatrix[7][114] , \sigMatrix[7][113] , 
        \sigMatrix[7][112] , \sigMatrix[7][111] , \sigMatrix[7][110] , 
        \sigMatrix[7][109] , \sigMatrix[7][108] , \sigMatrix[7][107] , 
        \sigMatrix[7][106] , \sigMatrix[7][105] , \sigMatrix[7][104] , 
        \sigMatrix[7][103] , \sigMatrix[7][102] , \sigMatrix[7][101] , 
        \sigMatrix[7][100] , \sigMatrix[7][99] , \sigMatrix[7][98] , 
        \sigMatrix[7][97] , \sigMatrix[7][96] , \sigMatrix[7][95] , 
        \sigMatrix[7][94] , \sigMatrix[7][93] , \sigMatrix[7][92] , 
        \sigMatrix[7][91] , \sigMatrix[7][90] , \sigMatrix[7][89] , 
        \sigMatrix[7][88] , \sigMatrix[7][87] , \sigMatrix[7][86] , 
        \sigMatrix[7][85] , \sigMatrix[7][84] , \sigMatrix[7][83] , 
        \sigMatrix[7][82] , \sigMatrix[7][81] , \sigMatrix[7][80] , 
        \sigMatrix[7][79] , \sigMatrix[7][78] , \sigMatrix[7][77] , 
        \sigMatrix[7][76] , \sigMatrix[7][75] , \sigMatrix[7][74] , 
        \sigMatrix[7][73] , \sigMatrix[7][72] , \sigMatrix[7][71] , 
        \sigMatrix[7][70] , \sigMatrix[7][69] , \sigMatrix[7][68] , 
        \sigMatrix[7][67] , \sigMatrix[7][66] , \sigMatrix[7][65] , 
        SYNOPSYS_UNCONNECTED__7}), .nextSum({\sigMatrix[7][63] , 
        \sigMatrix[7][62] , \sigMatrix[7][61] , \sigMatrix[7][60] , 
        \sigMatrix[7][59] , \sigMatrix[7][58] , \sigMatrix[7][57] , 
        \sigMatrix[7][56] , \sigMatrix[7][55] , \sigMatrix[7][54] , 
        \sigMatrix[7][53] , \sigMatrix[7][52] , \sigMatrix[7][51] , 
        \sigMatrix[7][50] , \sigMatrix[7][49] , \sigMatrix[7][48] , 
        \sigMatrix[7][47] , \sigMatrix[7][46] , \sigMatrix[7][45] , 
        \sigMatrix[7][44] , \sigMatrix[7][43] , \sigMatrix[7][42] , 
        \sigMatrix[7][41] , \sigMatrix[7][40] , \sigMatrix[7][39] , 
        \sigMatrix[7][38] , \sigMatrix[7][37] , \sigMatrix[7][36] , 
        \sigMatrix[7][35] , \sigMatrix[7][34] , \sigMatrix[7][33] , 
        \sigMatrix[7][32] , \sigMatrix[7][31] , \sigMatrix[7][30] , 
        \sigMatrix[7][29] , \sigMatrix[7][28] , \sigMatrix[7][27] , 
        \sigMatrix[7][26] , \sigMatrix[7][25] , \sigMatrix[7][24] , 
        \sigMatrix[7][23] , \sigMatrix[7][22] , \sigMatrix[7][21] , 
        \sigMatrix[7][20] , \sigMatrix[7][19] , \sigMatrix[7][18] , 
        \sigMatrix[7][17] , \sigMatrix[7][16] , \sigMatrix[7][15] , 
        \sigMatrix[7][14] , \sigMatrix[7][13] , \sigMatrix[7][12] , 
        \sigMatrix[7][11] , \sigMatrix[7][10] , \sigMatrix[7][9] , 
        \sigMatrix[7][8] , \sigMatrix[7][7] , \sigMatrix[7][6] , 
        \sigMatrix[7][5] , \sigMatrix[7][4] , \sigMatrix[7][3] , 
        \sigMatrix[7][2] , \sigMatrix[7][1] , \sigMatrix[7][0] }) );
  booth_mul_row_N64_RADIX3_8 booth_mul_row_1_8 ( .prevA({\sigMatrix[7][127] , 
        \sigMatrix[7][126] , \sigMatrix[7][125] , \sigMatrix[7][124] , 
        \sigMatrix[7][123] , \sigMatrix[7][122] , \sigMatrix[7][121] , 
        \sigMatrix[7][120] , \sigMatrix[7][119] , \sigMatrix[7][118] , 
        \sigMatrix[7][117] , \sigMatrix[7][116] , \sigMatrix[7][115] , 
        \sigMatrix[7][114] , \sigMatrix[7][113] , \sigMatrix[7][112] , 
        \sigMatrix[7][111] , \sigMatrix[7][110] , \sigMatrix[7][109] , 
        \sigMatrix[7][108] , \sigMatrix[7][107] , \sigMatrix[7][106] , 
        \sigMatrix[7][105] , \sigMatrix[7][104] , \sigMatrix[7][103] , 
        \sigMatrix[7][102] , \sigMatrix[7][101] , \sigMatrix[7][100] , 
        \sigMatrix[7][99] , \sigMatrix[7][98] , \sigMatrix[7][97] , 
        \sigMatrix[7][96] , \sigMatrix[7][95] , \sigMatrix[7][94] , 
        \sigMatrix[7][93] , \sigMatrix[7][92] , \sigMatrix[7][91] , 
        \sigMatrix[7][90] , \sigMatrix[7][89] , \sigMatrix[7][88] , 
        \sigMatrix[7][87] , \sigMatrix[7][86] , \sigMatrix[7][85] , 
        \sigMatrix[7][84] , \sigMatrix[7][83] , \sigMatrix[7][82] , 
        \sigMatrix[7][81] , \sigMatrix[7][80] , \sigMatrix[7][79] , 
        \sigMatrix[7][78] , \sigMatrix[7][77] , \sigMatrix[7][76] , 
        \sigMatrix[7][75] , \sigMatrix[7][74] , \sigMatrix[7][73] , 
        \sigMatrix[7][72] , \sigMatrix[7][71] , \sigMatrix[7][70] , 
        \sigMatrix[7][69] , \sigMatrix[7][68] , \sigMatrix[7][67] , 
        \sigMatrix[7][66] , \sigMatrix[7][65] , 1'b0}), .prevSum({
        \sigMatrix[7][63] , \sigMatrix[7][62] , \sigMatrix[7][61] , 
        \sigMatrix[7][60] , \sigMatrix[7][59] , \sigMatrix[7][58] , 
        \sigMatrix[7][57] , \sigMatrix[7][56] , \sigMatrix[7][55] , 
        \sigMatrix[7][54] , \sigMatrix[7][53] , \sigMatrix[7][52] , 
        \sigMatrix[7][51] , \sigMatrix[7][50] , \sigMatrix[7][49] , 
        \sigMatrix[7][48] , \sigMatrix[7][47] , \sigMatrix[7][46] , 
        \sigMatrix[7][45] , \sigMatrix[7][44] , \sigMatrix[7][43] , 
        \sigMatrix[7][42] , \sigMatrix[7][41] , \sigMatrix[7][40] , 
        \sigMatrix[7][39] , \sigMatrix[7][38] , \sigMatrix[7][37] , 
        \sigMatrix[7][36] , \sigMatrix[7][35] , \sigMatrix[7][34] , 
        \sigMatrix[7][33] , \sigMatrix[7][32] , \sigMatrix[7][31] , 
        \sigMatrix[7][30] , \sigMatrix[7][29] , \sigMatrix[7][28] , 
        \sigMatrix[7][27] , \sigMatrix[7][26] , \sigMatrix[7][25] , 
        \sigMatrix[7][24] , \sigMatrix[7][23] , \sigMatrix[7][22] , 
        \sigMatrix[7][21] , \sigMatrix[7][20] , \sigMatrix[7][19] , 
        \sigMatrix[7][18] , \sigMatrix[7][17] , \sigMatrix[7][16] , 
        \sigMatrix[7][15] , \sigMatrix[7][14] , \sigMatrix[7][13] , 
        \sigMatrix[7][12] , \sigMatrix[7][11] , \sigMatrix[7][10] , 
        \sigMatrix[7][9] , \sigMatrix[7][8] , \sigMatrix[7][7] , 
        \sigMatrix[7][6] , \sigMatrix[7][5] , \sigMatrix[7][4] , 
        \sigMatrix[7][3] , \sigMatrix[7][2] , \sigMatrix[7][1] , 
        \sigMatrix[7][0] }), .encoderIn(B_out_s[17:15]), .nextA({
        \sigMatrix[8][127] , \sigMatrix[8][126] , \sigMatrix[8][125] , 
        \sigMatrix[8][124] , \sigMatrix[8][123] , \sigMatrix[8][122] , 
        \sigMatrix[8][121] , \sigMatrix[8][120] , \sigMatrix[8][119] , 
        \sigMatrix[8][118] , \sigMatrix[8][117] , \sigMatrix[8][116] , 
        \sigMatrix[8][115] , \sigMatrix[8][114] , \sigMatrix[8][113] , 
        \sigMatrix[8][112] , \sigMatrix[8][111] , \sigMatrix[8][110] , 
        \sigMatrix[8][109] , \sigMatrix[8][108] , \sigMatrix[8][107] , 
        \sigMatrix[8][106] , \sigMatrix[8][105] , \sigMatrix[8][104] , 
        \sigMatrix[8][103] , \sigMatrix[8][102] , \sigMatrix[8][101] , 
        \sigMatrix[8][100] , \sigMatrix[8][99] , \sigMatrix[8][98] , 
        \sigMatrix[8][97] , \sigMatrix[8][96] , \sigMatrix[8][95] , 
        \sigMatrix[8][94] , \sigMatrix[8][93] , \sigMatrix[8][92] , 
        \sigMatrix[8][91] , \sigMatrix[8][90] , \sigMatrix[8][89] , 
        \sigMatrix[8][88] , \sigMatrix[8][87] , \sigMatrix[8][86] , 
        \sigMatrix[8][85] , \sigMatrix[8][84] , \sigMatrix[8][83] , 
        \sigMatrix[8][82] , \sigMatrix[8][81] , \sigMatrix[8][80] , 
        \sigMatrix[8][79] , \sigMatrix[8][78] , \sigMatrix[8][77] , 
        \sigMatrix[8][76] , \sigMatrix[8][75] , \sigMatrix[8][74] , 
        \sigMatrix[8][73] , \sigMatrix[8][72] , \sigMatrix[8][71] , 
        \sigMatrix[8][70] , \sigMatrix[8][69] , \sigMatrix[8][68] , 
        \sigMatrix[8][67] , \sigMatrix[8][66] , \sigMatrix[8][65] , 
        SYNOPSYS_UNCONNECTED__8}), .nextSum({\sigMatrix[8][63] , 
        \sigMatrix[8][62] , \sigMatrix[8][61] , \sigMatrix[8][60] , 
        \sigMatrix[8][59] , \sigMatrix[8][58] , \sigMatrix[8][57] , 
        \sigMatrix[8][56] , \sigMatrix[8][55] , \sigMatrix[8][54] , 
        \sigMatrix[8][53] , \sigMatrix[8][52] , \sigMatrix[8][51] , 
        \sigMatrix[8][50] , \sigMatrix[8][49] , \sigMatrix[8][48] , 
        \sigMatrix[8][47] , \sigMatrix[8][46] , \sigMatrix[8][45] , 
        \sigMatrix[8][44] , \sigMatrix[8][43] , \sigMatrix[8][42] , 
        \sigMatrix[8][41] , \sigMatrix[8][40] , \sigMatrix[8][39] , 
        \sigMatrix[8][38] , \sigMatrix[8][37] , \sigMatrix[8][36] , 
        \sigMatrix[8][35] , \sigMatrix[8][34] , \sigMatrix[8][33] , 
        \sigMatrix[8][32] , \sigMatrix[8][31] , \sigMatrix[8][30] , 
        \sigMatrix[8][29] , \sigMatrix[8][28] , \sigMatrix[8][27] , 
        \sigMatrix[8][26] , \sigMatrix[8][25] , \sigMatrix[8][24] , 
        \sigMatrix[8][23] , \sigMatrix[8][22] , \sigMatrix[8][21] , 
        \sigMatrix[8][20] , \sigMatrix[8][19] , \sigMatrix[8][18] , 
        \sigMatrix[8][17] , \sigMatrix[8][16] , \sigMatrix[8][15] , 
        \sigMatrix[8][14] , \sigMatrix[8][13] , \sigMatrix[8][12] , 
        \sigMatrix[8][11] , \sigMatrix[8][10] , \sigMatrix[8][9] , 
        \sigMatrix[8][8] , \sigMatrix[8][7] , \sigMatrix[8][6] , 
        \sigMatrix[8][5] , \sigMatrix[8][4] , \sigMatrix[8][3] , 
        \sigMatrix[8][2] , \sigMatrix[8][1] , \sigMatrix[8][0] }) );
  booth_mul_row_N64_RADIX3_7 booth_mul_row_1_9 ( .prevA({\sigMatrix[8][127] , 
        \sigMatrix[8][126] , \sigMatrix[8][125] , \sigMatrix[8][124] , 
        \sigMatrix[8][123] , \sigMatrix[8][122] , \sigMatrix[8][121] , 
        \sigMatrix[8][120] , \sigMatrix[8][119] , \sigMatrix[8][118] , 
        \sigMatrix[8][117] , \sigMatrix[8][116] , \sigMatrix[8][115] , 
        \sigMatrix[8][114] , \sigMatrix[8][113] , \sigMatrix[8][112] , 
        \sigMatrix[8][111] , \sigMatrix[8][110] , \sigMatrix[8][109] , 
        \sigMatrix[8][108] , \sigMatrix[8][107] , \sigMatrix[8][106] , 
        \sigMatrix[8][105] , \sigMatrix[8][104] , \sigMatrix[8][103] , 
        \sigMatrix[8][102] , \sigMatrix[8][101] , \sigMatrix[8][100] , 
        \sigMatrix[8][99] , \sigMatrix[8][98] , \sigMatrix[8][97] , 
        \sigMatrix[8][96] , \sigMatrix[8][95] , \sigMatrix[8][94] , 
        \sigMatrix[8][93] , \sigMatrix[8][92] , \sigMatrix[8][91] , 
        \sigMatrix[8][90] , \sigMatrix[8][89] , \sigMatrix[8][88] , 
        \sigMatrix[8][87] , \sigMatrix[8][86] , \sigMatrix[8][85] , 
        \sigMatrix[8][84] , \sigMatrix[8][83] , \sigMatrix[8][82] , 
        \sigMatrix[8][81] , \sigMatrix[8][80] , \sigMatrix[8][79] , 
        \sigMatrix[8][78] , \sigMatrix[8][77] , \sigMatrix[8][76] , 
        \sigMatrix[8][75] , \sigMatrix[8][74] , \sigMatrix[8][73] , 
        \sigMatrix[8][72] , \sigMatrix[8][71] , \sigMatrix[8][70] , 
        \sigMatrix[8][69] , \sigMatrix[8][68] , \sigMatrix[8][67] , 
        \sigMatrix[8][66] , \sigMatrix[8][65] , 1'b0}), .prevSum({
        \sigMatrix[8][63] , \sigMatrix[8][62] , \sigMatrix[8][61] , 
        \sigMatrix[8][60] , \sigMatrix[8][59] , \sigMatrix[8][58] , 
        \sigMatrix[8][57] , \sigMatrix[8][56] , \sigMatrix[8][55] , 
        \sigMatrix[8][54] , \sigMatrix[8][53] , \sigMatrix[8][52] , 
        \sigMatrix[8][51] , \sigMatrix[8][50] , \sigMatrix[8][49] , 
        \sigMatrix[8][48] , \sigMatrix[8][47] , \sigMatrix[8][46] , 
        \sigMatrix[8][45] , \sigMatrix[8][44] , \sigMatrix[8][43] , 
        \sigMatrix[8][42] , \sigMatrix[8][41] , \sigMatrix[8][40] , 
        \sigMatrix[8][39] , \sigMatrix[8][38] , \sigMatrix[8][37] , 
        \sigMatrix[8][36] , \sigMatrix[8][35] , \sigMatrix[8][34] , 
        \sigMatrix[8][33] , \sigMatrix[8][32] , \sigMatrix[8][31] , 
        \sigMatrix[8][30] , \sigMatrix[8][29] , \sigMatrix[8][28] , 
        \sigMatrix[8][27] , \sigMatrix[8][26] , \sigMatrix[8][25] , 
        \sigMatrix[8][24] , \sigMatrix[8][23] , \sigMatrix[8][22] , 
        \sigMatrix[8][21] , \sigMatrix[8][20] , \sigMatrix[8][19] , 
        \sigMatrix[8][18] , \sigMatrix[8][17] , \sigMatrix[8][16] , 
        \sigMatrix[8][15] , \sigMatrix[8][14] , \sigMatrix[8][13] , 
        \sigMatrix[8][12] , \sigMatrix[8][11] , \sigMatrix[8][10] , 
        \sigMatrix[8][9] , \sigMatrix[8][8] , \sigMatrix[8][7] , 
        \sigMatrix[8][6] , \sigMatrix[8][5] , \sigMatrix[8][4] , 
        \sigMatrix[8][3] , \sigMatrix[8][2] , \sigMatrix[8][1] , 
        \sigMatrix[8][0] }), .encoderIn(B_out_s[19:17]), .nextA({
        \sigMatrix[9][127] , \sigMatrix[9][126] , \sigMatrix[9][125] , 
        \sigMatrix[9][124] , \sigMatrix[9][123] , \sigMatrix[9][122] , 
        \sigMatrix[9][121] , \sigMatrix[9][120] , \sigMatrix[9][119] , 
        \sigMatrix[9][118] , \sigMatrix[9][117] , \sigMatrix[9][116] , 
        \sigMatrix[9][115] , \sigMatrix[9][114] , \sigMatrix[9][113] , 
        \sigMatrix[9][112] , \sigMatrix[9][111] , \sigMatrix[9][110] , 
        \sigMatrix[9][109] , \sigMatrix[9][108] , \sigMatrix[9][107] , 
        \sigMatrix[9][106] , \sigMatrix[9][105] , \sigMatrix[9][104] , 
        \sigMatrix[9][103] , \sigMatrix[9][102] , \sigMatrix[9][101] , 
        \sigMatrix[9][100] , \sigMatrix[9][99] , \sigMatrix[9][98] , 
        \sigMatrix[9][97] , \sigMatrix[9][96] , \sigMatrix[9][95] , 
        \sigMatrix[9][94] , \sigMatrix[9][93] , \sigMatrix[9][92] , 
        \sigMatrix[9][91] , \sigMatrix[9][90] , \sigMatrix[9][89] , 
        \sigMatrix[9][88] , \sigMatrix[9][87] , \sigMatrix[9][86] , 
        \sigMatrix[9][85] , \sigMatrix[9][84] , \sigMatrix[9][83] , 
        \sigMatrix[9][82] , \sigMatrix[9][81] , \sigMatrix[9][80] , 
        \sigMatrix[9][79] , \sigMatrix[9][78] , \sigMatrix[9][77] , 
        \sigMatrix[9][76] , \sigMatrix[9][75] , \sigMatrix[9][74] , 
        \sigMatrix[9][73] , \sigMatrix[9][72] , \sigMatrix[9][71] , 
        \sigMatrix[9][70] , \sigMatrix[9][69] , \sigMatrix[9][68] , 
        \sigMatrix[9][67] , \sigMatrix[9][66] , \sigMatrix[9][65] , 
        SYNOPSYS_UNCONNECTED__9}), .nextSum({\sigMatrix[9][63] , 
        \sigMatrix[9][62] , \sigMatrix[9][61] , \sigMatrix[9][60] , 
        \sigMatrix[9][59] , \sigMatrix[9][58] , \sigMatrix[9][57] , 
        \sigMatrix[9][56] , \sigMatrix[9][55] , \sigMatrix[9][54] , 
        \sigMatrix[9][53] , \sigMatrix[9][52] , \sigMatrix[9][51] , 
        \sigMatrix[9][50] , \sigMatrix[9][49] , \sigMatrix[9][48] , 
        \sigMatrix[9][47] , \sigMatrix[9][46] , \sigMatrix[9][45] , 
        \sigMatrix[9][44] , \sigMatrix[9][43] , \sigMatrix[9][42] , 
        \sigMatrix[9][41] , \sigMatrix[9][40] , \sigMatrix[9][39] , 
        \sigMatrix[9][38] , \sigMatrix[9][37] , \sigMatrix[9][36] , 
        \sigMatrix[9][35] , \sigMatrix[9][34] , \sigMatrix[9][33] , 
        \sigMatrix[9][32] , \sigMatrix[9][31] , \sigMatrix[9][30] , 
        \sigMatrix[9][29] , \sigMatrix[9][28] , \sigMatrix[9][27] , 
        \sigMatrix[9][26] , \sigMatrix[9][25] , \sigMatrix[9][24] , 
        \sigMatrix[9][23] , \sigMatrix[9][22] , \sigMatrix[9][21] , 
        \sigMatrix[9][20] , \sigMatrix[9][19] , \sigMatrix[9][18] , 
        \sigMatrix[9][17] , \sigMatrix[9][16] , \sigMatrix[9][15] , 
        \sigMatrix[9][14] , \sigMatrix[9][13] , \sigMatrix[9][12] , 
        \sigMatrix[9][11] , \sigMatrix[9][10] , \sigMatrix[9][9] , 
        \sigMatrix[9][8] , \sigMatrix[9][7] , \sigMatrix[9][6] , 
        \sigMatrix[9][5] , \sigMatrix[9][4] , \sigMatrix[9][3] , 
        \sigMatrix[9][2] , \sigMatrix[9][1] , \sigMatrix[9][0] }) );
  booth_mul_row_N64_RADIX3_6 booth_mul_row_1_10 ( .prevA({\sigMatrix[9][127] , 
        \sigMatrix[9][126] , \sigMatrix[9][125] , \sigMatrix[9][124] , 
        \sigMatrix[9][123] , \sigMatrix[9][122] , \sigMatrix[9][121] , 
        \sigMatrix[9][120] , \sigMatrix[9][119] , \sigMatrix[9][118] , 
        \sigMatrix[9][117] , \sigMatrix[9][116] , \sigMatrix[9][115] , 
        \sigMatrix[9][114] , \sigMatrix[9][113] , \sigMatrix[9][112] , 
        \sigMatrix[9][111] , \sigMatrix[9][110] , \sigMatrix[9][109] , 
        \sigMatrix[9][108] , \sigMatrix[9][107] , \sigMatrix[9][106] , 
        \sigMatrix[9][105] , \sigMatrix[9][104] , \sigMatrix[9][103] , 
        \sigMatrix[9][102] , \sigMatrix[9][101] , \sigMatrix[9][100] , 
        \sigMatrix[9][99] , \sigMatrix[9][98] , \sigMatrix[9][97] , 
        \sigMatrix[9][96] , \sigMatrix[9][95] , \sigMatrix[9][94] , 
        \sigMatrix[9][93] , \sigMatrix[9][92] , \sigMatrix[9][91] , 
        \sigMatrix[9][90] , \sigMatrix[9][89] , \sigMatrix[9][88] , 
        \sigMatrix[9][87] , \sigMatrix[9][86] , \sigMatrix[9][85] , 
        \sigMatrix[9][84] , \sigMatrix[9][83] , \sigMatrix[9][82] , 
        \sigMatrix[9][81] , \sigMatrix[9][80] , \sigMatrix[9][79] , 
        \sigMatrix[9][78] , \sigMatrix[9][77] , \sigMatrix[9][76] , 
        \sigMatrix[9][75] , \sigMatrix[9][74] , \sigMatrix[9][73] , 
        \sigMatrix[9][72] , \sigMatrix[9][71] , \sigMatrix[9][70] , 
        \sigMatrix[9][69] , \sigMatrix[9][68] , \sigMatrix[9][67] , 
        \sigMatrix[9][66] , \sigMatrix[9][65] , 1'b0}), .prevSum({
        \sigMatrix[9][63] , \sigMatrix[9][62] , \sigMatrix[9][61] , 
        \sigMatrix[9][60] , \sigMatrix[9][59] , \sigMatrix[9][58] , 
        \sigMatrix[9][57] , \sigMatrix[9][56] , \sigMatrix[9][55] , 
        \sigMatrix[9][54] , \sigMatrix[9][53] , \sigMatrix[9][52] , 
        \sigMatrix[9][51] , \sigMatrix[9][50] , \sigMatrix[9][49] , 
        \sigMatrix[9][48] , \sigMatrix[9][47] , \sigMatrix[9][46] , 
        \sigMatrix[9][45] , \sigMatrix[9][44] , \sigMatrix[9][43] , 
        \sigMatrix[9][42] , \sigMatrix[9][41] , \sigMatrix[9][40] , 
        \sigMatrix[9][39] , \sigMatrix[9][38] , \sigMatrix[9][37] , 
        \sigMatrix[9][36] , \sigMatrix[9][35] , \sigMatrix[9][34] , 
        \sigMatrix[9][33] , \sigMatrix[9][32] , \sigMatrix[9][31] , 
        \sigMatrix[9][30] , \sigMatrix[9][29] , \sigMatrix[9][28] , 
        \sigMatrix[9][27] , \sigMatrix[9][26] , \sigMatrix[9][25] , 
        \sigMatrix[9][24] , \sigMatrix[9][23] , \sigMatrix[9][22] , 
        \sigMatrix[9][21] , \sigMatrix[9][20] , \sigMatrix[9][19] , 
        \sigMatrix[9][18] , \sigMatrix[9][17] , \sigMatrix[9][16] , 
        \sigMatrix[9][15] , \sigMatrix[9][14] , \sigMatrix[9][13] , 
        \sigMatrix[9][12] , \sigMatrix[9][11] , \sigMatrix[9][10] , 
        \sigMatrix[9][9] , \sigMatrix[9][8] , \sigMatrix[9][7] , 
        \sigMatrix[9][6] , \sigMatrix[9][5] , \sigMatrix[9][4] , 
        \sigMatrix[9][3] , \sigMatrix[9][2] , \sigMatrix[9][1] , 
        \sigMatrix[9][0] }), .encoderIn(B_out_s[21:19]), .nextA({
        \sigMatrix[10][127] , \sigMatrix[10][126] , \sigMatrix[10][125] , 
        \sigMatrix[10][124] , \sigMatrix[10][123] , \sigMatrix[10][122] , 
        \sigMatrix[10][121] , \sigMatrix[10][120] , \sigMatrix[10][119] , 
        \sigMatrix[10][118] , \sigMatrix[10][117] , \sigMatrix[10][116] , 
        \sigMatrix[10][115] , \sigMatrix[10][114] , \sigMatrix[10][113] , 
        \sigMatrix[10][112] , \sigMatrix[10][111] , \sigMatrix[10][110] , 
        \sigMatrix[10][109] , \sigMatrix[10][108] , \sigMatrix[10][107] , 
        \sigMatrix[10][106] , \sigMatrix[10][105] , \sigMatrix[10][104] , 
        \sigMatrix[10][103] , \sigMatrix[10][102] , \sigMatrix[10][101] , 
        \sigMatrix[10][100] , \sigMatrix[10][99] , \sigMatrix[10][98] , 
        \sigMatrix[10][97] , \sigMatrix[10][96] , \sigMatrix[10][95] , 
        \sigMatrix[10][94] , \sigMatrix[10][93] , \sigMatrix[10][92] , 
        \sigMatrix[10][91] , \sigMatrix[10][90] , \sigMatrix[10][89] , 
        \sigMatrix[10][88] , \sigMatrix[10][87] , \sigMatrix[10][86] , 
        \sigMatrix[10][85] , \sigMatrix[10][84] , \sigMatrix[10][83] , 
        \sigMatrix[10][82] , \sigMatrix[10][81] , \sigMatrix[10][80] , 
        \sigMatrix[10][79] , \sigMatrix[10][78] , \sigMatrix[10][77] , 
        \sigMatrix[10][76] , \sigMatrix[10][75] , \sigMatrix[10][74] , 
        \sigMatrix[10][73] , \sigMatrix[10][72] , \sigMatrix[10][71] , 
        \sigMatrix[10][70] , \sigMatrix[10][69] , \sigMatrix[10][68] , 
        \sigMatrix[10][67] , \sigMatrix[10][66] , \sigMatrix[10][65] , 
        SYNOPSYS_UNCONNECTED__10}), .nextSum({\sigMatrix[10][63] , 
        \sigMatrix[10][62] , \sigMatrix[10][61] , \sigMatrix[10][60] , 
        \sigMatrix[10][59] , \sigMatrix[10][58] , \sigMatrix[10][57] , 
        \sigMatrix[10][56] , \sigMatrix[10][55] , \sigMatrix[10][54] , 
        \sigMatrix[10][53] , \sigMatrix[10][52] , \sigMatrix[10][51] , 
        \sigMatrix[10][50] , \sigMatrix[10][49] , \sigMatrix[10][48] , 
        \sigMatrix[10][47] , \sigMatrix[10][46] , \sigMatrix[10][45] , 
        \sigMatrix[10][44] , \sigMatrix[10][43] , \sigMatrix[10][42] , 
        \sigMatrix[10][41] , \sigMatrix[10][40] , \sigMatrix[10][39] , 
        \sigMatrix[10][38] , \sigMatrix[10][37] , \sigMatrix[10][36] , 
        \sigMatrix[10][35] , \sigMatrix[10][34] , \sigMatrix[10][33] , 
        \sigMatrix[10][32] , \sigMatrix[10][31] , \sigMatrix[10][30] , 
        \sigMatrix[10][29] , \sigMatrix[10][28] , \sigMatrix[10][27] , 
        \sigMatrix[10][26] , \sigMatrix[10][25] , \sigMatrix[10][24] , 
        \sigMatrix[10][23] , \sigMatrix[10][22] , \sigMatrix[10][21] , 
        \sigMatrix[10][20] , \sigMatrix[10][19] , \sigMatrix[10][18] , 
        \sigMatrix[10][17] , \sigMatrix[10][16] , \sigMatrix[10][15] , 
        \sigMatrix[10][14] , \sigMatrix[10][13] , \sigMatrix[10][12] , 
        \sigMatrix[10][11] , \sigMatrix[10][10] , \sigMatrix[10][9] , 
        \sigMatrix[10][8] , \sigMatrix[10][7] , \sigMatrix[10][6] , 
        \sigMatrix[10][5] , \sigMatrix[10][4] , \sigMatrix[10][3] , 
        \sigMatrix[10][2] , \sigMatrix[10][1] , \sigMatrix[10][0] }) );
  booth_mul_row_N64_RADIX3_5 booth_mul_row_1_11 ( .prevA({\sigMatrix[10][127] , 
        \sigMatrix[10][126] , \sigMatrix[10][125] , \sigMatrix[10][124] , 
        \sigMatrix[10][123] , \sigMatrix[10][122] , \sigMatrix[10][121] , 
        \sigMatrix[10][120] , \sigMatrix[10][119] , \sigMatrix[10][118] , 
        \sigMatrix[10][117] , \sigMatrix[10][116] , \sigMatrix[10][115] , 
        \sigMatrix[10][114] , \sigMatrix[10][113] , \sigMatrix[10][112] , 
        \sigMatrix[10][111] , \sigMatrix[10][110] , \sigMatrix[10][109] , 
        \sigMatrix[10][108] , \sigMatrix[10][107] , \sigMatrix[10][106] , 
        \sigMatrix[10][105] , \sigMatrix[10][104] , \sigMatrix[10][103] , 
        \sigMatrix[10][102] , \sigMatrix[10][101] , \sigMatrix[10][100] , 
        \sigMatrix[10][99] , \sigMatrix[10][98] , \sigMatrix[10][97] , 
        \sigMatrix[10][96] , \sigMatrix[10][95] , \sigMatrix[10][94] , 
        \sigMatrix[10][93] , \sigMatrix[10][92] , \sigMatrix[10][91] , 
        \sigMatrix[10][90] , \sigMatrix[10][89] , \sigMatrix[10][88] , 
        \sigMatrix[10][87] , \sigMatrix[10][86] , \sigMatrix[10][85] , 
        \sigMatrix[10][84] , \sigMatrix[10][83] , \sigMatrix[10][82] , 
        \sigMatrix[10][81] , \sigMatrix[10][80] , \sigMatrix[10][79] , 
        \sigMatrix[10][78] , \sigMatrix[10][77] , \sigMatrix[10][76] , 
        \sigMatrix[10][75] , \sigMatrix[10][74] , \sigMatrix[10][73] , 
        \sigMatrix[10][72] , \sigMatrix[10][71] , \sigMatrix[10][70] , 
        \sigMatrix[10][69] , \sigMatrix[10][68] , \sigMatrix[10][67] , 
        \sigMatrix[10][66] , \sigMatrix[10][65] , 1'b0}), .prevSum({
        \sigMatrix[10][63] , \sigMatrix[10][62] , \sigMatrix[10][61] , 
        \sigMatrix[10][60] , \sigMatrix[10][59] , \sigMatrix[10][58] , 
        \sigMatrix[10][57] , \sigMatrix[10][56] , \sigMatrix[10][55] , 
        \sigMatrix[10][54] , \sigMatrix[10][53] , \sigMatrix[10][52] , 
        \sigMatrix[10][51] , \sigMatrix[10][50] , \sigMatrix[10][49] , 
        \sigMatrix[10][48] , \sigMatrix[10][47] , \sigMatrix[10][46] , 
        \sigMatrix[10][45] , \sigMatrix[10][44] , \sigMatrix[10][43] , 
        \sigMatrix[10][42] , \sigMatrix[10][41] , \sigMatrix[10][40] , 
        \sigMatrix[10][39] , \sigMatrix[10][38] , \sigMatrix[10][37] , 
        \sigMatrix[10][36] , \sigMatrix[10][35] , \sigMatrix[10][34] , 
        \sigMatrix[10][33] , \sigMatrix[10][32] , \sigMatrix[10][31] , 
        \sigMatrix[10][30] , \sigMatrix[10][29] , \sigMatrix[10][28] , 
        \sigMatrix[10][27] , \sigMatrix[10][26] , \sigMatrix[10][25] , 
        \sigMatrix[10][24] , \sigMatrix[10][23] , \sigMatrix[10][22] , 
        \sigMatrix[10][21] , \sigMatrix[10][20] , \sigMatrix[10][19] , 
        \sigMatrix[10][18] , \sigMatrix[10][17] , \sigMatrix[10][16] , 
        \sigMatrix[10][15] , \sigMatrix[10][14] , \sigMatrix[10][13] , 
        \sigMatrix[10][12] , \sigMatrix[10][11] , \sigMatrix[10][10] , 
        \sigMatrix[10][9] , \sigMatrix[10][8] , \sigMatrix[10][7] , 
        \sigMatrix[10][6] , \sigMatrix[10][5] , \sigMatrix[10][4] , 
        \sigMatrix[10][3] , \sigMatrix[10][2] , \sigMatrix[10][1] , 
        \sigMatrix[10][0] }), .encoderIn(B_out_s[23:21]), .nextA({
        \sigMatrix[11][127] , \sigMatrix[11][126] , \sigMatrix[11][125] , 
        \sigMatrix[11][124] , \sigMatrix[11][123] , \sigMatrix[11][122] , 
        \sigMatrix[11][121] , \sigMatrix[11][120] , \sigMatrix[11][119] , 
        \sigMatrix[11][118] , \sigMatrix[11][117] , \sigMatrix[11][116] , 
        \sigMatrix[11][115] , \sigMatrix[11][114] , \sigMatrix[11][113] , 
        \sigMatrix[11][112] , \sigMatrix[11][111] , \sigMatrix[11][110] , 
        \sigMatrix[11][109] , \sigMatrix[11][108] , \sigMatrix[11][107] , 
        \sigMatrix[11][106] , \sigMatrix[11][105] , \sigMatrix[11][104] , 
        \sigMatrix[11][103] , \sigMatrix[11][102] , \sigMatrix[11][101] , 
        \sigMatrix[11][100] , \sigMatrix[11][99] , \sigMatrix[11][98] , 
        \sigMatrix[11][97] , \sigMatrix[11][96] , \sigMatrix[11][95] , 
        \sigMatrix[11][94] , \sigMatrix[11][93] , \sigMatrix[11][92] , 
        \sigMatrix[11][91] , \sigMatrix[11][90] , \sigMatrix[11][89] , 
        \sigMatrix[11][88] , \sigMatrix[11][87] , \sigMatrix[11][86] , 
        \sigMatrix[11][85] , \sigMatrix[11][84] , \sigMatrix[11][83] , 
        \sigMatrix[11][82] , \sigMatrix[11][81] , \sigMatrix[11][80] , 
        \sigMatrix[11][79] , \sigMatrix[11][78] , \sigMatrix[11][77] , 
        \sigMatrix[11][76] , \sigMatrix[11][75] , \sigMatrix[11][74] , 
        \sigMatrix[11][73] , \sigMatrix[11][72] , \sigMatrix[11][71] , 
        \sigMatrix[11][70] , \sigMatrix[11][69] , \sigMatrix[11][68] , 
        \sigMatrix[11][67] , \sigMatrix[11][66] , \sigMatrix[11][65] , 
        SYNOPSYS_UNCONNECTED__11}), .nextSum({\sigMatrix[11][63] , 
        \sigMatrix[11][62] , \sigMatrix[11][61] , \sigMatrix[11][60] , 
        \sigMatrix[11][59] , \sigMatrix[11][58] , \sigMatrix[11][57] , 
        \sigMatrix[11][56] , \sigMatrix[11][55] , \sigMatrix[11][54] , 
        \sigMatrix[11][53] , \sigMatrix[11][52] , \sigMatrix[11][51] , 
        \sigMatrix[11][50] , \sigMatrix[11][49] , \sigMatrix[11][48] , 
        \sigMatrix[11][47] , \sigMatrix[11][46] , \sigMatrix[11][45] , 
        \sigMatrix[11][44] , \sigMatrix[11][43] , \sigMatrix[11][42] , 
        \sigMatrix[11][41] , \sigMatrix[11][40] , \sigMatrix[11][39] , 
        \sigMatrix[11][38] , \sigMatrix[11][37] , \sigMatrix[11][36] , 
        \sigMatrix[11][35] , \sigMatrix[11][34] , \sigMatrix[11][33] , 
        \sigMatrix[11][32] , \sigMatrix[11][31] , \sigMatrix[11][30] , 
        \sigMatrix[11][29] , \sigMatrix[11][28] , \sigMatrix[11][27] , 
        \sigMatrix[11][26] , \sigMatrix[11][25] , \sigMatrix[11][24] , 
        \sigMatrix[11][23] , \sigMatrix[11][22] , \sigMatrix[11][21] , 
        \sigMatrix[11][20] , \sigMatrix[11][19] , \sigMatrix[11][18] , 
        \sigMatrix[11][17] , \sigMatrix[11][16] , \sigMatrix[11][15] , 
        \sigMatrix[11][14] , \sigMatrix[11][13] , \sigMatrix[11][12] , 
        \sigMatrix[11][11] , \sigMatrix[11][10] , \sigMatrix[11][9] , 
        \sigMatrix[11][8] , \sigMatrix[11][7] , \sigMatrix[11][6] , 
        \sigMatrix[11][5] , \sigMatrix[11][4] , \sigMatrix[11][3] , 
        \sigMatrix[11][2] , \sigMatrix[11][1] , \sigMatrix[11][0] }) );
  booth_mul_row_N64_RADIX3_4 booth_mul_row_1_12 ( .prevA({\sigMatrix[11][127] , 
        \sigMatrix[11][126] , \sigMatrix[11][125] , \sigMatrix[11][124] , 
        \sigMatrix[11][123] , \sigMatrix[11][122] , \sigMatrix[11][121] , 
        \sigMatrix[11][120] , \sigMatrix[11][119] , \sigMatrix[11][118] , 
        \sigMatrix[11][117] , \sigMatrix[11][116] , \sigMatrix[11][115] , 
        \sigMatrix[11][114] , \sigMatrix[11][113] , \sigMatrix[11][112] , 
        \sigMatrix[11][111] , \sigMatrix[11][110] , \sigMatrix[11][109] , 
        \sigMatrix[11][108] , \sigMatrix[11][107] , \sigMatrix[11][106] , 
        \sigMatrix[11][105] , \sigMatrix[11][104] , \sigMatrix[11][103] , 
        \sigMatrix[11][102] , \sigMatrix[11][101] , \sigMatrix[11][100] , 
        \sigMatrix[11][99] , \sigMatrix[11][98] , \sigMatrix[11][97] , 
        \sigMatrix[11][96] , \sigMatrix[11][95] , \sigMatrix[11][94] , 
        \sigMatrix[11][93] , \sigMatrix[11][92] , \sigMatrix[11][91] , 
        \sigMatrix[11][90] , \sigMatrix[11][89] , \sigMatrix[11][88] , 
        \sigMatrix[11][87] , \sigMatrix[11][86] , \sigMatrix[11][85] , 
        \sigMatrix[11][84] , \sigMatrix[11][83] , \sigMatrix[11][82] , 
        \sigMatrix[11][81] , \sigMatrix[11][80] , \sigMatrix[11][79] , 
        \sigMatrix[11][78] , \sigMatrix[11][77] , \sigMatrix[11][76] , 
        \sigMatrix[11][75] , \sigMatrix[11][74] , \sigMatrix[11][73] , 
        \sigMatrix[11][72] , \sigMatrix[11][71] , \sigMatrix[11][70] , 
        \sigMatrix[11][69] , \sigMatrix[11][68] , \sigMatrix[11][67] , 
        \sigMatrix[11][66] , \sigMatrix[11][65] , 1'b0}), .prevSum({
        \sigMatrix[11][63] , \sigMatrix[11][62] , \sigMatrix[11][61] , 
        \sigMatrix[11][60] , \sigMatrix[11][59] , \sigMatrix[11][58] , 
        \sigMatrix[11][57] , \sigMatrix[11][56] , \sigMatrix[11][55] , 
        \sigMatrix[11][54] , \sigMatrix[11][53] , \sigMatrix[11][52] , 
        \sigMatrix[11][51] , \sigMatrix[11][50] , \sigMatrix[11][49] , 
        \sigMatrix[11][48] , \sigMatrix[11][47] , \sigMatrix[11][46] , 
        \sigMatrix[11][45] , \sigMatrix[11][44] , \sigMatrix[11][43] , 
        \sigMatrix[11][42] , \sigMatrix[11][41] , \sigMatrix[11][40] , 
        \sigMatrix[11][39] , \sigMatrix[11][38] , \sigMatrix[11][37] , 
        \sigMatrix[11][36] , \sigMatrix[11][35] , \sigMatrix[11][34] , 
        \sigMatrix[11][33] , \sigMatrix[11][32] , \sigMatrix[11][31] , 
        \sigMatrix[11][30] , \sigMatrix[11][29] , \sigMatrix[11][28] , 
        \sigMatrix[11][27] , \sigMatrix[11][26] , \sigMatrix[11][25] , 
        \sigMatrix[11][24] , \sigMatrix[11][23] , \sigMatrix[11][22] , 
        \sigMatrix[11][21] , \sigMatrix[11][20] , \sigMatrix[11][19] , 
        \sigMatrix[11][18] , \sigMatrix[11][17] , \sigMatrix[11][16] , 
        \sigMatrix[11][15] , \sigMatrix[11][14] , \sigMatrix[11][13] , 
        \sigMatrix[11][12] , \sigMatrix[11][11] , \sigMatrix[11][10] , 
        \sigMatrix[11][9] , \sigMatrix[11][8] , \sigMatrix[11][7] , 
        \sigMatrix[11][6] , \sigMatrix[11][5] , \sigMatrix[11][4] , 
        \sigMatrix[11][3] , \sigMatrix[11][2] , \sigMatrix[11][1] , 
        \sigMatrix[11][0] }), .encoderIn(B_out_s[25:23]), .nextA({
        \sigMatrix[12][127] , \sigMatrix[12][126] , \sigMatrix[12][125] , 
        \sigMatrix[12][124] , \sigMatrix[12][123] , \sigMatrix[12][122] , 
        \sigMatrix[12][121] , \sigMatrix[12][120] , \sigMatrix[12][119] , 
        \sigMatrix[12][118] , \sigMatrix[12][117] , \sigMatrix[12][116] , 
        \sigMatrix[12][115] , \sigMatrix[12][114] , \sigMatrix[12][113] , 
        \sigMatrix[12][112] , \sigMatrix[12][111] , \sigMatrix[12][110] , 
        \sigMatrix[12][109] , \sigMatrix[12][108] , \sigMatrix[12][107] , 
        \sigMatrix[12][106] , \sigMatrix[12][105] , \sigMatrix[12][104] , 
        \sigMatrix[12][103] , \sigMatrix[12][102] , \sigMatrix[12][101] , 
        \sigMatrix[12][100] , \sigMatrix[12][99] , \sigMatrix[12][98] , 
        \sigMatrix[12][97] , \sigMatrix[12][96] , \sigMatrix[12][95] , 
        \sigMatrix[12][94] , \sigMatrix[12][93] , \sigMatrix[12][92] , 
        \sigMatrix[12][91] , \sigMatrix[12][90] , \sigMatrix[12][89] , 
        \sigMatrix[12][88] , \sigMatrix[12][87] , \sigMatrix[12][86] , 
        \sigMatrix[12][85] , \sigMatrix[12][84] , \sigMatrix[12][83] , 
        \sigMatrix[12][82] , \sigMatrix[12][81] , \sigMatrix[12][80] , 
        \sigMatrix[12][79] , \sigMatrix[12][78] , \sigMatrix[12][77] , 
        \sigMatrix[12][76] , \sigMatrix[12][75] , \sigMatrix[12][74] , 
        \sigMatrix[12][73] , \sigMatrix[12][72] , \sigMatrix[12][71] , 
        \sigMatrix[12][70] , \sigMatrix[12][69] , \sigMatrix[12][68] , 
        \sigMatrix[12][67] , \sigMatrix[12][66] , \sigMatrix[12][65] , 
        SYNOPSYS_UNCONNECTED__12}), .nextSum({\sigMatrix[12][63] , 
        \sigMatrix[12][62] , \sigMatrix[12][61] , \sigMatrix[12][60] , 
        \sigMatrix[12][59] , \sigMatrix[12][58] , \sigMatrix[12][57] , 
        \sigMatrix[12][56] , \sigMatrix[12][55] , \sigMatrix[12][54] , 
        \sigMatrix[12][53] , \sigMatrix[12][52] , \sigMatrix[12][51] , 
        \sigMatrix[12][50] , \sigMatrix[12][49] , \sigMatrix[12][48] , 
        \sigMatrix[12][47] , \sigMatrix[12][46] , \sigMatrix[12][45] , 
        \sigMatrix[12][44] , \sigMatrix[12][43] , \sigMatrix[12][42] , 
        \sigMatrix[12][41] , \sigMatrix[12][40] , \sigMatrix[12][39] , 
        \sigMatrix[12][38] , \sigMatrix[12][37] , \sigMatrix[12][36] , 
        \sigMatrix[12][35] , \sigMatrix[12][34] , \sigMatrix[12][33] , 
        \sigMatrix[12][32] , \sigMatrix[12][31] , \sigMatrix[12][30] , 
        \sigMatrix[12][29] , \sigMatrix[12][28] , \sigMatrix[12][27] , 
        \sigMatrix[12][26] , \sigMatrix[12][25] , \sigMatrix[12][24] , 
        \sigMatrix[12][23] , \sigMatrix[12][22] , \sigMatrix[12][21] , 
        \sigMatrix[12][20] , \sigMatrix[12][19] , \sigMatrix[12][18] , 
        \sigMatrix[12][17] , \sigMatrix[12][16] , \sigMatrix[12][15] , 
        \sigMatrix[12][14] , \sigMatrix[12][13] , \sigMatrix[12][12] , 
        \sigMatrix[12][11] , \sigMatrix[12][10] , \sigMatrix[12][9] , 
        \sigMatrix[12][8] , \sigMatrix[12][7] , \sigMatrix[12][6] , 
        \sigMatrix[12][5] , \sigMatrix[12][4] , \sigMatrix[12][3] , 
        \sigMatrix[12][2] , \sigMatrix[12][1] , \sigMatrix[12][0] }) );
  booth_mul_row_N64_RADIX3_3 booth_mul_row_1_13 ( .prevA({\sigMatrix[12][127] , 
        \sigMatrix[12][126] , \sigMatrix[12][125] , \sigMatrix[12][124] , 
        \sigMatrix[12][123] , \sigMatrix[12][122] , \sigMatrix[12][121] , 
        \sigMatrix[12][120] , \sigMatrix[12][119] , \sigMatrix[12][118] , 
        \sigMatrix[12][117] , \sigMatrix[12][116] , \sigMatrix[12][115] , 
        \sigMatrix[12][114] , \sigMatrix[12][113] , \sigMatrix[12][112] , 
        \sigMatrix[12][111] , \sigMatrix[12][110] , \sigMatrix[12][109] , 
        \sigMatrix[12][108] , \sigMatrix[12][107] , \sigMatrix[12][106] , 
        \sigMatrix[12][105] , \sigMatrix[12][104] , \sigMatrix[12][103] , 
        \sigMatrix[12][102] , \sigMatrix[12][101] , \sigMatrix[12][100] , 
        \sigMatrix[12][99] , \sigMatrix[12][98] , \sigMatrix[12][97] , 
        \sigMatrix[12][96] , \sigMatrix[12][95] , \sigMatrix[12][94] , 
        \sigMatrix[12][93] , \sigMatrix[12][92] , \sigMatrix[12][91] , 
        \sigMatrix[12][90] , \sigMatrix[12][89] , \sigMatrix[12][88] , 
        \sigMatrix[12][87] , \sigMatrix[12][86] , \sigMatrix[12][85] , 
        \sigMatrix[12][84] , \sigMatrix[12][83] , \sigMatrix[12][82] , 
        \sigMatrix[12][81] , \sigMatrix[12][80] , \sigMatrix[12][79] , 
        \sigMatrix[12][78] , \sigMatrix[12][77] , \sigMatrix[12][76] , 
        \sigMatrix[12][75] , \sigMatrix[12][74] , \sigMatrix[12][73] , 
        \sigMatrix[12][72] , \sigMatrix[12][71] , \sigMatrix[12][70] , 
        \sigMatrix[12][69] , \sigMatrix[12][68] , \sigMatrix[12][67] , 
        \sigMatrix[12][66] , \sigMatrix[12][65] , 1'b0}), .prevSum({
        \sigMatrix[12][63] , \sigMatrix[12][62] , \sigMatrix[12][61] , 
        \sigMatrix[12][60] , \sigMatrix[12][59] , \sigMatrix[12][58] , 
        \sigMatrix[12][57] , \sigMatrix[12][56] , \sigMatrix[12][55] , 
        \sigMatrix[12][54] , \sigMatrix[12][53] , \sigMatrix[12][52] , 
        \sigMatrix[12][51] , \sigMatrix[12][50] , \sigMatrix[12][49] , 
        \sigMatrix[12][48] , \sigMatrix[12][47] , \sigMatrix[12][46] , 
        \sigMatrix[12][45] , \sigMatrix[12][44] , \sigMatrix[12][43] , 
        \sigMatrix[12][42] , \sigMatrix[12][41] , \sigMatrix[12][40] , 
        \sigMatrix[12][39] , \sigMatrix[12][38] , \sigMatrix[12][37] , 
        \sigMatrix[12][36] , \sigMatrix[12][35] , \sigMatrix[12][34] , 
        \sigMatrix[12][33] , \sigMatrix[12][32] , \sigMatrix[12][31] , 
        \sigMatrix[12][30] , \sigMatrix[12][29] , \sigMatrix[12][28] , 
        \sigMatrix[12][27] , \sigMatrix[12][26] , \sigMatrix[12][25] , 
        \sigMatrix[12][24] , \sigMatrix[12][23] , \sigMatrix[12][22] , 
        \sigMatrix[12][21] , \sigMatrix[12][20] , \sigMatrix[12][19] , 
        \sigMatrix[12][18] , \sigMatrix[12][17] , \sigMatrix[12][16] , 
        \sigMatrix[12][15] , \sigMatrix[12][14] , \sigMatrix[12][13] , 
        \sigMatrix[12][12] , \sigMatrix[12][11] , \sigMatrix[12][10] , 
        \sigMatrix[12][9] , \sigMatrix[12][8] , \sigMatrix[12][7] , 
        \sigMatrix[12][6] , \sigMatrix[12][5] , \sigMatrix[12][4] , 
        \sigMatrix[12][3] , \sigMatrix[12][2] , \sigMatrix[12][1] , 
        \sigMatrix[12][0] }), .encoderIn(B_out_s[27:25]), .nextA({
        \sigMatrix[13][127] , \sigMatrix[13][126] , \sigMatrix[13][125] , 
        \sigMatrix[13][124] , \sigMatrix[13][123] , \sigMatrix[13][122] , 
        \sigMatrix[13][121] , \sigMatrix[13][120] , \sigMatrix[13][119] , 
        \sigMatrix[13][118] , \sigMatrix[13][117] , \sigMatrix[13][116] , 
        \sigMatrix[13][115] , \sigMatrix[13][114] , \sigMatrix[13][113] , 
        \sigMatrix[13][112] , \sigMatrix[13][111] , \sigMatrix[13][110] , 
        \sigMatrix[13][109] , \sigMatrix[13][108] , \sigMatrix[13][107] , 
        \sigMatrix[13][106] , \sigMatrix[13][105] , \sigMatrix[13][104] , 
        \sigMatrix[13][103] , \sigMatrix[13][102] , \sigMatrix[13][101] , 
        \sigMatrix[13][100] , \sigMatrix[13][99] , \sigMatrix[13][98] , 
        \sigMatrix[13][97] , \sigMatrix[13][96] , \sigMatrix[13][95] , 
        \sigMatrix[13][94] , \sigMatrix[13][93] , \sigMatrix[13][92] , 
        \sigMatrix[13][91] , \sigMatrix[13][90] , \sigMatrix[13][89] , 
        \sigMatrix[13][88] , \sigMatrix[13][87] , \sigMatrix[13][86] , 
        \sigMatrix[13][85] , \sigMatrix[13][84] , \sigMatrix[13][83] , 
        \sigMatrix[13][82] , \sigMatrix[13][81] , \sigMatrix[13][80] , 
        \sigMatrix[13][79] , \sigMatrix[13][78] , \sigMatrix[13][77] , 
        \sigMatrix[13][76] , \sigMatrix[13][75] , \sigMatrix[13][74] , 
        \sigMatrix[13][73] , \sigMatrix[13][72] , \sigMatrix[13][71] , 
        \sigMatrix[13][70] , \sigMatrix[13][69] , \sigMatrix[13][68] , 
        \sigMatrix[13][67] , \sigMatrix[13][66] , \sigMatrix[13][65] , 
        SYNOPSYS_UNCONNECTED__13}), .nextSum({\sigMatrix[13][63] , 
        \sigMatrix[13][62] , \sigMatrix[13][61] , \sigMatrix[13][60] , 
        \sigMatrix[13][59] , \sigMatrix[13][58] , \sigMatrix[13][57] , 
        \sigMatrix[13][56] , \sigMatrix[13][55] , \sigMatrix[13][54] , 
        \sigMatrix[13][53] , \sigMatrix[13][52] , \sigMatrix[13][51] , 
        \sigMatrix[13][50] , \sigMatrix[13][49] , \sigMatrix[13][48] , 
        \sigMatrix[13][47] , \sigMatrix[13][46] , \sigMatrix[13][45] , 
        \sigMatrix[13][44] , \sigMatrix[13][43] , \sigMatrix[13][42] , 
        \sigMatrix[13][41] , \sigMatrix[13][40] , \sigMatrix[13][39] , 
        \sigMatrix[13][38] , \sigMatrix[13][37] , \sigMatrix[13][36] , 
        \sigMatrix[13][35] , \sigMatrix[13][34] , \sigMatrix[13][33] , 
        \sigMatrix[13][32] , \sigMatrix[13][31] , \sigMatrix[13][30] , 
        \sigMatrix[13][29] , \sigMatrix[13][28] , \sigMatrix[13][27] , 
        \sigMatrix[13][26] , \sigMatrix[13][25] , \sigMatrix[13][24] , 
        \sigMatrix[13][23] , \sigMatrix[13][22] , \sigMatrix[13][21] , 
        \sigMatrix[13][20] , \sigMatrix[13][19] , \sigMatrix[13][18] , 
        \sigMatrix[13][17] , \sigMatrix[13][16] , \sigMatrix[13][15] , 
        \sigMatrix[13][14] , \sigMatrix[13][13] , \sigMatrix[13][12] , 
        \sigMatrix[13][11] , \sigMatrix[13][10] , \sigMatrix[13][9] , 
        \sigMatrix[13][8] , \sigMatrix[13][7] , \sigMatrix[13][6] , 
        \sigMatrix[13][5] , \sigMatrix[13][4] , \sigMatrix[13][3] , 
        \sigMatrix[13][2] , \sigMatrix[13][1] , \sigMatrix[13][0] }) );
  booth_mul_row_N64_RADIX3_2 booth_mul_row_1_14 ( .prevA({\sigMatrix[13][127] , 
        \sigMatrix[13][126] , \sigMatrix[13][125] , \sigMatrix[13][124] , 
        \sigMatrix[13][123] , \sigMatrix[13][122] , \sigMatrix[13][121] , 
        \sigMatrix[13][120] , \sigMatrix[13][119] , \sigMatrix[13][118] , 
        \sigMatrix[13][117] , \sigMatrix[13][116] , \sigMatrix[13][115] , 
        \sigMatrix[13][114] , \sigMatrix[13][113] , \sigMatrix[13][112] , 
        \sigMatrix[13][111] , \sigMatrix[13][110] , \sigMatrix[13][109] , 
        \sigMatrix[13][108] , \sigMatrix[13][107] , \sigMatrix[13][106] , 
        \sigMatrix[13][105] , \sigMatrix[13][104] , \sigMatrix[13][103] , 
        \sigMatrix[13][102] , \sigMatrix[13][101] , \sigMatrix[13][100] , 
        \sigMatrix[13][99] , \sigMatrix[13][98] , \sigMatrix[13][97] , 
        \sigMatrix[13][96] , \sigMatrix[13][95] , \sigMatrix[13][94] , 
        \sigMatrix[13][93] , \sigMatrix[13][92] , \sigMatrix[13][91] , 
        \sigMatrix[13][90] , \sigMatrix[13][89] , \sigMatrix[13][88] , 
        \sigMatrix[13][87] , \sigMatrix[13][86] , \sigMatrix[13][85] , 
        \sigMatrix[13][84] , \sigMatrix[13][83] , \sigMatrix[13][82] , 
        \sigMatrix[13][81] , \sigMatrix[13][80] , \sigMatrix[13][79] , 
        \sigMatrix[13][78] , \sigMatrix[13][77] , \sigMatrix[13][76] , 
        \sigMatrix[13][75] , \sigMatrix[13][74] , \sigMatrix[13][73] , 
        \sigMatrix[13][72] , \sigMatrix[13][71] , \sigMatrix[13][70] , 
        \sigMatrix[13][69] , \sigMatrix[13][68] , \sigMatrix[13][67] , 
        \sigMatrix[13][66] , \sigMatrix[13][65] , 1'b0}), .prevSum({
        \sigMatrix[13][63] , \sigMatrix[13][62] , \sigMatrix[13][61] , 
        \sigMatrix[13][60] , \sigMatrix[13][59] , \sigMatrix[13][58] , 
        \sigMatrix[13][57] , \sigMatrix[13][56] , \sigMatrix[13][55] , 
        \sigMatrix[13][54] , \sigMatrix[13][53] , \sigMatrix[13][52] , 
        \sigMatrix[13][51] , \sigMatrix[13][50] , \sigMatrix[13][49] , 
        \sigMatrix[13][48] , \sigMatrix[13][47] , \sigMatrix[13][46] , 
        \sigMatrix[13][45] , \sigMatrix[13][44] , \sigMatrix[13][43] , 
        \sigMatrix[13][42] , \sigMatrix[13][41] , \sigMatrix[13][40] , 
        \sigMatrix[13][39] , \sigMatrix[13][38] , \sigMatrix[13][37] , 
        \sigMatrix[13][36] , \sigMatrix[13][35] , \sigMatrix[13][34] , 
        \sigMatrix[13][33] , \sigMatrix[13][32] , \sigMatrix[13][31] , 
        \sigMatrix[13][30] , \sigMatrix[13][29] , \sigMatrix[13][28] , 
        \sigMatrix[13][27] , \sigMatrix[13][26] , \sigMatrix[13][25] , 
        \sigMatrix[13][24] , \sigMatrix[13][23] , \sigMatrix[13][22] , 
        \sigMatrix[13][21] , \sigMatrix[13][20] , \sigMatrix[13][19] , 
        \sigMatrix[13][18] , \sigMatrix[13][17] , \sigMatrix[13][16] , 
        \sigMatrix[13][15] , \sigMatrix[13][14] , \sigMatrix[13][13] , 
        \sigMatrix[13][12] , \sigMatrix[13][11] , \sigMatrix[13][10] , 
        \sigMatrix[13][9] , \sigMatrix[13][8] , \sigMatrix[13][7] , 
        \sigMatrix[13][6] , \sigMatrix[13][5] , \sigMatrix[13][4] , 
        \sigMatrix[13][3] , \sigMatrix[13][2] , \sigMatrix[13][1] , 
        \sigMatrix[13][0] }), .encoderIn(B_out_s[29:27]), .nextA({
        \sigMatrix[14][127] , \sigMatrix[14][126] , \sigMatrix[14][125] , 
        \sigMatrix[14][124] , \sigMatrix[14][123] , \sigMatrix[14][122] , 
        \sigMatrix[14][121] , \sigMatrix[14][120] , \sigMatrix[14][119] , 
        \sigMatrix[14][118] , \sigMatrix[14][117] , \sigMatrix[14][116] , 
        \sigMatrix[14][115] , \sigMatrix[14][114] , \sigMatrix[14][113] , 
        \sigMatrix[14][112] , \sigMatrix[14][111] , \sigMatrix[14][110] , 
        \sigMatrix[14][109] , \sigMatrix[14][108] , \sigMatrix[14][107] , 
        \sigMatrix[14][106] , \sigMatrix[14][105] , \sigMatrix[14][104] , 
        \sigMatrix[14][103] , \sigMatrix[14][102] , \sigMatrix[14][101] , 
        \sigMatrix[14][100] , \sigMatrix[14][99] , \sigMatrix[14][98] , 
        \sigMatrix[14][97] , \sigMatrix[14][96] , \sigMatrix[14][95] , 
        \sigMatrix[14][94] , \sigMatrix[14][93] , \sigMatrix[14][92] , 
        \sigMatrix[14][91] , \sigMatrix[14][90] , \sigMatrix[14][89] , 
        \sigMatrix[14][88] , \sigMatrix[14][87] , \sigMatrix[14][86] , 
        \sigMatrix[14][85] , \sigMatrix[14][84] , \sigMatrix[14][83] , 
        \sigMatrix[14][82] , \sigMatrix[14][81] , \sigMatrix[14][80] , 
        \sigMatrix[14][79] , \sigMatrix[14][78] , \sigMatrix[14][77] , 
        \sigMatrix[14][76] , \sigMatrix[14][75] , \sigMatrix[14][74] , 
        \sigMatrix[14][73] , \sigMatrix[14][72] , \sigMatrix[14][71] , 
        \sigMatrix[14][70] , \sigMatrix[14][69] , \sigMatrix[14][68] , 
        \sigMatrix[14][67] , \sigMatrix[14][66] , \sigMatrix[14][65] , 
        SYNOPSYS_UNCONNECTED__14}), .nextSum({\sigMatrix[14][63] , 
        \sigMatrix[14][62] , \sigMatrix[14][61] , \sigMatrix[14][60] , 
        \sigMatrix[14][59] , \sigMatrix[14][58] , \sigMatrix[14][57] , 
        \sigMatrix[14][56] , \sigMatrix[14][55] , \sigMatrix[14][54] , 
        \sigMatrix[14][53] , \sigMatrix[14][52] , \sigMatrix[14][51] , 
        \sigMatrix[14][50] , \sigMatrix[14][49] , \sigMatrix[14][48] , 
        \sigMatrix[14][47] , \sigMatrix[14][46] , \sigMatrix[14][45] , 
        \sigMatrix[14][44] , \sigMatrix[14][43] , \sigMatrix[14][42] , 
        \sigMatrix[14][41] , \sigMatrix[14][40] , \sigMatrix[14][39] , 
        \sigMatrix[14][38] , \sigMatrix[14][37] , \sigMatrix[14][36] , 
        \sigMatrix[14][35] , \sigMatrix[14][34] , \sigMatrix[14][33] , 
        \sigMatrix[14][32] , \sigMatrix[14][31] , \sigMatrix[14][30] , 
        \sigMatrix[14][29] , \sigMatrix[14][28] , \sigMatrix[14][27] , 
        \sigMatrix[14][26] , \sigMatrix[14][25] , \sigMatrix[14][24] , 
        \sigMatrix[14][23] , \sigMatrix[14][22] , \sigMatrix[14][21] , 
        \sigMatrix[14][20] , \sigMatrix[14][19] , \sigMatrix[14][18] , 
        \sigMatrix[14][17] , \sigMatrix[14][16] , \sigMatrix[14][15] , 
        \sigMatrix[14][14] , \sigMatrix[14][13] , \sigMatrix[14][12] , 
        \sigMatrix[14][11] , \sigMatrix[14][10] , \sigMatrix[14][9] , 
        \sigMatrix[14][8] , \sigMatrix[14][7] , \sigMatrix[14][6] , 
        \sigMatrix[14][5] , \sigMatrix[14][4] , \sigMatrix[14][3] , 
        \sigMatrix[14][2] , \sigMatrix[14][1] , \sigMatrix[14][0] }) );
  booth_mul_row_N64_RADIX3_1 booth_mul_row_1_15 ( .prevA({\sigMatrix[14][127] , 
        \sigMatrix[14][126] , \sigMatrix[14][125] , \sigMatrix[14][124] , 
        \sigMatrix[14][123] , \sigMatrix[14][122] , \sigMatrix[14][121] , 
        \sigMatrix[14][120] , \sigMatrix[14][119] , \sigMatrix[14][118] , 
        \sigMatrix[14][117] , \sigMatrix[14][116] , \sigMatrix[14][115] , 
        \sigMatrix[14][114] , \sigMatrix[14][113] , \sigMatrix[14][112] , 
        \sigMatrix[14][111] , \sigMatrix[14][110] , \sigMatrix[14][109] , 
        \sigMatrix[14][108] , \sigMatrix[14][107] , \sigMatrix[14][106] , 
        \sigMatrix[14][105] , \sigMatrix[14][104] , \sigMatrix[14][103] , 
        \sigMatrix[14][102] , \sigMatrix[14][101] , \sigMatrix[14][100] , 
        \sigMatrix[14][99] , \sigMatrix[14][98] , \sigMatrix[14][97] , 
        \sigMatrix[14][96] , \sigMatrix[14][95] , \sigMatrix[14][94] , 
        \sigMatrix[14][93] , \sigMatrix[14][92] , \sigMatrix[14][91] , 
        \sigMatrix[14][90] , \sigMatrix[14][89] , \sigMatrix[14][88] , 
        \sigMatrix[14][87] , \sigMatrix[14][86] , \sigMatrix[14][85] , 
        \sigMatrix[14][84] , \sigMatrix[14][83] , \sigMatrix[14][82] , 
        \sigMatrix[14][81] , \sigMatrix[14][80] , \sigMatrix[14][79] , 
        \sigMatrix[14][78] , \sigMatrix[14][77] , \sigMatrix[14][76] , 
        \sigMatrix[14][75] , \sigMatrix[14][74] , \sigMatrix[14][73] , 
        \sigMatrix[14][72] , \sigMatrix[14][71] , \sigMatrix[14][70] , 
        \sigMatrix[14][69] , \sigMatrix[14][68] , \sigMatrix[14][67] , 
        \sigMatrix[14][66] , \sigMatrix[14][65] , 1'b0}), .prevSum({
        \sigMatrix[14][63] , \sigMatrix[14][62] , \sigMatrix[14][61] , 
        \sigMatrix[14][60] , \sigMatrix[14][59] , \sigMatrix[14][58] , 
        \sigMatrix[14][57] , \sigMatrix[14][56] , \sigMatrix[14][55] , 
        \sigMatrix[14][54] , \sigMatrix[14][53] , \sigMatrix[14][52] , 
        \sigMatrix[14][51] , \sigMatrix[14][50] , \sigMatrix[14][49] , 
        \sigMatrix[14][48] , \sigMatrix[14][47] , \sigMatrix[14][46] , 
        \sigMatrix[14][45] , \sigMatrix[14][44] , \sigMatrix[14][43] , 
        \sigMatrix[14][42] , \sigMatrix[14][41] , \sigMatrix[14][40] , 
        \sigMatrix[14][39] , \sigMatrix[14][38] , \sigMatrix[14][37] , 
        \sigMatrix[14][36] , \sigMatrix[14][35] , \sigMatrix[14][34] , 
        \sigMatrix[14][33] , \sigMatrix[14][32] , \sigMatrix[14][31] , 
        \sigMatrix[14][30] , \sigMatrix[14][29] , \sigMatrix[14][28] , 
        \sigMatrix[14][27] , \sigMatrix[14][26] , \sigMatrix[14][25] , 
        \sigMatrix[14][24] , \sigMatrix[14][23] , \sigMatrix[14][22] , 
        \sigMatrix[14][21] , \sigMatrix[14][20] , \sigMatrix[14][19] , 
        \sigMatrix[14][18] , \sigMatrix[14][17] , \sigMatrix[14][16] , 
        \sigMatrix[14][15] , \sigMatrix[14][14] , \sigMatrix[14][13] , 
        \sigMatrix[14][12] , \sigMatrix[14][11] , \sigMatrix[14][10] , 
        \sigMatrix[14][9] , \sigMatrix[14][8] , \sigMatrix[14][7] , 
        \sigMatrix[14][6] , \sigMatrix[14][5] , \sigMatrix[14][4] , 
        \sigMatrix[14][3] , \sigMatrix[14][2] , \sigMatrix[14][1] , 
        \sigMatrix[14][0] }), .encoderIn(B_out_s[31:29]), .nextSum(P_s) );
  registers_N32_1 regs_out ( .Clk(Clk), .Rst(Rst), .A(P_s[63:32]), .B(
        P_s[31:0]), .A_out(P[63:32]), .B_out(P[31:0]) );
  BUF_X2 U2 ( .A(n8), .Z(n12) );
  BUF_X2 U3 ( .A(n9), .Z(n13) );
  BUF_X2 U4 ( .A(n9), .Z(n14) );
  BUF_X2 U5 ( .A(n8), .Z(n11) );
  BUF_X2 U6 ( .A(n8), .Z(n10) );
  BUF_X1 U7 ( .A(n9), .Z(n15) );
  BUF_X1 U9 ( .A(A_out_s[31]), .Z(n8) );
  BUF_X1 U10 ( .A(A_out_s[31]), .Z(n9) );
endmodule

