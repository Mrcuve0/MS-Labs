
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_register_file is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_register_file;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_register_file.all;

entity register_file is

   port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
         std_logic_vector (63 downto 0);  OUT1, OUT2 : out std_logic_vector (63
         downto 0));

end register_file;

architecture SYN_beh of register_file is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal OUT2_63_port, OUT2_62_port, OUT2_61_port, OUT2_60_port, OUT2_59_port,
      OUT2_58_port, OUT2_57_port, OUT2_56_port, OUT2_55_port, OUT2_54_port, 
      OUT2_53_port, OUT2_52_port, OUT2_51_port, OUT2_50_port, OUT2_49_port, 
      OUT2_48_port, OUT2_47_port, OUT2_46_port, OUT2_45_port, OUT2_44_port, 
      OUT2_43_port, OUT2_42_port, OUT2_41_port, OUT2_40_port, OUT2_39_port, 
      OUT2_38_port, OUT2_37_port, OUT2_36_port, OUT2_35_port, OUT2_34_port, 
      OUT2_33_port, OUT2_32_port, OUT2_31_port, OUT2_30_port, OUT2_29_port, 
      OUT2_28_port, OUT2_27_port, OUT2_26_port, OUT2_25_port, OUT2_24_port, 
      OUT2_23_port, OUT2_22_port, OUT2_21_port, OUT2_20_port, OUT2_19_port, 
      OUT2_18_port, OUT2_17_port, OUT2_16_port, OUT2_15_port, OUT2_14_port, 
      OUT2_13_port, OUT2_12_port, OUT2_11_port, OUT2_10_port, OUT2_9_port, 
      OUT2_8_port, OUT2_7_port, OUT2_6_port, OUT2_5_port, OUT2_4_port, 
      OUT2_3_port, OUT2_2_port, OUT2_1_port, OUT2_0_port, n77, n78, n79, n80, 
      n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95
      , n96, n97, n98, n99, n833, n834, n835, n836, n837, n838, n839, n840, 
      n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, 
      n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, 
      n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, 
      n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, 
      n889, n890, n891, n892, n893, n894, n895, n896, n4932, n4933, n4934, 
      n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, 
      n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, 
      n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, 
      n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, 
      n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, 
      n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, 
      n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, 
      n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, 
      n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, 
      n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, 
      n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, 
      n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, 
      n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, 
      n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, 
      n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, 
      n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, 
      n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, 
      n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, 
      n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, 
      n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, 
      n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, 
      n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, 
      n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, 
      n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, 
      n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, 
      n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, 
      n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, 
      n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, 
      n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, 
      n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, 
      n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, 
      n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, 
      n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, 
      n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, 
      n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, 
      n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, 
      n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, 
      n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, 
      n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, 
      n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, 
      n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, 
      n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, 
      n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, 
      n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, 
      n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, 
      n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, 
      n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, 
      n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, 
      n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, 
      n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, 
      n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, 
      n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, 
      n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, 
      n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, 
      n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, 
      n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, 
      n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, 
      n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, 
      n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, 
      n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, 
      n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, 
      n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, 
      n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, 
      n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, 
      n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, 
      n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, 
      n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, 
      n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, 
      n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, 
      n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, 
      n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, 
      n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, 
      n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, 
      n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, 
      n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, 
      n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, 
      n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, 
      n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, 
      n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, 
      n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, 
      n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, 
      n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, 
      n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, 
      n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, 
      n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, 
      n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, 
      n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, 
      n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, 
      n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, 
      n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, 
      n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, 
      n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, 
      n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, 
      n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, 
      n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, 
      n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, 
      n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, 
      n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, 
      n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, 
      n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, 
      n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, 
      n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, 
      n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, 
      n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, 
      n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, 
      n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, 
      n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, 
      n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, 
      n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, 
      n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, 
      n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, 
      n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, 
      n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, 
      n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, 
      n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, 
      n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, 
      n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, 
      n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, 
      n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, 
      n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, 
      n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, 
      n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, 
      n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, 
      n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, 
      n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, 
      n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, 
      n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, 
      n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, 
      n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, 
      n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, 
      n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, 
      n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, 
      n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, 
      n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, 
      n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, 
      n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, 
      n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, 
      n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, 
      n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, 
      n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, 
      n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, 
      n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, 
      n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, 
      n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, 
      n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, 
      n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, 
      n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, 
      n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, 
      n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, 
      n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, 
      n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, 
      n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, 
      n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, 
      n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, 
      n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, 
      n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, 
      n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, 
      n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, 
      n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, 
      n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, 
      n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, 
      n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, 
      n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, 
      n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, 
      n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, 
      n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, 
      n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, 
      n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, 
      n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, 
      n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, 
      n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, 
      n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, 
      n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, 
      n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, 
      n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, 
      n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, 
      n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, 
      n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, 
      n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, 
      n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, 
      n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, 
      n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, 
      n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, 
      n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, 
      n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, 
      n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, 
      n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, 
      n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, 
      n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, 
      n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, 
      n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, 
      n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, 
      n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, 
      n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, 
      n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, 
      n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, 
      n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, 
      n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, 
      n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, 
      n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, 
      n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, 
      n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, 
      n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, 
      n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, 
      n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, 
      n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, 
      n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, 
      n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, 
      n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, 
      n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, 
      n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, 
      n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, 
      n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, 
      n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, 
      n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, 
      n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, 
      n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, 
      n7105, n7106, n7107, n7300, n7301, n7302, n7303, n7304, n7305, n7306, 
      n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, 
      n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, 
      n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, 
      n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, 
      n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, 
      n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, 
      n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, 
      n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, 
      n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, 
      n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, 
      n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, 
      n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, 
      n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, 
      n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, 
      n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, 
      n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, 
      n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, 
      n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, 
      n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, 
      n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, 
      n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, 
      n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, 
      n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, 
      n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, 
      n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7646, 
      n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, 
      n7657, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, 
      n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, 
      n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, 
      n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, 
      n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, 
      n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, 
      n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, 
      n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, 
      n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, 
      n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, 
      n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, 
      n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, 
      n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, 
      n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, 
      n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, 
      n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8222, n8223, 
      n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, 
      n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, 
      n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, 
      n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, 
      n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, 
      n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, 
      n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, 
      n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, 
      n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, 
      n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, 
      n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, 
      n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, 
      n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, 
      n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, 
      n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, 
      n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, 
      n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, 
      n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, 
      n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, 
      n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, 
      n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, 
      n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, 
      n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, 
      n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, 
      n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, 
      n8538, n8539, n8540, n8541, n8606, n8607, n8608, n8609, n8610, n8611, 
      n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, 
      n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, 
      n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, 
      n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, 
      n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, 
      n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, 
      n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, 
      n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, 
      n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, 
      n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, 
      n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, 
      n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, 
      n8732, n8733, n8735, n8737, n8739, n8741, n8743, n8745, n8747, n8749, 
      n8751, n8753, n8755, n8757, n8759, n8761, n8763, n8765, n8767, n8769, 
      n8771, n8773, n8775, n8777, n8779, n8781, n8783, n8785, n8787, n8789, 
      n8791, n8793, n8795, n8797, n8799, n8801, n8803, n8805, n8807, n8809, 
      n8811, n8813, n8815, n8817, n8819, n8821, n8823, n8825, n8827, n8829, 
      n8831, n8833, n8835, n8837, n8839, n8841, n8843, n8845, n8847, n8849, 
      n8851, n8853, n8855, n8857, n8859, n8861, n8862, n8863, n8864, n8865, 
      n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, 
      n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, 
      n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, 
      n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, 
      n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, 
      n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, 
      n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, 
      n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, 
      n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, 
      n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, 
      n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, 
      n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, 
      n8986, n8987, n8988, n8989, n8990, n8992, n8994, n8996, n8998, n9000, 
      n9002, n9004, n9006, n9008, n9010, n9012, n9014, n9016, n9018, n9020, 
      n9022, n9024, n9026, n9028, n9030, n9032, n9034, n9036, n9038, n9040, 
      n9042, n9044, n9046, n9048, n9050, n9052, n9054, n9056, n9058, n9060, 
      n9062, n9064, n9066, n9068, n9070, n9072, n9074, n9076, n9078, n9080, 
      n9082, n9084, n9086, n9088, n9090, n9092, n9094, n9096, n9098, n9100, 
      n9102, n9104, n9106, n9108, n9110, n9112, n9114, n9116, n9118, n9119, 
      n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, 
      n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, 
      n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, 
      n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, 
      n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, 
      n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, 
      n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, 
      n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, 
      n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, 
      n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, 
      n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, 
      n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, 
      n9240, n9241, n9242, n9243, n9244, n9245, n11783, n11784, n11785, n11786,
      n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795, 
      n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804, 
      n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813, 
      n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822, 
      n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831, 
      n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840, 
      n11841, n11842, n11843, n11844, n11845, n11846, n17221, n17224, n17227, 
      n17230, n17233, n17236, n17239, n17242, n17245, n17248, n17251, n17254, 
      n17257, n17260, n17263, n17266, n17269, n17272, n17275, n17278, n17281, 
      n17284, n17287, n17290, n17293, n17296, n17299, n17302, n17305, n17308, 
      n17311, n17314, n17317, n17320, n17323, n17326, n17329, n17332, n17335, 
      n17338, n17341, n17344, n17347, n17350, n17353, n17356, n17359, n17362, 
      n17365, n17368, n17371, n17374, n17377, n17380, n17383, n17386, n17389, 
      n17392, n17395, n17398, n17401, n17404, n17407, n17410, n17471, n17472, 
      n17474, n17475, n17477, n17478, n17480, n17481, n17483, n17484, n17486, 
      n17487, n17489, n17490, n17492, n17493, n17495, n17496, n17498, n17499, 
      n17501, n17502, n17504, n17505, n17507, n17508, n17510, n17511, n17513, 
      n17514, n17516, n17517, n17519, n17520, n17522, n17523, n17525, n17526, 
      n17528, n17529, n17531, n17532, n17534, n17535, n17537, n17538, n17540, 
      n17541, n17543, n17544, n17546, n17547, n17549, n17550, n17552, n17553, 
      n17555, n17556, n17558, n17559, n17561, n17562, n17564, n17565, n17567, 
      n17568, n17570, n17571, n17573, n17574, n17576, n17577, n17579, n17580, 
      n17582, n17583, n17585, n17586, n17588, n17589, n17591, n17592, n17594, 
      n17595, n17597, n17598, n17600, n17601, n17603, n17604, n17606, n17607, 
      n17609, n17610, n17612, n17613, n17615, n17616, n17618, n17619, n17621, 
      n17622, n17624, n17625, n17627, n17628, n17630, n17631, n17633, n17634, 
      n17636, n17637, n17639, n17640, n17642, n17643, n17645, n17646, n17648, 
      n17649, n17651, n17652, n17654, n17655, n17657, n17658, n17660, n17661, 
      n19189, n19190, n19191, n19192, n19193, n19194, n19195, n19196, n19197, 
      n19198, n19199, n19200, n19201, n19202, n19203, n19204, n19205, n19206, 
      n19207, n19208, n19209, n19210, n19211, n19212, n19213, n19214, n19215, 
      n19216, n19217, n19218, n19219, n19220, n19221, n19222, n19223, n19224, 
      n19225, n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233, 
      n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241, n19242, 
      n19243, n19244, n19245, n19246, n19247, n19248, n19249, n19250, n19251, 
      n19252, n19253, n19254, n19255, n19256, n19257, n19258, n19259, n19260, 
      n19261, n19262, n19263, n19264, n19265, n19266, n19267, n19268, n19269, 
      n19270, n19271, n19272, n19273, n19274, n19275, n19276, n19277, n19278, 
      n19279, n19280, n19281, n19282, n19283, n19284, n19285, n19286, n19287, 
      n19288, n19289, n19290, n19291, n19292, n19293, n19294, n19295, n19296, 
      n19297, n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305, 
      n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313, n19314, 
      n19315, n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19323, 
      n19324, n19325, n19326, n19327, n19328, n19329, n19330, n19331, n19332, 
      n19333, n19334, n19335, n19336, n19337, n19338, n19339, n19340, n19341, 
      n19342, n19343, n19344, n19345, n19346, n19347, n19348, n19349, n19350, 
      n19351, n19352, n19353, n19354, n19355, n19356, n19357, n19358, n19359, 
      n19360, n19361, n19362, n19363, n19364, n19365, n19366, n19367, n19368, 
      n19369, n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377, 
      n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385, n19386, 
      n19387, n19388, n19389, n19390, n19391, n19392, n19393, n19394, n19395, 
      n19396, n19397, n19398, n19399, n19460, n19461, n19462, n19463, n19464, 
      n19465, n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473, 
      n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481, n19482, 
      n19483, n19484, n19485, n19486, n19487, n19488, n19489, n19490, n19491, 
      n19492, n19493, n19494, n19495, n19496, n19497, n19498, n19499, n19500, 
      n19501, n19502, n19503, n19504, n19505, n19506, n19507, n19508, n19509, 
      n19510, n19511, n19512, n19513, n19514, n19515, n19516, n19517, n19518, 
      n19519, n19520, n19521, n19522, n19523, n19524, n19525, n19526, n19527, 
      n19528, n19529, n19530, n19531, n19532, n19533, n19534, n19535, n19536, 
      n19537, n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545, 
      n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553, n19554, 
      n19555, n19556, n19557, n19558, n19559, n19560, n19561, n19562, n19563, 
      n19564, n19565, n19566, n19567, n19568, n19569, n19570, n19571, n19572, 
      n19573, n19574, n19575, n19576, n19577, n19578, n19579, n19580, n19581, 
      n19582, n19583, n19584, n19585, n19586, n19587, n19588, n19589, n19590, 
      n19591, n19592, n19593, n19594, n19595, n19596, n19597, n19598, n19599, 
      n19600, n19601, n19602, n19603, n19604, n19605, n19606, n19607, n19608, 
      n19609, n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617, 
      n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625, n19626, 
      n19627, n19628, n19629, n19630, n19631, n19632, n19633, n19634, n19635, 
      n19636, n19637, n19638, n19639, n19640, n19641, n19642, n19643, n19644, 
      n19645, n19646, n19647, n19648, n19649, n19650, n19651, n19652, n19653, 
      n19654, n19655, n19656, n19657, n19658, n19659, n19660, n19661, n19662, 
      n19663, n19664, n19665, n19666, n19667, n19668, n19669, n19670, n19671, 
      n19672, n19673, n19674, n19675, n19676, n19677, n19678, n19679, n19680, 
      n19681, n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689, 
      n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697, n19698, 
      n19699, n19700, n19701, n19702, n19703, n19704, n19705, n19706, n19707, 
      n19708, n19709, n19710, n19711, n19712, n19713, n19714, n19715, n19716, 
      n19717, n19718, n19719, n19720, n19721, n19722, n19723, n19724, n19725, 
      n19726, n19727, n19728, n19729, n19730, n19731, n19732, n19733, n19734, 
      n19735, n19736, n19737, n19802, n19803, n19804, n19805, n19806, n19807, 
      n19808, n19809, n19810, n19811, n19812, n19813, n19814, n19815, n19816, 
      n19817, n19822, n19823, n19824, n19825, n19826, n19827, n19828, n19829, 
      n19830, n19831, n19832, n19833, n19834, n19835, n19836, n19837, n19838, 
      n19839, n19840, n19841, n19842, n19843, n19844, n19845, n19846, n19847, 
      n19848, n19849, n19850, n19851, n19852, n19853, n19854, n19855, n19856, 
      n19857, n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865, 
      n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873, n19874, 
      n19875, n19876, n19877, n19878, n19879, n19880, n19881, n19882, n19883, 
      n19884, n19885, n19886, n19887, n19888, n19889, n19890, n19891, n19892, 
      n19893, n19894, n19895, n19896, n19897, n19898, n19899, n19900, n19901, 
      n19902, n19903, n19904, n19905, n19906, n19907, n19908, n19909, n19910, 
      n19911, n19912, n19913, n19914, n19915, n19916, n19917, n19918, n19919, 
      n19920, n19921, n19922, n19923, n19924, n19925, n19926, n19927, n19928, 
      n19929, n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009, 
      n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017, n20018, 
      n20019, n20020, n20021, n20022, n20023, n20024, n20025, n20026, n20027, 
      n20028, n20029, n20030, n20031, n20032, n20033, n20034, n20035, n20036, 
      n20037, n20038, n20039, n20040, n20041, n20042, n20043, n20044, n20045, 
      n20046, n20047, n20048, n20049, n20050, n20051, n20052, n20053, n20054, 
      n20055, n20056, n20057, n20058, n20059, n20060, n20061, n20062, n20063, 
      n20064, n20065, n20066, n20067, n20068, n20069, n20070, n20071, n20072, 
      n20073, n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129, 
      n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137, n20138, 
      n20139, n20140, n20141, n20142, n20143, n20144, n20145, n20146, n20147, 
      n20148, n20149, n20150, n20151, n20152, n20153, n20154, n20155, n20156, 
      n20157, n20158, n20159, n20160, n20161, n20162, n20163, n20164, n20165, 
      n20166, n20167, n20168, n20169, n20170, n20171, n20172, n20173, n20174, 
      n20175, n20176, n20177, n20178, n20179, n20180, n20181, n20182, n20183, 
      n20184, n20185, n20186, n20187, n20188, n20189, n20190, n20191, n20192, 
      n20193, n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201, 
      n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209, n20210, 
      n20211, n20212, n20213, n20214, n20215, n20216, n20217, n20218, n20219, 
      n20220, n20221, n20222, n20223, n20224, n20225, n20226, n20227, n20228, 
      n20229, n20230, n20231, n20232, n20233, n20234, n20235, n20236, n20237, 
      n20238, n20239, n20240, n20241, n20242, n20243, n20244, n20245, n20246, 
      n20247, n20248, n20249, n20250, n20251, n20252, n20253, n20254, n20255, 
      n20256, n20257, n20258, n20259, n20260, n20261, n20262, n20263, n20264, 
      n20265, n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273, 
      n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281, n20282, 
      n20283, n20284, n20285, n20286, n20287, n20288, n20289, n20290, n20291, 
      n20292, n20293, n20294, n20295, n20296, n20297, n20298, n20299, n20300, 
      n20301, n20302, n20303, n20304, n20305, n20306, n20307, n20308, n20309, 
      n20310, n20311, n20312, n20313, n20314, n20315, n20316, n20317, n20318, 
      n20319, n20320, n20321, n20322, n20323, n20324, n20325, n20326, n20327, 
      n20328, n20329, n20330, n20331, n20332, n20333, n20334, n20335, n20336, 
      n20337, n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345, 
      n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353, n20354, 
      n20355, n20356, n20357, n20358, n20359, n20360, n20361, n20362, n20363, 
      n20364, n20365, n20366, n20367, n20368, n20369, n20370, n20371, n20372, 
      n20373, n20374, n20375, n20376, n20377, n20378, n20379, n20380, n20381, 
      n20382, n20383, n20384, n20385, n20386, n20387, n20388, n20389, n20390, 
      n20391, n20392, n20393, n20394, n20395, n20396, n20397, n20398, n20399, 
      n20400, n20401, n20402, n20403, n20404, n20405, n20406, n20407, n20408, 
      n20409, n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417, 
      n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425, n20426, 
      n20427, n20428, n20429, n20430, n20431, n20432, n20433, n20434, n20435, 
      n20436, n20437, n20438, n20439, n20440, n20441, n20442, n20443, n20444, 
      n20445, n20446, n20447, n20448, n20449, n20450, n20451, n20452, n20453, 
      n20454, n20455, n20456, n20457, n20458, n20459, n20460, n20461, n20462, 
      n20463, n20464, n20465, n20466, n20467, n20468, n20469, n20470, n20471, 
      n20472, n20473, n20474, n20475, n20476, n20477, n20478, n20479, n20480, 
      n20481, n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489, 
      n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497, n20498, 
      n20499, n20500, n20501, n20502, n20503, n20504, n20505, n20506, n20507, 
      n20508, n20509, n20510, n20511, n20512, n20513, n20514, n20515, n20516, 
      n20517, n20518, n20519, n20520, n20521, n20522, n20523, n20524, n20525, 
      n20526, n20527, n20528, n20529, n20530, n20531, n20532, n20533, n20534, 
      n20535, n20536, n20537, n20538, n20539, n20540, n20541, n20542, n20543, 
      n20544, n20545, n20546, n20547, n20548, n20549, n20550, n20551, n20552, 
      n20553, n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561, 
      n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569, n20570, 
      n20571, n20572, n20573, n20574, n20575, n20576, n20577, n20578, n20579, 
      n20580, n20581, n20582, n20583, n20584, n20585, n20586, n20587, n20588, 
      n20589, n20590, n20591, n20592, n20593, n20594, n20595, n20596, n20597, 
      n20598, n20599, n20600, n20601, n20602, n20603, n20604, n20605, n20606, 
      n20607, n20608, n20609, n20610, n20611, n20612, n20613, n20614, n20615, 
      n20616, n20617, n20618, n20619, n20620, n20621, n20622, n20623, n20624, 
      n20625, n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633, 
      n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641, n20642, 
      n20643, n20644, n20645, n20646, n20647, n20648, n20649, n20650, n20651, 
      n20652, n20653, n20654, n20655, n20656, n20657, n20658, n20659, n20660, 
      n20661, n20662, n20663, n20664, n20665, n20666, n20667, n20668, n20669, 
      n20670, n20671, n20672, n20673, n20674, n20675, n20676, n20677, n20678, 
      n20679, n20680, n20681, n20682, n20683, n20684, n20685, n20686, n20687, 
      n20688, n20689, n20690, n20691, n20692, n20693, n20694, n20695, n20696, 
      n20697, n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705, 
      n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713, n20714, 
      n20715, n20716, n20717, n20718, n20719, n20720, n20721, n20722, n20723, 
      n20724, n20725, n20726, n20727, n20728, n20729, n20730, n20731, n20732, 
      n20733, n20734, n20735, n20736, n20737, n20738, n20739, n20740, n20741, 
      n20742, n20743, n20744, n20745, n20746, n20747, n20748, n20749, n20750, 
      n20751, n20752, n20753, n20754, n20755, n20756, n20757, n20758, n20759, 
      n20760, n20761, n20762, n20763, n20764, n20765, n20766, n20767, n20768, 
      n20769, n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777, 
      n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785, n20786, 
      n20787, n20788, n20789, n20790, n20791, n20792, n20793, n20794, n20795, 
      n20796, n20797, n20798, n20799, n20800, n20801, n20802, n20803, n20804, 
      n20805, n20806, n20807, n20808, n20809, n20810, n20811, n20812, n20813, 
      n20814, n20815, n20816, n20817, n20818, n20819, n20820, n20821, n20822, 
      n20823, n20824, n20825, n20826, n20827, n20828, n20829, n20830, n20831, 
      n20832, n20833, n20834, n20835, n20836, n20837, n20838, n20839, n20840, 
      n20841, n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849, 
      n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857, n20858, 
      n20859, n20860, n20861, n20862, n20863, n20864, n20865, n20866, n20867, 
      n20868, n20869, n20870, n20871, n20872, n20873, n20874, n20875, n20876, 
      n20877, n20878, n20879, n20880, n20881, n20882, n20883, n20884, n20885, 
      n20886, n20887, n20888, n20889, n20890, n20891, n20892, n20893, n20894, 
      n20895, n20896, n20897, n20898, n20899, n20900, n20901, n20902, n20903, 
      n20904, n20905, n20906, n20907, n20908, n20909, n20910, n20911, n20912, 
      n20913, n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921, 
      n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929, n20930, 
      n20931, n20932, n20933, n20934, n20935, n20936, n20937, n20938, n20939, 
      n20940, n20941, n20942, n20943, n20944, n20945, n20946, n20947, n20948, 
      n20949, n20950, n20951, n20952, n20953, n20954, n20955, n20956, n20957, 
      n20958, n20959, n20960, n20961, n20962, n20963, n20964, n20965, n20966, 
      n20967, n20968, n20969, n20970, n20971, n20972, n20973, n20974, n20975, 
      n20976, n20977, n20978, n20979, n20980, n20981, n20982, n20983, n20984, 
      n20985, n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993, 
      n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001, n21002, 
      n21003, n21004, n21005, n21006, n21007, n21008, n21009, n21010, n21011, 
      n21012, n21013, n21014, n21015, n21016, n21017, n21018, n21019, n21020, 
      n21021, n21022, n21023, n21024, n21025, n21026, n21027, n21028, n21029, 
      n21030, n21031, n21032, n21033, n21034, n21035, n21036, n21037, n21038, 
      n21039, n21040, n21041, n21042, n21043, n21044, n21045, n21046, n21047, 
      n21048, n21049, n21050, n21051, n21052, n21053, n21054, n21055, n21056, 
      n21057, n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065, 
      n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073, n21074, 
      n21075, n21076, n21077, n21078, n21079, n21080, n21081, n21082, n21083, 
      n21084, n21085, n21086, n21087, n21088, n21089, n21090, n21091, n21092, 
      n21093, n21094, n21095, n21096, n21097, n21098, n21099, n21100, n21101, 
      n21102, n21103, n21104, n21105, n21106, n21107, n21108, n21109, n21110, 
      n21111, n21112, n21113, n21114, n21115, n21116, n21117, n21118, n21119, 
      n21120, n21121, n21122, n21123, n21124, n21125, n21126, n21127, n21128, 
      n21129, n21130, n21131, n21132, n21133, n21134, n21135, n21136, n21137, 
      n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145, n21146, 
      n21147, n21148, n21149, n21150, n21151, n21152, n21153, n21154, n21155, 
      n21156, n21157, n21158, n21159, n21160, n21161, n21162, n21163, n21164, 
      n21165, n21166, n21167, n21168, n21169, n21170, n21171, n21172, n21173, 
      n21174, n21175, n21176, n21177, n21178, n21179, n21180, n21181, n21182, 
      n21183, n21184, n21185, n21186, n21187, n21188, n21189, n21190, n21191, 
      n21192, n21193, n21194, n21195, n21196, n21197, n21198, n21199, n21200, 
      n21201, n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209, 
      n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217, n21218, 
      n21219, n21220, n21221, n21222, n21223, n21224, n21225, n21226, n21227, 
      n21228, n21229, n21230, n21231, n21232, n21233, n21234, n21235, n21236, 
      n21237, n21238, n21239, n21240, n21241, n21242, n21243, n21244, n21245, 
      n21246, n21247, n21248, n21249, n21250, n21251, n21252, n21253, n21254, 
      n21255, n21256, n21257, n21258, n21259, n21260, n21261, n21262, n21263, 
      n21264, n21265, n21266, n21267, n21268, n21269, n21270, n21271, n21272, 
      n21273, n21274, n21275, n21276, n21277, n21278, n21279, n21280, n21281, 
      n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289, n21290, 
      n21291, n21292, n21293, n21294, n21295, n21296, n21297, n21298, n21299, 
      n21300, n21301, n21302, n21303, n21304, n21305, n21306, n21307, n21308, 
      n21309, n21310, n21311, n21312, n21313, n21314, n21315, n21316, n21317, 
      n21318, n21319, n21320, n21321, n21322, n21323, n21324, n21325, n21326, 
      n21327, n21328, n21329, n21330, n21331, n21332, n21333, n21334, n21335, 
      n21336, n21337, n21338, n21339, n21340, n21341, n21342, n21343, n21344, 
      n21345, n21346, n21347, n21348, n21349, n21350, n21351, n21352, n21353, 
      n21354, n21355, n21356, n21357, n21358, n21359, n21360, n21361, n21362, 
      n21363, n21364, n21365, n21366, n21367, n21368, n21369, n21370, n21371, 
      n21372, n21373, n21374, n21375, n21376, n21377, n21378, n21379, n21380, 
      n21381, n21382, n21383, n21384, n21385, n21386, n21387, n21388, n21389, 
      n21390, n21391, n21392, n21393, n21394, n21395, n21396, n21397, n21398, 
      n21399, n21400, n21401, n21402, n21403, n21404, n21405, n21406, n21407, 
      n21408, n21409, n21410, n21411, n21412, n21413, n21414, n21415, n21416, 
      n21417, n21418, n21419, n21420, n21421, n21422, n21423, n21424, n21425, 
      n21426, n21427, n21428, n21429, n21430, n21431, n21432, n21433, n21434, 
      n21435, n21436, n21437, n21438, n21439, n21440, n21441, n21442, n21443, 
      n21444, n21445, n21446, n21447, n21448, n21449, n21450, n21451, n21452, 
      n21453, n21454, n21455, n21456, n21457, n21458, n21459, n21460, n21461, 
      n21462, n21463, n21464, n21465, n21466, n21467, n21468, n21469, n21470, 
      n21471, n21472, n21473, n21474, n21475, n21476, n21477, n21478, n21479, 
      n21480, n21481, n21482, n21483, n21484, n21485, n21486, n21487, n21488, 
      n21489, n21490, n21491, n21492, n21493, n21494, n21495, n21496, n21497, 
      n21498, n21499, n21500, n21501, n21502, n21503, n21504, n21505, n21506, 
      n21507, n21508, n21509, n21510, n21511, n21512, n21513, n21514, n21515, 
      n21516, n21517, n21518, n21519, n21520, n21521, n21522, n21523, n21524, 
      n21525, n21526, n21527, n21528, n21529, n21530, n21531, n21532, n21533, 
      n21534, n21535, n21536, n21537, n21538, n21539, n21540, n21541, n21542, 
      n21543, n21544, n21545, n21546, n21547, n21548, n21549, n21550, n21551, 
      n21552, n21553, n21554, n21555, n21556, n21557, n21558, n21559, n21560, 
      n21561, n21562, n21563, n21564, n21565, n21566, n21567, n21568, n21569, 
      n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577, n21578, 
      n21579, n21580, n21581, n21582, n21583, n21584, n21585, n21586, n21587, 
      n21588, n21589, n21590, n21591, n21592, n21593, n21594, n21595, n21596, 
      n21597, n21598, n21599, n21600, n21601, n21602, n21603, n21604, n21605, 
      n21606, n21607, n21608, n21609, n21610, n21611, n21612, n21613, n21614, 
      n21615, n21616, n21617, n21618, n21619, n21620, n21621, n21622, n21623, 
      n21624, n21625, n21626, n21627, n21628, n21629, n21630, n21631, n21632, 
      n21633, n21634, n21635, n21636, n21637, n21638, n21639, n21640, n21641, 
      n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649, n21650, 
      n21651, n21652, n21653, n21654, n21655, n21656, n21657, n21658, n21659, 
      n21660, n21661, n21662, n21663, n21664, n21665, n21666, n21667, n21668, 
      n21669, n21670, n21671, n21672, n21673, n21674, n21675, n21676, n21677, 
      n21678, n21679, n21680, n21681, n21682, n21683, n21684, n21685, n21686, 
      n21687, n21688, n21689, n21690, n21691, n21692, n21693, n21694, n21695, 
      n21696, n21697, n21698, n21699, n21700, n21701, n21702, n21703, n21704, 
      n21705, n21706, n21707, n21708, n21709, n21710, n21711, n21712, n21713, 
      n21714, n21715, n21716, n21717, n21718, n21719, n21720, n21721, n21722, 
      n21723, n21724, n21725, n21726, n21727, n21728, n21729, n21730, n21731, 
      n21732, n21733, n21734, n21735, n21736, n21737, n21738, n21739, n21740, 
      n21741, n21742, n21743, n21744, n21745, n21746, n21747, n21748, n21749, 
      n21750, n21751, n21752, n21753, n21754, n21755, n21756, n21757, n21758, 
      n21759, n21760, n21761, n21762, n21763, n21764, n21765, n21766, n21767, 
      n21768, n21769, n21770, n21771, n21772, n21773, n21774, n21775, n21776, 
      n21777, n21778, n21779, n21780, n21781, n21782, n21783, n21784, n21785, 
      n21786, n21787, n21788, n21789, n21790, n21791, n21792, n21793, n21794, 
      n21795, n21796, n21797, n21798, n21799, n21800, n21801, n21802, n21803, 
      n21804, n21805, n21806, n21807, n21808, n21809, n21810, n21811, n21812, 
      n21813, n21814, n21815, n21816, n21817, n21818, n21819, n21820, n21821, 
      n21822, n21823, n21824, n21825, n21826, n21827, n21828, n21829, n21830, 
      n21831, n21832, n21833, n21834, n21835, n21836, n21837, n21838, n21839, 
      n21840, n21841, n21842, n21843, n21844, n21845, n21846, n21847, n21848, 
      n21849, n21850, n21851, n21852, n21853, n21854, n21855, n21856, n21857, 
      n21858, n21859, n21860, n21861, n21862, n21863, n21864, n21865, n21866, 
      n21867, n21868, n21869, n21870, n21871, n21872, n21873, n21874, n21875, 
      n21876, n21877, n21878, n21879, n21880, n21881, n21882, n21883, n21884, 
      n21885, n21886, n21887, n21888, n21889, n21890, n21891, n21892, n21893, 
      n21894, n21895, n21896, n21897, n21898, n21899, n21900, n21901, n21902, 
      n21903, n21904, n21905, n21906, n21907, n21908, n21909, n21910, n21911, 
      n21912, n21913, n21914, n21915, n21916, n21917, n21918, n21919, n21920, 
      n21921, n21922, n21923, n21924, n21925, n21926, n21927, n21928, n21929, 
      n21930, n21931, n21932, n21933, n21934, n21935, n21936, n21937, n21938, 
      n21939, n21940, n21941, n21942, n21943, n21944, n21945, n21946, n21947, 
      n21948, n21949, n21950, n21951, n21952, n21953, n21954, n21955, n21956, 
      n21957, n21958, n21959, n21960, n21961, n21962, n21963, n21964, n21965, 
      n21966, n21967, n21968, n21969, n21970, n21971, n21972, n21973, n21974, 
      n21975, n21976, n21977, n21978, n21979, n21980, n21981, n21982, n21983, 
      n21984, n21985, n21986, n21987, n21988, n21989, n21990, n21991, n21992, 
      n21993, n21994, n21995, n21996, n21997, n21998, n21999, n22000, n22001, 
      n22002, n22003, n22004, n22005, n22006, n22007, n22008, n22009, n22010, 
      n22011, n22012, n22013, n22014, n22015, n22016, n22017, n22018, n22019, 
      n22020, n22021, n22022, n22023, n22024, n22025, n22026, n22027, n22028, 
      n22029, n22030, n22031, n22032, n22033, n22034, n22035, n22036, n22037, 
      n22038, n22039, n22040, n22041, n22042, n22043, n22044, n22045, n22046, 
      n22047, n22048, n22049, n22050, n22051, n22052, n22053, n22054, n22055, 
      n22056, n22057, n22058, n22059, n22060, n22061, n22062, n22063, n22064, 
      n22065, n22066, n22067, n22068, n22069, n22070, n22071, n22072, n22073, 
      n22074, n22075, n22076, n22077, n22078, n22079, n22080, n22081, n22082, 
      n22083, n22084, n22085, n22086, n22087, n22088, n22089, n22090, n22091, 
      n22092, n22093, n22094, n22095, n22096, n22097, n22098, n22099, n22100, 
      n22101, n22102, n22103, n22104, n22105, n22106, n22107, n22108, n22109, 
      n22110, n22111, n22112, n22113, n22114, n22115, n22116, n22117, n22118, 
      n22119, n22120, n22121, n22122, n22123, n22124, n22125, n22126, n22127, 
      n22128, n22129, n22130, n22131, n22132, n22133, n22134, n22135, n22136, 
      n22137, n22138, n22139, n22140, n22141, n22142, n22143, n22144, n22145, 
      n22146, n22147, n22148, n22149, n22150, n22151, n22152, n22153, n22154, 
      n22155, n22156, n22157, n22158, n22159, n22160, n22161, n22162, n22163, 
      n22164, n22165, n22166, n22167, n22168, n22169, n22170, n22171, n22172, 
      n22173, n22174, n22175, n22176, n22177, n22178, n22179, n22180, n22181, 
      n22182, n22183, n22184, n22185, n22186, n22187, n22188, n22189, n22190, 
      n22191, n22192, n22193, n22194, n22195, n22196, n22197, n22198, n22199, 
      n22200, n22201, n22202, n22203, n22204, n22205, n22206, n22207, n22208, 
      n22209, n22210, n22211, n22212, n22213, n22214, n22215, n22216, n22217, 
      n22218, n22219, n22220, n22221, n22222, n22223, n22224, n22225, n22226, 
      n22227, n22228, n22229, n22230, n22231, n22232, n22233, n22234, n22235, 
      n22236, n22237, n22238, n22239, n22240, n22241, n22242, n22243, n22244, 
      n22245, n22246, n22247, n22248, n22249, n22250, n22251, n22252, n22253, 
      n22254, n22255, n22256, n22257, n22258, n22259, n22260, n22261, n22262, 
      n22263, n22264, n22265, n22266, n22267, n22268, n22269, n22270, n22271, 
      n22272, n22273, n22274, n22275, n22276, n22277, n22278, n22279, n22280, 
      n22281, n22282, n22283, n22284, n22285, n22286, n22287, n22288, n22289, 
      n22290, n22291, n22292, n22293, n22294, n22295, n22296, n22297, n22298, 
      n22299, n22300, n22301, n22302, n22303, n22304, n22305, n22306, n22307, 
      n22308, n22309, n22310, n22311, n22312, n22313, n22314, n22315, n22316, 
      n22317, n22318, n22319, n22320, n22321, n22322, n22323, n22324, n22325, 
      n22326, n22327, n22328, n22329, n22330, n22331, n22332, n22333, n22334, 
      n22335, n22336, n22337, n22338, n22339, n22340, n22341, n22342, n22343, 
      n22344, n22345, n22346, n22347, n22348, n22349, n22350, n22351, n22352, 
      n22353, n22354, n22355, n22356, n22357, n22358, n22359, n22360, n22361, 
      n22362, n22363, n22364, n22365, n22366, n22367, n22368, n22369, n22370, 
      n22371, n22372, n22373, n22374, n22375, n22376, n22377, n22378, n22379, 
      n22380, n22381, n22382, n22383, n22384, n22385, n22386, n22387, n22388, 
      n22389, n22390, n22391, n22392, n22393, n22394, n22395, n22396, n22397, 
      n22398, n22399, n22400, n22401, n22402, n22403, n22404, n22405, n22406, 
      n22407, n22408, n22409, n22410, n22411, n22412, n22413, n22414, n22415, 
      n22416, n22417, n22418, n22419, n22420, n22421, n22422, n22423, n22424, 
      n22425, n22426, n22427, n22428, n22429, n22430, n22431, n22432, n22433, 
      n22434, n22435, n22436, n22437, n22438, n22439, n22440, n22441, n22442, 
      n22443, n22444, n22445, n22446, n22447, n22448, n22449, n22450, n22451, 
      n22452, n22453, n22454, n22455, n22456, n22457, n22458, n22459, n22460, 
      n22461, n22462, n22463, n22464, n22465, n22466, n22467, n22468, n22469, 
      n22470, n22471, n22472, n22473, n22474, n22475, n22476, n22477, n22478, 
      n22479, n22480, n22481, n22482, n22483, n22484, n22485, n22486, n22487, 
      n22488, n22489, n22490, n22491, n22492, n22493, n22494, n22495, n22496, 
      n22497, n22498, n22499, n22500, n22501, n22502, n22503, n22504, n22505, 
      n22506, n22507, n22508, n22509, n22510, n22511, n22512, n22513, n22514, 
      n22515, n22516, n22517, n22518, n22519, n22520, n22521, n22522, n22523, 
      n22524, n22525, n22526, n22527, n22528, n22529, n22530, n22531, n22532, 
      n22533, n22534, n22535, n22536, n22537, n22538, n22539, n22540, n22541, 
      n22542, n22543, n22544, n22545, n22546, n22547, n22548, n22549, n22550, 
      n22551, n22552, n22553, n22554, n22555, n22556, n22557, n22558, n22559, 
      n22560, n22561, n22562, n22563, n22564, n22565, n22566, n22567, n22568, 
      n22569, n22570, n22571, n22572, n22573, n22574, n22575, n22576, n22577, 
      n22578, n22579, n22580, n22581, n22582, n22583, n22584, n22585, n22586, 
      n22587, n22588, n22589, n22590, n22591, n22592, n22593, n22594, n22595, 
      n22596, n22597, n22598, n22599, n22600, n22601, n22602, n22603, n22604, 
      n22605, n22606, n22607, n22608, n22609, n22610, n22611, n22612, n22613, 
      n22614, n22615, n22616, n22617, n22618, n22619, n22620, n22621, n22622, 
      n22623, n22624, n22625, n22626, n22627, n22628, n22629, n22630, n22631, 
      n22632, n22633, n22634, n22635, n22636, n22637, n22638, n22639, n22640, 
      n22641, n22642, n22643, n22644, n22645, n22646, n22647, n22648, n22649, 
      n22650, n22651, n22652, n22653, n22654, n22655, n22656, n22657, n22658, 
      n22659, n22660, n22661, n22662, n22663, n22664, n22665, n22666, n22667, 
      n22668, n22669, n22670, n22671, n22672, n22673, n22674, n22675, n22676, 
      n22677, n22678, n22679, n22680, n22681, n22682, n22683, n22684, n22685, 
      n22686, n22687, n22688, n22689, n22690, n22691, n22692, n22693, n22694, 
      n22695, n22696, n22697, n22698, n22699, n22700, n22701, n22702, n22703, 
      n22704, n22705, n22706, n22707, n22708, n22709, n22710, n22711, n22712, 
      n22713, n22714, n22715, n22716, n22717, n22718, n22719, n22720, n22721, 
      n22722, n22723, n22724, n22725, n22726, n22727, n22728, n22729, n22730, 
      n22731, n22732, n22733, n22734, n22735, n22736, n22737, n22738, n22739, 
      n22740, n22741, n22742, n22743, n22744, n22745, n22746, n22747, n22748, 
      n22749, n22750, n22751, n22752, n22753, n22754, n22755, n22756, n22757, 
      n22758, n22759, n22760, n22761, n22762, n22763, n22764, n22765, n22766, 
      n22767, n22768, n22769, n22770, n22771, n22772, n22773, n22774, n22775, 
      n22776, n22777, n22778, n22779, n22780, n22781, n22782, n22783, n22784, 
      n22785, n22786, n22787, n22788, n22789, n22790, n22791, n22792, n22793, 
      n22794, n22795, n22796, n22797, n22798, n22799, n22800, n22801, n22802, 
      n22803, n22804, n22805, n22806, n22807, n22808, n22809, n22810, n22811, 
      n22812, n22813, n22814, n22815, n22816, n22817, n22818, n22819, n22820, 
      n22821, n22822, n22823, n22824, n22825, n22826, n22827, n22828, n22829, 
      n22830, n22831, n22832, n22833, n22834, n22835, n22836, n22837, n22838, 
      n22839, n22840, n22841, n22842, n22843, n22844, n22845, n22846, n22847, 
      n22848, n22849, n22850, n22851, n22852, n22853, n22854, n22855, n22856, 
      n22857, n22858, n22859, n22860, n22861, n22862, n22863, n22864, n22865, 
      n22866, n22867, n22868, n22869, n22870, n22871, n22872, n22873, n22874, 
      n22875, n22876, n22877, n22878, n22879, n22880, n22881, n22882, n22883, 
      n22884, n22885, n22886, n22887, n22888, n22889, n22890, n22891, n22892, 
      n22893, n22894, n22895, n22896, n22897, n22898, n22899, n22900, n22901, 
      n22902, n22903, n22904, n22905, n22906, n22907, n22908, n22909, n22910, 
      n22911, n22912, n22913, n22914, n22915, n22916, n22917, n22918, n22919, 
      n22920, n22921, n22922, n22923, n22924, n22925, n22926, n22927, n22928, 
      n22929, n22930, n22931, n22932, n22933, n22934, n22935, n22936, n22937, 
      n22938, n22939, n22940, n22941, n22942, n22943, n22944, n22945, n22946, 
      n22947, n22948, n22949, n22950, n22951, n22952, n22953, n22954, n22955, 
      n22956, n22957, n22958, n22959, n22960, n22961, n22962, n22963, n22964, 
      n22965, n22966, n22967, n22968, n22969, n22970, n22971, n22972, n22973, 
      n22974, n22975, n22976, n22977, n22978, n22979, n22980, n22981, n22982, 
      n22983, n22984, n22985, n22986, n22987, n22988, n22989, n22990, n22991, 
      n22992, n22993, n22994, n22995, n22996, n22997, n22998, n22999, n23000, 
      n23001, n23002, n23003, n23004, n23005, n23006, n23007, n23008, n23009, 
      n23010, n23011, n23012, n23013, n23014, n23015, n23016, n23017, n23018, 
      n23019, n23020, n23021, n23022, n23023, n23024, n23025, n23026, n23027, 
      n23028, n23029, n23030, n23031, n23032, n23033, n23034, n23035, n23036, 
      n23037, n23038, n23039, n23040, n23041, n23042, n23043, n23044, n23045, 
      n23046, n23047, n23048, n23049, n23050, n23051, n23052, n23053, n23054, 
      n23055, n23056, n23057, n23058, n23059, n23060, n23061, n23062, n23063, 
      n23064, n23065, n23066, n23067, n23068, n23069, n23070, n23071, n23072, 
      n23073, n23074, n23075, n23076, n23077, n23078, n23079, n23080, n23081, 
      n23082, n23083, n23084, n23085, n23086, n23087, n23088, n23089, n23090, 
      n23091, n23092, n23093, n23094, n23095, n23096, n23097, n23098, n23099, 
      n23100, n23101, n23102, n23103, n23104, n23105, n23106, n23107, n23108, 
      n23109, n23110, n23111, n23112, n23113, n23114, n23115, n23116, n23117, 
      n23118, n23119, n23120, n23121, n23122, n23123, n23124, n23125, n23126, 
      n23127, n23128, n23129, n23130, n23131, n23132, n23133, n23134, n23135, 
      n23136, n23137, n23138, n23139, n23140, n23141, n23142, n23143, n23144, 
      n23145, n23146, n23147, n23148, n23149, n23150, n23151, n23152, n23153, 
      n23154, n23155, n23156, n23157, n23158, n23159, n23160, n23161, n23162, 
      n23163, n23164, n23165, n23166, n23167, n23168, n23169, n23170, n23171, 
      n23172, n23173, n23174, n23175, n23176, n23177, n23178, n23179, n23180, 
      n23181, n23182, n23183, n23184, n23185, n23186, n23187, n23188, n23189, 
      n23190, n23191, n23192, n23193, n23194, n23195, n23196, n23197, n23198, 
      n23199, n23200, n23201, n23202, n23203, n23204, n23205, n23206, n23207, 
      n23208, n23209, n23210, n23211, n23212, n23213, n23214, n23215, n23216, 
      n23217, n23218, n23219, n23220, n23221, n23222, n23223, n23224, n23225, 
      n23226, n23227, n23228, n23229, n23230, n23231, n23232, n23233, n23234, 
      n23235, n23236, n23237, n23238, n23239, n23240, n23241, n23242, n23243, 
      n23244, n23245, n23246, n23247, n23248, n23249, n23250, n23251, n23252, 
      n23253, n23254, n23255, n23256, n23257, n23258, n23259, n23260, n23261, 
      n23262, n23263, n23264, n23265, n23266, n23267, n23268, n23269, n23270, 
      n23271, n23272, n23273, n23274, n23275, n23276, n23277, n23278, n23279, 
      n23280, n23281, n23282, n23283, n23284, n23285, n23286, n23287, n23288, 
      n23289, n23290, n23291, n23292, n23293, n23294, n23295, n23296, n23297, 
      n23298, n23299, n23300, n23301, n23302, n23303, n23304, n23305, n23306, 
      n23307, n23308, n23309, n23310, n23311, n23312, n23313, n23314, n23315, 
      n23316, n23317, n23318, n23319, n23320, n23321, n23322, n23323, n23324, 
      n23325, n23326, n23327, n23328, n23329, n23330, n23331, n23332, n23333, 
      n23334, n23335, n23336, n23337, n23338, n23339, n23340, n23341, n23342, 
      n23343, n23344, n23345, n23346, n23347, n23348, n23349, n23350, n23351, 
      n23352, n23353, n23354, n23355, n23356, n23357, n23358, n23359, n23360, 
      n23361, n23362, n23363, n23364, n23365, n23366, n23367, n23368, n23369, 
      n23370, n23371, n23372, n23373, n23374, n23375, n23376, n23377, n23378, 
      n23379, n23380, n23381, n23382, n23383, n23384, n23385, n23386, n23387, 
      n23388, n23389, n23390, n23391, n23392, n23393, n23394, n23395, n23396, 
      n23397, n23398, n23399, n23400, n23401, n23402, n23403, n23404, n23405, 
      n23406, n23407, n23408, n23409, n23410, n23411, n23412, n23413, n23414, 
      n23415, n23416, n23417, n23418, n23419, n23420, n23421, n23422, n23423, 
      n23424, n23425, n23426, n23427, n23428, n23429, n23430, n23431, n23432, 
      n23433, n23434, n23435, n23436, n23437, n23438, n23439, n23440, n23441, 
      n23442, n23443, n23444, n23445, n23446, n23447, n23448, n23449, n23450, 
      n23451, n23452, n23453, n23454, n23455, n23456, n23457, n23458, n23459, 
      n23460, n23461, n23462, n23463, n23464, n23465, n23466, n23467, n23468, 
      n23469, n23470, n23471, n23472, n23473, n23474, n23475, n23476, n23477, 
      n23478, n23479, n23480, n23481, n23482, n23483, n23484, n23485, n23486, 
      n23487, n23488, n23489, n23490, n23491, n23492, n23493, n23494, n23495, 
      n23496, n23497, n23498, n23499, n23500, n23501, n23502, n23503, n23504, 
      n23505, n23506, n23507, n23508, n23509, n23510, n23511, n23512, n23513, 
      n23514, n23515, n23516, n23517, n23518, n23519, n23520, n23521, n23522, 
      n23523, n23524, n23525, n23526, n23527, n23528, n23529, n23530, n23531, 
      n23532, n23533, n23534, n23535, n23536, n23537, n23538, n23539, n23540, 
      n23541, n23542, n23543, n23544, n23545, n23546, n23547, n23548, n23549, 
      n23550, n23551, n23552, n23553, n23554, n23555, n23556, n23557, n23558, 
      n23559, n23560, n23561, n23562, n23563, n23564, n23565, n23566, n23567, 
      n23568, n23569, n23570, n23571, n23572, n23573, n23574, n23575, n23576, 
      n23577, n23578, n23579, n23580, n23581, n23582, n23583, n23584, n23585, 
      n23586, n23587, n23588, n23589, n23590, n23591, n23592, n23593, n23594, 
      n23595, n23596, n23597, n23598, n23599, n23600, n23601, n23602, n23603, 
      n23604, n23605, n23606, n23607, n23608, n23609, n23610, n23611, n23612, 
      n23613, n23614, n23615, n23616, n23617, n23618, n23619, n23620, n23621, 
      n23622, n23623, n23624, n23625, n23626, n23627, n23628, n23629, n23630, 
      n23631, n23632, n23633, n23634, n23635, n23636, n23637, n23638, n23639, 
      n23640, n23641, n23642, n23643, n23644, n23645, n23646, n23647, n23648, 
      n23649, n23650, n23651, n23652, n23653, n23654, n23655, n23656, n23657, 
      n23658, n23659, n23660, n23661, n23662, n23663, n23664, n23665, n23666, 
      n23667, n23668, n23669, n23670, n23671, n23672, n23673, n23674, n23675, 
      n23676, n23677, n23678, n23679, n23680, n23681, n23682, n23683, n23684, 
      n23685, n23686, n23687, n23688, n23689, n23690, n23691, n23692, n23693, 
      n23694, n23695, n23696, n23697, n23698, n23699, n23700, n23701, n23702, 
      n23703, n23704, n23705, n23706, n23707, n23708, n23709, n23710, n23711, 
      n23712, n23713, n23714, n23715, n23716, n23717, n23718, n23719, n23720, 
      n23721, n23722, n23723, n23724, n23725, n23726, n23727, n23728, n23729, 
      n23730, n23731, n23732, n23733, n23734, n23735, n23736, n23737, n23738, 
      n23739, n23740, n23741, n23742, n23743, n23744, n23745, n23746, n23747, 
      n23748, n23749, n23750, n23751, n23752, n23753, n23754, n23755, n23756, 
      n23757, n23758, n23759, n23760, n23761, n23762, n23763, n23856, n23858, 
      n23860, n23862, n23864, n23866, n23868, n23870, n23872, n23874, n23876, 
      n23878, n23880, n23882, n23884, n23886, n23888, n23890, n23892, n23894, 
      n23896, n23898, n23900, n23902, n23904, n23906, n23908, n23910, n23912, 
      n23914, n23916, n23918, n23920, n23922, n23924, n23926, n23928, n23930, 
      n23932, n23934, n23936, n23938, n23940, n23942, n23944, n23946, n23948, 
      n23950, n23952, n23953, n23954, n23955, n23956, n23957, n23958, n23959, 
      n23960, n23961, n23962, n23963, n23964, n23965, n23966, n23967, n23968, 
      n23969, n23970, n23971, n23972, n23973, n23974, n23975, n23976, n23977, 
      n23978, n23979, n23980, n23981, n23982, n23983, n23984, n23985, n23986, 
      n23987, n23988, n23989, n23990, n23991, n23992, n23993, n23994, n23995, 
      n23996, n23997, n23998, n23999, n24000, n24001, n24002, n24003, n24004, 
      n24005, n24006, n24007, n24008, n24009, n24010, n24011, n24012, n24013, 
      n24014, n24015, n24016, n24017, n24018, n24019, n24020, n24021, n24022, 
      n24023, n24024, n24025, n24026, n24027, n24028, n24029, n24030, n24031, 
      n24148, n24149, n24150, n24151, n24152, n24153, n24154, n24155, n24156, 
      n24157, n24158, n24159, n24160, n24161, n24162, n24163, n24164, n24165, 
      n24166, n24167, n24168, n24169, n24170, n24171, n24172, n24173, n24174, 
      n24175, n24176, n24177, n24178, n24179, n24180, n24181, n24182, n24183, 
      n24184, n24185, n24186, n24187, n24188, n24189, n24190, n24191, n24192, 
      n24193, n24194, n24195, n24196, n24197, n24198, n24199, n24200, n24201, 
      n24202, n24203, n24204, n24205, n24206, n24207, n24208, n24209, n24210, 
      n24211, n24212, n24213, n24214, n24215, n24216, n24217, n24218, n24219, 
      n24220, n24221, n24222, n24223, n24224, n24225, n24226, n24227, n24228, 
      n24229, n24230, n24231, n24232, n24233, n24234, n24235, n24236, n24237, 
      n24238, n24239, n24240, n24241, n24242, n24243, n24244, n24245, n24246, 
      n24247, n24248, n24249, n24250, n24251, n24252, n24253, n24254, n24255, 
      n24256, n24257, n24258, n24259, n24260, n24261, n24262, n24263, n24264, 
      n24265, n24266, n24267, n24268, n24269, n24270, n24271, n24272, n24273, 
      n24274, n24275, n24276, n24277, n24278, n24279, n24280, n24281, n24282, 
      n24283, n24284, n24285, n24286, n24287, n24288, n24289, n24290, n24291, 
      n24292, n24293, n24294, n24295, n24296, n24297, n24298, n24299, n24300, 
      n24301, n24302, n24303, n24304, n24305, n24306, n24307, n24308, n24309, 
      n24310, n24311, n24312, n24313, n24314, n24315, n24316, n24317, n24318, 
      n24319, n24320, n24321, n24322, n24323, n24324, n24325, n24326, n24327, 
      n24328, n24329, n24330, n24331, n24332, n24333, n24334, n24335, n24336, 
      n24337, n24338, n24339, n24340, n24341, n24342, n24343, n24344, n24345, 
      n24346, n24347, n24348, n24349, n24350, n24351, n24352, n24353, n24354, 
      n24355, n24356, n24357, n24358, n24359, n24360, n24361, n24362, n24363, 
      n24364, n24365, n24366, n24367, n24368, n24369, n24370, n24371, n24372, 
      n24373, n24374, n24375, n24376, n24377, n24378, n24379, n24380, n24381, 
      n24382, n24383, n24384, n24385, n24386, n24387, n24388, n24389, n24390, 
      n24391, n24392, n24393, n24394, n24395, n24396, n24397, n24398, n24399, 
      n24400, n24401, n24402, n24403, n24404, n24405, n24406, n24407, n24408, 
      n24409, n24410, n24411, n24412, n24413, n24414, n24415, n24416, n24417, 
      n24418, n24419, n24420, n24421, n24422, n24423, n24424, n24425, n24426, 
      n24427, n24428, n24429, n24430, n24431, n24432, n24433, n24434, n24435, 
      n24436, n24437, n24438, n24439, n24440, n24441, n24442, n24443, n24444, 
      n24445, n24446, n24447, n24448, n24449, n24450, n24451, n24452, n24453, 
      n24454, n24455, n24456, n24457, n24458, n24459, n24460, n24461, n24462, 
      n24463, n24464, n24465, n24466, n24467, n24468, n24469, n24470, n24471, 
      n24472, n24473, n24474, n24475, n24476, n24477, n24478, n24479, n24480, 
      n24481, n24482, n24483, n24484, n24485, n24486, n24487, n24488, n24489, 
      n24490, n24491, n24492, n24493, n24494, n24495, n24496, n24497, n24498, 
      n24499, n24500, n24501, n24502, n24503, n24504, n24505, n24506, n24507, 
      n24508, n24509, n24510, n24511, n24512, n24513, n24514, n24515, n24516, 
      n24517, n24518, n24519, n24520, n24521, n24522, n24523, n24524, n24525, 
      n24526, n24527, n24528, n24529, n24530, n24531, n24532, n24533, n24534, 
      n24535, n24536, n24537, n24538, n24539, n24540, n24541, n24542, n24543, 
      n24544, n24545, n24546, n24547, n24548, n24549, n24550, n24551, n24552, 
      n24553, n24554, n24555, n24556, n24557, n24558, n24559, n24560, n24561, 
      n24562, n24563, n24564, n24565, n24566, n24567, n24568, n24569, n24570, 
      n24571, n24572, n24573, n24574, n24575, n24576, n24577, n24578, n24579, 
      n24580, n24581, n24582, n24583, n24584, n24585, n24586, n24587, n24588, 
      n24589, n24590, n24591, n24592, n24593, n24594, n24595, n24596, n24597, 
      n24598, n24599, n24600, n24601, n24602, n24603, n24604, n24605, n24606, 
      n24607, n24608, n24609, n24610, n24611, n24612, n24613, n24614, n24615, 
      n24616, n24617, n24618, n24619, n24620, n24621, n24622, n24623, n24624, 
      n24625, n24626, n24627, n24628, n24629, n24630, n24631, n24632, n24633, 
      n24634, n24635, n24636, n24637, n24638, n24639, n24640, n24641, n24642, 
      n24643, n24644, n24645, n24646, n24647, n24648, n24649, n24650, n24651, 
      n24652, n24653, n24654, n24655, n24656, n24657, n24658, n24659, n24660, 
      n24661, n24662, n24663, n24664, n24665, n24666, n24667, n24668, n24669, 
      n24670, n24671, n24672, n24673, n24674, n24675, n24676, n24677, n24678, 
      n24679, n24680, n24681, n24682, n24683, n24684, n24685, n24686, n24687, 
      n24688, n24689, n24690, n24691, n24692, n24693, n24694, n24695, n24696, 
      n24697, n24698, n24699, n24700, n24701, n24702, n24703, n24704, n24705, 
      n24706, n24707, n24708, n24709, n24710, n24711, n24712, n24713, n24714, 
      n24715, n24716, n24717, n24718, n24719, n24720, n24721, n24722, n24723, 
      n24724, n24725, n24726, n24727, n24728, n24729, n24730, n24731, n24732, 
      n24733, n24734, n24735, n24736, n24737, n24738, n24739, n24740, n24741, 
      n24742, n24743, n24744, n24745, n24746, n24747, n24748, n24749, n24750, 
      n24751, n24752, n24753, n24754, n24755, n24756, n24757, n24758, n24759, 
      n24760, n24761, n24762, n24763, n24764, n24765, n24766, n24767, n24768, 
      n24769, n24770, n24771, n24772, n24773, n24774, n24775, n24776, n24777, 
      n24778, n24779, n24780, n24781, n24782, n24783, n24784, n24785, n24786, 
      n24787, n24788, n24789, n24790, n24791, n24792, n24793, n24794, n24795, 
      n24796, n24797, n24798, n24799, n24800, n24801, n24802, n24803, n24804, 
      n24805, n24806, n24807, n24808, n24809, n24810, n24811, n24812, n24813, 
      n24814, n24815, n24816, n24817, n24818, n24819, n24820, n24821, n24822, 
      n24823, n24824, n24825, n24826, n24827, n24828, n24829, n24830, n24831, 
      n24832, n24833, n24834, n24835, n24836, n24837, n24838, n24839, n24840, 
      n24841, n24842, n24843, n24844, n24845, n24846, n24847, n24848, n24849, 
      n24850, n24851, n24852, n24853, n24854, n24855, n24856, n24857, n24858, 
      n24859, n24860, n24861, n24862, n24863, n24864, n24865, n24866, n24867, 
      n24868, n24869, n24870, n24871, n24872, n24873, n24874, n24875, n24876, 
      n24877, n24878, n24879, n24880, n24881, n24882, n24883, n24884, n24885, 
      n24886, n24887, n24888, n24889, n24890, n24891, n24892, n24893, n24894, 
      n24895, n24896, n24897, n24898, n24899, n24900, n24901, n24902, n24903, 
      n24904, n24905, n24906, n24907, n24908, n24909, n24910, n24911, n24912, 
      n24913, n24914, n24915, n24916, n24917, n24918, n24919, n24920, n24921, 
      n24922, n24923, n24924, n24925, n24926, n24927, n24928, n24929, n24930, 
      n24931, n24932, n24933, n24934, n24935, n24936, n24937, n24938, n24939, 
      n24940, n24941, n24942, n24943, n24944, n24945, n24946, n24947, n24948, 
      n24949, n24950, n24951, n24952, n24953, n24954, n24955, n24956, n24957, 
      n24958, n24959, n24960, n24961, n24962, n24963, n24964, n24965, n24966, 
      n24967, n24968, n24969, n24970, n24971, n24972, n24973, n24974, n24975, 
      n24976, n24977, n24978, n24979, n24980, n24981, n24982, n24983, n24984, 
      n24985, n24986, n24987, n24988, n24989, n24990, n24991, n24992, n24993, 
      n24994, n24995, n24996, n24997, n24998, n24999, n25000, n25001, n25002, 
      n25003, n25004, n25005, n25006, n25007, n25008, n25009, n25010, n25011, 
      n25012, n25013, n25014, n25015, n25016, n25017, n25018, n25019, n25020, 
      n25021, n25022, n25023, n25024, n25025, n25026, n25027, n25028, n25029, 
      n25030, n25031, n25032, n25033, n25034, n25035, n25036, n25037, n25038, 
      n25039, n25040, n25041, n25042, n25043, n25044, n25045, n25046, n25047, 
      n25048, n25049, n25050, n25051, n25052, n25053, n25054, n25055, n25056, 
      n25057, n25058, n25059, n25060, n25061, n25062, n25063, n25064, n25065, 
      n25066, n25067, n25068, n25069, n25070, n25071, n25072, n25073, n25074, 
      n25075, n25076, n25077, n25078, n25079, n25080, n25081, n25082, n25083, 
      n25084, n25085, n25086, n25087, n25088, n25089, n25090, n25091, n25092, 
      n25093, n25094, n25095, n25096, n25097, n25098, n25099, n25100, n25101, 
      n25102, n25103, n25104, n25105, n25106, n25107, n25108, n25109, n25110, 
      n25111, n25112, n25113, n25114, n25115, n25116, n25117, n25118, n25119, 
      n25120, n25121, n25122, n25123, n25124, n25125, n25126, n25127, n25128, 
      n25129, n25130, n25131, n25132, n25133, n25134, n25135, n25136, n25137, 
      n25138, n25139, n25140, n25141, n25142, n25143, n25144, n25145, n25146, 
      n25147, n25148, n25149, n25150, n25151, n25152, n25153, n25154, n25155, 
      n25156, n25157, n25158, n25159, n25160, n25161, n25162, n25163, n25164, 
      n25165, n25166, n25167, n25168, n25169, n25170, n25171, n25172, n25173, 
      n25174, n25175, n25176, n25177, n25178, n25179, n25180, n25181, n25182, 
      n25183, n25184, n25185, n25186, n25187, n25188, n25189, n25190, n25191, 
      n25192, n25193, n25194, n25195, n25196, n25197, n25198, n25199, n25200, 
      n25201, n25202, n25203, n25204, n25205, n25206, n25207, n25208, n25209, 
      n25210, n25211, n25212, n25213, n25214, n25215, n25216, n25217, n25218, 
      n25219, n25220, n25221, n25222, n25223, n25224, n25225, n25226, n25227, 
      n25228, n25229, n25230, n25231, n25232, n25233, n25234, n25235, n25236, 
      n25237, n25238, n25239, n25240, n25241, n25242, n25243, n25244, n25245, 
      n25246, n25247, n25248, n25249, n25250, n25251, n25252, n25253, n25254, 
      n25255, n25256, n25257, n25258, n25259, n25260, n25261, n25262, n25263, 
      n25264, n25265, n25266, n25267, n25268, n25269, n25270, n25271, n25272, 
      n25273, n25274, n25275, n25276, n25277, n25278, n25279, n25280, n25281, 
      n25282, n25283, n25284, n25285, n25286, n25287, n25288, n25289, n25290, 
      n25291, n25292, n25293, n25294, n25295, n25296, n25297, n25298, n25299, 
      n25300, n25301, n25302, n25303, n25304, n25305, n25306, n25307, n25308, 
      n25309, n25310, n25311, n25312, n25313, n25314, n25315, n25316, n25317, 
      n25318, n25319, n25320, n25321, n25322, n25323, n25324, n25325, n25326, 
      n25327, n25328, n25329, n25330, n25331, n25332, n25333, n25334, n25335, 
      n25336, n25337, n25338, n25339, n25340, n25341, n25342, n25343, n25344, 
      n25345, n25346, n25347, n25348, n25349, n25350, n25351, n25352, n25353, 
      n25354, n25355, n25356, n25357, n25358, n25359, n25360, n25361, n25362, 
      n25363, n25364, n25365, n25366, n25367, n25368, n25369, n25370, n25371, 
      n25372, n25373, n25374, n25375, n25376, n25377, n25378, n25379, n25380, 
      n25381, n25382, n25383, n25384, n25385, n25386, n25387, n25388, n25389, 
      n25390, n25391, n25392, n25393, n25394, n25395, n25396, n25397, n25398, 
      n25399, n25400, n25401, n25402, n25403, n25404, n25405, n25406, n25407, 
      n25408, n25409, n25410, n25411, n25412, n25413, n25414, n25415, n25416, 
      n25417, n25418, n25419, n25420, n25421, n25422, n25423, n25424, n25425, 
      n25426, n25427, n25428, n25429, n25430, n25431, n25432, n25433, n25434, 
      n25435, n25436, n25437, n25438, n25439, n25440, n25441, n25442, n25443, 
      n25444, n25445, n25446, n25447, n25448, n25449, n25450, n25451, n25452, 
      n25453, n25454, n25455, n25456, n25457, n25458, n25459, n25460, n25461, 
      n25462, n25463, n25464, n25465, n25466, n25467, n25468, n25469, n25470, 
      n25471, n25472, n25473, n25474, n25475, n25476, n25477, n25478, n25479, 
      n25480, n25481, n25482, n25483, n25484, n25485, n25486, n25487, n25488, 
      n25489, n25490, n25491, n25492, n25493, n25494, n25495, n25496, n25497, 
      n25498, n25499, n25500, n25501, n25502, n25503, n25504, n25505, n25506, 
      n25507, n25508, n25509, n25510, n25511, n25512, n25513, n25514, n25515, 
      n25516, n25517, n25518, n25519, n25520, n25521, n25522, n25523, n25524, 
      n25525, n25526, n25527, n25528, n25529, n25530, n25531, n25532, n25533, 
      n25534, n25535, n25536, n25537, n25538, n25539, n25540, n25541, n25542, 
      n25543, n25544, n25545, n25546, n25547, n25548, n25549, n25550, n25551, 
      n25552, n25553, n25554, n25555, n25556, n25557, n25558, n25559, n25560, 
      n25561, n25562, n25563, n25564, n_1000, n_1001, n_1002, n_1003, n_1004, 
      n_1005, n_1006, n_1007, n_1008, n_1009, n_1010, n_1011, n_1012, n_1013, 
      n_1014, n_1015, n_1016, n_1017, n_1018, n_1019, n_1020, n_1021, n_1022, 
      n_1023, n_1024, n_1025, n_1026, n_1027, n_1028, n_1029, n_1030, n_1031, 
      n_1032, n_1033, n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, 
      n_1041, n_1042, n_1043, n_1044, n_1045, n_1046, n_1047, n_1048, n_1049, 
      n_1050, n_1051, n_1052, n_1053, n_1054, n_1055, n_1056, n_1057, n_1058, 
      n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, 
      n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, n_1076, 
      n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, n_1085, 
      n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, n_1092, n_1093, n_1094, 
      n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, n_1103, 
      n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, 
      n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, 
      n_1122, n_1123, n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, n_1130, 
      n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, n_1137, n_1138, n_1139, 
      n_1140, n_1141, n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, n_1148, 
      n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, n_1155, n_1156, n_1157, 
      n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, 
      n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, n_1175, 
      n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, n_1182, n_1183, n_1184, 
      n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, 
      n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, 
      n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, 
      n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, 
      n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, 
      n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, 
      n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, 
      n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, n_1256, 
      n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, 
      n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, 
      n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, 
      n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, 
      n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, 
      n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, 
      n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, n_1317, n_1318, n_1319, 
      n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, n_1326, n_1327, n_1328, 
      n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, n_1335, n_1336, n_1337, 
      n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, 
      n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, n_1353, n_1354, n_1355, 
      n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, n_1364, 
      n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, n_1373, 
      n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, n_1380, n_1381, n_1382, 
      n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, n_1389, n_1390, n_1391, 
      n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, n_1400, 
      n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, n_1407, n_1408, n_1409, 
      n_1410, n_1411, n_1412, n_1413, n_1414, n_1415, n_1416, n_1417, n_1418, 
      n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, 
      n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, 
      n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, n_1445, 
      n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, n_1452, n_1453, n_1454, 
      n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, n_1461, n_1462, n_1463, 
      n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, n_1470, n_1471, n_1472, 
      n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, n_1479, n_1480, n_1481, 
      n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, n_1488, n_1489, n_1490, 
      n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, n_1497, n_1498, n_1499, 
      n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, n_1506, n_1507, n_1508, 
      n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, n_1515, n_1516, n_1517, 
      n_1518, n_1519, n_1520, n_1521, n_1522, n_1523, n_1524, n_1525, n_1526, 
      n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, n_1533, n_1534, n_1535, 
      n_1536, n_1537, n_1538, n_1539, n_1540, n_1541, n_1542, n_1543, n_1544, 
      n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, n_1551, n_1552, n_1553, 
      n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, n_1560, n_1561, n_1562, 
      n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, n_1569, n_1570, n_1571, 
      n_1572, n_1573, n_1574, n_1575, n_1576, n_1577, n_1578, n_1579, n_1580, 
      n_1581, n_1582, n_1583, n_1584, n_1585, n_1586, n_1587, n_1588, n_1589, 
      n_1590, n_1591, n_1592, n_1593, n_1594, n_1595, n_1596, n_1597, n_1598, 
      n_1599, n_1600, n_1601, n_1602, n_1603, n_1604, n_1605, n_1606, n_1607, 
      n_1608, n_1609, n_1610, n_1611, n_1612, n_1613, n_1614, n_1615, n_1616, 
      n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, n_1623, n_1624, n_1625, 
      n_1626, n_1627, n_1628, n_1629, n_1630, n_1631, n_1632, n_1633, n_1634, 
      n_1635, n_1636, n_1637, n_1638, n_1639 : std_logic;

begin
   OUT2 <= ( OUT2_63_port, OUT2_62_port, OUT2_61_port, OUT2_60_port, 
      OUT2_59_port, OUT2_58_port, OUT2_57_port, OUT2_56_port, OUT2_55_port, 
      OUT2_54_port, OUT2_53_port, OUT2_52_port, OUT2_51_port, OUT2_50_port, 
      OUT2_49_port, OUT2_48_port, OUT2_47_port, OUT2_46_port, OUT2_45_port, 
      OUT2_44_port, OUT2_43_port, OUT2_42_port, OUT2_41_port, OUT2_40_port, 
      OUT2_39_port, OUT2_38_port, OUT2_37_port, OUT2_36_port, OUT2_35_port, 
      OUT2_34_port, OUT2_33_port, OUT2_32_port, OUT2_31_port, OUT2_30_port, 
      OUT2_29_port, OUT2_28_port, OUT2_27_port, OUT2_26_port, OUT2_25_port, 
      OUT2_24_port, OUT2_23_port, OUT2_22_port, OUT2_21_port, OUT2_20_port, 
      OUT2_19_port, OUT2_18_port, OUT2_17_port, OUT2_16_port, OUT2_15_port, 
      OUT2_14_port, OUT2_13_port, OUT2_12_port, OUT2_11_port, OUT2_10_port, 
      OUT2_9_port, OUT2_8_port, OUT2_7_port, OUT2_6_port, OUT2_5_port, 
      OUT2_4_port, OUT2_3_port, OUT2_2_port, OUT2_1_port, OUT2_0_port );
   
   REGISTERS_reg_11_63_inst : DFF_X1 port map( D => n6403, CK => CLK, Q => 
                           n19396, QN => n9118);
   REGISTERS_reg_11_62_inst : DFF_X1 port map( D => n6402, CK => CLK, Q => 
                           n19397, QN => n9120);
   REGISTERS_reg_11_61_inst : DFF_X1 port map( D => n6401, CK => CLK, Q => 
                           n19398, QN => n9122);
   REGISTERS_reg_11_60_inst : DFF_X1 port map( D => n6400, CK => CLK, Q => 
                           n19399, QN => n9124);
   REGISTERS_reg_11_59_inst : DFF_X1 port map( D => n6399, CK => CLK, Q => 
                           n24331, QN => n9126);
   REGISTERS_reg_11_58_inst : DFF_X1 port map( D => n6398, CK => CLK, Q => 
                           n24330, QN => n9128);
   REGISTERS_reg_11_57_inst : DFF_X1 port map( D => n6397, CK => CLK, Q => 
                           n24329, QN => n9130);
   REGISTERS_reg_11_56_inst : DFF_X1 port map( D => n6396, CK => CLK, Q => 
                           n24328, QN => n9132);
   REGISTERS_reg_11_55_inst : DFF_X1 port map( D => n6395, CK => CLK, Q => 
                           n24327, QN => n9134);
   REGISTERS_reg_11_54_inst : DFF_X1 port map( D => n6394, CK => CLK, Q => 
                           n24326, QN => n9136);
   REGISTERS_reg_11_53_inst : DFF_X1 port map( D => n6393, CK => CLK, Q => 
                           n24325, QN => n9138);
   REGISTERS_reg_11_52_inst : DFF_X1 port map( D => n6392, CK => CLK, Q => 
                           n24324, QN => n9140);
   REGISTERS_reg_11_51_inst : DFF_X1 port map( D => n6391, CK => CLK, Q => 
                           n24323, QN => n9142);
   REGISTERS_reg_11_50_inst : DFF_X1 port map( D => n6390, CK => CLK, Q => 
                           n24322, QN => n9144);
   REGISTERS_reg_11_49_inst : DFF_X1 port map( D => n6389, CK => CLK, Q => 
                           n24321, QN => n9146);
   REGISTERS_reg_11_48_inst : DFF_X1 port map( D => n6388, CK => CLK, Q => 
                           n24320, QN => n9148);
   REGISTERS_reg_11_47_inst : DFF_X1 port map( D => n6387, CK => CLK, Q => 
                           n24319, QN => n9150);
   REGISTERS_reg_11_46_inst : DFF_X1 port map( D => n6386, CK => CLK, Q => 
                           n24318, QN => n9152);
   REGISTERS_reg_11_45_inst : DFF_X1 port map( D => n6385, CK => CLK, Q => 
                           n24317, QN => n9154);
   REGISTERS_reg_11_44_inst : DFF_X1 port map( D => n6384, CK => CLK, Q => 
                           n24316, QN => n9156);
   REGISTERS_reg_11_43_inst : DFF_X1 port map( D => n6383, CK => CLK, Q => 
                           n24315, QN => n9158);
   REGISTERS_reg_11_42_inst : DFF_X1 port map( D => n6382, CK => CLK, Q => 
                           n24314, QN => n9160);
   REGISTERS_reg_11_41_inst : DFF_X1 port map( D => n6381, CK => CLK, Q => 
                           n24313, QN => n9162);
   REGISTERS_reg_11_40_inst : DFF_X1 port map( D => n6380, CK => CLK, Q => 
                           n24312, QN => n9164);
   REGISTERS_reg_11_39_inst : DFF_X1 port map( D => n6379, CK => CLK, Q => 
                           n24311, QN => n9166);
   REGISTERS_reg_11_38_inst : DFF_X1 port map( D => n6378, CK => CLK, Q => 
                           n24310, QN => n9168);
   REGISTERS_reg_11_37_inst : DFF_X1 port map( D => n6377, CK => CLK, Q => 
                           n24309, QN => n9170);
   REGISTERS_reg_11_36_inst : DFF_X1 port map( D => n6376, CK => CLK, Q => 
                           n24308, QN => n9172);
   REGISTERS_reg_11_35_inst : DFF_X1 port map( D => n6375, CK => CLK, Q => 
                           n24307, QN => n9174);
   REGISTERS_reg_11_34_inst : DFF_X1 port map( D => n6374, CK => CLK, Q => 
                           n24306, QN => n9176);
   REGISTERS_reg_11_33_inst : DFF_X1 port map( D => n6373, CK => CLK, Q => 
                           n24305, QN => n9178);
   REGISTERS_reg_11_32_inst : DFF_X1 port map( D => n6372, CK => CLK, Q => 
                           n24304, QN => n9180);
   REGISTERS_reg_11_31_inst : DFF_X1 port map( D => n6371, CK => CLK, Q => 
                           n24303, QN => n9182);
   REGISTERS_reg_11_30_inst : DFF_X1 port map( D => n6370, CK => CLK, Q => 
                           n24302, QN => n9184);
   REGISTERS_reg_11_29_inst : DFF_X1 port map( D => n6369, CK => CLK, Q => 
                           n24301, QN => n9186);
   REGISTERS_reg_11_28_inst : DFF_X1 port map( D => n6368, CK => CLK, Q => 
                           n24300, QN => n9188);
   REGISTERS_reg_11_27_inst : DFF_X1 port map( D => n6367, CK => CLK, Q => 
                           n24299, QN => n9190);
   REGISTERS_reg_11_26_inst : DFF_X1 port map( D => n6366, CK => CLK, Q => 
                           n24298, QN => n9192);
   REGISTERS_reg_11_25_inst : DFF_X1 port map( D => n6365, CK => CLK, Q => 
                           n24297, QN => n9194);
   REGISTERS_reg_11_24_inst : DFF_X1 port map( D => n6364, CK => CLK, Q => 
                           n24296, QN => n9196);
   REGISTERS_reg_11_23_inst : DFF_X1 port map( D => n6363, CK => CLK, Q => 
                           n24295, QN => n9198);
   REGISTERS_reg_11_22_inst : DFF_X1 port map( D => n6362, CK => CLK, Q => 
                           n24294, QN => n9200);
   REGISTERS_reg_11_21_inst : DFF_X1 port map( D => n6361, CK => CLK, Q => 
                           n24293, QN => n9202);
   REGISTERS_reg_11_20_inst : DFF_X1 port map( D => n6360, CK => CLK, Q => 
                           n24292, QN => n9204);
   REGISTERS_reg_11_19_inst : DFF_X1 port map( D => n6359, CK => CLK, Q => 
                           n24291, QN => n9206);
   REGISTERS_reg_11_18_inst : DFF_X1 port map( D => n6358, CK => CLK, Q => 
                           n24290, QN => n9208);
   REGISTERS_reg_11_17_inst : DFF_X1 port map( D => n6357, CK => CLK, Q => 
                           n24289, QN => n9210);
   REGISTERS_reg_11_16_inst : DFF_X1 port map( D => n6356, CK => CLK, Q => 
                           n24288, QN => n9212);
   REGISTERS_reg_11_15_inst : DFF_X1 port map( D => n6355, CK => CLK, Q => 
                           n24287, QN => n9214);
   REGISTERS_reg_11_14_inst : DFF_X1 port map( D => n6354, CK => CLK, Q => 
                           n24286, QN => n9216);
   REGISTERS_reg_11_13_inst : DFF_X1 port map( D => n6353, CK => CLK, Q => 
                           n24285, QN => n9218);
   REGISTERS_reg_11_12_inst : DFF_X1 port map( D => n6352, CK => CLK, Q => 
                           n24284, QN => n9220);
   REGISTERS_reg_11_11_inst : DFF_X1 port map( D => n6351, CK => CLK, Q => 
                           n24283, QN => n9222);
   REGISTERS_reg_11_10_inst : DFF_X1 port map( D => n6350, CK => CLK, Q => 
                           n24282, QN => n9224);
   REGISTERS_reg_11_9_inst : DFF_X1 port map( D => n6349, CK => CLK, Q => 
                           n24281, QN => n9226);
   REGISTERS_reg_11_8_inst : DFF_X1 port map( D => n6348, CK => CLK, Q => 
                           n24280, QN => n9228);
   REGISTERS_reg_11_7_inst : DFF_X1 port map( D => n6347, CK => CLK, Q => 
                           n24279, QN => n9230);
   REGISTERS_reg_11_6_inst : DFF_X1 port map( D => n6346, CK => CLK, Q => 
                           n24278, QN => n9232);
   REGISTERS_reg_11_5_inst : DFF_X1 port map( D => n6345, CK => CLK, Q => 
                           n24277, QN => n9234);
   REGISTERS_reg_11_4_inst : DFF_X1 port map( D => n6344, CK => CLK, Q => 
                           n24276, QN => n9236);
   REGISTERS_reg_11_3_inst : DFF_X1 port map( D => n6343, CK => CLK, Q => 
                           n24275, QN => n9238);
   REGISTERS_reg_11_2_inst : DFF_X1 port map( D => n6342, CK => CLK, Q => 
                           n24274, QN => n9240);
   REGISTERS_reg_11_1_inst : DFF_X1 port map( D => n6341, CK => CLK, Q => 
                           n24273, QN => n9242);
   REGISTERS_reg_11_0_inst : DFF_X1 port map( D => n6340, CK => CLK, Q => 
                           n24272, QN => n9244);
   REGISTERS_reg_13_63_inst : DFF_X1 port map( D => n6275, CK => CLK, Q => 
                           n_1000, QN => n833);
   REGISTERS_reg_13_62_inst : DFF_X1 port map( D => n6274, CK => CLK, Q => 
                           n_1001, QN => n834);
   REGISTERS_reg_13_61_inst : DFF_X1 port map( D => n6273, CK => CLK, Q => 
                           n_1002, QN => n835);
   REGISTERS_reg_13_60_inst : DFF_X1 port map( D => n6272, CK => CLK, Q => 
                           n_1003, QN => n836);
   REGISTERS_reg_13_59_inst : DFF_X1 port map( D => n6271, CK => CLK, Q => 
                           n_1004, QN => n837);
   REGISTERS_reg_13_58_inst : DFF_X1 port map( D => n6270, CK => CLK, Q => 
                           n_1005, QN => n838);
   REGISTERS_reg_13_57_inst : DFF_X1 port map( D => n6269, CK => CLK, Q => 
                           n_1006, QN => n839);
   REGISTERS_reg_13_56_inst : DFF_X1 port map( D => n6268, CK => CLK, Q => 
                           n_1007, QN => n840);
   REGISTERS_reg_13_55_inst : DFF_X1 port map( D => n6267, CK => CLK, Q => 
                           n_1008, QN => n841);
   REGISTERS_reg_13_54_inst : DFF_X1 port map( D => n6266, CK => CLK, Q => 
                           n_1009, QN => n842);
   REGISTERS_reg_13_53_inst : DFF_X1 port map( D => n6265, CK => CLK, Q => 
                           n_1010, QN => n843);
   REGISTERS_reg_13_52_inst : DFF_X1 port map( D => n6264, CK => CLK, Q => 
                           n_1011, QN => n844);
   REGISTERS_reg_13_51_inst : DFF_X1 port map( D => n6263, CK => CLK, Q => 
                           n_1012, QN => n845);
   REGISTERS_reg_13_50_inst : DFF_X1 port map( D => n6262, CK => CLK, Q => 
                           n_1013, QN => n846);
   REGISTERS_reg_13_49_inst : DFF_X1 port map( D => n6261, CK => CLK, Q => 
                           n_1014, QN => n847);
   REGISTERS_reg_13_48_inst : DFF_X1 port map( D => n6260, CK => CLK, Q => 
                           n_1015, QN => n848);
   REGISTERS_reg_13_47_inst : DFF_X1 port map( D => n6259, CK => CLK, Q => 
                           n_1016, QN => n849);
   REGISTERS_reg_13_46_inst : DFF_X1 port map( D => n6258, CK => CLK, Q => 
                           n_1017, QN => n850);
   REGISTERS_reg_13_45_inst : DFF_X1 port map( D => n6257, CK => CLK, Q => 
                           n_1018, QN => n851);
   REGISTERS_reg_13_44_inst : DFF_X1 port map( D => n6256, CK => CLK, Q => 
                           n_1019, QN => n852);
   REGISTERS_reg_13_43_inst : DFF_X1 port map( D => n6255, CK => CLK, Q => 
                           n_1020, QN => n853);
   REGISTERS_reg_13_42_inst : DFF_X1 port map( D => n6254, CK => CLK, Q => 
                           n_1021, QN => n854);
   REGISTERS_reg_13_41_inst : DFF_X1 port map( D => n6253, CK => CLK, Q => 
                           n_1022, QN => n855);
   REGISTERS_reg_13_40_inst : DFF_X1 port map( D => n6252, CK => CLK, Q => 
                           n_1023, QN => n856);
   REGISTERS_reg_13_39_inst : DFF_X1 port map( D => n6251, CK => CLK, Q => 
                           n_1024, QN => n857);
   REGISTERS_reg_13_38_inst : DFF_X1 port map( D => n6250, CK => CLK, Q => 
                           n_1025, QN => n858);
   REGISTERS_reg_13_37_inst : DFF_X1 port map( D => n6249, CK => CLK, Q => 
                           n_1026, QN => n859);
   REGISTERS_reg_13_36_inst : DFF_X1 port map( D => n6248, CK => CLK, Q => 
                           n_1027, QN => n860);
   REGISTERS_reg_13_35_inst : DFF_X1 port map( D => n6247, CK => CLK, Q => 
                           n_1028, QN => n861);
   REGISTERS_reg_13_34_inst : DFF_X1 port map( D => n6246, CK => CLK, Q => 
                           n_1029, QN => n862);
   REGISTERS_reg_13_33_inst : DFF_X1 port map( D => n6245, CK => CLK, Q => 
                           n_1030, QN => n863);
   REGISTERS_reg_13_32_inst : DFF_X1 port map( D => n6244, CK => CLK, Q => 
                           n_1031, QN => n864);
   REGISTERS_reg_13_31_inst : DFF_X1 port map( D => n6243, CK => CLK, Q => 
                           n_1032, QN => n865);
   REGISTERS_reg_13_30_inst : DFF_X1 port map( D => n6242, CK => CLK, Q => 
                           n_1033, QN => n866);
   REGISTERS_reg_13_29_inst : DFF_X1 port map( D => n6241, CK => CLK, Q => 
                           n_1034, QN => n867);
   REGISTERS_reg_13_28_inst : DFF_X1 port map( D => n6240, CK => CLK, Q => 
                           n_1035, QN => n868);
   REGISTERS_reg_13_27_inst : DFF_X1 port map( D => n6239, CK => CLK, Q => 
                           n_1036, QN => n869);
   REGISTERS_reg_13_26_inst : DFF_X1 port map( D => n6238, CK => CLK, Q => 
                           n_1037, QN => n870);
   REGISTERS_reg_13_25_inst : DFF_X1 port map( D => n6237, CK => CLK, Q => 
                           n_1038, QN => n871);
   REGISTERS_reg_13_24_inst : DFF_X1 port map( D => n6236, CK => CLK, Q => 
                           n_1039, QN => n872);
   REGISTERS_reg_13_23_inst : DFF_X1 port map( D => n6235, CK => CLK, Q => 
                           n_1040, QN => n873);
   REGISTERS_reg_13_22_inst : DFF_X1 port map( D => n6234, CK => CLK, Q => 
                           n_1041, QN => n874);
   REGISTERS_reg_13_21_inst : DFF_X1 port map( D => n6233, CK => CLK, Q => 
                           n_1042, QN => n875);
   REGISTERS_reg_13_20_inst : DFF_X1 port map( D => n6232, CK => CLK, Q => 
                           n_1043, QN => n876);
   REGISTERS_reg_13_19_inst : DFF_X1 port map( D => n6231, CK => CLK, Q => 
                           n_1044, QN => n877);
   REGISTERS_reg_13_18_inst : DFF_X1 port map( D => n6230, CK => CLK, Q => 
                           n_1045, QN => n878);
   REGISTERS_reg_13_17_inst : DFF_X1 port map( D => n6229, CK => CLK, Q => 
                           n_1046, QN => n879);
   REGISTERS_reg_13_16_inst : DFF_X1 port map( D => n6228, CK => CLK, Q => 
                           n_1047, QN => n880);
   REGISTERS_reg_13_15_inst : DFF_X1 port map( D => n6227, CK => CLK, Q => 
                           n_1048, QN => n881);
   REGISTERS_reg_13_14_inst : DFF_X1 port map( D => n6226, CK => CLK, Q => 
                           n_1049, QN => n882);
   REGISTERS_reg_13_13_inst : DFF_X1 port map( D => n6225, CK => CLK, Q => 
                           n_1050, QN => n883);
   REGISTERS_reg_13_12_inst : DFF_X1 port map( D => n6224, CK => CLK, Q => 
                           n_1051, QN => n884);
   REGISTERS_reg_13_11_inst : DFF_X1 port map( D => n6223, CK => CLK, Q => 
                           n_1052, QN => n885);
   REGISTERS_reg_13_10_inst : DFF_X1 port map( D => n6222, CK => CLK, Q => 
                           n_1053, QN => n886);
   REGISTERS_reg_13_9_inst : DFF_X1 port map( D => n6221, CK => CLK, Q => 
                           n_1054, QN => n887);
   REGISTERS_reg_13_8_inst : DFF_X1 port map( D => n6220, CK => CLK, Q => 
                           n_1055, QN => n888);
   REGISTERS_reg_13_7_inst : DFF_X1 port map( D => n6219, CK => CLK, Q => 
                           n_1056, QN => n889);
   REGISTERS_reg_13_6_inst : DFF_X1 port map( D => n6218, CK => CLK, Q => 
                           n_1057, QN => n890);
   REGISTERS_reg_13_5_inst : DFF_X1 port map( D => n6217, CK => CLK, Q => 
                           n_1058, QN => n891);
   REGISTERS_reg_13_4_inst : DFF_X1 port map( D => n6216, CK => CLK, Q => 
                           n_1059, QN => n892);
   REGISTERS_reg_13_3_inst : DFF_X1 port map( D => n6215, CK => CLK, Q => 
                           n_1060, QN => n893);
   REGISTERS_reg_13_2_inst : DFF_X1 port map( D => n6214, CK => CLK, Q => 
                           n_1061, QN => n894);
   REGISTERS_reg_13_1_inst : DFF_X1 port map( D => n6213, CK => CLK, Q => 
                           n_1062, QN => n895);
   REGISTERS_reg_13_0_inst : DFF_X1 port map( D => n6212, CK => CLK, Q => 
                           n_1063, QN => n896);
   REGISTERS_reg_23_59_inst : DFF_X1 port map( D => n5631, CK => CLK, Q => 
                           n19588, QN => n9127);
   REGISTERS_reg_23_58_inst : DFF_X1 port map( D => n5630, CK => CLK, Q => 
                           n19589, QN => n9129);
   REGISTERS_reg_23_57_inst : DFF_X1 port map( D => n5629, CK => CLK, Q => 
                           n19590, QN => n9131);
   REGISTERS_reg_23_56_inst : DFF_X1 port map( D => n5628, CK => CLK, Q => 
                           n19591, QN => n9133);
   REGISTERS_reg_23_55_inst : DFF_X1 port map( D => n5627, CK => CLK, Q => 
                           n19592, QN => n9135);
   REGISTERS_reg_23_54_inst : DFF_X1 port map( D => n5626, CK => CLK, Q => 
                           n19593, QN => n9137);
   REGISTERS_reg_23_53_inst : DFF_X1 port map( D => n5625, CK => CLK, Q => 
                           n19594, QN => n9139);
   REGISTERS_reg_23_52_inst : DFF_X1 port map( D => n5624, CK => CLK, Q => 
                           n19595, QN => n9141);
   REGISTERS_reg_23_51_inst : DFF_X1 port map( D => n5623, CK => CLK, Q => 
                           n19596, QN => n9143);
   REGISTERS_reg_23_50_inst : DFF_X1 port map( D => n5622, CK => CLK, Q => 
                           n19597, QN => n9145);
   REGISTERS_reg_23_49_inst : DFF_X1 port map( D => n5621, CK => CLK, Q => 
                           n19598, QN => n9147);
   REGISTERS_reg_23_48_inst : DFF_X1 port map( D => n5620, CK => CLK, Q => 
                           n19599, QN => n9149);
   REGISTERS_reg_23_47_inst : DFF_X1 port map( D => n5619, CK => CLK, Q => 
                           n19600, QN => n9151);
   REGISTERS_reg_23_46_inst : DFF_X1 port map( D => n5618, CK => CLK, Q => 
                           n19601, QN => n9153);
   REGISTERS_reg_23_45_inst : DFF_X1 port map( D => n5617, CK => CLK, Q => 
                           n19602, QN => n9155);
   REGISTERS_reg_23_44_inst : DFF_X1 port map( D => n5616, CK => CLK, Q => 
                           n19603, QN => n9157);
   REGISTERS_reg_23_43_inst : DFF_X1 port map( D => n5615, CK => CLK, Q => 
                           n19604, QN => n9159);
   REGISTERS_reg_23_42_inst : DFF_X1 port map( D => n5614, CK => CLK, Q => 
                           n19605, QN => n9161);
   REGISTERS_reg_23_41_inst : DFF_X1 port map( D => n5613, CK => CLK, Q => 
                           n19606, QN => n9163);
   REGISTERS_reg_23_40_inst : DFF_X1 port map( D => n5612, CK => CLK, Q => 
                           n19607, QN => n9165);
   REGISTERS_reg_23_39_inst : DFF_X1 port map( D => n5611, CK => CLK, Q => 
                           n19608, QN => n9167);
   REGISTERS_reg_23_38_inst : DFF_X1 port map( D => n5610, CK => CLK, Q => 
                           n19609, QN => n9169);
   REGISTERS_reg_23_37_inst : DFF_X1 port map( D => n5609, CK => CLK, Q => 
                           n19610, QN => n9171);
   REGISTERS_reg_23_36_inst : DFF_X1 port map( D => n5608, CK => CLK, Q => 
                           n19611, QN => n9173);
   REGISTERS_reg_23_35_inst : DFF_X1 port map( D => n5607, CK => CLK, Q => 
                           n19612, QN => n9175);
   REGISTERS_reg_23_34_inst : DFF_X1 port map( D => n5606, CK => CLK, Q => 
                           n19613, QN => n9177);
   REGISTERS_reg_23_33_inst : DFF_X1 port map( D => n5605, CK => CLK, Q => 
                           n19614, QN => n9179);
   REGISTERS_reg_23_32_inst : DFF_X1 port map( D => n5604, CK => CLK, Q => 
                           n19615, QN => n9181);
   REGISTERS_reg_23_31_inst : DFF_X1 port map( D => n5603, CK => CLK, Q => 
                           n19616, QN => n9183);
   REGISTERS_reg_23_30_inst : DFF_X1 port map( D => n5602, CK => CLK, Q => 
                           n19617, QN => n9185);
   REGISTERS_reg_23_29_inst : DFF_X1 port map( D => n5601, CK => CLK, Q => 
                           n19618, QN => n9187);
   REGISTERS_reg_23_28_inst : DFF_X1 port map( D => n5600, CK => CLK, Q => 
                           n19619, QN => n9189);
   REGISTERS_reg_23_27_inst : DFF_X1 port map( D => n5599, CK => CLK, Q => 
                           n19620, QN => n9191);
   REGISTERS_reg_23_26_inst : DFF_X1 port map( D => n5598, CK => CLK, Q => 
                           n19621, QN => n9193);
   REGISTERS_reg_23_25_inst : DFF_X1 port map( D => n5597, CK => CLK, Q => 
                           n19622, QN => n9195);
   REGISTERS_reg_23_24_inst : DFF_X1 port map( D => n5596, CK => CLK, Q => 
                           n19623, QN => n9197);
   REGISTERS_reg_23_23_inst : DFF_X1 port map( D => n5595, CK => CLK, Q => 
                           n19624, QN => n9199);
   REGISTERS_reg_23_22_inst : DFF_X1 port map( D => n5594, CK => CLK, Q => 
                           n19625, QN => n9201);
   REGISTERS_reg_23_21_inst : DFF_X1 port map( D => n5593, CK => CLK, Q => 
                           n19626, QN => n9203);
   REGISTERS_reg_23_20_inst : DFF_X1 port map( D => n5592, CK => CLK, Q => 
                           n19627, QN => n9205);
   REGISTERS_reg_23_19_inst : DFF_X1 port map( D => n5591, CK => CLK, Q => 
                           n19628, QN => n9207);
   REGISTERS_reg_23_18_inst : DFF_X1 port map( D => n5590, CK => CLK, Q => 
                           n19629, QN => n9209);
   REGISTERS_reg_23_17_inst : DFF_X1 port map( D => n5589, CK => CLK, Q => 
                           n19630, QN => n9211);
   REGISTERS_reg_23_16_inst : DFF_X1 port map( D => n5588, CK => CLK, Q => 
                           n19631, QN => n9213);
   REGISTERS_reg_23_15_inst : DFF_X1 port map( D => n5587, CK => CLK, Q => 
                           n19632, QN => n9215);
   REGISTERS_reg_23_14_inst : DFF_X1 port map( D => n5586, CK => CLK, Q => 
                           n19633, QN => n9217);
   REGISTERS_reg_23_13_inst : DFF_X1 port map( D => n5585, CK => CLK, Q => 
                           n19634, QN => n9219);
   REGISTERS_reg_23_12_inst : DFF_X1 port map( D => n5584, CK => CLK, Q => 
                           n19635, QN => n9221);
   REGISTERS_reg_23_11_inst : DFF_X1 port map( D => n5583, CK => CLK, Q => 
                           n19636, QN => n9223);
   REGISTERS_reg_23_10_inst : DFF_X1 port map( D => n5582, CK => CLK, Q => 
                           n19637, QN => n9225);
   REGISTERS_reg_23_9_inst : DFF_X1 port map( D => n5581, CK => CLK, Q => 
                           n19638, QN => n9227);
   REGISTERS_reg_23_8_inst : DFF_X1 port map( D => n5580, CK => CLK, Q => 
                           n19639, QN => n9229);
   REGISTERS_reg_23_7_inst : DFF_X1 port map( D => n5579, CK => CLK, Q => 
                           n19640, QN => n9231);
   REGISTERS_reg_23_6_inst : DFF_X1 port map( D => n5578, CK => CLK, Q => 
                           n19641, QN => n9233);
   REGISTERS_reg_23_5_inst : DFF_X1 port map( D => n5577, CK => CLK, Q => 
                           n19642, QN => n9235);
   REGISTERS_reg_23_4_inst : DFF_X1 port map( D => n5576, CK => CLK, Q => 
                           n19643, QN => n9237);
   REGISTERS_reg_23_3_inst : DFF_X1 port map( D => n5575, CK => CLK, Q => 
                           n19644, QN => n9239);
   REGISTERS_reg_23_2_inst : DFF_X1 port map( D => n5574, CK => CLK, Q => 
                           n19645, QN => n9241);
   REGISTERS_reg_23_1_inst : DFF_X1 port map( D => n5573, CK => CLK, Q => 
                           n19646, QN => n9243);
   REGISTERS_reg_23_0_inst : DFF_X1 port map( D => n5572, CK => CLK, Q => 
                           n19647, QN => n9245);
   REGISTERS_reg_25_62_inst : DFF_X1 port map( D => n5506, CK => CLK, Q => 
                           n_1064, QN => n7303);
   REGISTERS_reg_25_61_inst : DFF_X1 port map( D => n5505, CK => CLK, Q => 
                           n_1065, QN => n7305);
   REGISTERS_reg_25_60_inst : DFF_X1 port map( D => n5504, CK => CLK, Q => 
                           n_1066, QN => n7307);
   REGISTERS_reg_25_59_inst : DFF_X1 port map( D => n5503, CK => CLK, Q => 
                           n_1067, QN => n7309);
   REGISTERS_reg_25_58_inst : DFF_X1 port map( D => n5502, CK => CLK, Q => 
                           n_1068, QN => n7311);
   REGISTERS_reg_25_57_inst : DFF_X1 port map( D => n5501, CK => CLK, Q => 
                           n_1069, QN => n7313);
   REGISTERS_reg_25_56_inst : DFF_X1 port map( D => n5500, CK => CLK, Q => 
                           n_1070, QN => n7315);
   REGISTERS_reg_25_55_inst : DFF_X1 port map( D => n5499, CK => CLK, Q => 
                           n_1071, QN => n7317);
   REGISTERS_reg_25_54_inst : DFF_X1 port map( D => n5498, CK => CLK, Q => 
                           n_1072, QN => n7319);
   REGISTERS_reg_25_53_inst : DFF_X1 port map( D => n5497, CK => CLK, Q => 
                           n_1073, QN => n7321);
   REGISTERS_reg_25_52_inst : DFF_X1 port map( D => n5496, CK => CLK, Q => 
                           n_1074, QN => n7323);
   REGISTERS_reg_25_51_inst : DFF_X1 port map( D => n5495, CK => CLK, Q => 
                           n_1075, QN => n7325);
   REGISTERS_reg_25_50_inst : DFF_X1 port map( D => n5494, CK => CLK, Q => 
                           n_1076, QN => n7327);
   REGISTERS_reg_25_49_inst : DFF_X1 port map( D => n5493, CK => CLK, Q => 
                           n_1077, QN => n7329);
   REGISTERS_reg_25_48_inst : DFF_X1 port map( D => n5492, CK => CLK, Q => 
                           n_1078, QN => n7331);
   REGISTERS_reg_25_47_inst : DFF_X1 port map( D => n5491, CK => CLK, Q => 
                           n_1079, QN => n7333);
   REGISTERS_reg_25_46_inst : DFF_X1 port map( D => n5490, CK => CLK, Q => 
                           n_1080, QN => n7335);
   REGISTERS_reg_25_45_inst : DFF_X1 port map( D => n5489, CK => CLK, Q => 
                           n_1081, QN => n7337);
   REGISTERS_reg_25_44_inst : DFF_X1 port map( D => n5488, CK => CLK, Q => 
                           n_1082, QN => n7339);
   REGISTERS_reg_25_43_inst : DFF_X1 port map( D => n5487, CK => CLK, Q => 
                           n_1083, QN => n7341);
   REGISTERS_reg_25_42_inst : DFF_X1 port map( D => n5486, CK => CLK, Q => 
                           n_1084, QN => n7343);
   REGISTERS_reg_25_41_inst : DFF_X1 port map( D => n5485, CK => CLK, Q => 
                           n_1085, QN => n7345);
   REGISTERS_reg_25_40_inst : DFF_X1 port map( D => n5484, CK => CLK, Q => 
                           n_1086, QN => n7347);
   REGISTERS_reg_25_39_inst : DFF_X1 port map( D => n5483, CK => CLK, Q => 
                           n_1087, QN => n7349);
   REGISTERS_reg_25_38_inst : DFF_X1 port map( D => n5482, CK => CLK, Q => 
                           n_1088, QN => n7351);
   REGISTERS_reg_25_37_inst : DFF_X1 port map( D => n5481, CK => CLK, Q => 
                           n_1089, QN => n7353);
   REGISTERS_reg_25_36_inst : DFF_X1 port map( D => n5480, CK => CLK, Q => 
                           n_1090, QN => n7355);
   REGISTERS_reg_25_35_inst : DFF_X1 port map( D => n5479, CK => CLK, Q => 
                           n_1091, QN => n7357);
   REGISTERS_reg_25_34_inst : DFF_X1 port map( D => n5478, CK => CLK, Q => 
                           n_1092, QN => n7359);
   REGISTERS_reg_25_33_inst : DFF_X1 port map( D => n5477, CK => CLK, Q => 
                           n_1093, QN => n7361);
   REGISTERS_reg_25_32_inst : DFF_X1 port map( D => n5476, CK => CLK, Q => 
                           n_1094, QN => n7363);
   REGISTERS_reg_25_31_inst : DFF_X1 port map( D => n5475, CK => CLK, Q => 
                           n_1095, QN => n7365);
   REGISTERS_reg_25_30_inst : DFF_X1 port map( D => n5474, CK => CLK, Q => 
                           n_1096, QN => n7367);
   REGISTERS_reg_25_29_inst : DFF_X1 port map( D => n5473, CK => CLK, Q => 
                           n_1097, QN => n7369);
   REGISTERS_reg_25_28_inst : DFF_X1 port map( D => n5472, CK => CLK, Q => 
                           n_1098, QN => n7371);
   REGISTERS_reg_25_27_inst : DFF_X1 port map( D => n5471, CK => CLK, Q => 
                           n_1099, QN => n7373);
   REGISTERS_reg_25_26_inst : DFF_X1 port map( D => n5470, CK => CLK, Q => 
                           n_1100, QN => n7375);
   REGISTERS_reg_25_25_inst : DFF_X1 port map( D => n5469, CK => CLK, Q => 
                           n_1101, QN => n7377);
   REGISTERS_reg_25_24_inst : DFF_X1 port map( D => n5468, CK => CLK, Q => 
                           n_1102, QN => n7379);
   REGISTERS_reg_25_23_inst : DFF_X1 port map( D => n5467, CK => CLK, Q => 
                           n_1103, QN => n7381);
   REGISTERS_reg_25_22_inst : DFF_X1 port map( D => n5466, CK => CLK, Q => 
                           n_1104, QN => n7383);
   REGISTERS_reg_25_21_inst : DFF_X1 port map( D => n5465, CK => CLK, Q => 
                           n_1105, QN => n7385);
   REGISTERS_reg_25_20_inst : DFF_X1 port map( D => n5464, CK => CLK, Q => 
                           n_1106, QN => n7387);
   REGISTERS_reg_25_19_inst : DFF_X1 port map( D => n5463, CK => CLK, Q => 
                           n_1107, QN => n7389);
   REGISTERS_reg_25_18_inst : DFF_X1 port map( D => n5462, CK => CLK, Q => 
                           n_1108, QN => n7391);
   REGISTERS_reg_25_17_inst : DFF_X1 port map( D => n5461, CK => CLK, Q => 
                           n_1109, QN => n7393);
   REGISTERS_reg_25_16_inst : DFF_X1 port map( D => n5460, CK => CLK, Q => 
                           n_1110, QN => n7395);
   REGISTERS_reg_25_15_inst : DFF_X1 port map( D => n5459, CK => CLK, Q => 
                           n_1111, QN => n7397);
   REGISTERS_reg_25_14_inst : DFF_X1 port map( D => n5458, CK => CLK, Q => 
                           n_1112, QN => n7399);
   REGISTERS_reg_25_13_inst : DFF_X1 port map( D => n5457, CK => CLK, Q => 
                           n_1113, QN => n7401);
   REGISTERS_reg_25_12_inst : DFF_X1 port map( D => n5456, CK => CLK, Q => 
                           n_1114, QN => n7403);
   REGISTERS_reg_25_11_inst : DFF_X1 port map( D => n5455, CK => CLK, Q => 
                           n_1115, QN => n7405);
   REGISTERS_reg_25_10_inst : DFF_X1 port map( D => n5454, CK => CLK, Q => 
                           n_1116, QN => n7407);
   REGISTERS_reg_25_9_inst : DFF_X1 port map( D => n5453, CK => CLK, Q => 
                           n_1117, QN => n7409);
   REGISTERS_reg_25_8_inst : DFF_X1 port map( D => n5452, CK => CLK, Q => 
                           n_1118, QN => n7411);
   REGISTERS_reg_25_7_inst : DFF_X1 port map( D => n5451, CK => CLK, Q => 
                           n_1119, QN => n7413);
   REGISTERS_reg_25_6_inst : DFF_X1 port map( D => n5450, CK => CLK, Q => 
                           n_1120, QN => n7415);
   REGISTERS_reg_25_5_inst : DFF_X1 port map( D => n5449, CK => CLK, Q => 
                           n_1121, QN => n7417);
   REGISTERS_reg_25_4_inst : DFF_X1 port map( D => n5448, CK => CLK, Q => 
                           n_1122, QN => n7419);
   REGISTERS_reg_25_3_inst : DFF_X1 port map( D => n5447, CK => CLK, Q => 
                           n_1123, QN => n7421);
   REGISTERS_reg_25_2_inst : DFF_X1 port map( D => n5446, CK => CLK, Q => 
                           n_1124, QN => n7423);
   REGISTERS_reg_25_1_inst : DFF_X1 port map( D => n5445, CK => CLK, Q => 
                           n_1125, QN => n7425);
   REGISTERS_reg_25_0_inst : DFF_X1 port map( D => n5444, CK => CLK, Q => 
                           n_1126, QN => n7427);
   REGISTERS_reg_29_63_inst : DFF_X1 port map( D => n5251, CK => CLK, Q => 
                           n24355, QN => n8862);
   REGISTERS_reg_29_62_inst : DFF_X1 port map( D => n5250, CK => CLK, Q => 
                           n24354, QN => n8864);
   REGISTERS_reg_29_61_inst : DFF_X1 port map( D => n5249, CK => CLK, Q => 
                           n24353, QN => n8866);
   REGISTERS_reg_29_60_inst : DFF_X1 port map( D => n5248, CK => CLK, Q => 
                           n24352, QN => n8868);
   REGISTERS_reg_29_59_inst : DFF_X1 port map( D => n5247, CK => CLK, Q => 
                           n24351, QN => n8870);
   REGISTERS_reg_29_58_inst : DFF_X1 port map( D => n5246, CK => CLK, Q => 
                           n24350, QN => n8872);
   REGISTERS_reg_29_57_inst : DFF_X1 port map( D => n5245, CK => CLK, Q => 
                           n24349, QN => n8874);
   REGISTERS_reg_29_56_inst : DFF_X1 port map( D => n5244, CK => CLK, Q => 
                           n24348, QN => n8876);
   REGISTERS_reg_29_55_inst : DFF_X1 port map( D => n5243, CK => CLK, Q => 
                           n24347, QN => n8878);
   REGISTERS_reg_29_54_inst : DFF_X1 port map( D => n5242, CK => CLK, Q => 
                           n24346, QN => n8880);
   REGISTERS_reg_29_53_inst : DFF_X1 port map( D => n5241, CK => CLK, Q => 
                           n24345, QN => n8882);
   REGISTERS_reg_29_52_inst : DFF_X1 port map( D => n5240, CK => CLK, Q => 
                           n24344, QN => n8884);
   REGISTERS_reg_29_51_inst : DFF_X1 port map( D => n5239, CK => CLK, Q => 
                           n24343, QN => n8886);
   REGISTERS_reg_29_50_inst : DFF_X1 port map( D => n5238, CK => CLK, Q => 
                           n24342, QN => n8888);
   REGISTERS_reg_29_49_inst : DFF_X1 port map( D => n5237, CK => CLK, Q => 
                           n24341, QN => n8890);
   REGISTERS_reg_29_48_inst : DFF_X1 port map( D => n5236, CK => CLK, Q => 
                           n24340, QN => n8892);
   REGISTERS_reg_29_47_inst : DFF_X1 port map( D => n5235, CK => CLK, Q => 
                           n24339, QN => n8894);
   REGISTERS_reg_29_46_inst : DFF_X1 port map( D => n5234, CK => CLK, Q => 
                           n24338, QN => n8896);
   REGISTERS_reg_29_45_inst : DFF_X1 port map( D => n5233, CK => CLK, Q => 
                           n24337, QN => n8898);
   REGISTERS_reg_29_44_inst : DFF_X1 port map( D => n5232, CK => CLK, Q => 
                           n24336, QN => n8900);
   REGISTERS_reg_29_43_inst : DFF_X1 port map( D => n5231, CK => CLK, Q => 
                           n24335, QN => n8902);
   REGISTERS_reg_29_42_inst : DFF_X1 port map( D => n5230, CK => CLK, Q => 
                           n24334, QN => n8904);
   REGISTERS_reg_29_41_inst : DFF_X1 port map( D => n5229, CK => CLK, Q => 
                           n24333, QN => n8906);
   REGISTERS_reg_29_40_inst : DFF_X1 port map( D => n5228, CK => CLK, Q => 
                           n24332, QN => n8908);
   REGISTERS_reg_29_39_inst : DFF_X1 port map( D => n5227, CK => CLK, Q => 
                           n24395, QN => n8910);
   REGISTERS_reg_29_38_inst : DFF_X1 port map( D => n5226, CK => CLK, Q => 
                           n24394, QN => n8912);
   REGISTERS_reg_29_37_inst : DFF_X1 port map( D => n5225, CK => CLK, Q => 
                           n24393, QN => n8914);
   REGISTERS_reg_29_36_inst : DFF_X1 port map( D => n5224, CK => CLK, Q => 
                           n24392, QN => n8916);
   REGISTERS_reg_29_35_inst : DFF_X1 port map( D => n5223, CK => CLK, Q => 
                           n24391, QN => n8918);
   REGISTERS_reg_29_34_inst : DFF_X1 port map( D => n5222, CK => CLK, Q => 
                           n24390, QN => n8920);
   REGISTERS_reg_29_33_inst : DFF_X1 port map( D => n5221, CK => CLK, Q => 
                           n24389, QN => n8922);
   REGISTERS_reg_29_32_inst : DFF_X1 port map( D => n5220, CK => CLK, Q => 
                           n24388, QN => n8924);
   REGISTERS_reg_29_31_inst : DFF_X1 port map( D => n5219, CK => CLK, Q => 
                           n24387, QN => n8926);
   REGISTERS_reg_29_30_inst : DFF_X1 port map( D => n5218, CK => CLK, Q => 
                           n24386, QN => n8928);
   REGISTERS_reg_29_29_inst : DFF_X1 port map( D => n5217, CK => CLK, Q => 
                           n24385, QN => n8930);
   REGISTERS_reg_29_28_inst : DFF_X1 port map( D => n5216, CK => CLK, Q => 
                           n24384, QN => n8932);
   REGISTERS_reg_29_27_inst : DFF_X1 port map( D => n5215, CK => CLK, Q => 
                           n24383, QN => n8934);
   REGISTERS_reg_29_26_inst : DFF_X1 port map( D => n5214, CK => CLK, Q => 
                           n24382, QN => n8936);
   REGISTERS_reg_29_25_inst : DFF_X1 port map( D => n5213, CK => CLK, Q => 
                           n24381, QN => n8938);
   REGISTERS_reg_29_24_inst : DFF_X1 port map( D => n5212, CK => CLK, Q => 
                           n24380, QN => n8940);
   REGISTERS_reg_29_23_inst : DFF_X1 port map( D => n5211, CK => CLK, Q => 
                           n24379, QN => n8942);
   REGISTERS_reg_29_22_inst : DFF_X1 port map( D => n5210, CK => CLK, Q => 
                           n24378, QN => n8944);
   REGISTERS_reg_29_21_inst : DFF_X1 port map( D => n5209, CK => CLK, Q => 
                           n24377, QN => n8946);
   REGISTERS_reg_29_20_inst : DFF_X1 port map( D => n5208, CK => CLK, Q => 
                           n24376, QN => n8948);
   REGISTERS_reg_29_19_inst : DFF_X1 port map( D => n5207, CK => CLK, Q => 
                           n24375, QN => n8950);
   REGISTERS_reg_29_18_inst : DFF_X1 port map( D => n5206, CK => CLK, Q => 
                           n24374, QN => n8952);
   REGISTERS_reg_29_17_inst : DFF_X1 port map( D => n5205, CK => CLK, Q => 
                           n24373, QN => n8954);
   REGISTERS_reg_29_16_inst : DFF_X1 port map( D => n5204, CK => CLK, Q => 
                           n24372, QN => n8956);
   REGISTERS_reg_29_15_inst : DFF_X1 port map( D => n5203, CK => CLK, Q => 
                           n24371, QN => n8958);
   REGISTERS_reg_29_14_inst : DFF_X1 port map( D => n5202, CK => CLK, Q => 
                           n24370, QN => n8960);
   REGISTERS_reg_29_13_inst : DFF_X1 port map( D => n5201, CK => CLK, Q => 
                           n24369, QN => n8962);
   REGISTERS_reg_29_12_inst : DFF_X1 port map( D => n5200, CK => CLK, Q => 
                           n24368, QN => n8964);
   REGISTERS_reg_29_11_inst : DFF_X1 port map( D => n5199, CK => CLK, Q => 
                           n24367, QN => n8966);
   REGISTERS_reg_29_10_inst : DFF_X1 port map( D => n5198, CK => CLK, Q => 
                           n24366, QN => n8968);
   REGISTERS_reg_29_9_inst : DFF_X1 port map( D => n5197, CK => CLK, Q => 
                           n24365, QN => n8970);
   REGISTERS_reg_29_8_inst : DFF_X1 port map( D => n5196, CK => CLK, Q => 
                           n24364, QN => n8972);
   REGISTERS_reg_29_7_inst : DFF_X1 port map( D => n5195, CK => CLK, Q => 
                           n24363, QN => n8974);
   REGISTERS_reg_29_6_inst : DFF_X1 port map( D => n5194, CK => CLK, Q => 
                           n24362, QN => n8976);
   REGISTERS_reg_29_5_inst : DFF_X1 port map( D => n5193, CK => CLK, Q => 
                           n24361, QN => n8978);
   REGISTERS_reg_29_4_inst : DFF_X1 port map( D => n5192, CK => CLK, Q => 
                           n24360, QN => n8980);
   REGISTERS_reg_29_3_inst : DFF_X1 port map( D => n5191, CK => CLK, Q => 
                           n24359, QN => n8982);
   REGISTERS_reg_29_2_inst : DFF_X1 port map( D => n5190, CK => CLK, Q => 
                           n24358, QN => n8984);
   REGISTERS_reg_29_1_inst : DFF_X1 port map( D => n5189, CK => CLK, Q => 
                           n24357, QN => n8986);
   REGISTERS_reg_29_0_inst : DFF_X1 port map( D => n5188, CK => CLK, Q => 
                           n24356, QN => n8988);
   OUT1_reg_63_inst : DFF_X1 port map( D => n5059, CK => CLK, Q => OUT1(63), QN
                           => n11846);
   OUT1_reg_62_inst : DFF_X1 port map( D => n5058, CK => CLK, Q => OUT1(62), QN
                           => n11845);
   OUT1_reg_61_inst : DFF_X1 port map( D => n5057, CK => CLK, Q => OUT1(61), QN
                           => n11844);
   OUT1_reg_60_inst : DFF_X1 port map( D => n5056, CK => CLK, Q => OUT1(60), QN
                           => n11843);
   OUT1_reg_59_inst : DFF_X1 port map( D => n5055, CK => CLK, Q => OUT1(59), QN
                           => n11842);
   OUT1_reg_58_inst : DFF_X1 port map( D => n5054, CK => CLK, Q => OUT1(58), QN
                           => n11841);
   OUT1_reg_57_inst : DFF_X1 port map( D => n5053, CK => CLK, Q => OUT1(57), QN
                           => n11840);
   OUT1_reg_56_inst : DFF_X1 port map( D => n5052, CK => CLK, Q => OUT1(56), QN
                           => n11839);
   OUT1_reg_55_inst : DFF_X1 port map( D => n5051, CK => CLK, Q => OUT1(55), QN
                           => n11838);
   OUT1_reg_54_inst : DFF_X1 port map( D => n5050, CK => CLK, Q => OUT1(54), QN
                           => n11837);
   OUT1_reg_53_inst : DFF_X1 port map( D => n5049, CK => CLK, Q => OUT1(53), QN
                           => n11836);
   OUT1_reg_52_inst : DFF_X1 port map( D => n5048, CK => CLK, Q => OUT1(52), QN
                           => n11835);
   OUT1_reg_51_inst : DFF_X1 port map( D => n5047, CK => CLK, Q => OUT1(51), QN
                           => n11834);
   OUT1_reg_50_inst : DFF_X1 port map( D => n5046, CK => CLK, Q => OUT1(50), QN
                           => n11833);
   OUT1_reg_49_inst : DFF_X1 port map( D => n5045, CK => CLK, Q => OUT1(49), QN
                           => n11832);
   OUT1_reg_48_inst : DFF_X1 port map( D => n5044, CK => CLK, Q => OUT1(48), QN
                           => n11831);
   OUT1_reg_47_inst : DFF_X1 port map( D => n5043, CK => CLK, Q => OUT1(47), QN
                           => n11830);
   OUT1_reg_46_inst : DFF_X1 port map( D => n5042, CK => CLK, Q => OUT1(46), QN
                           => n11829);
   OUT1_reg_45_inst : DFF_X1 port map( D => n5041, CK => CLK, Q => OUT1(45), QN
                           => n11828);
   OUT1_reg_44_inst : DFF_X1 port map( D => n5040, CK => CLK, Q => OUT1(44), QN
                           => n11827);
   OUT1_reg_43_inst : DFF_X1 port map( D => n5039, CK => CLK, Q => OUT1(43), QN
                           => n11826);
   OUT1_reg_42_inst : DFF_X1 port map( D => n5038, CK => CLK, Q => OUT1(42), QN
                           => n11825);
   OUT1_reg_41_inst : DFF_X1 port map( D => n5037, CK => CLK, Q => OUT1(41), QN
                           => n11824);
   OUT1_reg_40_inst : DFF_X1 port map( D => n5036, CK => CLK, Q => OUT1(40), QN
                           => n11823);
   OUT1_reg_39_inst : DFF_X1 port map( D => n5035, CK => CLK, Q => OUT1(39), QN
                           => n11822);
   OUT1_reg_38_inst : DFF_X1 port map( D => n5034, CK => CLK, Q => OUT1(38), QN
                           => n11821);
   OUT1_reg_37_inst : DFF_X1 port map( D => n5033, CK => CLK, Q => OUT1(37), QN
                           => n11820);
   OUT1_reg_36_inst : DFF_X1 port map( D => n5032, CK => CLK, Q => OUT1(36), QN
                           => n11819);
   OUT1_reg_35_inst : DFF_X1 port map( D => n5031, CK => CLK, Q => OUT1(35), QN
                           => n11818);
   OUT1_reg_34_inst : DFF_X1 port map( D => n5030, CK => CLK, Q => OUT1(34), QN
                           => n11817);
   OUT1_reg_33_inst : DFF_X1 port map( D => n5029, CK => CLK, Q => OUT1(33), QN
                           => n11816);
   OUT1_reg_32_inst : DFF_X1 port map( D => n5028, CK => CLK, Q => OUT1(32), QN
                           => n11815);
   OUT1_reg_31_inst : DFF_X1 port map( D => n5027, CK => CLK, Q => OUT1(31), QN
                           => n11814);
   OUT1_reg_30_inst : DFF_X1 port map( D => n5026, CK => CLK, Q => OUT1(30), QN
                           => n11813);
   OUT1_reg_29_inst : DFF_X1 port map( D => n5025, CK => CLK, Q => OUT1(29), QN
                           => n11812);
   OUT1_reg_28_inst : DFF_X1 port map( D => n5024, CK => CLK, Q => OUT1(28), QN
                           => n11811);
   OUT1_reg_27_inst : DFF_X1 port map( D => n5023, CK => CLK, Q => OUT1(27), QN
                           => n11810);
   OUT1_reg_26_inst : DFF_X1 port map( D => n5022, CK => CLK, Q => OUT1(26), QN
                           => n11809);
   OUT1_reg_25_inst : DFF_X1 port map( D => n5021, CK => CLK, Q => OUT1(25), QN
                           => n11808);
   OUT1_reg_24_inst : DFF_X1 port map( D => n5020, CK => CLK, Q => OUT1(24), QN
                           => n11807);
   OUT1_reg_23_inst : DFF_X1 port map( D => n5019, CK => CLK, Q => OUT1(23), QN
                           => n11806);
   OUT1_reg_22_inst : DFF_X1 port map( D => n5018, CK => CLK, Q => OUT1(22), QN
                           => n11805);
   OUT1_reg_21_inst : DFF_X1 port map( D => n5017, CK => CLK, Q => OUT1(21), QN
                           => n11804);
   OUT1_reg_20_inst : DFF_X1 port map( D => n5016, CK => CLK, Q => OUT1(20), QN
                           => n11803);
   OUT1_reg_19_inst : DFF_X1 port map( D => n5015, CK => CLK, Q => OUT1(19), QN
                           => n11802);
   OUT1_reg_18_inst : DFF_X1 port map( D => n5014, CK => CLK, Q => OUT1(18), QN
                           => n11801);
   OUT1_reg_17_inst : DFF_X1 port map( D => n5013, CK => CLK, Q => OUT1(17), QN
                           => n11800);
   OUT1_reg_16_inst : DFF_X1 port map( D => n5012, CK => CLK, Q => OUT1(16), QN
                           => n11799);
   OUT1_reg_15_inst : DFF_X1 port map( D => n5011, CK => CLK, Q => OUT1(15), QN
                           => n11798);
   OUT1_reg_14_inst : DFF_X1 port map( D => n5010, CK => CLK, Q => OUT1(14), QN
                           => n11797);
   OUT1_reg_13_inst : DFF_X1 port map( D => n5009, CK => CLK, Q => OUT1(13), QN
                           => n11796);
   OUT1_reg_12_inst : DFF_X1 port map( D => n5008, CK => CLK, Q => OUT1(12), QN
                           => n11795);
   OUT1_reg_11_inst : DFF_X1 port map( D => n5007, CK => CLK, Q => OUT1(11), QN
                           => n11794);
   OUT1_reg_10_inst : DFF_X1 port map( D => n5006, CK => CLK, Q => OUT1(10), QN
                           => n11793);
   OUT1_reg_9_inst : DFF_X1 port map( D => n5005, CK => CLK, Q => OUT1(9), QN 
                           => n11792);
   OUT1_reg_8_inst : DFF_X1 port map( D => n5004, CK => CLK, Q => OUT1(8), QN 
                           => n11791);
   OUT1_reg_7_inst : DFF_X1 port map( D => n5003, CK => CLK, Q => OUT1(7), QN 
                           => n11790);
   OUT1_reg_6_inst : DFF_X1 port map( D => n5002, CK => CLK, Q => OUT1(6), QN 
                           => n11789);
   OUT1_reg_5_inst : DFF_X1 port map( D => n5001, CK => CLK, Q => OUT1(5), QN 
                           => n11788);
   OUT1_reg_4_inst : DFF_X1 port map( D => n5000, CK => CLK, Q => OUT1(4), QN 
                           => n11787);
   OUT1_reg_3_inst : DFF_X1 port map( D => n4999, CK => CLK, Q => OUT1(3), QN 
                           => n11786);
   OUT1_reg_2_inst : DFF_X1 port map( D => n4998, CK => CLK, Q => OUT1(2), QN 
                           => n11785);
   OUT1_reg_1_inst : DFF_X1 port map( D => n4997, CK => CLK, Q => OUT1(1), QN 
                           => n11784);
   OUT1_reg_0_inst : DFF_X1 port map( D => n4996, CK => CLK, Q => OUT1(0), QN 
                           => n11783);
   OUT2_reg_39_inst : DFF_X1 port map( D => n4971, CK => CLK, Q => OUT2_39_port
                           , QN => n_1127);
   OUT2_reg_38_inst : DFF_X1 port map( D => n4970, CK => CLK, Q => OUT2_38_port
                           , QN => n_1128);
   OUT2_reg_37_inst : DFF_X1 port map( D => n4969, CK => CLK, Q => OUT2_37_port
                           , QN => n_1129);
   OUT2_reg_36_inst : DFF_X1 port map( D => n4968, CK => CLK, Q => OUT2_36_port
                           , QN => n_1130);
   OUT2_reg_35_inst : DFF_X1 port map( D => n4967, CK => CLK, Q => OUT2_35_port
                           , QN => n_1131);
   OUT2_reg_34_inst : DFF_X1 port map( D => n4966, CK => CLK, Q => OUT2_34_port
                           , QN => n_1132);
   OUT2_reg_33_inst : DFF_X1 port map( D => n4965, CK => CLK, Q => OUT2_33_port
                           , QN => n_1133);
   OUT2_reg_32_inst : DFF_X1 port map( D => n4964, CK => CLK, Q => OUT2_32_port
                           , QN => n_1134);
   OUT2_reg_31_inst : DFF_X1 port map( D => n4963, CK => CLK, Q => OUT2_31_port
                           , QN => n_1135);
   OUT2_reg_30_inst : DFF_X1 port map( D => n4962, CK => CLK, Q => OUT2_30_port
                           , QN => n_1136);
   OUT2_reg_29_inst : DFF_X1 port map( D => n4961, CK => CLK, Q => OUT2_29_port
                           , QN => n_1137);
   OUT2_reg_28_inst : DFF_X1 port map( D => n4960, CK => CLK, Q => OUT2_28_port
                           , QN => n_1138);
   OUT2_reg_27_inst : DFF_X1 port map( D => n4959, CK => CLK, Q => OUT2_27_port
                           , QN => n_1139);
   OUT2_reg_26_inst : DFF_X1 port map( D => n4958, CK => CLK, Q => OUT2_26_port
                           , QN => n_1140);
   OUT2_reg_25_inst : DFF_X1 port map( D => n4957, CK => CLK, Q => OUT2_25_port
                           , QN => n_1141);
   OUT2_reg_24_inst : DFF_X1 port map( D => n4956, CK => CLK, Q => OUT2_24_port
                           , QN => n_1142);
   OUT2_reg_23_inst : DFF_X1 port map( D => n4955, CK => CLK, Q => OUT2_23_port
                           , QN => n_1143);
   OUT2_reg_22_inst : DFF_X1 port map( D => n4954, CK => CLK, Q => OUT2_22_port
                           , QN => n_1144);
   OUT2_reg_21_inst : DFF_X1 port map( D => n4953, CK => CLK, Q => OUT2_21_port
                           , QN => n_1145);
   OUT2_reg_20_inst : DFF_X1 port map( D => n4952, CK => CLK, Q => OUT2_20_port
                           , QN => n_1146);
   OUT2_reg_19_inst : DFF_X1 port map( D => n4951, CK => CLK, Q => OUT2_19_port
                           , QN => n_1147);
   OUT2_reg_18_inst : DFF_X1 port map( D => n4950, CK => CLK, Q => OUT2_18_port
                           , QN => n_1148);
   OUT2_reg_17_inst : DFF_X1 port map( D => n4949, CK => CLK, Q => OUT2_17_port
                           , QN => n_1149);
   OUT2_reg_16_inst : DFF_X1 port map( D => n4948, CK => CLK, Q => OUT2_16_port
                           , QN => n_1150);
   OUT2_reg_15_inst : DFF_X1 port map( D => n4947, CK => CLK, Q => OUT2_15_port
                           , QN => n_1151);
   OUT2_reg_14_inst : DFF_X1 port map( D => n4946, CK => CLK, Q => OUT2_14_port
                           , QN => n_1152);
   OUT2_reg_13_inst : DFF_X1 port map( D => n4945, CK => CLK, Q => OUT2_13_port
                           , QN => n_1153);
   OUT2_reg_12_inst : DFF_X1 port map( D => n4944, CK => CLK, Q => OUT2_12_port
                           , QN => n_1154);
   OUT2_reg_11_inst : DFF_X1 port map( D => n4943, CK => CLK, Q => OUT2_11_port
                           , QN => n_1155);
   OUT2_reg_10_inst : DFF_X1 port map( D => n4942, CK => CLK, Q => OUT2_10_port
                           , QN => n_1156);
   OUT2_reg_9_inst : DFF_X1 port map( D => n4941, CK => CLK, Q => OUT2_9_port, 
                           QN => n_1157);
   OUT2_reg_8_inst : DFF_X1 port map( D => n4940, CK => CLK, Q => OUT2_8_port, 
                           QN => n_1158);
   OUT2_reg_7_inst : DFF_X1 port map( D => n4939, CK => CLK, Q => OUT2_7_port, 
                           QN => n_1159);
   OUT2_reg_6_inst : DFF_X1 port map( D => n4938, CK => CLK, Q => OUT2_6_port, 
                           QN => n_1160);
   OUT2_reg_5_inst : DFF_X1 port map( D => n4937, CK => CLK, Q => OUT2_5_port, 
                           QN => n_1161);
   OUT2_reg_4_inst : DFF_X1 port map( D => n4936, CK => CLK, Q => OUT2_4_port, 
                           QN => n_1162);
   OUT2_reg_3_inst : DFF_X1 port map( D => n4935, CK => CLK, Q => OUT2_3_port, 
                           QN => n_1163);
   OUT2_reg_2_inst : DFF_X1 port map( D => n4934, CK => CLK, Q => OUT2_2_port, 
                           QN => n_1164);
   OUT2_reg_1_inst : DFF_X1 port map( D => n4933, CK => CLK, Q => OUT2_1_port, 
                           QN => n_1165);
   OUT2_reg_0_inst : DFF_X1 port map( D => n4932, CK => CLK, Q => OUT2_0_port, 
                           QN => n_1166);
   REGISTERS_reg_19_63_inst : DFF_X1 port map( D => n5891, CK => CLK, Q => 
                           n19802, QN => n8863);
   REGISTERS_reg_19_62_inst : DFF_X1 port map( D => n5890, CK => CLK, Q => 
                           n19803, QN => n8865);
   REGISTERS_reg_19_61_inst : DFF_X1 port map( D => n5889, CK => CLK, Q => 
                           n19804, QN => n8867);
   REGISTERS_reg_19_60_inst : DFF_X1 port map( D => n5888, CK => CLK, Q => 
                           n19805, QN => n8869);
   REGISTERS_reg_15_63_inst : DFF_X1 port map( D => n6147, CK => CLK, Q => 
                           n19810, QN => n7300);
   REGISTERS_reg_15_62_inst : DFF_X1 port map( D => n6146, CK => CLK, Q => 
                           n19811, QN => n7302);
   REGISTERS_reg_15_61_inst : DFF_X1 port map( D => n6145, CK => CLK, Q => 
                           n19812, QN => n7304);
   REGISTERS_reg_15_60_inst : DFF_X1 port map( D => n6144, CK => CLK, Q => 
                           n19813, QN => n7306);
   REGISTERS_reg_10_63_inst : DFF_X1 port map( D => n6467, CK => CLK, Q => 
                           n19814, QN => n7428);
   REGISTERS_reg_10_62_inst : DFF_X1 port map( D => n6466, CK => CLK, Q => 
                           n19815, QN => n7430);
   REGISTERS_reg_10_61_inst : DFF_X1 port map( D => n6465, CK => CLK, Q => 
                           n19816, QN => n7432);
   REGISTERS_reg_10_60_inst : DFF_X1 port map( D => n6464, CK => CLK, Q => 
                           n19817, QN => n7434);
   REGISTERS_reg_5_63_inst : DFF_X1 port map( D => n6787, CK => CLK, Q => 
                           n24211, QN => n17221);
   REGISTERS_reg_5_62_inst : DFF_X1 port map( D => n6786, CK => CLK, Q => 
                           n24210, QN => n17224);
   REGISTERS_reg_5_61_inst : DFF_X1 port map( D => n6785, CK => CLK, Q => 
                           n24209, QN => n17227);
   REGISTERS_reg_5_60_inst : DFF_X1 port map( D => n6784, CK => CLK, Q => 
                           n24208, QN => n17230);
   REGISTERS_reg_19_59_inst : DFF_X1 port map( D => n5887, CK => CLK, Q => 
                           n19822, QN => n8871);
   REGISTERS_reg_19_58_inst : DFF_X1 port map( D => n5886, CK => CLK, Q => 
                           n19823, QN => n8873);
   REGISTERS_reg_19_57_inst : DFF_X1 port map( D => n5885, CK => CLK, Q => 
                           n19824, QN => n8875);
   REGISTERS_reg_19_56_inst : DFF_X1 port map( D => n5884, CK => CLK, Q => 
                           n19825, QN => n8877);
   REGISTERS_reg_19_55_inst : DFF_X1 port map( D => n5883, CK => CLK, Q => 
                           n19826, QN => n8879);
   REGISTERS_reg_19_54_inst : DFF_X1 port map( D => n5882, CK => CLK, Q => 
                           n19827, QN => n8881);
   REGISTERS_reg_19_53_inst : DFF_X1 port map( D => n5881, CK => CLK, Q => 
                           n19828, QN => n8883);
   REGISTERS_reg_19_52_inst : DFF_X1 port map( D => n5880, CK => CLK, Q => 
                           n19829, QN => n8885);
   REGISTERS_reg_19_51_inst : DFF_X1 port map( D => n5879, CK => CLK, Q => 
                           n19830, QN => n8887);
   REGISTERS_reg_19_50_inst : DFF_X1 port map( D => n5878, CK => CLK, Q => 
                           n19831, QN => n8889);
   REGISTERS_reg_19_49_inst : DFF_X1 port map( D => n5877, CK => CLK, Q => 
                           n19832, QN => n8891);
   REGISTERS_reg_19_48_inst : DFF_X1 port map( D => n5876, CK => CLK, Q => 
                           n19833, QN => n8893);
   REGISTERS_reg_19_47_inst : DFF_X1 port map( D => n5875, CK => CLK, Q => 
                           n19834, QN => n8895);
   REGISTERS_reg_19_46_inst : DFF_X1 port map( D => n5874, CK => CLK, Q => 
                           n19835, QN => n8897);
   REGISTERS_reg_19_45_inst : DFF_X1 port map( D => n5873, CK => CLK, Q => 
                           n19836, QN => n8899);
   REGISTERS_reg_19_44_inst : DFF_X1 port map( D => n5872, CK => CLK, Q => 
                           n19837, QN => n8901);
   REGISTERS_reg_19_43_inst : DFF_X1 port map( D => n5871, CK => CLK, Q => 
                           n19838, QN => n8903);
   REGISTERS_reg_19_42_inst : DFF_X1 port map( D => n5870, CK => CLK, Q => 
                           n19839, QN => n8905);
   REGISTERS_reg_19_41_inst : DFF_X1 port map( D => n5869, CK => CLK, Q => 
                           n19840, QN => n8907);
   REGISTERS_reg_19_40_inst : DFF_X1 port map( D => n5868, CK => CLK, Q => 
                           n19841, QN => n8909);
   REGISTERS_reg_19_39_inst : DFF_X1 port map( D => n5867, CK => CLK, Q => 
                           n19842, QN => n8911);
   REGISTERS_reg_19_38_inst : DFF_X1 port map( D => n5866, CK => CLK, Q => 
                           n19843, QN => n8913);
   REGISTERS_reg_19_37_inst : DFF_X1 port map( D => n5865, CK => CLK, Q => 
                           n19844, QN => n8915);
   REGISTERS_reg_19_36_inst : DFF_X1 port map( D => n5864, CK => CLK, Q => 
                           n19845, QN => n8917);
   REGISTERS_reg_19_35_inst : DFF_X1 port map( D => n5863, CK => CLK, Q => 
                           n19846, QN => n8919);
   REGISTERS_reg_19_34_inst : DFF_X1 port map( D => n5862, CK => CLK, Q => 
                           n19847, QN => n8921);
   REGISTERS_reg_19_33_inst : DFF_X1 port map( D => n5861, CK => CLK, Q => 
                           n19848, QN => n8923);
   REGISTERS_reg_19_32_inst : DFF_X1 port map( D => n5860, CK => CLK, Q => 
                           n19849, QN => n8925);
   REGISTERS_reg_19_31_inst : DFF_X1 port map( D => n5859, CK => CLK, Q => 
                           n19850, QN => n8927);
   REGISTERS_reg_19_30_inst : DFF_X1 port map( D => n5858, CK => CLK, Q => 
                           n19851, QN => n8929);
   REGISTERS_reg_19_29_inst : DFF_X1 port map( D => n5857, CK => CLK, Q => 
                           n19852, QN => n8931);
   REGISTERS_reg_19_28_inst : DFF_X1 port map( D => n5856, CK => CLK, Q => 
                           n19853, QN => n8933);
   REGISTERS_reg_19_27_inst : DFF_X1 port map( D => n5855, CK => CLK, Q => 
                           n19854, QN => n8935);
   REGISTERS_reg_19_26_inst : DFF_X1 port map( D => n5854, CK => CLK, Q => 
                           n19855, QN => n8937);
   REGISTERS_reg_19_25_inst : DFF_X1 port map( D => n5853, CK => CLK, Q => 
                           n19856, QN => n8939);
   REGISTERS_reg_19_24_inst : DFF_X1 port map( D => n5852, CK => CLK, Q => 
                           n19857, QN => n8941);
   REGISTERS_reg_15_59_inst : DFF_X1 port map( D => n6143, CK => CLK, Q => 
                           n19894, QN => n7308);
   REGISTERS_reg_15_58_inst : DFF_X1 port map( D => n6142, CK => CLK, Q => 
                           n19895, QN => n7310);
   REGISTERS_reg_15_57_inst : DFF_X1 port map( D => n6141, CK => CLK, Q => 
                           n19896, QN => n7312);
   REGISTERS_reg_15_56_inst : DFF_X1 port map( D => n6140, CK => CLK, Q => 
                           n19897, QN => n7314);
   REGISTERS_reg_15_55_inst : DFF_X1 port map( D => n6139, CK => CLK, Q => 
                           n19898, QN => n7316);
   REGISTERS_reg_15_54_inst : DFF_X1 port map( D => n6138, CK => CLK, Q => 
                           n19899, QN => n7318);
   REGISTERS_reg_15_53_inst : DFF_X1 port map( D => n6137, CK => CLK, Q => 
                           n19900, QN => n7320);
   REGISTERS_reg_15_52_inst : DFF_X1 port map( D => n6136, CK => CLK, Q => 
                           n19901, QN => n7322);
   REGISTERS_reg_15_51_inst : DFF_X1 port map( D => n6135, CK => CLK, Q => 
                           n19902, QN => n7324);
   REGISTERS_reg_15_50_inst : DFF_X1 port map( D => n6134, CK => CLK, Q => 
                           n19903, QN => n7326);
   REGISTERS_reg_15_49_inst : DFF_X1 port map( D => n6133, CK => CLK, Q => 
                           n19904, QN => n7328);
   REGISTERS_reg_15_48_inst : DFF_X1 port map( D => n6132, CK => CLK, Q => 
                           n19905, QN => n7330);
   REGISTERS_reg_15_47_inst : DFF_X1 port map( D => n6131, CK => CLK, Q => 
                           n19906, QN => n7332);
   REGISTERS_reg_15_46_inst : DFF_X1 port map( D => n6130, CK => CLK, Q => 
                           n19907, QN => n7334);
   REGISTERS_reg_15_45_inst : DFF_X1 port map( D => n6129, CK => CLK, Q => 
                           n19908, QN => n7336);
   REGISTERS_reg_15_44_inst : DFF_X1 port map( D => n6128, CK => CLK, Q => 
                           n19909, QN => n7338);
   REGISTERS_reg_15_43_inst : DFF_X1 port map( D => n6127, CK => CLK, Q => 
                           n19910, QN => n7340);
   REGISTERS_reg_15_42_inst : DFF_X1 port map( D => n6126, CK => CLK, Q => 
                           n19911, QN => n7342);
   REGISTERS_reg_15_41_inst : DFF_X1 port map( D => n6125, CK => CLK, Q => 
                           n19912, QN => n7344);
   REGISTERS_reg_15_40_inst : DFF_X1 port map( D => n6124, CK => CLK, Q => 
                           n19913, QN => n7346);
   REGISTERS_reg_15_39_inst : DFF_X1 port map( D => n6123, CK => CLK, Q => 
                           n19914, QN => n7348);
   REGISTERS_reg_15_38_inst : DFF_X1 port map( D => n6122, CK => CLK, Q => 
                           n19915, QN => n7350);
   REGISTERS_reg_15_37_inst : DFF_X1 port map( D => n6121, CK => CLK, Q => 
                           n19916, QN => n7352);
   REGISTERS_reg_15_36_inst : DFF_X1 port map( D => n6120, CK => CLK, Q => 
                           n19917, QN => n7354);
   REGISTERS_reg_15_35_inst : DFF_X1 port map( D => n6119, CK => CLK, Q => 
                           n19918, QN => n7356);
   REGISTERS_reg_15_34_inst : DFF_X1 port map( D => n6118, CK => CLK, Q => 
                           n19919, QN => n7358);
   REGISTERS_reg_15_33_inst : DFF_X1 port map( D => n6117, CK => CLK, Q => 
                           n19920, QN => n7360);
   REGISTERS_reg_15_32_inst : DFF_X1 port map( D => n6116, CK => CLK, Q => 
                           n19921, QN => n7362);
   REGISTERS_reg_15_31_inst : DFF_X1 port map( D => n6115, CK => CLK, Q => 
                           n19922, QN => n7364);
   REGISTERS_reg_15_30_inst : DFF_X1 port map( D => n6114, CK => CLK, Q => 
                           n19923, QN => n7366);
   REGISTERS_reg_15_29_inst : DFF_X1 port map( D => n6113, CK => CLK, Q => 
                           n19924, QN => n7368);
   REGISTERS_reg_15_28_inst : DFF_X1 port map( D => n6112, CK => CLK, Q => 
                           n19925, QN => n7370);
   REGISTERS_reg_15_27_inst : DFF_X1 port map( D => n6111, CK => CLK, Q => 
                           n19926, QN => n7372);
   REGISTERS_reg_15_26_inst : DFF_X1 port map( D => n6110, CK => CLK, Q => 
                           n19927, QN => n7374);
   REGISTERS_reg_15_25_inst : DFF_X1 port map( D => n6109, CK => CLK, Q => 
                           n19928, QN => n7376);
   REGISTERS_reg_15_24_inst : DFF_X1 port map( D => n6108, CK => CLK, Q => 
                           n19929, QN => n7378);
   REGISTERS_reg_10_59_inst : DFF_X1 port map( D => n6463, CK => CLK, Q => 
                           n24207, QN => n7436);
   REGISTERS_reg_10_58_inst : DFF_X1 port map( D => n6462, CK => CLK, Q => 
                           n24206, QN => n7438);
   REGISTERS_reg_10_57_inst : DFF_X1 port map( D => n6461, CK => CLK, Q => 
                           n24205, QN => n7440);
   REGISTERS_reg_10_56_inst : DFF_X1 port map( D => n6460, CK => CLK, Q => 
                           n24204, QN => n7442);
   REGISTERS_reg_10_55_inst : DFF_X1 port map( D => n6459, CK => CLK, Q => 
                           n24203, QN => n7444);
   REGISTERS_reg_10_54_inst : DFF_X1 port map( D => n6458, CK => CLK, Q => 
                           n24202, QN => n7446);
   REGISTERS_reg_10_53_inst : DFF_X1 port map( D => n6457, CK => CLK, Q => 
                           n24201, QN => n7448);
   REGISTERS_reg_10_52_inst : DFF_X1 port map( D => n6456, CK => CLK, Q => 
                           n24200, QN => n7450);
   REGISTERS_reg_10_51_inst : DFF_X1 port map( D => n6455, CK => CLK, Q => 
                           n24199, QN => n7452);
   REGISTERS_reg_10_50_inst : DFF_X1 port map( D => n6454, CK => CLK, Q => 
                           n24198, QN => n7454);
   REGISTERS_reg_10_49_inst : DFF_X1 port map( D => n6453, CK => CLK, Q => 
                           n24197, QN => n7456);
   REGISTERS_reg_10_48_inst : DFF_X1 port map( D => n6452, CK => CLK, Q => 
                           n24196, QN => n7458);
   REGISTERS_reg_10_47_inst : DFF_X1 port map( D => n6451, CK => CLK, Q => 
                           n24195, QN => n7460);
   REGISTERS_reg_10_46_inst : DFF_X1 port map( D => n6450, CK => CLK, Q => 
                           n24194, QN => n7462);
   REGISTERS_reg_10_45_inst : DFF_X1 port map( D => n6449, CK => CLK, Q => 
                           n24193, QN => n7464);
   REGISTERS_reg_10_44_inst : DFF_X1 port map( D => n6448, CK => CLK, Q => 
                           n24192, QN => n7466);
   REGISTERS_reg_10_43_inst : DFF_X1 port map( D => n6447, CK => CLK, Q => 
                           n24191, QN => n7468);
   REGISTERS_reg_10_42_inst : DFF_X1 port map( D => n6446, CK => CLK, Q => 
                           n24190, QN => n7470);
   REGISTERS_reg_10_41_inst : DFF_X1 port map( D => n6445, CK => CLK, Q => 
                           n24189, QN => n7472);
   REGISTERS_reg_10_40_inst : DFF_X1 port map( D => n6444, CK => CLK, Q => 
                           n24188, QN => n7474);
   REGISTERS_reg_10_39_inst : DFF_X1 port map( D => n6443, CK => CLK, Q => 
                           n24187, QN => n7476);
   REGISTERS_reg_10_38_inst : DFF_X1 port map( D => n6442, CK => CLK, Q => 
                           n24186, QN => n7478);
   REGISTERS_reg_10_37_inst : DFF_X1 port map( D => n6441, CK => CLK, Q => 
                           n24185, QN => n7480);
   REGISTERS_reg_10_36_inst : DFF_X1 port map( D => n6440, CK => CLK, Q => 
                           n24184, QN => n7482);
   REGISTERS_reg_10_35_inst : DFF_X1 port map( D => n6439, CK => CLK, Q => 
                           n24183, QN => n7484);
   REGISTERS_reg_10_34_inst : DFF_X1 port map( D => n6438, CK => CLK, Q => 
                           n24182, QN => n7486);
   REGISTERS_reg_10_33_inst : DFF_X1 port map( D => n6437, CK => CLK, Q => 
                           n24181, QN => n7488);
   REGISTERS_reg_10_32_inst : DFF_X1 port map( D => n6436, CK => CLK, Q => 
                           n24180, QN => n7490);
   REGISTERS_reg_10_31_inst : DFF_X1 port map( D => n6435, CK => CLK, Q => 
                           n24179, QN => n7492);
   REGISTERS_reg_10_30_inst : DFF_X1 port map( D => n6434, CK => CLK, Q => 
                           n24178, QN => n7494);
   REGISTERS_reg_10_29_inst : DFF_X1 port map( D => n6433, CK => CLK, Q => 
                           n24177, QN => n7496);
   REGISTERS_reg_10_28_inst : DFF_X1 port map( D => n6432, CK => CLK, Q => 
                           n24176, QN => n7498);
   REGISTERS_reg_10_27_inst : DFF_X1 port map( D => n6431, CK => CLK, Q => 
                           n24175, QN => n7500);
   REGISTERS_reg_10_26_inst : DFF_X1 port map( D => n6430, CK => CLK, Q => 
                           n24174, QN => n7502);
   REGISTERS_reg_10_25_inst : DFF_X1 port map( D => n6429, CK => CLK, Q => 
                           n24173, QN => n7504);
   REGISTERS_reg_10_24_inst : DFF_X1 port map( D => n6428, CK => CLK, Q => 
                           n24172, QN => n7506);
   REGISTERS_reg_5_59_inst : DFF_X1 port map( D => n6783, CK => CLK, Q => 
                           n24271, QN => n17233);
   REGISTERS_reg_5_58_inst : DFF_X1 port map( D => n6782, CK => CLK, Q => 
                           n24270, QN => n17236);
   REGISTERS_reg_5_57_inst : DFF_X1 port map( D => n6781, CK => CLK, Q => 
                           n24269, QN => n17239);
   REGISTERS_reg_5_56_inst : DFF_X1 port map( D => n6780, CK => CLK, Q => 
                           n24268, QN => n17242);
   REGISTERS_reg_5_55_inst : DFF_X1 port map( D => n6779, CK => CLK, Q => 
                           n24267, QN => n17245);
   REGISTERS_reg_5_54_inst : DFF_X1 port map( D => n6778, CK => CLK, Q => 
                           n24266, QN => n17248);
   REGISTERS_reg_5_53_inst : DFF_X1 port map( D => n6777, CK => CLK, Q => 
                           n24265, QN => n17251);
   REGISTERS_reg_5_52_inst : DFF_X1 port map( D => n6776, CK => CLK, Q => 
                           n24264, QN => n17254);
   REGISTERS_reg_5_51_inst : DFF_X1 port map( D => n6775, CK => CLK, Q => 
                           n24263, QN => n17257);
   REGISTERS_reg_5_50_inst : DFF_X1 port map( D => n6774, CK => CLK, Q => 
                           n24262, QN => n17260);
   REGISTERS_reg_5_49_inst : DFF_X1 port map( D => n6773, CK => CLK, Q => 
                           n24261, QN => n17263);
   REGISTERS_reg_5_48_inst : DFF_X1 port map( D => n6772, CK => CLK, Q => 
                           n24260, QN => n17266);
   REGISTERS_reg_5_47_inst : DFF_X1 port map( D => n6771, CK => CLK, Q => 
                           n24259, QN => n17269);
   REGISTERS_reg_5_46_inst : DFF_X1 port map( D => n6770, CK => CLK, Q => 
                           n24258, QN => n17272);
   REGISTERS_reg_5_45_inst : DFF_X1 port map( D => n6769, CK => CLK, Q => 
                           n24257, QN => n17275);
   REGISTERS_reg_5_44_inst : DFF_X1 port map( D => n6768, CK => CLK, Q => 
                           n24256, QN => n17278);
   REGISTERS_reg_5_43_inst : DFF_X1 port map( D => n6767, CK => CLK, Q => 
                           n24255, QN => n17281);
   REGISTERS_reg_5_42_inst : DFF_X1 port map( D => n6766, CK => CLK, Q => 
                           n24254, QN => n17284);
   REGISTERS_reg_5_41_inst : DFF_X1 port map( D => n6765, CK => CLK, Q => 
                           n24253, QN => n17287);
   REGISTERS_reg_5_40_inst : DFF_X1 port map( D => n6764, CK => CLK, Q => 
                           n24252, QN => n17290);
   REGISTERS_reg_5_39_inst : DFF_X1 port map( D => n6763, CK => CLK, Q => 
                           n24251, QN => n17293);
   REGISTERS_reg_5_38_inst : DFF_X1 port map( D => n6762, CK => CLK, Q => 
                           n24250, QN => n17296);
   REGISTERS_reg_5_37_inst : DFF_X1 port map( D => n6761, CK => CLK, Q => 
                           n24249, QN => n17299);
   REGISTERS_reg_5_36_inst : DFF_X1 port map( D => n6760, CK => CLK, Q => 
                           n24248, QN => n17302);
   REGISTERS_reg_5_35_inst : DFF_X1 port map( D => n6759, CK => CLK, Q => 
                           n24247, QN => n17305);
   REGISTERS_reg_5_34_inst : DFF_X1 port map( D => n6758, CK => CLK, Q => 
                           n24246, QN => n17308);
   REGISTERS_reg_5_33_inst : DFF_X1 port map( D => n6757, CK => CLK, Q => 
                           n24245, QN => n17311);
   REGISTERS_reg_5_32_inst : DFF_X1 port map( D => n6756, CK => CLK, Q => 
                           n24244, QN => n17314);
   REGISTERS_reg_5_31_inst : DFF_X1 port map( D => n6755, CK => CLK, Q => 
                           n24243, QN => n17317);
   REGISTERS_reg_5_30_inst : DFF_X1 port map( D => n6754, CK => CLK, Q => 
                           n24242, QN => n17320);
   REGISTERS_reg_5_29_inst : DFF_X1 port map( D => n6753, CK => CLK, Q => 
                           n24241, QN => n17323);
   REGISTERS_reg_5_28_inst : DFF_X1 port map( D => n6752, CK => CLK, Q => 
                           n24240, QN => n17326);
   REGISTERS_reg_5_27_inst : DFF_X1 port map( D => n6751, CK => CLK, Q => 
                           n24239, QN => n17329);
   REGISTERS_reg_5_26_inst : DFF_X1 port map( D => n6750, CK => CLK, Q => 
                           n24238, QN => n17332);
   REGISTERS_reg_5_25_inst : DFF_X1 port map( D => n6749, CK => CLK, Q => 
                           n24237, QN => n17335);
   REGISTERS_reg_5_24_inst : DFF_X1 port map( D => n6748, CK => CLK, Q => 
                           n24236, QN => n17338);
   REGISTERS_reg_19_23_inst : DFF_X1 port map( D => n5851, CK => CLK, Q => 
                           n20002, QN => n8943);
   REGISTERS_reg_19_22_inst : DFF_X1 port map( D => n5850, CK => CLK, Q => 
                           n20003, QN => n8945);
   REGISTERS_reg_19_21_inst : DFF_X1 port map( D => n5849, CK => CLK, Q => 
                           n20004, QN => n8947);
   REGISTERS_reg_19_20_inst : DFF_X1 port map( D => n5848, CK => CLK, Q => 
                           n20005, QN => n8949);
   REGISTERS_reg_19_19_inst : DFF_X1 port map( D => n5847, CK => CLK, Q => 
                           n20006, QN => n8951);
   REGISTERS_reg_19_18_inst : DFF_X1 port map( D => n5846, CK => CLK, Q => 
                           n20007, QN => n8953);
   REGISTERS_reg_19_17_inst : DFF_X1 port map( D => n5845, CK => CLK, Q => 
                           n20008, QN => n8955);
   REGISTERS_reg_19_16_inst : DFF_X1 port map( D => n5844, CK => CLK, Q => 
                           n20009, QN => n8957);
   REGISTERS_reg_19_15_inst : DFF_X1 port map( D => n5843, CK => CLK, Q => 
                           n20010, QN => n8959);
   REGISTERS_reg_19_14_inst : DFF_X1 port map( D => n5842, CK => CLK, Q => 
                           n20011, QN => n8961);
   REGISTERS_reg_19_13_inst : DFF_X1 port map( D => n5841, CK => CLK, Q => 
                           n20012, QN => n8963);
   REGISTERS_reg_19_12_inst : DFF_X1 port map( D => n5840, CK => CLK, Q => 
                           n20013, QN => n8965);
   REGISTERS_reg_19_11_inst : DFF_X1 port map( D => n5839, CK => CLK, Q => 
                           n20014, QN => n8967);
   REGISTERS_reg_19_10_inst : DFF_X1 port map( D => n5838, CK => CLK, Q => 
                           n20015, QN => n8969);
   REGISTERS_reg_19_9_inst : DFF_X1 port map( D => n5837, CK => CLK, Q => 
                           n20016, QN => n8971);
   REGISTERS_reg_19_8_inst : DFF_X1 port map( D => n5836, CK => CLK, Q => 
                           n20017, QN => n8973);
   REGISTERS_reg_19_7_inst : DFF_X1 port map( D => n5835, CK => CLK, Q => 
                           n20018, QN => n8975);
   REGISTERS_reg_19_6_inst : DFF_X1 port map( D => n5834, CK => CLK, Q => 
                           n20019, QN => n8977);
   REGISTERS_reg_19_5_inst : DFF_X1 port map( D => n5833, CK => CLK, Q => 
                           n20020, QN => n8979);
   REGISTERS_reg_19_4_inst : DFF_X1 port map( D => n5832, CK => CLK, Q => 
                           n20021, QN => n8981);
   REGISTERS_reg_19_3_inst : DFF_X1 port map( D => n5831, CK => CLK, Q => 
                           n20022, QN => n8983);
   REGISTERS_reg_19_2_inst : DFF_X1 port map( D => n5830, CK => CLK, Q => 
                           n20023, QN => n8985);
   REGISTERS_reg_19_1_inst : DFF_X1 port map( D => n5829, CK => CLK, Q => 
                           n20024, QN => n8987);
   REGISTERS_reg_19_0_inst : DFF_X1 port map( D => n5828, CK => CLK, Q => 
                           n20025, QN => n8989);
   REGISTERS_reg_15_23_inst : DFF_X1 port map( D => n6107, CK => CLK, Q => 
                           n20050, QN => n7380);
   REGISTERS_reg_15_22_inst : DFF_X1 port map( D => n6106, CK => CLK, Q => 
                           n20051, QN => n7382);
   REGISTERS_reg_15_21_inst : DFF_X1 port map( D => n6105, CK => CLK, Q => 
                           n20052, QN => n7384);
   REGISTERS_reg_15_20_inst : DFF_X1 port map( D => n6104, CK => CLK, Q => 
                           n20053, QN => n7386);
   REGISTERS_reg_15_19_inst : DFF_X1 port map( D => n6103, CK => CLK, Q => 
                           n20054, QN => n7388);
   REGISTERS_reg_15_18_inst : DFF_X1 port map( D => n6102, CK => CLK, Q => 
                           n20055, QN => n7390);
   REGISTERS_reg_15_17_inst : DFF_X1 port map( D => n6101, CK => CLK, Q => 
                           n20056, QN => n7392);
   REGISTERS_reg_15_16_inst : DFF_X1 port map( D => n6100, CK => CLK, Q => 
                           n20057, QN => n7394);
   REGISTERS_reg_15_15_inst : DFF_X1 port map( D => n6099, CK => CLK, Q => 
                           n20058, QN => n7396);
   REGISTERS_reg_15_14_inst : DFF_X1 port map( D => n6098, CK => CLK, Q => 
                           n20059, QN => n7398);
   REGISTERS_reg_15_13_inst : DFF_X1 port map( D => n6097, CK => CLK, Q => 
                           n20060, QN => n7400);
   REGISTERS_reg_15_12_inst : DFF_X1 port map( D => n6096, CK => CLK, Q => 
                           n20061, QN => n7402);
   REGISTERS_reg_15_11_inst : DFF_X1 port map( D => n6095, CK => CLK, Q => 
                           n20062, QN => n7404);
   REGISTERS_reg_15_10_inst : DFF_X1 port map( D => n6094, CK => CLK, Q => 
                           n20063, QN => n7406);
   REGISTERS_reg_15_9_inst : DFF_X1 port map( D => n6093, CK => CLK, Q => 
                           n20064, QN => n7408);
   REGISTERS_reg_15_8_inst : DFF_X1 port map( D => n6092, CK => CLK, Q => 
                           n20065, QN => n7410);
   REGISTERS_reg_15_7_inst : DFF_X1 port map( D => n6091, CK => CLK, Q => 
                           n20066, QN => n7412);
   REGISTERS_reg_15_6_inst : DFF_X1 port map( D => n6090, CK => CLK, Q => 
                           n20067, QN => n7414);
   REGISTERS_reg_15_5_inst : DFF_X1 port map( D => n6089, CK => CLK, Q => 
                           n20068, QN => n7416);
   REGISTERS_reg_15_4_inst : DFF_X1 port map( D => n6088, CK => CLK, Q => 
                           n20069, QN => n7418);
   REGISTERS_reg_15_3_inst : DFF_X1 port map( D => n6087, CK => CLK, Q => 
                           n20070, QN => n7420);
   REGISTERS_reg_15_2_inst : DFF_X1 port map( D => n6086, CK => CLK, Q => 
                           n20071, QN => n7422);
   REGISTERS_reg_15_1_inst : DFF_X1 port map( D => n6085, CK => CLK, Q => 
                           n20072, QN => n7424);
   REGISTERS_reg_15_0_inst : DFF_X1 port map( D => n6084, CK => CLK, Q => 
                           n20073, QN => n7426);
   REGISTERS_reg_10_23_inst : DFF_X1 port map( D => n6427, CK => CLK, Q => 
                           n24171, QN => n7508);
   REGISTERS_reg_10_22_inst : DFF_X1 port map( D => n6426, CK => CLK, Q => 
                           n24170, QN => n7510);
   REGISTERS_reg_10_21_inst : DFF_X1 port map( D => n6425, CK => CLK, Q => 
                           n24169, QN => n7512);
   REGISTERS_reg_10_20_inst : DFF_X1 port map( D => n6424, CK => CLK, Q => 
                           n24168, QN => n7514);
   REGISTERS_reg_10_19_inst : DFF_X1 port map( D => n6423, CK => CLK, Q => 
                           n24167, QN => n7516);
   REGISTERS_reg_10_18_inst : DFF_X1 port map( D => n6422, CK => CLK, Q => 
                           n24166, QN => n7518);
   REGISTERS_reg_10_17_inst : DFF_X1 port map( D => n6421, CK => CLK, Q => 
                           n24165, QN => n7520);
   REGISTERS_reg_10_16_inst : DFF_X1 port map( D => n6420, CK => CLK, Q => 
                           n24164, QN => n7522);
   REGISTERS_reg_10_15_inst : DFF_X1 port map( D => n6419, CK => CLK, Q => 
                           n24163, QN => n7524);
   REGISTERS_reg_10_14_inst : DFF_X1 port map( D => n6418, CK => CLK, Q => 
                           n24162, QN => n7526);
   REGISTERS_reg_10_13_inst : DFF_X1 port map( D => n6417, CK => CLK, Q => 
                           n24161, QN => n7528);
   REGISTERS_reg_10_12_inst : DFF_X1 port map( D => n6416, CK => CLK, Q => 
                           n24160, QN => n7530);
   REGISTERS_reg_10_11_inst : DFF_X1 port map( D => n6415, CK => CLK, Q => 
                           n24159, QN => n7532);
   REGISTERS_reg_10_10_inst : DFF_X1 port map( D => n6414, CK => CLK, Q => 
                           n24158, QN => n7534);
   REGISTERS_reg_10_9_inst : DFF_X1 port map( D => n6413, CK => CLK, Q => 
                           n24157, QN => n7536);
   REGISTERS_reg_10_8_inst : DFF_X1 port map( D => n6412, CK => CLK, Q => 
                           n24156, QN => n7538);
   REGISTERS_reg_10_7_inst : DFF_X1 port map( D => n6411, CK => CLK, Q => 
                           n24155, QN => n7540);
   REGISTERS_reg_10_6_inst : DFF_X1 port map( D => n6410, CK => CLK, Q => 
                           n24154, QN => n7542);
   REGISTERS_reg_10_5_inst : DFF_X1 port map( D => n6409, CK => CLK, Q => 
                           n24153, QN => n7544);
   REGISTERS_reg_10_4_inst : DFF_X1 port map( D => n6408, CK => CLK, Q => 
                           n24152, QN => n7546);
   REGISTERS_reg_10_3_inst : DFF_X1 port map( D => n6407, CK => CLK, Q => 
                           n24151, QN => n7548);
   REGISTERS_reg_10_2_inst : DFF_X1 port map( D => n6406, CK => CLK, Q => 
                           n24150, QN => n7550);
   REGISTERS_reg_10_1_inst : DFF_X1 port map( D => n6405, CK => CLK, Q => 
                           n24149, QN => n7552);
   REGISTERS_reg_10_0_inst : DFF_X1 port map( D => n6404, CK => CLK, Q => 
                           n24148, QN => n7554);
   REGISTERS_reg_5_23_inst : DFF_X1 port map( D => n6747, CK => CLK, Q => 
                           n24235, QN => n17341);
   REGISTERS_reg_5_22_inst : DFF_X1 port map( D => n6746, CK => CLK, Q => 
                           n24234, QN => n17344);
   REGISTERS_reg_5_21_inst : DFF_X1 port map( D => n6745, CK => CLK, Q => 
                           n24233, QN => n17347);
   REGISTERS_reg_5_20_inst : DFF_X1 port map( D => n6744, CK => CLK, Q => 
                           n24232, QN => n17350);
   REGISTERS_reg_5_19_inst : DFF_X1 port map( D => n6743, CK => CLK, Q => 
                           n24231, QN => n17353);
   REGISTERS_reg_5_18_inst : DFF_X1 port map( D => n6742, CK => CLK, Q => 
                           n24230, QN => n17356);
   REGISTERS_reg_5_17_inst : DFF_X1 port map( D => n6741, CK => CLK, Q => 
                           n24229, QN => n17359);
   REGISTERS_reg_5_16_inst : DFF_X1 port map( D => n6740, CK => CLK, Q => 
                           n24228, QN => n17362);
   REGISTERS_reg_5_15_inst : DFF_X1 port map( D => n6739, CK => CLK, Q => 
                           n24227, QN => n17365);
   REGISTERS_reg_5_14_inst : DFF_X1 port map( D => n6738, CK => CLK, Q => 
                           n24226, QN => n17368);
   REGISTERS_reg_5_13_inst : DFF_X1 port map( D => n6737, CK => CLK, Q => 
                           n24225, QN => n17371);
   REGISTERS_reg_5_12_inst : DFF_X1 port map( D => n6736, CK => CLK, Q => 
                           n24224, QN => n17374);
   REGISTERS_reg_5_11_inst : DFF_X1 port map( D => n6735, CK => CLK, Q => 
                           n24223, QN => n17377);
   REGISTERS_reg_5_10_inst : DFF_X1 port map( D => n6734, CK => CLK, Q => 
                           n24222, QN => n17380);
   REGISTERS_reg_5_9_inst : DFF_X1 port map( D => n6733, CK => CLK, Q => n24221
                           , QN => n17383);
   REGISTERS_reg_5_8_inst : DFF_X1 port map( D => n6732, CK => CLK, Q => n24220
                           , QN => n17386);
   REGISTERS_reg_5_7_inst : DFF_X1 port map( D => n6731, CK => CLK, Q => n24219
                           , QN => n17389);
   REGISTERS_reg_5_6_inst : DFF_X1 port map( D => n6730, CK => CLK, Q => n24218
                           , QN => n17392);
   REGISTERS_reg_5_5_inst : DFF_X1 port map( D => n6729, CK => CLK, Q => n24217
                           , QN => n17395);
   REGISTERS_reg_5_4_inst : DFF_X1 port map( D => n6728, CK => CLK, Q => n24216
                           , QN => n17398);
   REGISTERS_reg_5_3_inst : DFF_X1 port map( D => n6727, CK => CLK, Q => n24215
                           , QN => n17401);
   REGISTERS_reg_5_2_inst : DFF_X1 port map( D => n6726, CK => CLK, Q => n24214
                           , QN => n17404);
   REGISTERS_reg_5_1_inst : DFF_X1 port map( D => n6725, CK => CLK, Q => n24213
                           , QN => n17407);
   REGISTERS_reg_5_0_inst : DFF_X1 port map( D => n6724, CK => CLK, Q => n24212
                           , QN => n17410);
   REGISTERS_reg_1_51_inst : DFF_X1 port map( D => n7031, CK => CLK, Q => 
                           n20122, QN => n77);
   REGISTERS_reg_1_50_inst : DFF_X1 port map( D => n7030, CK => CLK, Q => 
                           n20123, QN => n78);
   REGISTERS_reg_1_49_inst : DFF_X1 port map( D => n7029, CK => CLK, Q => 
                           n20124, QN => n79);
   REGISTERS_reg_1_48_inst : DFF_X1 port map( D => n7028, CK => CLK, Q => 
                           n20125, QN => n80);
   REGISTERS_reg_1_47_inst : DFF_X1 port map( D => n7027, CK => CLK, Q => 
                           n20126, QN => n81);
   REGISTERS_reg_1_46_inst : DFF_X1 port map( D => n7026, CK => CLK, Q => 
                           n20127, QN => n82);
   REGISTERS_reg_1_45_inst : DFF_X1 port map( D => n7025, CK => CLK, Q => 
                           n20128, QN => n83);
   REGISTERS_reg_1_44_inst : DFF_X1 port map( D => n7024, CK => CLK, Q => 
                           n20129, QN => n84);
   REGISTERS_reg_1_43_inst : DFF_X1 port map( D => n7023, CK => CLK, Q => 
                           n20130, QN => n85);
   REGISTERS_reg_1_41_inst : DFF_X1 port map( D => n7021, CK => CLK, Q => 
                           n20131, QN => n87);
   REGISTERS_reg_1_39_inst : DFF_X1 port map( D => n7019, CK => CLK, Q => 
                           n20132, QN => n89);
   REGISTERS_reg_1_35_inst : DFF_X1 port map( D => n7015, CK => CLK, Q => 
                           n20133, QN => n93);
   REGISTERS_reg_1_42_inst : DFF_X1 port map( D => n7022, CK => CLK, Q => 
                           n20134, QN => n86);
   REGISTERS_reg_1_40_inst : DFF_X1 port map( D => n7020, CK => CLK, Q => 
                           n20135, QN => n88);
   REGISTERS_reg_1_38_inst : DFF_X1 port map( D => n7018, CK => CLK, Q => 
                           n20136, QN => n90);
   REGISTERS_reg_1_37_inst : DFF_X1 port map( D => n7017, CK => CLK, Q => 
                           n20137, QN => n91);
   REGISTERS_reg_1_36_inst : DFF_X1 port map( D => n7016, CK => CLK, Q => 
                           n20138, QN => n92);
   REGISTERS_reg_1_34_inst : DFF_X1 port map( D => n7014, CK => CLK, Q => 
                           n20139, QN => n94);
   REGISTERS_reg_1_33_inst : DFF_X1 port map( D => n7013, CK => CLK, Q => 
                           n20140, QN => n95);
   REGISTERS_reg_1_32_inst : DFF_X1 port map( D => n7012, CK => CLK, Q => 
                           n20141, QN => n96);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n7011, CK => CLK, Q => 
                           n20142, QN => n97);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n7010, CK => CLK, Q => 
                           n20143, QN => n98);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n7009, CK => CLK, Q => 
                           n20144, QN => n99);
   REGISTERS_reg_23_63_inst : DFF_X1 port map( D => n5635, CK => CLK, Q => 
                           n20153, QN => n9119);
   REGISTERS_reg_23_62_inst : DFF_X1 port map( D => n5634, CK => CLK, Q => 
                           n20154, QN => n9121);
   REGISTERS_reg_23_61_inst : DFF_X1 port map( D => n5633, CK => CLK, Q => 
                           n20155, QN => n9123);
   REGISTERS_reg_23_60_inst : DFF_X1 port map( D => n5632, CK => CLK, Q => 
                           n20156, QN => n9125);
   U18613 : NAND3_X1 port map( A1 => n19192, A2 => n19191, A3 => n21269, ZN => 
                           n21253);
   U18614 : NAND3_X1 port map( A1 => n21269, A2 => n19191, A3 => ADD_WR(3), ZN 
                           => n21271);
   U18615 : NAND3_X1 port map( A1 => n21269, A2 => n19192, A3 => ADD_WR(4), ZN 
                           => n21280);
   U18616 : NAND3_X1 port map( A1 => n19194, A2 => n19193, A3 => n19195, ZN => 
                           n21254);
   U18617 : NAND3_X1 port map( A1 => n19194, A2 => n19193, A3 => ADD_WR(0), ZN 
                           => n21256);
   U18618 : NAND3_X1 port map( A1 => n19195, A2 => n19193, A3 => ADD_WR(1), ZN 
                           => n21258);
   U18619 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n19193, A3 => ADD_WR(1), 
                           ZN => n21260);
   U18620 : NAND3_X1 port map( A1 => n19195, A2 => n19194, A3 => ADD_WR(2), ZN 
                           => n21262);
   U18621 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n19194, A3 => ADD_WR(2), 
                           ZN => n21264);
   U18622 : NAND3_X1 port map( A1 => ADD_WR(1), A2 => n19195, A3 => ADD_WR(2), 
                           ZN => n21266);
   U18623 : NAND3_X1 port map( A1 => ADD_WR(3), A2 => n21269, A3 => ADD_WR(4), 
                           ZN => n21289);
   U18624 : NAND3_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(0), A3 => 
                           ADD_WR(2), ZN => n21268);
   REGISTERS_reg_22_63_inst : DFF_X1 port map( D => n5699, CK => CLK, Q => 
                           n19524, QN => n7429);
   REGISTERS_reg_22_62_inst : DFF_X1 port map( D => n5698, CK => CLK, Q => 
                           n19525, QN => n7431);
   REGISTERS_reg_22_61_inst : DFF_X1 port map( D => n5697, CK => CLK, Q => 
                           n19526, QN => n7433);
   REGISTERS_reg_22_60_inst : DFF_X1 port map( D => n5696, CK => CLK, Q => 
                           n19527, QN => n7435);
   REGISTERS_reg_18_63_inst : DFF_X1 port map( D => n5955, CK => CLK, Q => 
                           n19806, QN => n8735);
   REGISTERS_reg_18_62_inst : DFF_X1 port map( D => n5954, CK => CLK, Q => 
                           n19807, QN => n8737);
   REGISTERS_reg_18_61_inst : DFF_X1 port map( D => n5953, CK => CLK, Q => 
                           n19808, QN => n8739);
   REGISTERS_reg_18_60_inst : DFF_X1 port map( D => n5952, CK => CLK, Q => 
                           n19809, QN => n8741);
   REGISTERS_reg_14_63_inst : DFF_X1 port map( D => n6211, CK => CLK, Q => 
                           n19460, QN => n8990);
   REGISTERS_reg_14_62_inst : DFF_X1 port map( D => n6210, CK => CLK, Q => 
                           n19461, QN => n8992);
   REGISTERS_reg_14_61_inst : DFF_X1 port map( D => n6209, CK => CLK, Q => 
                           n19462, QN => n8994);
   REGISTERS_reg_14_60_inst : DFF_X1 port map( D => n6208, CK => CLK, Q => 
                           n19463, QN => n8996);
   REGISTERS_reg_22_59_inst : DFF_X1 port map( D => n5695, CK => CLK, Q => 
                           n19528, QN => n7437);
   REGISTERS_reg_22_58_inst : DFF_X1 port map( D => n5694, CK => CLK, Q => 
                           n19529, QN => n7439);
   REGISTERS_reg_22_57_inst : DFF_X1 port map( D => n5693, CK => CLK, Q => 
                           n19530, QN => n7441);
   REGISTERS_reg_22_56_inst : DFF_X1 port map( D => n5692, CK => CLK, Q => 
                           n19531, QN => n7443);
   REGISTERS_reg_22_55_inst : DFF_X1 port map( D => n5691, CK => CLK, Q => 
                           n19532, QN => n7445);
   REGISTERS_reg_22_54_inst : DFF_X1 port map( D => n5690, CK => CLK, Q => 
                           n19533, QN => n7447);
   REGISTERS_reg_22_53_inst : DFF_X1 port map( D => n5689, CK => CLK, Q => 
                           n19534, QN => n7449);
   REGISTERS_reg_22_52_inst : DFF_X1 port map( D => n5688, CK => CLK, Q => 
                           n19535, QN => n7451);
   REGISTERS_reg_22_51_inst : DFF_X1 port map( D => n5687, CK => CLK, Q => 
                           n19536, QN => n7453);
   REGISTERS_reg_22_50_inst : DFF_X1 port map( D => n5686, CK => CLK, Q => 
                           n19537, QN => n7455);
   REGISTERS_reg_22_49_inst : DFF_X1 port map( D => n5685, CK => CLK, Q => 
                           n19538, QN => n7457);
   REGISTERS_reg_22_48_inst : DFF_X1 port map( D => n5684, CK => CLK, Q => 
                           n19539, QN => n7459);
   REGISTERS_reg_22_47_inst : DFF_X1 port map( D => n5683, CK => CLK, Q => 
                           n19540, QN => n7461);
   REGISTERS_reg_22_46_inst : DFF_X1 port map( D => n5682, CK => CLK, Q => 
                           n19541, QN => n7463);
   REGISTERS_reg_22_45_inst : DFF_X1 port map( D => n5681, CK => CLK, Q => 
                           n19542, QN => n7465);
   REGISTERS_reg_22_44_inst : DFF_X1 port map( D => n5680, CK => CLK, Q => 
                           n19543, QN => n7467);
   REGISTERS_reg_22_43_inst : DFF_X1 port map( D => n5679, CK => CLK, Q => 
                           n19544, QN => n7469);
   REGISTERS_reg_22_42_inst : DFF_X1 port map( D => n5678, CK => CLK, Q => 
                           n19545, QN => n7471);
   REGISTERS_reg_22_41_inst : DFF_X1 port map( D => n5677, CK => CLK, Q => 
                           n19546, QN => n7473);
   REGISTERS_reg_22_40_inst : DFF_X1 port map( D => n5676, CK => CLK, Q => 
                           n19547, QN => n7475);
   REGISTERS_reg_22_39_inst : DFF_X1 port map( D => n5675, CK => CLK, Q => 
                           n19548, QN => n7477);
   REGISTERS_reg_22_38_inst : DFF_X1 port map( D => n5674, CK => CLK, Q => 
                           n19549, QN => n7479);
   REGISTERS_reg_22_37_inst : DFF_X1 port map( D => n5673, CK => CLK, Q => 
                           n19550, QN => n7481);
   REGISTERS_reg_22_36_inst : DFF_X1 port map( D => n5672, CK => CLK, Q => 
                           n19551, QN => n7483);
   REGISTERS_reg_22_35_inst : DFF_X1 port map( D => n5671, CK => CLK, Q => 
                           n19552, QN => n7485);
   REGISTERS_reg_22_34_inst : DFF_X1 port map( D => n5670, CK => CLK, Q => 
                           n19553, QN => n7487);
   REGISTERS_reg_22_33_inst : DFF_X1 port map( D => n5669, CK => CLK, Q => 
                           n19554, QN => n7489);
   REGISTERS_reg_22_32_inst : DFF_X1 port map( D => n5668, CK => CLK, Q => 
                           n19555, QN => n7491);
   REGISTERS_reg_22_31_inst : DFF_X1 port map( D => n5667, CK => CLK, Q => 
                           n19556, QN => n7493);
   REGISTERS_reg_22_30_inst : DFF_X1 port map( D => n5666, CK => CLK, Q => 
                           n19557, QN => n7495);
   REGISTERS_reg_22_29_inst : DFF_X1 port map( D => n5665, CK => CLK, Q => 
                           n19558, QN => n7497);
   REGISTERS_reg_22_28_inst : DFF_X1 port map( D => n5664, CK => CLK, Q => 
                           n19559, QN => n7499);
   REGISTERS_reg_22_27_inst : DFF_X1 port map( D => n5663, CK => CLK, Q => 
                           n19560, QN => n7501);
   REGISTERS_reg_22_26_inst : DFF_X1 port map( D => n5662, CK => CLK, Q => 
                           n19561, QN => n7503);
   REGISTERS_reg_22_25_inst : DFF_X1 port map( D => n5661, CK => CLK, Q => 
                           n19562, QN => n7505);
   REGISTERS_reg_22_24_inst : DFF_X1 port map( D => n5660, CK => CLK, Q => 
                           n19563, QN => n7507);
   REGISTERS_reg_18_59_inst : DFF_X1 port map( D => n5951, CK => CLK, Q => 
                           n19858, QN => n8743);
   REGISTERS_reg_18_58_inst : DFF_X1 port map( D => n5950, CK => CLK, Q => 
                           n19859, QN => n8745);
   REGISTERS_reg_18_57_inst : DFF_X1 port map( D => n5949, CK => CLK, Q => 
                           n19860, QN => n8747);
   REGISTERS_reg_18_56_inst : DFF_X1 port map( D => n5948, CK => CLK, Q => 
                           n19861, QN => n8749);
   REGISTERS_reg_18_55_inst : DFF_X1 port map( D => n5947, CK => CLK, Q => 
                           n19862, QN => n8751);
   REGISTERS_reg_18_54_inst : DFF_X1 port map( D => n5946, CK => CLK, Q => 
                           n19863, QN => n8753);
   REGISTERS_reg_18_53_inst : DFF_X1 port map( D => n5945, CK => CLK, Q => 
                           n19864, QN => n8755);
   REGISTERS_reg_18_52_inst : DFF_X1 port map( D => n5944, CK => CLK, Q => 
                           n19865, QN => n8757);
   REGISTERS_reg_18_51_inst : DFF_X1 port map( D => n5943, CK => CLK, Q => 
                           n19866, QN => n8759);
   REGISTERS_reg_18_50_inst : DFF_X1 port map( D => n5942, CK => CLK, Q => 
                           n19867, QN => n8761);
   REGISTERS_reg_18_49_inst : DFF_X1 port map( D => n5941, CK => CLK, Q => 
                           n19868, QN => n8763);
   REGISTERS_reg_18_48_inst : DFF_X1 port map( D => n5940, CK => CLK, Q => 
                           n19869, QN => n8765);
   REGISTERS_reg_18_47_inst : DFF_X1 port map( D => n5939, CK => CLK, Q => 
                           n19870, QN => n8767);
   REGISTERS_reg_18_46_inst : DFF_X1 port map( D => n5938, CK => CLK, Q => 
                           n19871, QN => n8769);
   REGISTERS_reg_18_45_inst : DFF_X1 port map( D => n5937, CK => CLK, Q => 
                           n19872, QN => n8771);
   REGISTERS_reg_18_44_inst : DFF_X1 port map( D => n5936, CK => CLK, Q => 
                           n19873, QN => n8773);
   REGISTERS_reg_18_43_inst : DFF_X1 port map( D => n5935, CK => CLK, Q => 
                           n19874, QN => n8775);
   REGISTERS_reg_18_42_inst : DFF_X1 port map( D => n5934, CK => CLK, Q => 
                           n19875, QN => n8777);
   REGISTERS_reg_18_41_inst : DFF_X1 port map( D => n5933, CK => CLK, Q => 
                           n19876, QN => n8779);
   REGISTERS_reg_18_40_inst : DFF_X1 port map( D => n5932, CK => CLK, Q => 
                           n19877, QN => n8781);
   REGISTERS_reg_18_39_inst : DFF_X1 port map( D => n5931, CK => CLK, Q => 
                           n19878, QN => n8783);
   REGISTERS_reg_18_38_inst : DFF_X1 port map( D => n5930, CK => CLK, Q => 
                           n19879, QN => n8785);
   REGISTERS_reg_18_37_inst : DFF_X1 port map( D => n5929, CK => CLK, Q => 
                           n19880, QN => n8787);
   REGISTERS_reg_18_36_inst : DFF_X1 port map( D => n5928, CK => CLK, Q => 
                           n19881, QN => n8789);
   REGISTERS_reg_18_35_inst : DFF_X1 port map( D => n5927, CK => CLK, Q => 
                           n19882, QN => n8791);
   REGISTERS_reg_18_34_inst : DFF_X1 port map( D => n5926, CK => CLK, Q => 
                           n19883, QN => n8793);
   REGISTERS_reg_18_33_inst : DFF_X1 port map( D => n5925, CK => CLK, Q => 
                           n19884, QN => n8795);
   REGISTERS_reg_18_32_inst : DFF_X1 port map( D => n5924, CK => CLK, Q => 
                           n19885, QN => n8797);
   REGISTERS_reg_18_31_inst : DFF_X1 port map( D => n5923, CK => CLK, Q => 
                           n19886, QN => n8799);
   REGISTERS_reg_18_30_inst : DFF_X1 port map( D => n5922, CK => CLK, Q => 
                           n19887, QN => n8801);
   REGISTERS_reg_18_29_inst : DFF_X1 port map( D => n5921, CK => CLK, Q => 
                           n19888, QN => n8803);
   REGISTERS_reg_18_28_inst : DFF_X1 port map( D => n5920, CK => CLK, Q => 
                           n19889, QN => n8805);
   REGISTERS_reg_18_27_inst : DFF_X1 port map( D => n5919, CK => CLK, Q => 
                           n19890, QN => n8807);
   REGISTERS_reg_18_26_inst : DFF_X1 port map( D => n5918, CK => CLK, Q => 
                           n19891, QN => n8809);
   REGISTERS_reg_18_25_inst : DFF_X1 port map( D => n5917, CK => CLK, Q => 
                           n19892, QN => n8811);
   REGISTERS_reg_18_24_inst : DFF_X1 port map( D => n5916, CK => CLK, Q => 
                           n19893, QN => n8813);
   REGISTERS_reg_14_59_inst : DFF_X1 port map( D => n6207, CK => CLK, Q => 
                           n19464, QN => n8998);
   REGISTERS_reg_14_58_inst : DFF_X1 port map( D => n6206, CK => CLK, Q => 
                           n19465, QN => n9000);
   REGISTERS_reg_14_57_inst : DFF_X1 port map( D => n6205, CK => CLK, Q => 
                           n19466, QN => n9002);
   REGISTERS_reg_14_56_inst : DFF_X1 port map( D => n6204, CK => CLK, Q => 
                           n19467, QN => n9004);
   REGISTERS_reg_14_55_inst : DFF_X1 port map( D => n6203, CK => CLK, Q => 
                           n19468, QN => n9006);
   REGISTERS_reg_14_54_inst : DFF_X1 port map( D => n6202, CK => CLK, Q => 
                           n19469, QN => n9008);
   REGISTERS_reg_14_53_inst : DFF_X1 port map( D => n6201, CK => CLK, Q => 
                           n19470, QN => n9010);
   REGISTERS_reg_14_52_inst : DFF_X1 port map( D => n6200, CK => CLK, Q => 
                           n19471, QN => n9012);
   REGISTERS_reg_14_51_inst : DFF_X1 port map( D => n6199, CK => CLK, Q => 
                           n19472, QN => n9014);
   REGISTERS_reg_14_50_inst : DFF_X1 port map( D => n6198, CK => CLK, Q => 
                           n19473, QN => n9016);
   REGISTERS_reg_14_49_inst : DFF_X1 port map( D => n6197, CK => CLK, Q => 
                           n19474, QN => n9018);
   REGISTERS_reg_14_48_inst : DFF_X1 port map( D => n6196, CK => CLK, Q => 
                           n19475, QN => n9020);
   REGISTERS_reg_14_47_inst : DFF_X1 port map( D => n6195, CK => CLK, Q => 
                           n19476, QN => n9022);
   REGISTERS_reg_14_46_inst : DFF_X1 port map( D => n6194, CK => CLK, Q => 
                           n19477, QN => n9024);
   REGISTERS_reg_14_45_inst : DFF_X1 port map( D => n6193, CK => CLK, Q => 
                           n19478, QN => n9026);
   REGISTERS_reg_14_44_inst : DFF_X1 port map( D => n6192, CK => CLK, Q => 
                           n19479, QN => n9028);
   REGISTERS_reg_14_43_inst : DFF_X1 port map( D => n6191, CK => CLK, Q => 
                           n19480, QN => n9030);
   REGISTERS_reg_14_42_inst : DFF_X1 port map( D => n6190, CK => CLK, Q => 
                           n19481, QN => n9032);
   REGISTERS_reg_14_41_inst : DFF_X1 port map( D => n6189, CK => CLK, Q => 
                           n19482, QN => n9034);
   REGISTERS_reg_14_40_inst : DFF_X1 port map( D => n6188, CK => CLK, Q => 
                           n19483, QN => n9036);
   REGISTERS_reg_14_39_inst : DFF_X1 port map( D => n6187, CK => CLK, Q => 
                           n19484, QN => n9038);
   REGISTERS_reg_14_38_inst : DFF_X1 port map( D => n6186, CK => CLK, Q => 
                           n19485, QN => n9040);
   REGISTERS_reg_14_37_inst : DFF_X1 port map( D => n6185, CK => CLK, Q => 
                           n19486, QN => n9042);
   REGISTERS_reg_14_36_inst : DFF_X1 port map( D => n6184, CK => CLK, Q => 
                           n19487, QN => n9044);
   REGISTERS_reg_14_35_inst : DFF_X1 port map( D => n6183, CK => CLK, Q => 
                           n19488, QN => n9046);
   REGISTERS_reg_14_34_inst : DFF_X1 port map( D => n6182, CK => CLK, Q => 
                           n19489, QN => n9048);
   REGISTERS_reg_14_33_inst : DFF_X1 port map( D => n6181, CK => CLK, Q => 
                           n19490, QN => n9050);
   REGISTERS_reg_14_32_inst : DFF_X1 port map( D => n6180, CK => CLK, Q => 
                           n19491, QN => n9052);
   REGISTERS_reg_14_31_inst : DFF_X1 port map( D => n6179, CK => CLK, Q => 
                           n19492, QN => n9054);
   REGISTERS_reg_14_30_inst : DFF_X1 port map( D => n6178, CK => CLK, Q => 
                           n19493, QN => n9056);
   REGISTERS_reg_14_29_inst : DFF_X1 port map( D => n6177, CK => CLK, Q => 
                           n19494, QN => n9058);
   REGISTERS_reg_14_28_inst : DFF_X1 port map( D => n6176, CK => CLK, Q => 
                           n19495, QN => n9060);
   REGISTERS_reg_14_27_inst : DFF_X1 port map( D => n6175, CK => CLK, Q => 
                           n19496, QN => n9062);
   REGISTERS_reg_14_26_inst : DFF_X1 port map( D => n6174, CK => CLK, Q => 
                           n19497, QN => n9064);
   REGISTERS_reg_14_25_inst : DFF_X1 port map( D => n6173, CK => CLK, Q => 
                           n19498, QN => n9066);
   REGISTERS_reg_14_24_inst : DFF_X1 port map( D => n6172, CK => CLK, Q => 
                           n19499, QN => n9068);
   REGISTERS_reg_22_23_inst : DFF_X1 port map( D => n5659, CK => CLK, Q => 
                           n19564, QN => n7509);
   REGISTERS_reg_22_22_inst : DFF_X1 port map( D => n5658, CK => CLK, Q => 
                           n19565, QN => n7511);
   REGISTERS_reg_22_21_inst : DFF_X1 port map( D => n5657, CK => CLK, Q => 
                           n19566, QN => n7513);
   REGISTERS_reg_22_20_inst : DFF_X1 port map( D => n5656, CK => CLK, Q => 
                           n19567, QN => n7515);
   REGISTERS_reg_22_19_inst : DFF_X1 port map( D => n5655, CK => CLK, Q => 
                           n19568, QN => n7517);
   REGISTERS_reg_22_18_inst : DFF_X1 port map( D => n5654, CK => CLK, Q => 
                           n19569, QN => n7519);
   REGISTERS_reg_22_17_inst : DFF_X1 port map( D => n5653, CK => CLK, Q => 
                           n19570, QN => n7521);
   REGISTERS_reg_22_16_inst : DFF_X1 port map( D => n5652, CK => CLK, Q => 
                           n19571, QN => n7523);
   REGISTERS_reg_22_15_inst : DFF_X1 port map( D => n5651, CK => CLK, Q => 
                           n19572, QN => n7525);
   REGISTERS_reg_22_14_inst : DFF_X1 port map( D => n5650, CK => CLK, Q => 
                           n19573, QN => n7527);
   REGISTERS_reg_22_13_inst : DFF_X1 port map( D => n5649, CK => CLK, Q => 
                           n19574, QN => n7529);
   REGISTERS_reg_22_12_inst : DFF_X1 port map( D => n5648, CK => CLK, Q => 
                           n19575, QN => n7531);
   REGISTERS_reg_22_11_inst : DFF_X1 port map( D => n5647, CK => CLK, Q => 
                           n19576, QN => n7533);
   REGISTERS_reg_22_10_inst : DFF_X1 port map( D => n5646, CK => CLK, Q => 
                           n19577, QN => n7535);
   REGISTERS_reg_22_9_inst : DFF_X1 port map( D => n5645, CK => CLK, Q => 
                           n19578, QN => n7537);
   REGISTERS_reg_22_8_inst : DFF_X1 port map( D => n5644, CK => CLK, Q => 
                           n19579, QN => n7539);
   REGISTERS_reg_22_7_inst : DFF_X1 port map( D => n5643, CK => CLK, Q => 
                           n19580, QN => n7541);
   REGISTERS_reg_22_6_inst : DFF_X1 port map( D => n5642, CK => CLK, Q => 
                           n19581, QN => n7543);
   REGISTERS_reg_22_5_inst : DFF_X1 port map( D => n5641, CK => CLK, Q => 
                           n19582, QN => n7545);
   REGISTERS_reg_22_4_inst : DFF_X1 port map( D => n5640, CK => CLK, Q => 
                           n19583, QN => n7547);
   REGISTERS_reg_22_3_inst : DFF_X1 port map( D => n5639, CK => CLK, Q => 
                           n19584, QN => n7549);
   REGISTERS_reg_22_2_inst : DFF_X1 port map( D => n5638, CK => CLK, Q => 
                           n19585, QN => n7551);
   REGISTERS_reg_22_1_inst : DFF_X1 port map( D => n5637, CK => CLK, Q => 
                           n19586, QN => n7553);
   REGISTERS_reg_22_0_inst : DFF_X1 port map( D => n5636, CK => CLK, Q => 
                           n19587, QN => n7555);
   REGISTERS_reg_18_23_inst : DFF_X1 port map( D => n5915, CK => CLK, Q => 
                           n20026, QN => n8815);
   REGISTERS_reg_18_22_inst : DFF_X1 port map( D => n5914, CK => CLK, Q => 
                           n20027, QN => n8817);
   REGISTERS_reg_18_21_inst : DFF_X1 port map( D => n5913, CK => CLK, Q => 
                           n20028, QN => n8819);
   REGISTERS_reg_18_20_inst : DFF_X1 port map( D => n5912, CK => CLK, Q => 
                           n20029, QN => n8821);
   REGISTERS_reg_18_19_inst : DFF_X1 port map( D => n5911, CK => CLK, Q => 
                           n20030, QN => n8823);
   REGISTERS_reg_18_18_inst : DFF_X1 port map( D => n5910, CK => CLK, Q => 
                           n20031, QN => n8825);
   REGISTERS_reg_18_17_inst : DFF_X1 port map( D => n5909, CK => CLK, Q => 
                           n20032, QN => n8827);
   REGISTERS_reg_18_16_inst : DFF_X1 port map( D => n5908, CK => CLK, Q => 
                           n20033, QN => n8829);
   REGISTERS_reg_18_15_inst : DFF_X1 port map( D => n5907, CK => CLK, Q => 
                           n20034, QN => n8831);
   REGISTERS_reg_18_14_inst : DFF_X1 port map( D => n5906, CK => CLK, Q => 
                           n20035, QN => n8833);
   REGISTERS_reg_18_13_inst : DFF_X1 port map( D => n5905, CK => CLK, Q => 
                           n20036, QN => n8835);
   REGISTERS_reg_18_12_inst : DFF_X1 port map( D => n5904, CK => CLK, Q => 
                           n20037, QN => n8837);
   REGISTERS_reg_18_11_inst : DFF_X1 port map( D => n5903, CK => CLK, Q => 
                           n20038, QN => n8839);
   REGISTERS_reg_18_10_inst : DFF_X1 port map( D => n5902, CK => CLK, Q => 
                           n20039, QN => n8841);
   REGISTERS_reg_18_9_inst : DFF_X1 port map( D => n5901, CK => CLK, Q => 
                           n20040, QN => n8843);
   REGISTERS_reg_18_8_inst : DFF_X1 port map( D => n5900, CK => CLK, Q => 
                           n20041, QN => n8845);
   REGISTERS_reg_18_7_inst : DFF_X1 port map( D => n5899, CK => CLK, Q => 
                           n20042, QN => n8847);
   REGISTERS_reg_18_6_inst : DFF_X1 port map( D => n5898, CK => CLK, Q => 
                           n20043, QN => n8849);
   REGISTERS_reg_18_5_inst : DFF_X1 port map( D => n5897, CK => CLK, Q => 
                           n20044, QN => n8851);
   REGISTERS_reg_18_4_inst : DFF_X1 port map( D => n5896, CK => CLK, Q => 
                           n20045, QN => n8853);
   REGISTERS_reg_18_3_inst : DFF_X1 port map( D => n5895, CK => CLK, Q => 
                           n20046, QN => n8855);
   REGISTERS_reg_18_2_inst : DFF_X1 port map( D => n5894, CK => CLK, Q => 
                           n20047, QN => n8857);
   REGISTERS_reg_18_1_inst : DFF_X1 port map( D => n5893, CK => CLK, Q => 
                           n20048, QN => n8859);
   REGISTERS_reg_18_0_inst : DFF_X1 port map( D => n5892, CK => CLK, Q => 
                           n20049, QN => n8861);
   REGISTERS_reg_14_23_inst : DFF_X1 port map( D => n6171, CK => CLK, Q => 
                           n19500, QN => n9070);
   REGISTERS_reg_14_22_inst : DFF_X1 port map( D => n6170, CK => CLK, Q => 
                           n19501, QN => n9072);
   REGISTERS_reg_14_21_inst : DFF_X1 port map( D => n6169, CK => CLK, Q => 
                           n19502, QN => n9074);
   REGISTERS_reg_14_20_inst : DFF_X1 port map( D => n6168, CK => CLK, Q => 
                           n19503, QN => n9076);
   REGISTERS_reg_14_19_inst : DFF_X1 port map( D => n6167, CK => CLK, Q => 
                           n19504, QN => n9078);
   REGISTERS_reg_14_18_inst : DFF_X1 port map( D => n6166, CK => CLK, Q => 
                           n19505, QN => n9080);
   REGISTERS_reg_14_17_inst : DFF_X1 port map( D => n6165, CK => CLK, Q => 
                           n19506, QN => n9082);
   REGISTERS_reg_14_16_inst : DFF_X1 port map( D => n6164, CK => CLK, Q => 
                           n19507, QN => n9084);
   REGISTERS_reg_14_15_inst : DFF_X1 port map( D => n6163, CK => CLK, Q => 
                           n19508, QN => n9086);
   REGISTERS_reg_14_14_inst : DFF_X1 port map( D => n6162, CK => CLK, Q => 
                           n19509, QN => n9088);
   REGISTERS_reg_14_13_inst : DFF_X1 port map( D => n6161, CK => CLK, Q => 
                           n19510, QN => n9090);
   REGISTERS_reg_14_12_inst : DFF_X1 port map( D => n6160, CK => CLK, Q => 
                           n19511, QN => n9092);
   REGISTERS_reg_14_11_inst : DFF_X1 port map( D => n6159, CK => CLK, Q => 
                           n19512, QN => n9094);
   REGISTERS_reg_14_10_inst : DFF_X1 port map( D => n6158, CK => CLK, Q => 
                           n19513, QN => n9096);
   REGISTERS_reg_14_9_inst : DFF_X1 port map( D => n6157, CK => CLK, Q => 
                           n19514, QN => n9098);
   REGISTERS_reg_14_8_inst : DFF_X1 port map( D => n6156, CK => CLK, Q => 
                           n19515, QN => n9100);
   REGISTERS_reg_14_7_inst : DFF_X1 port map( D => n6155, CK => CLK, Q => 
                           n19516, QN => n9102);
   REGISTERS_reg_14_6_inst : DFF_X1 port map( D => n6154, CK => CLK, Q => 
                           n19517, QN => n9104);
   REGISTERS_reg_14_5_inst : DFF_X1 port map( D => n6153, CK => CLK, Q => 
                           n19518, QN => n9106);
   REGISTERS_reg_14_4_inst : DFF_X1 port map( D => n6152, CK => CLK, Q => 
                           n19519, QN => n9108);
   REGISTERS_reg_14_3_inst : DFF_X1 port map( D => n6151, CK => CLK, Q => 
                           n19520, QN => n9110);
   REGISTERS_reg_14_2_inst : DFF_X1 port map( D => n6150, CK => CLK, Q => 
                           n19521, QN => n9112);
   REGISTERS_reg_14_1_inst : DFF_X1 port map( D => n6149, CK => CLK, Q => 
                           n19522, QN => n9114);
   REGISTERS_reg_14_0_inst : DFF_X1 port map( D => n6148, CK => CLK, Q => 
                           n19523, QN => n9116);
   REGISTERS_reg_25_63_inst : DFF_X1 port map( D => n5507, CK => CLK, Q => 
                           n_1167, QN => n7301);
   REGISTERS_reg_31_3_inst : DFF_X1 port map( D => n5063, CK => CLK, Q => n8282
                           , QN => n20187);
   REGISTERS_reg_31_2_inst : DFF_X1 port map( D => n5062, CK => CLK, Q => n8283
                           , QN => n20188);
   REGISTERS_reg_31_1_inst : DFF_X1 port map( D => n5061, CK => CLK, Q => n8284
                           , QN => n20189);
   REGISTERS_reg_31_0_inst : DFF_X1 port map( D => n5060, CK => CLK, Q => n8285
                           , QN => n20526);
   REGISTERS_reg_31_39_inst : DFF_X1 port map( D => n5099, CK => CLK, Q => 
                           n8246, QN => n20214);
   REGISTERS_reg_31_38_inst : DFF_X1 port map( D => n5098, CK => CLK, Q => 
                           n8247, QN => n20215);
   REGISTERS_reg_31_37_inst : DFF_X1 port map( D => n5097, CK => CLK, Q => 
                           n8248, QN => n20216);
   REGISTERS_reg_31_36_inst : DFF_X1 port map( D => n5096, CK => CLK, Q => 
                           n8249, QN => n20217);
   REGISTERS_reg_31_35_inst : DFF_X1 port map( D => n5095, CK => CLK, Q => 
                           n8250, QN => n20218);
   REGISTERS_reg_31_34_inst : DFF_X1 port map( D => n5094, CK => CLK, Q => 
                           n8251, QN => n20219);
   REGISTERS_reg_31_33_inst : DFF_X1 port map( D => n5093, CK => CLK, Q => 
                           n8252, QN => n20220);
   REGISTERS_reg_31_32_inst : DFF_X1 port map( D => n5092, CK => CLK, Q => 
                           n8253, QN => n20221);
   REGISTERS_reg_31_31_inst : DFF_X1 port map( D => n5091, CK => CLK, Q => 
                           n8254, QN => n20222);
   REGISTERS_reg_31_30_inst : DFF_X1 port map( D => n5090, CK => CLK, Q => 
                           n8255, QN => n20223);
   REGISTERS_reg_31_29_inst : DFF_X1 port map( D => n5089, CK => CLK, Q => 
                           n8256, QN => n20224);
   REGISTERS_reg_31_28_inst : DFF_X1 port map( D => n5088, CK => CLK, Q => 
                           n8257, QN => n20225);
   REGISTERS_reg_31_27_inst : DFF_X1 port map( D => n5087, CK => CLK, Q => 
                           n8258, QN => n20226);
   REGISTERS_reg_31_26_inst : DFF_X1 port map( D => n5086, CK => CLK, Q => 
                           n8259, QN => n20227);
   REGISTERS_reg_31_25_inst : DFF_X1 port map( D => n5085, CK => CLK, Q => 
                           n8260, QN => n20228);
   REGISTERS_reg_31_24_inst : DFF_X1 port map( D => n5084, CK => CLK, Q => 
                           n8261, QN => n20229);
   REGISTERS_reg_31_23_inst : DFF_X1 port map( D => n5083, CK => CLK, Q => 
                           n8262, QN => n20230);
   REGISTERS_reg_31_22_inst : DFF_X1 port map( D => n5082, CK => CLK, Q => 
                           n8263, QN => n20231);
   REGISTERS_reg_31_21_inst : DFF_X1 port map( D => n5081, CK => CLK, Q => 
                           n8264, QN => n20232);
   REGISTERS_reg_31_20_inst : DFF_X1 port map( D => n5080, CK => CLK, Q => 
                           n8265, QN => n20233);
   REGISTERS_reg_31_19_inst : DFF_X1 port map( D => n5079, CK => CLK, Q => 
                           n8266, QN => n20234);
   REGISTERS_reg_31_18_inst : DFF_X1 port map( D => n5078, CK => CLK, Q => 
                           n8267, QN => n20235);
   REGISTERS_reg_31_17_inst : DFF_X1 port map( D => n5077, CK => CLK, Q => 
                           n8268, QN => n20236);
   REGISTERS_reg_31_16_inst : DFF_X1 port map( D => n5076, CK => CLK, Q => 
                           n8269, QN => n20237);
   REGISTERS_reg_31_15_inst : DFF_X1 port map( D => n5075, CK => CLK, Q => 
                           n8270, QN => n20238);
   REGISTERS_reg_31_14_inst : DFF_X1 port map( D => n5074, CK => CLK, Q => 
                           n8271, QN => n20239);
   REGISTERS_reg_31_13_inst : DFF_X1 port map( D => n5073, CK => CLK, Q => 
                           n8272, QN => n20240);
   REGISTERS_reg_31_12_inst : DFF_X1 port map( D => n5072, CK => CLK, Q => 
                           n8273, QN => n20241);
   REGISTERS_reg_31_11_inst : DFF_X1 port map( D => n5071, CK => CLK, Q => 
                           n8274, QN => n20242);
   REGISTERS_reg_31_10_inst : DFF_X1 port map( D => n5070, CK => CLK, Q => 
                           n8275, QN => n20243);
   REGISTERS_reg_31_9_inst : DFF_X1 port map( D => n5069, CK => CLK, Q => n8276
                           , QN => n20244);
   REGISTERS_reg_31_8_inst : DFF_X1 port map( D => n5068, CK => CLK, Q => n8277
                           , QN => n20245);
   REGISTERS_reg_31_7_inst : DFF_X1 port map( D => n5067, CK => CLK, Q => n8278
                           , QN => n20246);
   REGISTERS_reg_31_6_inst : DFF_X1 port map( D => n5066, CK => CLK, Q => n8279
                           , QN => n20247);
   REGISTERS_reg_31_5_inst : DFF_X1 port map( D => n5065, CK => CLK, Q => n8280
                           , QN => n20248);
   REGISTERS_reg_31_4_inst : DFF_X1 port map( D => n5064, CK => CLK, Q => n8281
                           , QN => n20249);
   REGISTERS_reg_31_63_inst : DFF_X1 port map( D => n5123, CK => CLK, Q => 
                           n8222, QN => n20190);
   REGISTERS_reg_31_62_inst : DFF_X1 port map( D => n5122, CK => CLK, Q => 
                           n8223, QN => n20191);
   REGISTERS_reg_31_61_inst : DFF_X1 port map( D => n5121, CK => CLK, Q => 
                           n8224, QN => n20192);
   REGISTERS_reg_31_60_inst : DFF_X1 port map( D => n5120, CK => CLK, Q => 
                           n8225, QN => n20193);
   REGISTERS_reg_31_59_inst : DFF_X1 port map( D => n5119, CK => CLK, Q => 
                           n8226, QN => n20194);
   REGISTERS_reg_31_58_inst : DFF_X1 port map( D => n5118, CK => CLK, Q => 
                           n8227, QN => n20195);
   REGISTERS_reg_31_57_inst : DFF_X1 port map( D => n5117, CK => CLK, Q => 
                           n8228, QN => n20196);
   REGISTERS_reg_31_56_inst : DFF_X1 port map( D => n5116, CK => CLK, Q => 
                           n8229, QN => n20197);
   REGISTERS_reg_31_55_inst : DFF_X1 port map( D => n5115, CK => CLK, Q => 
                           n8230, QN => n20198);
   REGISTERS_reg_31_54_inst : DFF_X1 port map( D => n5114, CK => CLK, Q => 
                           n8231, QN => n20199);
   REGISTERS_reg_31_53_inst : DFF_X1 port map( D => n5113, CK => CLK, Q => 
                           n8232, QN => n20200);
   REGISTERS_reg_31_52_inst : DFF_X1 port map( D => n5112, CK => CLK, Q => 
                           n8233, QN => n20201);
   REGISTERS_reg_31_51_inst : DFF_X1 port map( D => n5111, CK => CLK, Q => 
                           n8234, QN => n20202);
   REGISTERS_reg_31_50_inst : DFF_X1 port map( D => n5110, CK => CLK, Q => 
                           n8235, QN => n20203);
   REGISTERS_reg_31_49_inst : DFF_X1 port map( D => n5109, CK => CLK, Q => 
                           n8236, QN => n20204);
   REGISTERS_reg_31_48_inst : DFF_X1 port map( D => n5108, CK => CLK, Q => 
                           n8237, QN => n20205);
   REGISTERS_reg_31_47_inst : DFF_X1 port map( D => n5107, CK => CLK, Q => 
                           n8238, QN => n20206);
   REGISTERS_reg_31_46_inst : DFF_X1 port map( D => n5106, CK => CLK, Q => 
                           n8239, QN => n20207);
   REGISTERS_reg_31_45_inst : DFF_X1 port map( D => n5105, CK => CLK, Q => 
                           n8240, QN => n20208);
   REGISTERS_reg_31_44_inst : DFF_X1 port map( D => n5104, CK => CLK, Q => 
                           n8241, QN => n20209);
   REGISTERS_reg_31_43_inst : DFF_X1 port map( D => n5103, CK => CLK, Q => 
                           n8242, QN => n20210);
   REGISTERS_reg_31_42_inst : DFF_X1 port map( D => n5102, CK => CLK, Q => 
                           n8243, QN => n20211);
   REGISTERS_reg_31_41_inst : DFF_X1 port map( D => n5101, CK => CLK, Q => 
                           n8244, QN => n20212);
   REGISTERS_reg_31_40_inst : DFF_X1 port map( D => n5100, CK => CLK, Q => 
                           n8245, QN => n20213);
   REGISTERS_reg_20_63_inst : DFF_X1 port map( D => n5827, CK => CLK, Q => 
                           n_1168, QN => n20514);
   REGISTERS_reg_20_62_inst : DFF_X1 port map( D => n5826, CK => CLK, Q => 
                           n_1169, QN => n20515);
   REGISTERS_reg_20_61_inst : DFF_X1 port map( D => n5825, CK => CLK, Q => 
                           n_1170, QN => n20516);
   REGISTERS_reg_20_60_inst : DFF_X1 port map( D => n5824, CK => CLK, Q => 
                           n_1171, QN => n20517);
   REGISTERS_reg_3_63_inst : DFF_X1 port map( D => n6915, CK => CLK, Q => 
                           n_1172, QN => n20250);
   REGISTERS_reg_3_62_inst : DFF_X1 port map( D => n6914, CK => CLK, Q => 
                           n_1173, QN => n20251);
   REGISTERS_reg_3_61_inst : DFF_X1 port map( D => n6913, CK => CLK, Q => 
                           n_1174, QN => n20252);
   REGISTERS_reg_3_60_inst : DFF_X1 port map( D => n6912, CK => CLK, Q => 
                           n_1175, QN => n20253);
   REGISTERS_reg_17_63_inst : DFF_X1 port map( D => n6019, CK => CLK, Q => 
                           n_1176, QN => n20262);
   REGISTERS_reg_17_62_inst : DFF_X1 port map( D => n6018, CK => CLK, Q => 
                           n_1177, QN => n20263);
   REGISTERS_reg_17_61_inst : DFF_X1 port map( D => n6017, CK => CLK, Q => 
                           n_1178, QN => n20264);
   REGISTERS_reg_17_60_inst : DFF_X1 port map( D => n6016, CK => CLK, Q => 
                           n_1179, QN => n20265);
   REGISTERS_reg_24_63_inst : DFF_X1 port map( D => n5571, CK => CLK, Q => 
                           n_1180, QN => n20149);
   REGISTERS_reg_24_62_inst : DFF_X1 port map( D => n5570, CK => CLK, Q => 
                           n_1181, QN => n20150);
   REGISTERS_reg_24_61_inst : DFF_X1 port map( D => n5569, CK => CLK, Q => 
                           n_1182, QN => n20151);
   REGISTERS_reg_24_60_inst : DFF_X1 port map( D => n5568, CK => CLK, Q => 
                           n_1183, QN => n20152);
   REGISTERS_reg_7_63_inst : DFF_X1 port map( D => n6659, CK => CLK, Q => 
                           n_1184, QN => n20539);
   REGISTERS_reg_7_62_inst : DFF_X1 port map( D => n6658, CK => CLK, Q => 
                           n_1185, QN => n20540);
   REGISTERS_reg_7_61_inst : DFF_X1 port map( D => n6657, CK => CLK, Q => 
                           n_1186, QN => n20541);
   REGISTERS_reg_7_60_inst : DFF_X1 port map( D => n6656, CK => CLK, Q => 
                           n_1187, QN => n20542);
   REGISTERS_reg_6_63_inst : DFF_X1 port map( D => n6723, CK => CLK, Q => 
                           n_1188, QN => n20522);
   REGISTERS_reg_6_62_inst : DFF_X1 port map( D => n6722, CK => CLK, Q => 
                           n_1189, QN => n20523);
   REGISTERS_reg_6_61_inst : DFF_X1 port map( D => n6721, CK => CLK, Q => 
                           n_1190, QN => n20524);
   REGISTERS_reg_6_60_inst : DFF_X1 port map( D => n6720, CK => CLK, Q => 
                           n_1191, QN => n20525);
   REGISTERS_reg_2_63_inst : DFF_X1 port map( D => n6979, CK => CLK, Q => 
                           n_1192, QN => n20258);
   REGISTERS_reg_2_62_inst : DFF_X1 port map( D => n6978, CK => CLK, Q => 
                           n_1193, QN => n20259);
   REGISTERS_reg_2_61_inst : DFF_X1 port map( D => n6977, CK => CLK, Q => 
                           n_1194, QN => n20260);
   REGISTERS_reg_2_60_inst : DFF_X1 port map( D => n6976, CK => CLK, Q => 
                           n_1195, QN => n20261);
   REGISTERS_reg_20_59_inst : DFF_X1 port map( D => n5823, CK => CLK, Q => 
                           n_1196, QN => n20619);
   REGISTERS_reg_20_58_inst : DFF_X1 port map( D => n5822, CK => CLK, Q => 
                           n_1197, QN => n20620);
   REGISTERS_reg_20_57_inst : DFF_X1 port map( D => n5821, CK => CLK, Q => 
                           n_1198, QN => n20621);
   REGISTERS_reg_20_56_inst : DFF_X1 port map( D => n5820, CK => CLK, Q => 
                           n_1199, QN => n20622);
   REGISTERS_reg_20_55_inst : DFF_X1 port map( D => n5819, CK => CLK, Q => 
                           n_1200, QN => n20623);
   REGISTERS_reg_20_54_inst : DFF_X1 port map( D => n5818, CK => CLK, Q => 
                           n_1201, QN => n20624);
   REGISTERS_reg_20_53_inst : DFF_X1 port map( D => n5817, CK => CLK, Q => 
                           n_1202, QN => n20625);
   REGISTERS_reg_20_52_inst : DFF_X1 port map( D => n5816, CK => CLK, Q => 
                           n_1203, QN => n20626);
   REGISTERS_reg_20_51_inst : DFF_X1 port map( D => n5815, CK => CLK, Q => 
                           n_1204, QN => n20627);
   REGISTERS_reg_20_50_inst : DFF_X1 port map( D => n5814, CK => CLK, Q => 
                           n_1205, QN => n20628);
   REGISTERS_reg_20_49_inst : DFF_X1 port map( D => n5813, CK => CLK, Q => 
                           n_1206, QN => n20629);
   REGISTERS_reg_20_48_inst : DFF_X1 port map( D => n5812, CK => CLK, Q => 
                           n_1207, QN => n20630);
   REGISTERS_reg_20_47_inst : DFF_X1 port map( D => n5811, CK => CLK, Q => 
                           n_1208, QN => n20631);
   REGISTERS_reg_20_46_inst : DFF_X1 port map( D => n5810, CK => CLK, Q => 
                           n_1209, QN => n20632);
   REGISTERS_reg_20_45_inst : DFF_X1 port map( D => n5809, CK => CLK, Q => 
                           n_1210, QN => n20633);
   REGISTERS_reg_20_44_inst : DFF_X1 port map( D => n5808, CK => CLK, Q => 
                           n_1211, QN => n20634);
   REGISTERS_reg_20_43_inst : DFF_X1 port map( D => n5807, CK => CLK, Q => 
                           n_1212, QN => n20635);
   REGISTERS_reg_20_42_inst : DFF_X1 port map( D => n5806, CK => CLK, Q => 
                           n_1213, QN => n20636);
   REGISTERS_reg_20_41_inst : DFF_X1 port map( D => n5805, CK => CLK, Q => 
                           n_1214, QN => n20637);
   REGISTERS_reg_20_40_inst : DFF_X1 port map( D => n5804, CK => CLK, Q => 
                           n_1215, QN => n20638);
   REGISTERS_reg_20_39_inst : DFF_X1 port map( D => n5803, CK => CLK, Q => 
                           n_1216, QN => n20639);
   REGISTERS_reg_20_38_inst : DFF_X1 port map( D => n5802, CK => CLK, Q => 
                           n_1217, QN => n20640);
   REGISTERS_reg_20_37_inst : DFF_X1 port map( D => n5801, CK => CLK, Q => 
                           n_1218, QN => n20641);
   REGISTERS_reg_20_36_inst : DFF_X1 port map( D => n5800, CK => CLK, Q => 
                           n_1219, QN => n20642);
   REGISTERS_reg_20_35_inst : DFF_X1 port map( D => n5799, CK => CLK, Q => 
                           n_1220, QN => n20643);
   REGISTERS_reg_20_34_inst : DFF_X1 port map( D => n5798, CK => CLK, Q => 
                           n_1221, QN => n20644);
   REGISTERS_reg_20_33_inst : DFF_X1 port map( D => n5797, CK => CLK, Q => 
                           n_1222, QN => n20645);
   REGISTERS_reg_20_32_inst : DFF_X1 port map( D => n5796, CK => CLK, Q => 
                           n_1223, QN => n20646);
   REGISTERS_reg_20_31_inst : DFF_X1 port map( D => n5795, CK => CLK, Q => 
                           n_1224, QN => n20647);
   REGISTERS_reg_20_30_inst : DFF_X1 port map( D => n5794, CK => CLK, Q => 
                           n_1225, QN => n20648);
   REGISTERS_reg_20_29_inst : DFF_X1 port map( D => n5793, CK => CLK, Q => 
                           n_1226, QN => n20649);
   REGISTERS_reg_20_28_inst : DFF_X1 port map( D => n5792, CK => CLK, Q => 
                           n_1227, QN => n20650);
   REGISTERS_reg_20_27_inst : DFF_X1 port map( D => n5791, CK => CLK, Q => 
                           n_1228, QN => n20651);
   REGISTERS_reg_20_26_inst : DFF_X1 port map( D => n5790, CK => CLK, Q => 
                           n_1229, QN => n20652);
   REGISTERS_reg_20_25_inst : DFF_X1 port map( D => n5789, CK => CLK, Q => 
                           n_1230, QN => n20653);
   REGISTERS_reg_20_24_inst : DFF_X1 port map( D => n5788, CK => CLK, Q => 
                           n_1231, QN => n20654);
   REGISTERS_reg_3_59_inst : DFF_X1 port map( D => n6911, CK => CLK, Q => 
                           n_1232, QN => n20266);
   REGISTERS_reg_3_58_inst : DFF_X1 port map( D => n6910, CK => CLK, Q => 
                           n_1233, QN => n20267);
   REGISTERS_reg_3_57_inst : DFF_X1 port map( D => n6909, CK => CLK, Q => 
                           n_1234, QN => n20268);
   REGISTERS_reg_3_56_inst : DFF_X1 port map( D => n6908, CK => CLK, Q => 
                           n_1235, QN => n20269);
   REGISTERS_reg_3_55_inst : DFF_X1 port map( D => n6907, CK => CLK, Q => 
                           n_1236, QN => n20270);
   REGISTERS_reg_3_54_inst : DFF_X1 port map( D => n6906, CK => CLK, Q => 
                           n_1237, QN => n20271);
   REGISTERS_reg_3_53_inst : DFF_X1 port map( D => n6905, CK => CLK, Q => 
                           n_1238, QN => n20272);
   REGISTERS_reg_3_52_inst : DFF_X1 port map( D => n6904, CK => CLK, Q => 
                           n_1239, QN => n20273);
   REGISTERS_reg_3_51_inst : DFF_X1 port map( D => n6903, CK => CLK, Q => 
                           n_1240, QN => n20274);
   REGISTERS_reg_3_50_inst : DFF_X1 port map( D => n6902, CK => CLK, Q => 
                           n_1241, QN => n20275);
   REGISTERS_reg_3_49_inst : DFF_X1 port map( D => n6901, CK => CLK, Q => 
                           n_1242, QN => n20276);
   REGISTERS_reg_3_48_inst : DFF_X1 port map( D => n6900, CK => CLK, Q => 
                           n_1243, QN => n20277);
   REGISTERS_reg_3_47_inst : DFF_X1 port map( D => n6899, CK => CLK, Q => 
                           n_1244, QN => n20278);
   REGISTERS_reg_3_46_inst : DFF_X1 port map( D => n6898, CK => CLK, Q => 
                           n_1245, QN => n20279);
   REGISTERS_reg_3_45_inst : DFF_X1 port map( D => n6897, CK => CLK, Q => 
                           n_1246, QN => n20280);
   REGISTERS_reg_3_44_inst : DFF_X1 port map( D => n6896, CK => CLK, Q => 
                           n_1247, QN => n20281);
   REGISTERS_reg_3_43_inst : DFF_X1 port map( D => n6895, CK => CLK, Q => 
                           n_1248, QN => n20282);
   REGISTERS_reg_3_42_inst : DFF_X1 port map( D => n6894, CK => CLK, Q => 
                           n_1249, QN => n20283);
   REGISTERS_reg_3_41_inst : DFF_X1 port map( D => n6893, CK => CLK, Q => 
                           n_1250, QN => n20284);
   REGISTERS_reg_3_40_inst : DFF_X1 port map( D => n6892, CK => CLK, Q => 
                           n_1251, QN => n20285);
   REGISTERS_reg_3_39_inst : DFF_X1 port map( D => n6891, CK => CLK, Q => 
                           n_1252, QN => n20286);
   REGISTERS_reg_3_38_inst : DFF_X1 port map( D => n6890, CK => CLK, Q => 
                           n_1253, QN => n20287);
   REGISTERS_reg_3_37_inst : DFF_X1 port map( D => n6889, CK => CLK, Q => 
                           n_1254, QN => n20288);
   REGISTERS_reg_3_36_inst : DFF_X1 port map( D => n6888, CK => CLK, Q => 
                           n_1255, QN => n20289);
   REGISTERS_reg_3_35_inst : DFF_X1 port map( D => n6887, CK => CLK, Q => 
                           n_1256, QN => n20290);
   REGISTERS_reg_3_34_inst : DFF_X1 port map( D => n6886, CK => CLK, Q => 
                           n_1257, QN => n20291);
   REGISTERS_reg_3_33_inst : DFF_X1 port map( D => n6885, CK => CLK, Q => 
                           n_1258, QN => n20292);
   REGISTERS_reg_3_32_inst : DFF_X1 port map( D => n6884, CK => CLK, Q => 
                           n_1259, QN => n20293);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n6883, CK => CLK, Q => 
                           n_1260, QN => n20294);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n6882, CK => CLK, Q => 
                           n_1261, QN => n20295);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n6881, CK => CLK, Q => 
                           n_1262, QN => n20296);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n6880, CK => CLK, Q => 
                           n_1263, QN => n20297);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n6879, CK => CLK, Q => 
                           n_1264, QN => n20298);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n6878, CK => CLK, Q => 
                           n_1265, QN => n20299);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n6877, CK => CLK, Q => 
                           n_1266, QN => n20300);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n6876, CK => CLK, Q => 
                           n_1267, QN => n20301);
   REGISTERS_reg_20_23_inst : DFF_X1 port map( D => n5787, CK => CLK, Q => 
                           n_1268, QN => n20775);
   REGISTERS_reg_20_22_inst : DFF_X1 port map( D => n5786, CK => CLK, Q => 
                           n_1269, QN => n20776);
   REGISTERS_reg_20_21_inst : DFF_X1 port map( D => n5785, CK => CLK, Q => 
                           n_1270, QN => n20777);
   REGISTERS_reg_20_20_inst : DFF_X1 port map( D => n5784, CK => CLK, Q => 
                           n_1271, QN => n20778);
   REGISTERS_reg_20_19_inst : DFF_X1 port map( D => n5783, CK => CLK, Q => 
                           n_1272, QN => n20779);
   REGISTERS_reg_20_18_inst : DFF_X1 port map( D => n5782, CK => CLK, Q => 
                           n_1273, QN => n20780);
   REGISTERS_reg_20_17_inst : DFF_X1 port map( D => n5781, CK => CLK, Q => 
                           n_1274, QN => n20781);
   REGISTERS_reg_20_16_inst : DFF_X1 port map( D => n5780, CK => CLK, Q => 
                           n_1275, QN => n20782);
   REGISTERS_reg_20_15_inst : DFF_X1 port map( D => n5779, CK => CLK, Q => 
                           n_1276, QN => n20783);
   REGISTERS_reg_20_14_inst : DFF_X1 port map( D => n5778, CK => CLK, Q => 
                           n_1277, QN => n20784);
   REGISTERS_reg_20_13_inst : DFF_X1 port map( D => n5777, CK => CLK, Q => 
                           n_1278, QN => n20785);
   REGISTERS_reg_20_12_inst : DFF_X1 port map( D => n5776, CK => CLK, Q => 
                           n_1279, QN => n20786);
   REGISTERS_reg_20_11_inst : DFF_X1 port map( D => n5775, CK => CLK, Q => 
                           n_1280, QN => n20787);
   REGISTERS_reg_20_10_inst : DFF_X1 port map( D => n5774, CK => CLK, Q => 
                           n_1281, QN => n20788);
   REGISTERS_reg_20_9_inst : DFF_X1 port map( D => n5773, CK => CLK, Q => 
                           n_1282, QN => n20789);
   REGISTERS_reg_20_8_inst : DFF_X1 port map( D => n5772, CK => CLK, Q => 
                           n_1283, QN => n20790);
   REGISTERS_reg_20_7_inst : DFF_X1 port map( D => n5771, CK => CLK, Q => 
                           n_1284, QN => n20791);
   REGISTERS_reg_20_6_inst : DFF_X1 port map( D => n5770, CK => CLK, Q => 
                           n_1285, QN => n20792);
   REGISTERS_reg_20_5_inst : DFF_X1 port map( D => n5769, CK => CLK, Q => 
                           n_1286, QN => n20793);
   REGISTERS_reg_20_4_inst : DFF_X1 port map( D => n5768, CK => CLK, Q => 
                           n_1287, QN => n20794);
   REGISTERS_reg_20_3_inst : DFF_X1 port map( D => n5767, CK => CLK, Q => 
                           n_1288, QN => n20795);
   REGISTERS_reg_20_2_inst : DFF_X1 port map( D => n5766, CK => CLK, Q => 
                           n_1289, QN => n20796);
   REGISTERS_reg_20_1_inst : DFF_X1 port map( D => n5765, CK => CLK, Q => 
                           n_1290, QN => n20797);
   REGISTERS_reg_20_0_inst : DFF_X1 port map( D => n5764, CK => CLK, Q => 
                           n_1291, QN => n20798);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n6875, CK => CLK, Q => 
                           n_1292, QN => n20374);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n6874, CK => CLK, Q => 
                           n_1293, QN => n20375);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n6873, CK => CLK, Q => 
                           n_1294, QN => n20376);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n6872, CK => CLK, Q => 
                           n_1295, QN => n20377);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n6871, CK => CLK, Q => 
                           n_1296, QN => n20378);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n6870, CK => CLK, Q => 
                           n_1297, QN => n20379);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n6869, CK => CLK, Q => 
                           n_1298, QN => n20380);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n6868, CK => CLK, Q => 
                           n_1299, QN => n20381);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n6867, CK => CLK, Q => 
                           n_1300, QN => n20382);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n6866, CK => CLK, Q => 
                           n_1301, QN => n20383);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n6865, CK => CLK, Q => 
                           n_1302, QN => n20384);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n6864, CK => CLK, Q => 
                           n_1303, QN => n20385);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n6863, CK => CLK, Q => 
                           n_1304, QN => n20386);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n6862, CK => CLK, Q => 
                           n_1305, QN => n20387);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n6861, CK => CLK, Q => n_1306
                           , QN => n20388);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n6860, CK => CLK, Q => n_1307
                           , QN => n20389);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n6859, CK => CLK, Q => n_1308
                           , QN => n20390);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n6858, CK => CLK, Q => n_1309
                           , QN => n20391);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n6857, CK => CLK, Q => n_1310
                           , QN => n20392);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n6856, CK => CLK, Q => n_1311
                           , QN => n20393);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n6855, CK => CLK, Q => n_1312
                           , QN => n20394);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n6854, CK => CLK, Q => n_1313
                           , QN => n20395);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n6853, CK => CLK, Q => n_1314
                           , QN => n20396);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n6852, CK => CLK, Q => n_1315
                           , QN => n20397);
   REGISTERS_reg_17_59_inst : DFF_X1 port map( D => n6015, CK => CLK, Q => 
                           n_1316, QN => n20446);
   REGISTERS_reg_17_58_inst : DFF_X1 port map( D => n6014, CK => CLK, Q => 
                           n_1317, QN => n20447);
   REGISTERS_reg_17_57_inst : DFF_X1 port map( D => n6013, CK => CLK, Q => 
                           n_1318, QN => n20448);
   REGISTERS_reg_17_56_inst : DFF_X1 port map( D => n6012, CK => CLK, Q => 
                           n_1319, QN => n20449);
   REGISTERS_reg_17_55_inst : DFF_X1 port map( D => n6011, CK => CLK, Q => 
                           n_1320, QN => n20450);
   REGISTERS_reg_17_54_inst : DFF_X1 port map( D => n6010, CK => CLK, Q => 
                           n_1321, QN => n20451);
   REGISTERS_reg_17_53_inst : DFF_X1 port map( D => n6009, CK => CLK, Q => 
                           n_1322, QN => n20452);
   REGISTERS_reg_17_52_inst : DFF_X1 port map( D => n6008, CK => CLK, Q => 
                           n_1323, QN => n20453);
   REGISTERS_reg_17_51_inst : DFF_X1 port map( D => n6007, CK => CLK, Q => 
                           n_1324, QN => n20454);
   REGISTERS_reg_17_50_inst : DFF_X1 port map( D => n6006, CK => CLK, Q => 
                           n_1325, QN => n20455);
   REGISTERS_reg_17_49_inst : DFF_X1 port map( D => n6005, CK => CLK, Q => 
                           n_1326, QN => n20456);
   REGISTERS_reg_17_48_inst : DFF_X1 port map( D => n6004, CK => CLK, Q => 
                           n_1327, QN => n20457);
   REGISTERS_reg_17_47_inst : DFF_X1 port map( D => n6003, CK => CLK, Q => 
                           n_1328, QN => n20458);
   REGISTERS_reg_17_46_inst : DFF_X1 port map( D => n6002, CK => CLK, Q => 
                           n_1329, QN => n20459);
   REGISTERS_reg_17_45_inst : DFF_X1 port map( D => n6001, CK => CLK, Q => 
                           n_1330, QN => n20460);
   REGISTERS_reg_17_44_inst : DFF_X1 port map( D => n6000, CK => CLK, Q => 
                           n_1331, QN => n20461);
   REGISTERS_reg_17_43_inst : DFF_X1 port map( D => n5999, CK => CLK, Q => 
                           n_1332, QN => n20462);
   REGISTERS_reg_17_42_inst : DFF_X1 port map( D => n5998, CK => CLK, Q => 
                           n_1333, QN => n20463);
   REGISTERS_reg_17_41_inst : DFF_X1 port map( D => n5997, CK => CLK, Q => 
                           n_1334, QN => n20464);
   REGISTERS_reg_17_40_inst : DFF_X1 port map( D => n5996, CK => CLK, Q => 
                           n_1335, QN => n20465);
   REGISTERS_reg_17_39_inst : DFF_X1 port map( D => n5995, CK => CLK, Q => 
                           n_1336, QN => n20466);
   REGISTERS_reg_17_38_inst : DFF_X1 port map( D => n5994, CK => CLK, Q => 
                           n_1337, QN => n20467);
   REGISTERS_reg_17_37_inst : DFF_X1 port map( D => n5993, CK => CLK, Q => 
                           n_1338, QN => n20468);
   REGISTERS_reg_17_36_inst : DFF_X1 port map( D => n5992, CK => CLK, Q => 
                           n_1339, QN => n20469);
   REGISTERS_reg_17_35_inst : DFF_X1 port map( D => n5991, CK => CLK, Q => 
                           n_1340, QN => n20470);
   REGISTERS_reg_17_34_inst : DFF_X1 port map( D => n5990, CK => CLK, Q => 
                           n_1341, QN => n20471);
   REGISTERS_reg_17_33_inst : DFF_X1 port map( D => n5989, CK => CLK, Q => 
                           n_1342, QN => n20472);
   REGISTERS_reg_17_32_inst : DFF_X1 port map( D => n5988, CK => CLK, Q => 
                           n_1343, QN => n20473);
   REGISTERS_reg_17_31_inst : DFF_X1 port map( D => n5987, CK => CLK, Q => 
                           n_1344, QN => n20474);
   REGISTERS_reg_17_30_inst : DFF_X1 port map( D => n5986, CK => CLK, Q => 
                           n_1345, QN => n20475);
   REGISTERS_reg_17_29_inst : DFF_X1 port map( D => n5985, CK => CLK, Q => 
                           n_1346, QN => n20476);
   REGISTERS_reg_17_28_inst : DFF_X1 port map( D => n5984, CK => CLK, Q => 
                           n_1347, QN => n20477);
   REGISTERS_reg_17_27_inst : DFF_X1 port map( D => n5983, CK => CLK, Q => 
                           n_1348, QN => n20478);
   REGISTERS_reg_17_26_inst : DFF_X1 port map( D => n5982, CK => CLK, Q => 
                           n_1349, QN => n20479);
   REGISTERS_reg_17_25_inst : DFF_X1 port map( D => n5981, CK => CLK, Q => 
                           n_1350, QN => n20480);
   REGISTERS_reg_17_24_inst : DFF_X1 port map( D => n5980, CK => CLK, Q => 
                           n_1351, QN => n20481);
   REGISTERS_reg_24_59_inst : DFF_X1 port map( D => n5567, CK => CLK, Q => 
                           n_1352, QN => n19648);
   REGISTERS_reg_24_58_inst : DFF_X1 port map( D => n5566, CK => CLK, Q => 
                           n_1353, QN => n19649);
   REGISTERS_reg_24_57_inst : DFF_X1 port map( D => n5565, CK => CLK, Q => 
                           n_1354, QN => n19650);
   REGISTERS_reg_24_56_inst : DFF_X1 port map( D => n5564, CK => CLK, Q => 
                           n_1355, QN => n19651);
   REGISTERS_reg_24_55_inst : DFF_X1 port map( D => n5563, CK => CLK, Q => 
                           n_1356, QN => n19652);
   REGISTERS_reg_24_54_inst : DFF_X1 port map( D => n5562, CK => CLK, Q => 
                           n_1357, QN => n19653);
   REGISTERS_reg_24_53_inst : DFF_X1 port map( D => n5561, CK => CLK, Q => 
                           n_1358, QN => n19654);
   REGISTERS_reg_24_52_inst : DFF_X1 port map( D => n5560, CK => CLK, Q => 
                           n_1359, QN => n19655);
   REGISTERS_reg_24_51_inst : DFF_X1 port map( D => n5559, CK => CLK, Q => 
                           n_1360, QN => n19656);
   REGISTERS_reg_24_50_inst : DFF_X1 port map( D => n5558, CK => CLK, Q => 
                           n_1361, QN => n19657);
   REGISTERS_reg_24_49_inst : DFF_X1 port map( D => n5557, CK => CLK, Q => 
                           n_1362, QN => n19658);
   REGISTERS_reg_24_48_inst : DFF_X1 port map( D => n5556, CK => CLK, Q => 
                           n_1363, QN => n19659);
   REGISTERS_reg_24_47_inst : DFF_X1 port map( D => n5555, CK => CLK, Q => 
                           n_1364, QN => n19660);
   REGISTERS_reg_24_46_inst : DFF_X1 port map( D => n5554, CK => CLK, Q => 
                           n_1365, QN => n19661);
   REGISTERS_reg_24_45_inst : DFF_X1 port map( D => n5553, CK => CLK, Q => 
                           n_1366, QN => n19662);
   REGISTERS_reg_24_44_inst : DFF_X1 port map( D => n5552, CK => CLK, Q => 
                           n_1367, QN => n19663);
   REGISTERS_reg_24_43_inst : DFF_X1 port map( D => n5551, CK => CLK, Q => 
                           n_1368, QN => n19664);
   REGISTERS_reg_24_42_inst : DFF_X1 port map( D => n5550, CK => CLK, Q => 
                           n_1369, QN => n19665);
   REGISTERS_reg_24_41_inst : DFF_X1 port map( D => n5549, CK => CLK, Q => 
                           n_1370, QN => n19666);
   REGISTERS_reg_24_40_inst : DFF_X1 port map( D => n5548, CK => CLK, Q => 
                           n_1371, QN => n19667);
   REGISTERS_reg_24_39_inst : DFF_X1 port map( D => n5547, CK => CLK, Q => 
                           n_1372, QN => n19668);
   REGISTERS_reg_24_38_inst : DFF_X1 port map( D => n5546, CK => CLK, Q => 
                           n_1373, QN => n19669);
   REGISTERS_reg_24_37_inst : DFF_X1 port map( D => n5545, CK => CLK, Q => 
                           n_1374, QN => n19670);
   REGISTERS_reg_24_36_inst : DFF_X1 port map( D => n5544, CK => CLK, Q => 
                           n_1375, QN => n19671);
   REGISTERS_reg_24_35_inst : DFF_X1 port map( D => n5543, CK => CLK, Q => 
                           n_1376, QN => n19672);
   REGISTERS_reg_24_34_inst : DFF_X1 port map( D => n5542, CK => CLK, Q => 
                           n_1377, QN => n19673);
   REGISTERS_reg_24_33_inst : DFF_X1 port map( D => n5541, CK => CLK, Q => 
                           n_1378, QN => n19674);
   REGISTERS_reg_24_32_inst : DFF_X1 port map( D => n5540, CK => CLK, Q => 
                           n_1379, QN => n19675);
   REGISTERS_reg_24_31_inst : DFF_X1 port map( D => n5539, CK => CLK, Q => 
                           n_1380, QN => n19676);
   REGISTERS_reg_24_30_inst : DFF_X1 port map( D => n5538, CK => CLK, Q => 
                           n_1381, QN => n19677);
   REGISTERS_reg_24_29_inst : DFF_X1 port map( D => n5537, CK => CLK, Q => 
                           n_1382, QN => n19678);
   REGISTERS_reg_24_28_inst : DFF_X1 port map( D => n5536, CK => CLK, Q => 
                           n_1383, QN => n19679);
   REGISTERS_reg_24_27_inst : DFF_X1 port map( D => n5535, CK => CLK, Q => 
                           n_1384, QN => n19680);
   REGISTERS_reg_24_26_inst : DFF_X1 port map( D => n5534, CK => CLK, Q => 
                           n_1385, QN => n19681);
   REGISTERS_reg_24_25_inst : DFF_X1 port map( D => n5533, CK => CLK, Q => 
                           n_1386, QN => n19682);
   REGISTERS_reg_24_24_inst : DFF_X1 port map( D => n5532, CK => CLK, Q => 
                           n_1387, QN => n19683);
   REGISTERS_reg_7_59_inst : DFF_X1 port map( D => n6655, CK => CLK, Q => 
                           n_1388, QN => n20979);
   REGISTERS_reg_7_58_inst : DFF_X1 port map( D => n6654, CK => CLK, Q => 
                           n_1389, QN => n20980);
   REGISTERS_reg_7_57_inst : DFF_X1 port map( D => n6653, CK => CLK, Q => 
                           n_1390, QN => n20981);
   REGISTERS_reg_7_56_inst : DFF_X1 port map( D => n6652, CK => CLK, Q => 
                           n_1391, QN => n20982);
   REGISTERS_reg_7_55_inst : DFF_X1 port map( D => n6651, CK => CLK, Q => 
                           n_1392, QN => n20983);
   REGISTERS_reg_7_54_inst : DFF_X1 port map( D => n6650, CK => CLK, Q => 
                           n_1393, QN => n20984);
   REGISTERS_reg_7_53_inst : DFF_X1 port map( D => n6649, CK => CLK, Q => 
                           n_1394, QN => n20985);
   REGISTERS_reg_7_52_inst : DFF_X1 port map( D => n6648, CK => CLK, Q => 
                           n_1395, QN => n20986);
   REGISTERS_reg_7_51_inst : DFF_X1 port map( D => n6647, CK => CLK, Q => 
                           n_1396, QN => n20987);
   REGISTERS_reg_7_50_inst : DFF_X1 port map( D => n6646, CK => CLK, Q => 
                           n_1397, QN => n20988);
   REGISTERS_reg_7_49_inst : DFF_X1 port map( D => n6645, CK => CLK, Q => 
                           n_1398, QN => n20989);
   REGISTERS_reg_7_48_inst : DFF_X1 port map( D => n6644, CK => CLK, Q => 
                           n_1399, QN => n20990);
   REGISTERS_reg_7_47_inst : DFF_X1 port map( D => n6643, CK => CLK, Q => 
                           n_1400, QN => n20991);
   REGISTERS_reg_7_46_inst : DFF_X1 port map( D => n6642, CK => CLK, Q => 
                           n_1401, QN => n20992);
   REGISTERS_reg_7_45_inst : DFF_X1 port map( D => n6641, CK => CLK, Q => 
                           n_1402, QN => n20993);
   REGISTERS_reg_7_44_inst : DFF_X1 port map( D => n6640, CK => CLK, Q => 
                           n_1403, QN => n20994);
   REGISTERS_reg_7_43_inst : DFF_X1 port map( D => n6639, CK => CLK, Q => 
                           n_1404, QN => n20995);
   REGISTERS_reg_7_42_inst : DFF_X1 port map( D => n6638, CK => CLK, Q => 
                           n_1405, QN => n20996);
   REGISTERS_reg_7_41_inst : DFF_X1 port map( D => n6637, CK => CLK, Q => 
                           n_1406, QN => n20997);
   REGISTERS_reg_7_40_inst : DFF_X1 port map( D => n6636, CK => CLK, Q => 
                           n_1407, QN => n20998);
   REGISTERS_reg_7_39_inst : DFF_X1 port map( D => n6635, CK => CLK, Q => 
                           n_1408, QN => n20999);
   REGISTERS_reg_7_38_inst : DFF_X1 port map( D => n6634, CK => CLK, Q => 
                           n_1409, QN => n21000);
   REGISTERS_reg_7_37_inst : DFF_X1 port map( D => n6633, CK => CLK, Q => 
                           n_1410, QN => n21001);
   REGISTERS_reg_7_36_inst : DFF_X1 port map( D => n6632, CK => CLK, Q => 
                           n_1411, QN => n21002);
   REGISTERS_reg_7_35_inst : DFF_X1 port map( D => n6631, CK => CLK, Q => 
                           n_1412, QN => n21003);
   REGISTERS_reg_7_34_inst : DFF_X1 port map( D => n6630, CK => CLK, Q => 
                           n_1413, QN => n21004);
   REGISTERS_reg_7_33_inst : DFF_X1 port map( D => n6629, CK => CLK, Q => 
                           n_1414, QN => n21005);
   REGISTERS_reg_7_32_inst : DFF_X1 port map( D => n6628, CK => CLK, Q => 
                           n_1415, QN => n21006);
   REGISTERS_reg_7_31_inst : DFF_X1 port map( D => n6627, CK => CLK, Q => 
                           n_1416, QN => n21007);
   REGISTERS_reg_7_30_inst : DFF_X1 port map( D => n6626, CK => CLK, Q => 
                           n_1417, QN => n21008);
   REGISTERS_reg_7_29_inst : DFF_X1 port map( D => n6625, CK => CLK, Q => 
                           n_1418, QN => n21009);
   REGISTERS_reg_7_28_inst : DFF_X1 port map( D => n6624, CK => CLK, Q => 
                           n_1419, QN => n21010);
   REGISTERS_reg_7_27_inst : DFF_X1 port map( D => n6623, CK => CLK, Q => 
                           n_1420, QN => n21011);
   REGISTERS_reg_7_26_inst : DFF_X1 port map( D => n6622, CK => CLK, Q => 
                           n_1421, QN => n21012);
   REGISTERS_reg_7_25_inst : DFF_X1 port map( D => n6621, CK => CLK, Q => 
                           n_1422, QN => n21013);
   REGISTERS_reg_7_24_inst : DFF_X1 port map( D => n6620, CK => CLK, Q => 
                           n_1423, QN => n21014);
   REGISTERS_reg_6_59_inst : DFF_X1 port map( D => n6719, CK => CLK, Q => 
                           n_1424, QN => n20691);
   REGISTERS_reg_6_58_inst : DFF_X1 port map( D => n6718, CK => CLK, Q => 
                           n_1425, QN => n20692);
   REGISTERS_reg_6_57_inst : DFF_X1 port map( D => n6717, CK => CLK, Q => 
                           n_1426, QN => n20693);
   REGISTERS_reg_6_56_inst : DFF_X1 port map( D => n6716, CK => CLK, Q => 
                           n_1427, QN => n20694);
   REGISTERS_reg_6_55_inst : DFF_X1 port map( D => n6715, CK => CLK, Q => 
                           n_1428, QN => n20695);
   REGISTERS_reg_6_54_inst : DFF_X1 port map( D => n6714, CK => CLK, Q => 
                           n_1429, QN => n20696);
   REGISTERS_reg_6_53_inst : DFF_X1 port map( D => n6713, CK => CLK, Q => 
                           n_1430, QN => n20697);
   REGISTERS_reg_6_52_inst : DFF_X1 port map( D => n6712, CK => CLK, Q => 
                           n_1431, QN => n20698);
   REGISTERS_reg_6_51_inst : DFF_X1 port map( D => n6711, CK => CLK, Q => 
                           n_1432, QN => n20699);
   REGISTERS_reg_6_50_inst : DFF_X1 port map( D => n6710, CK => CLK, Q => 
                           n_1433, QN => n20700);
   REGISTERS_reg_6_49_inst : DFF_X1 port map( D => n6709, CK => CLK, Q => 
                           n_1434, QN => n20701);
   REGISTERS_reg_6_48_inst : DFF_X1 port map( D => n6708, CK => CLK, Q => 
                           n_1435, QN => n20702);
   REGISTERS_reg_6_47_inst : DFF_X1 port map( D => n6707, CK => CLK, Q => 
                           n_1436, QN => n20703);
   REGISTERS_reg_6_46_inst : DFF_X1 port map( D => n6706, CK => CLK, Q => 
                           n_1437, QN => n20704);
   REGISTERS_reg_6_45_inst : DFF_X1 port map( D => n6705, CK => CLK, Q => 
                           n_1438, QN => n20705);
   REGISTERS_reg_6_44_inst : DFF_X1 port map( D => n6704, CK => CLK, Q => 
                           n_1439, QN => n20706);
   REGISTERS_reg_6_43_inst : DFF_X1 port map( D => n6703, CK => CLK, Q => 
                           n_1440, QN => n20707);
   REGISTERS_reg_6_42_inst : DFF_X1 port map( D => n6702, CK => CLK, Q => 
                           n_1441, QN => n20708);
   REGISTERS_reg_6_41_inst : DFF_X1 port map( D => n6701, CK => CLK, Q => 
                           n_1442, QN => n20709);
   REGISTERS_reg_6_40_inst : DFF_X1 port map( D => n6700, CK => CLK, Q => 
                           n_1443, QN => n20710);
   REGISTERS_reg_6_39_inst : DFF_X1 port map( D => n6699, CK => CLK, Q => 
                           n_1444, QN => n20711);
   REGISTERS_reg_6_38_inst : DFF_X1 port map( D => n6698, CK => CLK, Q => 
                           n_1445, QN => n20712);
   REGISTERS_reg_6_37_inst : DFF_X1 port map( D => n6697, CK => CLK, Q => 
                           n_1446, QN => n20713);
   REGISTERS_reg_6_36_inst : DFF_X1 port map( D => n6696, CK => CLK, Q => 
                           n_1447, QN => n20714);
   REGISTERS_reg_6_35_inst : DFF_X1 port map( D => n6695, CK => CLK, Q => 
                           n_1448, QN => n20715);
   REGISTERS_reg_6_34_inst : DFF_X1 port map( D => n6694, CK => CLK, Q => 
                           n_1449, QN => n20716);
   REGISTERS_reg_6_33_inst : DFF_X1 port map( D => n6693, CK => CLK, Q => 
                           n_1450, QN => n20717);
   REGISTERS_reg_6_32_inst : DFF_X1 port map( D => n6692, CK => CLK, Q => 
                           n_1451, QN => n20718);
   REGISTERS_reg_6_31_inst : DFF_X1 port map( D => n6691, CK => CLK, Q => 
                           n_1452, QN => n20719);
   REGISTERS_reg_6_30_inst : DFF_X1 port map( D => n6690, CK => CLK, Q => 
                           n_1453, QN => n20720);
   REGISTERS_reg_6_29_inst : DFF_X1 port map( D => n6689, CK => CLK, Q => 
                           n_1454, QN => n20721);
   REGISTERS_reg_6_28_inst : DFF_X1 port map( D => n6688, CK => CLK, Q => 
                           n_1455, QN => n20722);
   REGISTERS_reg_6_27_inst : DFF_X1 port map( D => n6687, CK => CLK, Q => 
                           n_1456, QN => n20723);
   REGISTERS_reg_6_26_inst : DFF_X1 port map( D => n6686, CK => CLK, Q => 
                           n_1457, QN => n20724);
   REGISTERS_reg_6_25_inst : DFF_X1 port map( D => n6685, CK => CLK, Q => 
                           n_1458, QN => n20725);
   REGISTERS_reg_6_24_inst : DFF_X1 port map( D => n6684, CK => CLK, Q => 
                           n_1459, QN => n20726);
   REGISTERS_reg_2_59_inst : DFF_X1 port map( D => n6975, CK => CLK, Q => 
                           n_1460, QN => n20338);
   REGISTERS_reg_2_58_inst : DFF_X1 port map( D => n6974, CK => CLK, Q => 
                           n_1461, QN => n20339);
   REGISTERS_reg_2_57_inst : DFF_X1 port map( D => n6973, CK => CLK, Q => 
                           n_1462, QN => n20340);
   REGISTERS_reg_2_56_inst : DFF_X1 port map( D => n6972, CK => CLK, Q => 
                           n_1463, QN => n20341);
   REGISTERS_reg_2_55_inst : DFF_X1 port map( D => n6971, CK => CLK, Q => 
                           n_1464, QN => n20342);
   REGISTERS_reg_2_54_inst : DFF_X1 port map( D => n6970, CK => CLK, Q => 
                           n_1465, QN => n20343);
   REGISTERS_reg_2_53_inst : DFF_X1 port map( D => n6969, CK => CLK, Q => 
                           n_1466, QN => n20344);
   REGISTERS_reg_2_52_inst : DFF_X1 port map( D => n6968, CK => CLK, Q => 
                           n_1467, QN => n20345);
   REGISTERS_reg_2_51_inst : DFF_X1 port map( D => n6967, CK => CLK, Q => 
                           n_1468, QN => n20346);
   REGISTERS_reg_2_50_inst : DFF_X1 port map( D => n6966, CK => CLK, Q => 
                           n_1469, QN => n20347);
   REGISTERS_reg_2_49_inst : DFF_X1 port map( D => n6965, CK => CLK, Q => 
                           n_1470, QN => n20348);
   REGISTERS_reg_2_48_inst : DFF_X1 port map( D => n6964, CK => CLK, Q => 
                           n_1471, QN => n20349);
   REGISTERS_reg_2_47_inst : DFF_X1 port map( D => n6963, CK => CLK, Q => 
                           n_1472, QN => n20350);
   REGISTERS_reg_2_46_inst : DFF_X1 port map( D => n6962, CK => CLK, Q => 
                           n_1473, QN => n20351);
   REGISTERS_reg_2_45_inst : DFF_X1 port map( D => n6961, CK => CLK, Q => 
                           n_1474, QN => n20352);
   REGISTERS_reg_2_44_inst : DFF_X1 port map( D => n6960, CK => CLK, Q => 
                           n_1475, QN => n20353);
   REGISTERS_reg_2_43_inst : DFF_X1 port map( D => n6959, CK => CLK, Q => 
                           n_1476, QN => n20354);
   REGISTERS_reg_2_42_inst : DFF_X1 port map( D => n6958, CK => CLK, Q => 
                           n_1477, QN => n20355);
   REGISTERS_reg_2_41_inst : DFF_X1 port map( D => n6957, CK => CLK, Q => 
                           n_1478, QN => n20356);
   REGISTERS_reg_2_40_inst : DFF_X1 port map( D => n6956, CK => CLK, Q => 
                           n_1479, QN => n20357);
   REGISTERS_reg_2_39_inst : DFF_X1 port map( D => n6955, CK => CLK, Q => 
                           n_1480, QN => n20358);
   REGISTERS_reg_2_38_inst : DFF_X1 port map( D => n6954, CK => CLK, Q => 
                           n_1481, QN => n20359);
   REGISTERS_reg_2_37_inst : DFF_X1 port map( D => n6953, CK => CLK, Q => 
                           n_1482, QN => n20360);
   REGISTERS_reg_2_36_inst : DFF_X1 port map( D => n6952, CK => CLK, Q => 
                           n_1483, QN => n20361);
   REGISTERS_reg_2_35_inst : DFF_X1 port map( D => n6951, CK => CLK, Q => 
                           n_1484, QN => n20362);
   REGISTERS_reg_2_34_inst : DFF_X1 port map( D => n6950, CK => CLK, Q => 
                           n_1485, QN => n20363);
   REGISTERS_reg_2_33_inst : DFF_X1 port map( D => n6949, CK => CLK, Q => 
                           n_1486, QN => n20364);
   REGISTERS_reg_2_32_inst : DFF_X1 port map( D => n6948, CK => CLK, Q => 
                           n_1487, QN => n20365);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n6947, CK => CLK, Q => 
                           n_1488, QN => n20366);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n6946, CK => CLK, Q => 
                           n_1489, QN => n20367);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n6945, CK => CLK, Q => 
                           n_1490, QN => n20368);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n6944, CK => CLK, Q => 
                           n_1491, QN => n20369);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n6943, CK => CLK, Q => 
                           n_1492, QN => n20370);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n6942, CK => CLK, Q => 
                           n_1493, QN => n20371);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n6941, CK => CLK, Q => 
                           n_1494, QN => n20372);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n6940, CK => CLK, Q => 
                           n_1495, QN => n20373);
   REGISTERS_reg_17_23_inst : DFF_X1 port map( D => n5979, CK => CLK, Q => 
                           n_1496, QN => n20482);
   REGISTERS_reg_17_22_inst : DFF_X1 port map( D => n5978, CK => CLK, Q => 
                           n_1497, QN => n20483);
   REGISTERS_reg_17_21_inst : DFF_X1 port map( D => n5977, CK => CLK, Q => 
                           n_1498, QN => n20484);
   REGISTERS_reg_17_20_inst : DFF_X1 port map( D => n5976, CK => CLK, Q => 
                           n_1499, QN => n20485);
   REGISTERS_reg_17_19_inst : DFF_X1 port map( D => n5975, CK => CLK, Q => 
                           n_1500, QN => n20486);
   REGISTERS_reg_17_18_inst : DFF_X1 port map( D => n5974, CK => CLK, Q => 
                           n_1501, QN => n20487);
   REGISTERS_reg_17_17_inst : DFF_X1 port map( D => n5973, CK => CLK, Q => 
                           n_1502, QN => n20488);
   REGISTERS_reg_17_16_inst : DFF_X1 port map( D => n5972, CK => CLK, Q => 
                           n_1503, QN => n20489);
   REGISTERS_reg_17_15_inst : DFF_X1 port map( D => n5971, CK => CLK, Q => 
                           n_1504, QN => n20490);
   REGISTERS_reg_17_14_inst : DFF_X1 port map( D => n5970, CK => CLK, Q => 
                           n_1505, QN => n20491);
   REGISTERS_reg_17_13_inst : DFF_X1 port map( D => n5969, CK => CLK, Q => 
                           n_1506, QN => n20492);
   REGISTERS_reg_17_12_inst : DFF_X1 port map( D => n5968, CK => CLK, Q => 
                           n_1507, QN => n20493);
   REGISTERS_reg_17_11_inst : DFF_X1 port map( D => n5967, CK => CLK, Q => 
                           n_1508, QN => n20494);
   REGISTERS_reg_17_10_inst : DFF_X1 port map( D => n5966, CK => CLK, Q => 
                           n_1509, QN => n20495);
   REGISTERS_reg_17_9_inst : DFF_X1 port map( D => n5965, CK => CLK, Q => 
                           n_1510, QN => n20496);
   REGISTERS_reg_17_8_inst : DFF_X1 port map( D => n5964, CK => CLK, Q => 
                           n_1511, QN => n20497);
   REGISTERS_reg_17_7_inst : DFF_X1 port map( D => n5963, CK => CLK, Q => 
                           n_1512, QN => n20498);
   REGISTERS_reg_17_6_inst : DFF_X1 port map( D => n5962, CK => CLK, Q => 
                           n_1513, QN => n20499);
   REGISTERS_reg_17_5_inst : DFF_X1 port map( D => n5961, CK => CLK, Q => 
                           n_1514, QN => n20500);
   REGISTERS_reg_17_4_inst : DFF_X1 port map( D => n5960, CK => CLK, Q => 
                           n_1515, QN => n20501);
   REGISTERS_reg_17_3_inst : DFF_X1 port map( D => n5959, CK => CLK, Q => 
                           n_1516, QN => n20502);
   REGISTERS_reg_17_2_inst : DFF_X1 port map( D => n5958, CK => CLK, Q => 
                           n_1517, QN => n20503);
   REGISTERS_reg_17_1_inst : DFF_X1 port map( D => n5957, CK => CLK, Q => 
                           n_1518, QN => n20504);
   REGISTERS_reg_17_0_inst : DFF_X1 port map( D => n5956, CK => CLK, Q => 
                           n_1519, QN => n20505);
   REGISTERS_reg_24_23_inst : DFF_X1 port map( D => n5531, CK => CLK, Q => 
                           n_1520, QN => n19684);
   REGISTERS_reg_24_22_inst : DFF_X1 port map( D => n5530, CK => CLK, Q => 
                           n_1521, QN => n19685);
   REGISTERS_reg_24_21_inst : DFF_X1 port map( D => n5529, CK => CLK, Q => 
                           n_1522, QN => n19686);
   REGISTERS_reg_24_20_inst : DFF_X1 port map( D => n5528, CK => CLK, Q => 
                           n_1523, QN => n19687);
   REGISTERS_reg_24_19_inst : DFF_X1 port map( D => n5527, CK => CLK, Q => 
                           n_1524, QN => n19688);
   REGISTERS_reg_24_18_inst : DFF_X1 port map( D => n5526, CK => CLK, Q => 
                           n_1525, QN => n19689);
   REGISTERS_reg_24_17_inst : DFF_X1 port map( D => n5525, CK => CLK, Q => 
                           n_1526, QN => n19690);
   REGISTERS_reg_24_16_inst : DFF_X1 port map( D => n5524, CK => CLK, Q => 
                           n_1527, QN => n19691);
   REGISTERS_reg_24_15_inst : DFF_X1 port map( D => n5523, CK => CLK, Q => 
                           n_1528, QN => n19692);
   REGISTERS_reg_24_14_inst : DFF_X1 port map( D => n5522, CK => CLK, Q => 
                           n_1529, QN => n19693);
   REGISTERS_reg_24_13_inst : DFF_X1 port map( D => n5521, CK => CLK, Q => 
                           n_1530, QN => n19694);
   REGISTERS_reg_24_12_inst : DFF_X1 port map( D => n5520, CK => CLK, Q => 
                           n_1531, QN => n19695);
   REGISTERS_reg_24_11_inst : DFF_X1 port map( D => n5519, CK => CLK, Q => 
                           n_1532, QN => n19696);
   REGISTERS_reg_24_10_inst : DFF_X1 port map( D => n5518, CK => CLK, Q => 
                           n_1533, QN => n19697);
   REGISTERS_reg_24_9_inst : DFF_X1 port map( D => n5517, CK => CLK, Q => 
                           n_1534, QN => n19698);
   REGISTERS_reg_24_8_inst : DFF_X1 port map( D => n5516, CK => CLK, Q => 
                           n_1535, QN => n19699);
   REGISTERS_reg_24_7_inst : DFF_X1 port map( D => n5515, CK => CLK, Q => 
                           n_1536, QN => n19700);
   REGISTERS_reg_24_6_inst : DFF_X1 port map( D => n5514, CK => CLK, Q => 
                           n_1537, QN => n19701);
   REGISTERS_reg_24_5_inst : DFF_X1 port map( D => n5513, CK => CLK, Q => 
                           n_1538, QN => n19702);
   REGISTERS_reg_24_4_inst : DFF_X1 port map( D => n5512, CK => CLK, Q => 
                           n_1539, QN => n19703);
   REGISTERS_reg_24_3_inst : DFF_X1 port map( D => n5511, CK => CLK, Q => 
                           n_1540, QN => n19704);
   REGISTERS_reg_24_2_inst : DFF_X1 port map( D => n5510, CK => CLK, Q => 
                           n_1541, QN => n19705);
   REGISTERS_reg_24_1_inst : DFF_X1 port map( D => n5509, CK => CLK, Q => 
                           n_1542, QN => n19706);
   REGISTERS_reg_24_0_inst : DFF_X1 port map( D => n5508, CK => CLK, Q => 
                           n_1543, QN => n19707);
   REGISTERS_reg_7_23_inst : DFF_X1 port map( D => n6619, CK => CLK, Q => 
                           n_1544, QN => n21099);
   REGISTERS_reg_7_22_inst : DFF_X1 port map( D => n6618, CK => CLK, Q => 
                           n_1545, QN => n21100);
   REGISTERS_reg_7_21_inst : DFF_X1 port map( D => n6617, CK => CLK, Q => 
                           n_1546, QN => n21101);
   REGISTERS_reg_7_20_inst : DFF_X1 port map( D => n6616, CK => CLK, Q => 
                           n_1547, QN => n21102);
   REGISTERS_reg_7_19_inst : DFF_X1 port map( D => n6615, CK => CLK, Q => 
                           n_1548, QN => n21103);
   REGISTERS_reg_7_18_inst : DFF_X1 port map( D => n6614, CK => CLK, Q => 
                           n_1549, QN => n21104);
   REGISTERS_reg_7_17_inst : DFF_X1 port map( D => n6613, CK => CLK, Q => 
                           n_1550, QN => n21105);
   REGISTERS_reg_7_16_inst : DFF_X1 port map( D => n6612, CK => CLK, Q => 
                           n_1551, QN => n21106);
   REGISTERS_reg_7_15_inst : DFF_X1 port map( D => n6611, CK => CLK, Q => 
                           n_1552, QN => n21107);
   REGISTERS_reg_7_14_inst : DFF_X1 port map( D => n6610, CK => CLK, Q => 
                           n_1553, QN => n21108);
   REGISTERS_reg_7_13_inst : DFF_X1 port map( D => n6609, CK => CLK, Q => 
                           n_1554, QN => n21109);
   REGISTERS_reg_7_12_inst : DFF_X1 port map( D => n6608, CK => CLK, Q => 
                           n_1555, QN => n21110);
   REGISTERS_reg_7_11_inst : DFF_X1 port map( D => n6607, CK => CLK, Q => 
                           n_1556, QN => n21111);
   REGISTERS_reg_7_10_inst : DFF_X1 port map( D => n6606, CK => CLK, Q => 
                           n_1557, QN => n21112);
   REGISTERS_reg_7_9_inst : DFF_X1 port map( D => n6605, CK => CLK, Q => n_1558
                           , QN => n21113);
   REGISTERS_reg_7_8_inst : DFF_X1 port map( D => n6604, CK => CLK, Q => n_1559
                           , QN => n21114);
   REGISTERS_reg_7_7_inst : DFF_X1 port map( D => n6603, CK => CLK, Q => n_1560
                           , QN => n21115);
   REGISTERS_reg_7_6_inst : DFF_X1 port map( D => n6602, CK => CLK, Q => n_1561
                           , QN => n21116);
   REGISTERS_reg_7_5_inst : DFF_X1 port map( D => n6601, CK => CLK, Q => n_1562
                           , QN => n21117);
   REGISTERS_reg_7_4_inst : DFF_X1 port map( D => n6600, CK => CLK, Q => n_1563
                           , QN => n21118);
   REGISTERS_reg_7_3_inst : DFF_X1 port map( D => n6599, CK => CLK, Q => n_1564
                           , QN => n21119);
   REGISTERS_reg_7_2_inst : DFF_X1 port map( D => n6598, CK => CLK, Q => n_1565
                           , QN => n21120);
   REGISTERS_reg_7_1_inst : DFF_X1 port map( D => n6597, CK => CLK, Q => n_1566
                           , QN => n21121);
   REGISTERS_reg_7_0_inst : DFF_X1 port map( D => n6596, CK => CLK, Q => n_1567
                           , QN => n21122);
   REGISTERS_reg_6_23_inst : DFF_X1 port map( D => n6683, CK => CLK, Q => 
                           n_1568, QN => n20823);
   REGISTERS_reg_6_22_inst : DFF_X1 port map( D => n6682, CK => CLK, Q => 
                           n_1569, QN => n20824);
   REGISTERS_reg_6_21_inst : DFF_X1 port map( D => n6681, CK => CLK, Q => 
                           n_1570, QN => n20825);
   REGISTERS_reg_6_20_inst : DFF_X1 port map( D => n6680, CK => CLK, Q => 
                           n_1571, QN => n20826);
   REGISTERS_reg_6_19_inst : DFF_X1 port map( D => n6679, CK => CLK, Q => 
                           n_1572, QN => n20827);
   REGISTERS_reg_6_18_inst : DFF_X1 port map( D => n6678, CK => CLK, Q => 
                           n_1573, QN => n20828);
   REGISTERS_reg_6_17_inst : DFF_X1 port map( D => n6677, CK => CLK, Q => 
                           n_1574, QN => n20829);
   REGISTERS_reg_6_16_inst : DFF_X1 port map( D => n6676, CK => CLK, Q => 
                           n_1575, QN => n20830);
   REGISTERS_reg_6_15_inst : DFF_X1 port map( D => n6675, CK => CLK, Q => 
                           n_1576, QN => n20831);
   REGISTERS_reg_6_14_inst : DFF_X1 port map( D => n6674, CK => CLK, Q => 
                           n_1577, QN => n20832);
   REGISTERS_reg_6_13_inst : DFF_X1 port map( D => n6673, CK => CLK, Q => 
                           n_1578, QN => n20833);
   REGISTERS_reg_6_12_inst : DFF_X1 port map( D => n6672, CK => CLK, Q => 
                           n_1579, QN => n20834);
   REGISTERS_reg_6_11_inst : DFF_X1 port map( D => n6671, CK => CLK, Q => 
                           n_1580, QN => n20835);
   REGISTERS_reg_6_10_inst : DFF_X1 port map( D => n6670, CK => CLK, Q => 
                           n_1581, QN => n20836);
   REGISTERS_reg_6_9_inst : DFF_X1 port map( D => n6669, CK => CLK, Q => n_1582
                           , QN => n20837);
   REGISTERS_reg_6_8_inst : DFF_X1 port map( D => n6668, CK => CLK, Q => n_1583
                           , QN => n20838);
   REGISTERS_reg_6_7_inst : DFF_X1 port map( D => n6667, CK => CLK, Q => n_1584
                           , QN => n20839);
   REGISTERS_reg_6_6_inst : DFF_X1 port map( D => n6666, CK => CLK, Q => n_1585
                           , QN => n20840);
   REGISTERS_reg_6_5_inst : DFF_X1 port map( D => n6665, CK => CLK, Q => n_1586
                           , QN => n20841);
   REGISTERS_reg_6_4_inst : DFF_X1 port map( D => n6664, CK => CLK, Q => n_1587
                           , QN => n20842);
   REGISTERS_reg_6_3_inst : DFF_X1 port map( D => n6663, CK => CLK, Q => n_1588
                           , QN => n20843);
   REGISTERS_reg_6_2_inst : DFF_X1 port map( D => n6662, CK => CLK, Q => n_1589
                           , QN => n20844);
   REGISTERS_reg_6_1_inst : DFF_X1 port map( D => n6661, CK => CLK, Q => n_1590
                           , QN => n20845);
   REGISTERS_reg_6_0_inst : DFF_X1 port map( D => n6660, CK => CLK, Q => n_1591
                           , QN => n20846);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n6939, CK => CLK, Q => 
                           n_1592, QN => n20422);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n6938, CK => CLK, Q => 
                           n_1593, QN => n20423);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n6937, CK => CLK, Q => 
                           n_1594, QN => n20424);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n6936, CK => CLK, Q => 
                           n_1595, QN => n20425);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n6935, CK => CLK, Q => 
                           n_1596, QN => n20426);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n6934, CK => CLK, Q => 
                           n_1597, QN => n20427);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n6933, CK => CLK, Q => 
                           n_1598, QN => n20428);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n6932, CK => CLK, Q => 
                           n_1599, QN => n20429);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n6931, CK => CLK, Q => 
                           n_1600, QN => n20430);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n6930, CK => CLK, Q => 
                           n_1601, QN => n20431);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n6929, CK => CLK, Q => 
                           n_1602, QN => n20432);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n6928, CK => CLK, Q => 
                           n_1603, QN => n20433);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n6927, CK => CLK, Q => 
                           n_1604, QN => n20434);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n6926, CK => CLK, Q => 
                           n_1605, QN => n20435);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n6925, CK => CLK, Q => n_1606
                           , QN => n20436);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n6924, CK => CLK, Q => n_1607
                           , QN => n20437);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n6923, CK => CLK, Q => n_1608
                           , QN => n20438);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n6922, CK => CLK, Q => n_1609
                           , QN => n20439);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n6921, CK => CLK, Q => n_1610
                           , QN => n20440);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n6920, CK => CLK, Q => n_1611
                           , QN => n20441);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n6919, CK => CLK, Q => n_1612
                           , QN => n20442);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n6918, CK => CLK, Q => n_1613
                           , QN => n20443);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n6917, CK => CLK, Q => n_1614
                           , QN => n20444);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n6916, CK => CLK, Q => n_1615
                           , QN => n20445);
   REGISTERS_reg_4_63_inst : DFF_X1 port map( D => n6851, CK => CLK, Q => 
                           n17661, QN => n19332);
   REGISTERS_reg_4_62_inst : DFF_X1 port map( D => n6850, CK => CLK, Q => 
                           n17658, QN => n19333);
   REGISTERS_reg_4_61_inst : DFF_X1 port map( D => n6849, CK => CLK, Q => 
                           n17655, QN => n19334);
   REGISTERS_reg_4_60_inst : DFF_X1 port map( D => n6848, CK => CLK, Q => 
                           n17652, QN => n19335);
   REGISTERS_reg_21_63_inst : DFF_X1 port map( D => n5763, CK => CLK, Q => 
                           n8478, QN => n20543);
   REGISTERS_reg_21_62_inst : DFF_X1 port map( D => n5762, CK => CLK, Q => 
                           n8479, QN => n20544);
   REGISTERS_reg_21_61_inst : DFF_X1 port map( D => n5761, CK => CLK, Q => 
                           n8480, QN => n20545);
   REGISTERS_reg_21_60_inst : DFF_X1 port map( D => n5760, CK => CLK, Q => 
                           n8481, QN => n20546);
   REGISTERS_reg_16_63_inst : DFF_X1 port map( D => n6083, CK => CLK, Q => 
                           n8606, QN => n20518);
   REGISTERS_reg_16_62_inst : DFF_X1 port map( D => n6082, CK => CLK, Q => 
                           n8607, QN => n20519);
   REGISTERS_reg_16_61_inst : DFF_X1 port map( D => n6081, CK => CLK, Q => 
                           n8608, QN => n20520);
   REGISTERS_reg_16_60_inst : DFF_X1 port map( D => n6080, CK => CLK, Q => 
                           n8609, QN => n20521);
   REGISTERS_reg_9_63_inst : DFF_X1 port map( D => n6531, CK => CLK, Q => 
                           n23967, QN => n20254);
   REGISTERS_reg_9_62_inst : DFF_X1 port map( D => n6530, CK => CLK, Q => 
                           n23966, QN => n20255);
   REGISTERS_reg_9_61_inst : DFF_X1 port map( D => n6529, CK => CLK, Q => 
                           n23965, QN => n20256);
   REGISTERS_reg_9_60_inst : DFF_X1 port map( D => n6528, CK => CLK, Q => 
                           n23964, QN => n20257);
   REGISTERS_reg_0_63_inst : DFF_X1 port map( D => n7107, CK => CLK, Q => 
                           n17660, QN => n19268);
   REGISTERS_reg_0_62_inst : DFF_X1 port map( D => n7106, CK => CLK, Q => 
                           n17657, QN => n19269);
   REGISTERS_reg_0_61_inst : DFF_X1 port map( D => n7105, CK => CLK, Q => 
                           n17654, QN => n19270);
   REGISTERS_reg_0_60_inst : DFF_X1 port map( D => n7104, CK => CLK, Q => 
                           n17651, QN => n19271);
   REGISTERS_reg_4_59_inst : DFF_X1 port map( D => n6847, CK => CLK, Q => 
                           n17649, QN => n19336);
   REGISTERS_reg_4_58_inst : DFF_X1 port map( D => n6846, CK => CLK, Q => 
                           n17646, QN => n19337);
   REGISTERS_reg_4_57_inst : DFF_X1 port map( D => n6845, CK => CLK, Q => 
                           n17643, QN => n19338);
   REGISTERS_reg_4_56_inst : DFF_X1 port map( D => n6844, CK => CLK, Q => 
                           n17640, QN => n19339);
   REGISTERS_reg_4_55_inst : DFF_X1 port map( D => n6843, CK => CLK, Q => 
                           n17637, QN => n19340);
   REGISTERS_reg_4_54_inst : DFF_X1 port map( D => n6842, CK => CLK, Q => 
                           n17634, QN => n19341);
   REGISTERS_reg_4_53_inst : DFF_X1 port map( D => n6841, CK => CLK, Q => 
                           n17631, QN => n19342);
   REGISTERS_reg_4_52_inst : DFF_X1 port map( D => n6840, CK => CLK, Q => 
                           n17628, QN => n19343);
   REGISTERS_reg_4_51_inst : DFF_X1 port map( D => n6839, CK => CLK, Q => 
                           n17538, QN => n19344);
   REGISTERS_reg_4_50_inst : DFF_X1 port map( D => n6838, CK => CLK, Q => 
                           n17535, QN => n19345);
   REGISTERS_reg_4_49_inst : DFF_X1 port map( D => n6837, CK => CLK, Q => 
                           n17532, QN => n19346);
   REGISTERS_reg_4_48_inst : DFF_X1 port map( D => n6836, CK => CLK, Q => 
                           n17529, QN => n19347);
   REGISTERS_reg_4_47_inst : DFF_X1 port map( D => n6835, CK => CLK, Q => 
                           n17526, QN => n19348);
   REGISTERS_reg_4_46_inst : DFF_X1 port map( D => n6834, CK => CLK, Q => 
                           n17523, QN => n19349);
   REGISTERS_reg_4_45_inst : DFF_X1 port map( D => n6833, CK => CLK, Q => 
                           n17520, QN => n19350);
   REGISTERS_reg_4_44_inst : DFF_X1 port map( D => n6832, CK => CLK, Q => 
                           n17517, QN => n19351);
   REGISTERS_reg_4_43_inst : DFF_X1 port map( D => n6831, CK => CLK, Q => 
                           n17514, QN => n19352);
   REGISTERS_reg_4_42_inst : DFF_X1 port map( D => n6830, CK => CLK, Q => 
                           n17511, QN => n19353);
   REGISTERS_reg_4_41_inst : DFF_X1 port map( D => n6829, CK => CLK, Q => 
                           n17508, QN => n19354);
   REGISTERS_reg_4_40_inst : DFF_X1 port map( D => n6828, CK => CLK, Q => 
                           n17505, QN => n19355);
   REGISTERS_reg_4_39_inst : DFF_X1 port map( D => n6827, CK => CLK, Q => 
                           n17502, QN => n19356);
   REGISTERS_reg_4_38_inst : DFF_X1 port map( D => n6826, CK => CLK, Q => 
                           n17499, QN => n19357);
   REGISTERS_reg_4_37_inst : DFF_X1 port map( D => n6825, CK => CLK, Q => 
                           n17496, QN => n19358);
   REGISTERS_reg_4_36_inst : DFF_X1 port map( D => n6824, CK => CLK, Q => 
                           n17493, QN => n19359);
   REGISTERS_reg_4_35_inst : DFF_X1 port map( D => n6823, CK => CLK, Q => 
                           n17490, QN => n19360);
   REGISTERS_reg_4_34_inst : DFF_X1 port map( D => n6822, CK => CLK, Q => 
                           n17487, QN => n19361);
   REGISTERS_reg_4_33_inst : DFF_X1 port map( D => n6821, CK => CLK, Q => 
                           n17484, QN => n19362);
   REGISTERS_reg_4_32_inst : DFF_X1 port map( D => n6820, CK => CLK, Q => 
                           n17481, QN => n19363);
   REGISTERS_reg_4_31_inst : DFF_X1 port map( D => n6819, CK => CLK, Q => 
                           n17478, QN => n19364);
   REGISTERS_reg_4_30_inst : DFF_X1 port map( D => n6818, CK => CLK, Q => 
                           n17475, QN => n19365);
   REGISTERS_reg_4_29_inst : DFF_X1 port map( D => n6817, CK => CLK, Q => 
                           n17472, QN => n19366);
   REGISTERS_reg_4_28_inst : DFF_X1 port map( D => n6816, CK => CLK, Q => 
                           n17625, QN => n19367);
   REGISTERS_reg_4_27_inst : DFF_X1 port map( D => n6815, CK => CLK, Q => 
                           n17622, QN => n19368);
   REGISTERS_reg_4_26_inst : DFF_X1 port map( D => n6814, CK => CLK, Q => 
                           n17619, QN => n19369);
   REGISTERS_reg_4_25_inst : DFF_X1 port map( D => n6813, CK => CLK, Q => 
                           n17616, QN => n19370);
   REGISTERS_reg_4_24_inst : DFF_X1 port map( D => n6812, CK => CLK, Q => 
                           n17613, QN => n19371);
   REGISTERS_reg_21_59_inst : DFF_X1 port map( D => n5759, CK => CLK, Q => 
                           n8482, QN => n21015);
   REGISTERS_reg_21_58_inst : DFF_X1 port map( D => n5758, CK => CLK, Q => 
                           n8483, QN => n21016);
   REGISTERS_reg_21_57_inst : DFF_X1 port map( D => n5757, CK => CLK, Q => 
                           n8484, QN => n21017);
   REGISTERS_reg_21_56_inst : DFF_X1 port map( D => n5756, CK => CLK, Q => 
                           n8485, QN => n21018);
   REGISTERS_reg_21_55_inst : DFF_X1 port map( D => n5755, CK => CLK, Q => 
                           n8486, QN => n21019);
   REGISTERS_reg_21_54_inst : DFF_X1 port map( D => n5754, CK => CLK, Q => 
                           n8487, QN => n21020);
   REGISTERS_reg_21_53_inst : DFF_X1 port map( D => n5753, CK => CLK, Q => 
                           n8488, QN => n21021);
   REGISTERS_reg_21_52_inst : DFF_X1 port map( D => n5752, CK => CLK, Q => 
                           n8489, QN => n21022);
   REGISTERS_reg_21_51_inst : DFF_X1 port map( D => n5751, CK => CLK, Q => 
                           n8490, QN => n21023);
   REGISTERS_reg_21_50_inst : DFF_X1 port map( D => n5750, CK => CLK, Q => 
                           n8491, QN => n21024);
   REGISTERS_reg_21_49_inst : DFF_X1 port map( D => n5749, CK => CLK, Q => 
                           n8492, QN => n21025);
   REGISTERS_reg_21_48_inst : DFF_X1 port map( D => n5748, CK => CLK, Q => 
                           n8493, QN => n21026);
   REGISTERS_reg_21_47_inst : DFF_X1 port map( D => n5747, CK => CLK, Q => 
                           n8494, QN => n21027);
   REGISTERS_reg_21_46_inst : DFF_X1 port map( D => n5746, CK => CLK, Q => 
                           n8495, QN => n21028);
   REGISTERS_reg_21_45_inst : DFF_X1 port map( D => n5745, CK => CLK, Q => 
                           n8496, QN => n21029);
   REGISTERS_reg_21_44_inst : DFF_X1 port map( D => n5744, CK => CLK, Q => 
                           n8497, QN => n21030);
   REGISTERS_reg_21_43_inst : DFF_X1 port map( D => n5743, CK => CLK, Q => 
                           n8498, QN => n21031);
   REGISTERS_reg_21_42_inst : DFF_X1 port map( D => n5742, CK => CLK, Q => 
                           n8499, QN => n21032);
   REGISTERS_reg_21_41_inst : DFF_X1 port map( D => n5741, CK => CLK, Q => 
                           n8500, QN => n21033);
   REGISTERS_reg_21_40_inst : DFF_X1 port map( D => n5740, CK => CLK, Q => 
                           n8501, QN => n21034);
   REGISTERS_reg_21_39_inst : DFF_X1 port map( D => n5739, CK => CLK, Q => 
                           n8502, QN => n21035);
   REGISTERS_reg_21_38_inst : DFF_X1 port map( D => n5738, CK => CLK, Q => 
                           n8503, QN => n21036);
   REGISTERS_reg_21_37_inst : DFF_X1 port map( D => n5737, CK => CLK, Q => 
                           n8504, QN => n21037);
   REGISTERS_reg_21_36_inst : DFF_X1 port map( D => n5736, CK => CLK, Q => 
                           n8505, QN => n21038);
   REGISTERS_reg_21_35_inst : DFF_X1 port map( D => n5735, CK => CLK, Q => 
                           n8506, QN => n21039);
   REGISTERS_reg_21_34_inst : DFF_X1 port map( D => n5734, CK => CLK, Q => 
                           n8507, QN => n21040);
   REGISTERS_reg_21_33_inst : DFF_X1 port map( D => n5733, CK => CLK, Q => 
                           n8508, QN => n21041);
   REGISTERS_reg_21_32_inst : DFF_X1 port map( D => n5732, CK => CLK, Q => 
                           n8509, QN => n21042);
   REGISTERS_reg_21_31_inst : DFF_X1 port map( D => n5731, CK => CLK, Q => 
                           n8510, QN => n21043);
   REGISTERS_reg_21_30_inst : DFF_X1 port map( D => n5730, CK => CLK, Q => 
                           n8511, QN => n21044);
   REGISTERS_reg_21_29_inst : DFF_X1 port map( D => n5729, CK => CLK, Q => 
                           n8512, QN => n21045);
   REGISTERS_reg_21_28_inst : DFF_X1 port map( D => n5728, CK => CLK, Q => 
                           n8513, QN => n21046);
   REGISTERS_reg_21_27_inst : DFF_X1 port map( D => n5727, CK => CLK, Q => 
                           n8514, QN => n21047);
   REGISTERS_reg_21_26_inst : DFF_X1 port map( D => n5726, CK => CLK, Q => 
                           n8515, QN => n21048);
   REGISTERS_reg_21_25_inst : DFF_X1 port map( D => n5725, CK => CLK, Q => 
                           n8516, QN => n21049);
   REGISTERS_reg_21_24_inst : DFF_X1 port map( D => n5724, CK => CLK, Q => 
                           n8517, QN => n21050);
   REGISTERS_reg_4_23_inst : DFF_X1 port map( D => n6811, CK => CLK, Q => 
                           n17610, QN => n19372);
   REGISTERS_reg_4_22_inst : DFF_X1 port map( D => n6810, CK => CLK, Q => 
                           n17607, QN => n19373);
   REGISTERS_reg_4_21_inst : DFF_X1 port map( D => n6809, CK => CLK, Q => 
                           n17604, QN => n19374);
   REGISTERS_reg_4_20_inst : DFF_X1 port map( D => n6808, CK => CLK, Q => 
                           n17601, QN => n19375);
   REGISTERS_reg_4_19_inst : DFF_X1 port map( D => n6807, CK => CLK, Q => 
                           n17598, QN => n19376);
   REGISTERS_reg_4_18_inst : DFF_X1 port map( D => n6806, CK => CLK, Q => 
                           n17595, QN => n19377);
   REGISTERS_reg_4_17_inst : DFF_X1 port map( D => n6805, CK => CLK, Q => 
                           n17592, QN => n19378);
   REGISTERS_reg_4_16_inst : DFF_X1 port map( D => n6804, CK => CLK, Q => 
                           n17589, QN => n19379);
   REGISTERS_reg_4_15_inst : DFF_X1 port map( D => n6803, CK => CLK, Q => 
                           n17586, QN => n19380);
   REGISTERS_reg_4_14_inst : DFF_X1 port map( D => n6802, CK => CLK, Q => 
                           n17583, QN => n19381);
   REGISTERS_reg_4_13_inst : DFF_X1 port map( D => n6801, CK => CLK, Q => 
                           n17580, QN => n19382);
   REGISTERS_reg_4_12_inst : DFF_X1 port map( D => n6800, CK => CLK, Q => 
                           n17577, QN => n19383);
   REGISTERS_reg_4_11_inst : DFF_X1 port map( D => n6799, CK => CLK, Q => 
                           n17574, QN => n19384);
   REGISTERS_reg_4_10_inst : DFF_X1 port map( D => n6798, CK => CLK, Q => 
                           n17571, QN => n19385);
   REGISTERS_reg_4_9_inst : DFF_X1 port map( D => n6797, CK => CLK, Q => n17568
                           , QN => n19386);
   REGISTERS_reg_4_8_inst : DFF_X1 port map( D => n6796, CK => CLK, Q => n17565
                           , QN => n19387);
   REGISTERS_reg_4_7_inst : DFF_X1 port map( D => n6795, CK => CLK, Q => n17562
                           , QN => n19388);
   REGISTERS_reg_4_6_inst : DFF_X1 port map( D => n6794, CK => CLK, Q => n17559
                           , QN => n19389);
   REGISTERS_reg_4_5_inst : DFF_X1 port map( D => n6793, CK => CLK, Q => n17556
                           , QN => n19390);
   REGISTERS_reg_4_4_inst : DFF_X1 port map( D => n6792, CK => CLK, Q => n17553
                           , QN => n19391);
   REGISTERS_reg_4_3_inst : DFF_X1 port map( D => n6791, CK => CLK, Q => n17550
                           , QN => n19392);
   REGISTERS_reg_4_2_inst : DFF_X1 port map( D => n6790, CK => CLK, Q => n17547
                           , QN => n19393);
   REGISTERS_reg_4_1_inst : DFF_X1 port map( D => n6789, CK => CLK, Q => n17544
                           , QN => n19394);
   REGISTERS_reg_4_0_inst : DFF_X1 port map( D => n6788, CK => CLK, Q => n17541
                           , QN => n19395);
   REGISTERS_reg_12_63_inst : DFF_X1 port map( D => n6339, CK => CLK, Q => 
                           n8286, QN => n20531);
   REGISTERS_reg_12_62_inst : DFF_X1 port map( D => n6338, CK => CLK, Q => 
                           n8287, QN => n20532);
   REGISTERS_reg_12_61_inst : DFF_X1 port map( D => n6337, CK => CLK, Q => 
                           n8288, QN => n20533);
   REGISTERS_reg_12_60_inst : DFF_X1 port map( D => n6336, CK => CLK, Q => 
                           n8289, QN => n20534);
   REGISTERS_reg_8_63_inst : DFF_X1 port map( D => n6595, CK => CLK, Q => n8030
                           , QN => n20535);
   REGISTERS_reg_8_62_inst : DFF_X1 port map( D => n6594, CK => CLK, Q => n8031
                           , QN => n20536);
   REGISTERS_reg_8_61_inst : DFF_X1 port map( D => n6593, CK => CLK, Q => n8032
                           , QN => n20537);
   REGISTERS_reg_8_60_inst : DFF_X1 port map( D => n6592, CK => CLK, Q => n8033
                           , QN => n20538);
   REGISTERS_reg_21_23_inst : DFF_X1 port map( D => n5723, CK => CLK, Q => 
                           n8518, QN => n21123);
   REGISTERS_reg_21_22_inst : DFF_X1 port map( D => n5722, CK => CLK, Q => 
                           n8519, QN => n21124);
   REGISTERS_reg_21_21_inst : DFF_X1 port map( D => n5721, CK => CLK, Q => 
                           n8520, QN => n21125);
   REGISTERS_reg_21_20_inst : DFF_X1 port map( D => n5720, CK => CLK, Q => 
                           n8521, QN => n21126);
   REGISTERS_reg_21_19_inst : DFF_X1 port map( D => n5719, CK => CLK, Q => 
                           n8522, QN => n21127);
   REGISTERS_reg_21_18_inst : DFF_X1 port map( D => n5718, CK => CLK, Q => 
                           n8523, QN => n21128);
   REGISTERS_reg_21_17_inst : DFF_X1 port map( D => n5717, CK => CLK, Q => 
                           n8524, QN => n21129);
   REGISTERS_reg_21_16_inst : DFF_X1 port map( D => n5716, CK => CLK, Q => 
                           n8525, QN => n21130);
   REGISTERS_reg_21_15_inst : DFF_X1 port map( D => n5715, CK => CLK, Q => 
                           n8526, QN => n21131);
   REGISTERS_reg_21_14_inst : DFF_X1 port map( D => n5714, CK => CLK, Q => 
                           n8527, QN => n21132);
   REGISTERS_reg_21_13_inst : DFF_X1 port map( D => n5713, CK => CLK, Q => 
                           n8528, QN => n21133);
   REGISTERS_reg_21_12_inst : DFF_X1 port map( D => n5712, CK => CLK, Q => 
                           n8529, QN => n21134);
   REGISTERS_reg_21_11_inst : DFF_X1 port map( D => n5711, CK => CLK, Q => 
                           n8530, QN => n21135);
   REGISTERS_reg_21_10_inst : DFF_X1 port map( D => n5710, CK => CLK, Q => 
                           n8531, QN => n21136);
   REGISTERS_reg_21_9_inst : DFF_X1 port map( D => n5709, CK => CLK, Q => n8532
                           , QN => n21137);
   REGISTERS_reg_21_8_inst : DFF_X1 port map( D => n5708, CK => CLK, Q => n8533
                           , QN => n21138);
   REGISTERS_reg_21_7_inst : DFF_X1 port map( D => n5707, CK => CLK, Q => n8534
                           , QN => n21139);
   REGISTERS_reg_21_6_inst : DFF_X1 port map( D => n5706, CK => CLK, Q => n8535
                           , QN => n21140);
   REGISTERS_reg_21_5_inst : DFF_X1 port map( D => n5705, CK => CLK, Q => n8536
                           , QN => n21141);
   REGISTERS_reg_21_4_inst : DFF_X1 port map( D => n5704, CK => CLK, Q => n8537
                           , QN => n21142);
   REGISTERS_reg_21_3_inst : DFF_X1 port map( D => n5703, CK => CLK, Q => n8538
                           , QN => n21143);
   REGISTERS_reg_21_2_inst : DFF_X1 port map( D => n5702, CK => CLK, Q => n8539
                           , QN => n21144);
   REGISTERS_reg_21_1_inst : DFF_X1 port map( D => n5701, CK => CLK, Q => n8540
                           , QN => n21145);
   REGISTERS_reg_21_0_inst : DFF_X1 port map( D => n5700, CK => CLK, Q => n8541
                           , QN => n21146);
   REGISTERS_reg_28_63_inst : DFF_X1 port map( D => n5315, CK => CLK, Q => 
                           n24031, QN => n20145);
   REGISTERS_reg_28_62_inst : DFF_X1 port map( D => n5314, CK => CLK, Q => 
                           n24030, QN => n20146);
   REGISTERS_reg_28_61_inst : DFF_X1 port map( D => n5313, CK => CLK, Q => 
                           n24029, QN => n20147);
   REGISTERS_reg_28_60_inst : DFF_X1 port map( D => n5312, CK => CLK, Q => 
                           n24028, QN => n20148);
   REGISTERS_reg_30_63_inst : DFF_X1 port map( D => n5187, CK => CLK, Q => 
                           n8670, QN => n20506);
   REGISTERS_reg_30_62_inst : DFF_X1 port map( D => n5186, CK => CLK, Q => 
                           n8671, QN => n20507);
   REGISTERS_reg_30_61_inst : DFF_X1 port map( D => n5185, CK => CLK, Q => 
                           n8672, QN => n20508);
   REGISTERS_reg_30_60_inst : DFF_X1 port map( D => n5184, CK => CLK, Q => 
                           n8673, QN => n20509);
   REGISTERS_reg_26_63_inst : DFF_X1 port map( D => n5443, CK => CLK, Q => 
                           n8350, QN => n20510);
   REGISTERS_reg_26_62_inst : DFF_X1 port map( D => n5442, CK => CLK, Q => 
                           n8351, QN => n20511);
   REGISTERS_reg_26_61_inst : DFF_X1 port map( D => n5441, CK => CLK, Q => 
                           n8352, QN => n20512);
   REGISTERS_reg_26_60_inst : DFF_X1 port map( D => n5440, CK => CLK, Q => 
                           n8353, QN => n20513);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n6981, CK => CLK, Q => n7708,
                           QN => n21147);
   REGISTERS_reg_16_59_inst : DFF_X1 port map( D => n6079, CK => CLK, Q => 
                           n8610, QN => n20655);
   REGISTERS_reg_16_58_inst : DFF_X1 port map( D => n6078, CK => CLK, Q => 
                           n8611, QN => n20656);
   REGISTERS_reg_16_57_inst : DFF_X1 port map( D => n6077, CK => CLK, Q => 
                           n8612, QN => n20657);
   REGISTERS_reg_16_56_inst : DFF_X1 port map( D => n6076, CK => CLK, Q => 
                           n8613, QN => n20658);
   REGISTERS_reg_16_55_inst : DFF_X1 port map( D => n6075, CK => CLK, Q => 
                           n8614, QN => n20659);
   REGISTERS_reg_16_54_inst : DFF_X1 port map( D => n6074, CK => CLK, Q => 
                           n8615, QN => n20660);
   REGISTERS_reg_16_53_inst : DFF_X1 port map( D => n6073, CK => CLK, Q => 
                           n8616, QN => n20661);
   REGISTERS_reg_16_52_inst : DFF_X1 port map( D => n6072, CK => CLK, Q => 
                           n8617, QN => n20662);
   REGISTERS_reg_16_51_inst : DFF_X1 port map( D => n6071, CK => CLK, Q => 
                           n8618, QN => n20663);
   REGISTERS_reg_16_50_inst : DFF_X1 port map( D => n6070, CK => CLK, Q => 
                           n8619, QN => n20664);
   REGISTERS_reg_16_49_inst : DFF_X1 port map( D => n6069, CK => CLK, Q => 
                           n8620, QN => n20665);
   REGISTERS_reg_16_48_inst : DFF_X1 port map( D => n6068, CK => CLK, Q => 
                           n8621, QN => n20666);
   REGISTERS_reg_16_47_inst : DFF_X1 port map( D => n6067, CK => CLK, Q => 
                           n8622, QN => n20667);
   REGISTERS_reg_16_46_inst : DFF_X1 port map( D => n6066, CK => CLK, Q => 
                           n8623, QN => n20668);
   REGISTERS_reg_16_45_inst : DFF_X1 port map( D => n6065, CK => CLK, Q => 
                           n8624, QN => n20669);
   REGISTERS_reg_16_44_inst : DFF_X1 port map( D => n6064, CK => CLK, Q => 
                           n8625, QN => n20670);
   REGISTERS_reg_16_43_inst : DFF_X1 port map( D => n6063, CK => CLK, Q => 
                           n8626, QN => n20671);
   REGISTERS_reg_16_42_inst : DFF_X1 port map( D => n6062, CK => CLK, Q => 
                           n8627, QN => n20672);
   REGISTERS_reg_16_41_inst : DFF_X1 port map( D => n6061, CK => CLK, Q => 
                           n8628, QN => n20673);
   REGISTERS_reg_16_40_inst : DFF_X1 port map( D => n6060, CK => CLK, Q => 
                           n8629, QN => n20674);
   REGISTERS_reg_16_39_inst : DFF_X1 port map( D => n6059, CK => CLK, Q => 
                           n8630, QN => n20675);
   REGISTERS_reg_16_38_inst : DFF_X1 port map( D => n6058, CK => CLK, Q => 
                           n8631, QN => n20676);
   REGISTERS_reg_16_37_inst : DFF_X1 port map( D => n6057, CK => CLK, Q => 
                           n8632, QN => n20677);
   REGISTERS_reg_16_36_inst : DFF_X1 port map( D => n6056, CK => CLK, Q => 
                           n8633, QN => n20678);
   REGISTERS_reg_16_35_inst : DFF_X1 port map( D => n6055, CK => CLK, Q => 
                           n8634, QN => n20679);
   REGISTERS_reg_16_34_inst : DFF_X1 port map( D => n6054, CK => CLK, Q => 
                           n8635, QN => n20680);
   REGISTERS_reg_16_33_inst : DFF_X1 port map( D => n6053, CK => CLK, Q => 
                           n8636, QN => n20681);
   REGISTERS_reg_16_32_inst : DFF_X1 port map( D => n6052, CK => CLK, Q => 
                           n8637, QN => n20682);
   REGISTERS_reg_16_31_inst : DFF_X1 port map( D => n6051, CK => CLK, Q => 
                           n8638, QN => n20683);
   REGISTERS_reg_16_30_inst : DFF_X1 port map( D => n6050, CK => CLK, Q => 
                           n8639, QN => n20684);
   REGISTERS_reg_16_29_inst : DFF_X1 port map( D => n6049, CK => CLK, Q => 
                           n8640, QN => n20685);
   REGISTERS_reg_16_28_inst : DFF_X1 port map( D => n6048, CK => CLK, Q => 
                           n8641, QN => n20686);
   REGISTERS_reg_16_27_inst : DFF_X1 port map( D => n6047, CK => CLK, Q => 
                           n8642, QN => n20687);
   REGISTERS_reg_16_26_inst : DFF_X1 port map( D => n6046, CK => CLK, Q => 
                           n8643, QN => n20688);
   REGISTERS_reg_16_25_inst : DFF_X1 port map( D => n6045, CK => CLK, Q => 
                           n8644, QN => n20689);
   REGISTERS_reg_16_24_inst : DFF_X1 port map( D => n6044, CK => CLK, Q => 
                           n8645, QN => n20690);
   REGISTERS_reg_9_59_inst : DFF_X1 port map( D => n6527, CK => CLK, Q => 
                           n23963, QN => n20302);
   REGISTERS_reg_9_58_inst : DFF_X1 port map( D => n6526, CK => CLK, Q => 
                           n23962, QN => n20303);
   REGISTERS_reg_9_57_inst : DFF_X1 port map( D => n6525, CK => CLK, Q => 
                           n23961, QN => n20304);
   REGISTERS_reg_9_56_inst : DFF_X1 port map( D => n6524, CK => CLK, Q => 
                           n23960, QN => n20305);
   REGISTERS_reg_9_55_inst : DFF_X1 port map( D => n6523, CK => CLK, Q => 
                           n23959, QN => n20306);
   REGISTERS_reg_9_54_inst : DFF_X1 port map( D => n6522, CK => CLK, Q => 
                           n23958, QN => n20307);
   REGISTERS_reg_9_53_inst : DFF_X1 port map( D => n6521, CK => CLK, Q => 
                           n23957, QN => n20308);
   REGISTERS_reg_9_52_inst : DFF_X1 port map( D => n6520, CK => CLK, Q => 
                           n23956, QN => n20309);
   REGISTERS_reg_9_51_inst : DFF_X1 port map( D => n6519, CK => CLK, Q => 
                           n23955, QN => n20310);
   REGISTERS_reg_9_50_inst : DFF_X1 port map( D => n6518, CK => CLK, Q => 
                           n23954, QN => n20311);
   REGISTERS_reg_9_49_inst : DFF_X1 port map( D => n6517, CK => CLK, Q => 
                           n23953, QN => n20312);
   REGISTERS_reg_9_48_inst : DFF_X1 port map( D => n6516, CK => CLK, Q => 
                           n23952, QN => n20313);
   REGISTERS_reg_9_47_inst : DFF_X1 port map( D => n6515, CK => CLK, Q => 
                           n23950, QN => n20314);
   REGISTERS_reg_9_46_inst : DFF_X1 port map( D => n6514, CK => CLK, Q => 
                           n23948, QN => n20315);
   REGISTERS_reg_9_45_inst : DFF_X1 port map( D => n6513, CK => CLK, Q => 
                           n23946, QN => n20316);
   REGISTERS_reg_9_44_inst : DFF_X1 port map( D => n6512, CK => CLK, Q => 
                           n23944, QN => n20317);
   REGISTERS_reg_9_43_inst : DFF_X1 port map( D => n6511, CK => CLK, Q => 
                           n23942, QN => n20318);
   REGISTERS_reg_9_42_inst : DFF_X1 port map( D => n6510, CK => CLK, Q => 
                           n23940, QN => n20319);
   REGISTERS_reg_9_41_inst : DFF_X1 port map( D => n6509, CK => CLK, Q => 
                           n23938, QN => n20320);
   REGISTERS_reg_9_40_inst : DFF_X1 port map( D => n6508, CK => CLK, Q => 
                           n23936, QN => n20321);
   REGISTERS_reg_9_39_inst : DFF_X1 port map( D => n6507, CK => CLK, Q => 
                           n23934, QN => n20322);
   REGISTERS_reg_9_38_inst : DFF_X1 port map( D => n6506, CK => CLK, Q => 
                           n23932, QN => n20323);
   REGISTERS_reg_9_37_inst : DFF_X1 port map( D => n6505, CK => CLK, Q => 
                           n23930, QN => n20324);
   REGISTERS_reg_9_36_inst : DFF_X1 port map( D => n6504, CK => CLK, Q => 
                           n23928, QN => n20325);
   REGISTERS_reg_9_35_inst : DFF_X1 port map( D => n6503, CK => CLK, Q => 
                           n23926, QN => n20326);
   REGISTERS_reg_9_34_inst : DFF_X1 port map( D => n6502, CK => CLK, Q => 
                           n23924, QN => n20327);
   REGISTERS_reg_9_33_inst : DFF_X1 port map( D => n6501, CK => CLK, Q => 
                           n23922, QN => n20328);
   REGISTERS_reg_9_32_inst : DFF_X1 port map( D => n6500, CK => CLK, Q => 
                           n23920, QN => n20329);
   REGISTERS_reg_9_31_inst : DFF_X1 port map( D => n6499, CK => CLK, Q => 
                           n23918, QN => n20330);
   REGISTERS_reg_9_30_inst : DFF_X1 port map( D => n6498, CK => CLK, Q => 
                           n23916, QN => n20331);
   REGISTERS_reg_9_29_inst : DFF_X1 port map( D => n6497, CK => CLK, Q => 
                           n23914, QN => n20332);
   REGISTERS_reg_9_28_inst : DFF_X1 port map( D => n6496, CK => CLK, Q => 
                           n23912, QN => n20333);
   REGISTERS_reg_9_27_inst : DFF_X1 port map( D => n6495, CK => CLK, Q => 
                           n23910, QN => n20334);
   REGISTERS_reg_9_26_inst : DFF_X1 port map( D => n6494, CK => CLK, Q => 
                           n23908, QN => n20335);
   REGISTERS_reg_9_25_inst : DFF_X1 port map( D => n6493, CK => CLK, Q => 
                           n23906, QN => n20336);
   REGISTERS_reg_9_24_inst : DFF_X1 port map( D => n6492, CK => CLK, Q => 
                           n23904, QN => n20337);
   REGISTERS_reg_16_23_inst : DFF_X1 port map( D => n6043, CK => CLK, Q => 
                           n8646, QN => n20799);
   REGISTERS_reg_16_22_inst : DFF_X1 port map( D => n6042, CK => CLK, Q => 
                           n8647, QN => n20800);
   REGISTERS_reg_16_21_inst : DFF_X1 port map( D => n6041, CK => CLK, Q => 
                           n8648, QN => n20801);
   REGISTERS_reg_16_20_inst : DFF_X1 port map( D => n6040, CK => CLK, Q => 
                           n8649, QN => n20802);
   REGISTERS_reg_16_19_inst : DFF_X1 port map( D => n6039, CK => CLK, Q => 
                           n8650, QN => n20803);
   REGISTERS_reg_16_18_inst : DFF_X1 port map( D => n6038, CK => CLK, Q => 
                           n8651, QN => n20804);
   REGISTERS_reg_16_17_inst : DFF_X1 port map( D => n6037, CK => CLK, Q => 
                           n8652, QN => n20805);
   REGISTERS_reg_16_16_inst : DFF_X1 port map( D => n6036, CK => CLK, Q => 
                           n8653, QN => n20806);
   REGISTERS_reg_16_15_inst : DFF_X1 port map( D => n6035, CK => CLK, Q => 
                           n8654, QN => n20807);
   REGISTERS_reg_16_14_inst : DFF_X1 port map( D => n6034, CK => CLK, Q => 
                           n8655, QN => n20808);
   REGISTERS_reg_16_13_inst : DFF_X1 port map( D => n6033, CK => CLK, Q => 
                           n8656, QN => n20809);
   REGISTERS_reg_16_12_inst : DFF_X1 port map( D => n6032, CK => CLK, Q => 
                           n8657, QN => n20810);
   REGISTERS_reg_16_11_inst : DFF_X1 port map( D => n6031, CK => CLK, Q => 
                           n8658, QN => n20811);
   REGISTERS_reg_16_10_inst : DFF_X1 port map( D => n6030, CK => CLK, Q => 
                           n8659, QN => n20812);
   REGISTERS_reg_16_9_inst : DFF_X1 port map( D => n6029, CK => CLK, Q => n8660
                           , QN => n20813);
   REGISTERS_reg_16_8_inst : DFF_X1 port map( D => n6028, CK => CLK, Q => n8661
                           , QN => n20814);
   REGISTERS_reg_16_7_inst : DFF_X1 port map( D => n6027, CK => CLK, Q => n8662
                           , QN => n20815);
   REGISTERS_reg_16_6_inst : DFF_X1 port map( D => n6026, CK => CLK, Q => n8663
                           , QN => n20816);
   REGISTERS_reg_16_5_inst : DFF_X1 port map( D => n6025, CK => CLK, Q => n8664
                           , QN => n20817);
   REGISTERS_reg_16_4_inst : DFF_X1 port map( D => n6024, CK => CLK, Q => n8665
                           , QN => n20818);
   REGISTERS_reg_16_3_inst : DFF_X1 port map( D => n6023, CK => CLK, Q => n8666
                           , QN => n20819);
   REGISTERS_reg_16_2_inst : DFF_X1 port map( D => n6022, CK => CLK, Q => n8667
                           , QN => n20820);
   REGISTERS_reg_16_1_inst : DFF_X1 port map( D => n6021, CK => CLK, Q => n8668
                           , QN => n20821);
   REGISTERS_reg_16_0_inst : DFF_X1 port map( D => n6020, CK => CLK, Q => n8669
                           , QN => n20822);
   REGISTERS_reg_0_59_inst : DFF_X1 port map( D => n7103, CK => CLK, Q => 
                           n17648, QN => n19272);
   REGISTERS_reg_0_58_inst : DFF_X1 port map( D => n7102, CK => CLK, Q => 
                           n17645, QN => n19273);
   REGISTERS_reg_0_57_inst : DFF_X1 port map( D => n7101, CK => CLK, Q => 
                           n17642, QN => n19274);
   REGISTERS_reg_0_56_inst : DFF_X1 port map( D => n7100, CK => CLK, Q => 
                           n17639, QN => n19275);
   REGISTERS_reg_0_55_inst : DFF_X1 port map( D => n7099, CK => CLK, Q => 
                           n17636, QN => n19276);
   REGISTERS_reg_0_54_inst : DFF_X1 port map( D => n7098, CK => CLK, Q => 
                           n17633, QN => n19277);
   REGISTERS_reg_0_53_inst : DFF_X1 port map( D => n7097, CK => CLK, Q => 
                           n17630, QN => n19278);
   REGISTERS_reg_0_52_inst : DFF_X1 port map( D => n7096, CK => CLK, Q => 
                           n17627, QN => n19279);
   REGISTERS_reg_0_51_inst : DFF_X1 port map( D => n7095, CK => CLK, Q => 
                           n17537, QN => n19280);
   REGISTERS_reg_0_50_inst : DFF_X1 port map( D => n7094, CK => CLK, Q => 
                           n17534, QN => n19281);
   REGISTERS_reg_0_49_inst : DFF_X1 port map( D => n7093, CK => CLK, Q => 
                           n17531, QN => n19282);
   REGISTERS_reg_0_48_inst : DFF_X1 port map( D => n7092, CK => CLK, Q => 
                           n17528, QN => n19283);
   REGISTERS_reg_0_47_inst : DFF_X1 port map( D => n7091, CK => CLK, Q => 
                           n17525, QN => n19284);
   REGISTERS_reg_0_46_inst : DFF_X1 port map( D => n7090, CK => CLK, Q => 
                           n17522, QN => n19285);
   REGISTERS_reg_0_45_inst : DFF_X1 port map( D => n7089, CK => CLK, Q => 
                           n17519, QN => n19286);
   REGISTERS_reg_0_44_inst : DFF_X1 port map( D => n7088, CK => CLK, Q => 
                           n17516, QN => n19287);
   REGISTERS_reg_0_43_inst : DFF_X1 port map( D => n7087, CK => CLK, Q => 
                           n17513, QN => n19288);
   REGISTERS_reg_0_42_inst : DFF_X1 port map( D => n7086, CK => CLK, Q => 
                           n17510, QN => n19289);
   REGISTERS_reg_0_41_inst : DFF_X1 port map( D => n7085, CK => CLK, Q => 
                           n17507, QN => n19290);
   REGISTERS_reg_0_40_inst : DFF_X1 port map( D => n7084, CK => CLK, Q => 
                           n17504, QN => n19291);
   REGISTERS_reg_0_39_inst : DFF_X1 port map( D => n7083, CK => CLK, Q => 
                           n17501, QN => n19292);
   REGISTERS_reg_0_38_inst : DFF_X1 port map( D => n7082, CK => CLK, Q => 
                           n17498, QN => n19293);
   REGISTERS_reg_0_37_inst : DFF_X1 port map( D => n7081, CK => CLK, Q => 
                           n17495, QN => n19294);
   REGISTERS_reg_0_36_inst : DFF_X1 port map( D => n7080, CK => CLK, Q => 
                           n17492, QN => n19295);
   REGISTERS_reg_0_35_inst : DFF_X1 port map( D => n7079, CK => CLK, Q => 
                           n17489, QN => n19296);
   REGISTERS_reg_0_34_inst : DFF_X1 port map( D => n7078, CK => CLK, Q => 
                           n17486, QN => n19297);
   REGISTERS_reg_0_33_inst : DFF_X1 port map( D => n7077, CK => CLK, Q => 
                           n17483, QN => n19298);
   REGISTERS_reg_0_32_inst : DFF_X1 port map( D => n7076, CK => CLK, Q => 
                           n17480, QN => n19299);
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n7075, CK => CLK, Q => 
                           n17477, QN => n19300);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n7074, CK => CLK, Q => 
                           n17474, QN => n19301);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n7073, CK => CLK, Q => 
                           n17471, QN => n19302);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n7072, CK => CLK, Q => 
                           n17624, QN => n19303);
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n7071, CK => CLK, Q => 
                           n17621, QN => n19304);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n7070, CK => CLK, Q => 
                           n17618, QN => n19305);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n7069, CK => CLK, Q => 
                           n17615, QN => n19306);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n7068, CK => CLK, Q => 
                           n17612, QN => n19307);
   REGISTERS_reg_9_23_inst : DFF_X1 port map( D => n6491, CK => CLK, Q => 
                           n23902, QN => n20398);
   REGISTERS_reg_9_22_inst : DFF_X1 port map( D => n6490, CK => CLK, Q => 
                           n23900, QN => n20399);
   REGISTERS_reg_9_21_inst : DFF_X1 port map( D => n6489, CK => CLK, Q => 
                           n23898, QN => n20400);
   REGISTERS_reg_9_20_inst : DFF_X1 port map( D => n6488, CK => CLK, Q => 
                           n23896, QN => n20401);
   REGISTERS_reg_9_19_inst : DFF_X1 port map( D => n6487, CK => CLK, Q => 
                           n23894, QN => n20402);
   REGISTERS_reg_9_18_inst : DFF_X1 port map( D => n6486, CK => CLK, Q => 
                           n23892, QN => n20403);
   REGISTERS_reg_9_17_inst : DFF_X1 port map( D => n6485, CK => CLK, Q => 
                           n23890, QN => n20404);
   REGISTERS_reg_9_16_inst : DFF_X1 port map( D => n6484, CK => CLK, Q => 
                           n23888, QN => n20405);
   REGISTERS_reg_9_15_inst : DFF_X1 port map( D => n6483, CK => CLK, Q => 
                           n23886, QN => n20406);
   REGISTERS_reg_9_14_inst : DFF_X1 port map( D => n6482, CK => CLK, Q => 
                           n23884, QN => n20407);
   REGISTERS_reg_9_13_inst : DFF_X1 port map( D => n6481, CK => CLK, Q => 
                           n23882, QN => n20408);
   REGISTERS_reg_9_12_inst : DFF_X1 port map( D => n6480, CK => CLK, Q => 
                           n23880, QN => n20409);
   REGISTERS_reg_9_11_inst : DFF_X1 port map( D => n6479, CK => CLK, Q => 
                           n23878, QN => n20410);
   REGISTERS_reg_9_10_inst : DFF_X1 port map( D => n6478, CK => CLK, Q => 
                           n23876, QN => n20411);
   REGISTERS_reg_9_9_inst : DFF_X1 port map( D => n6477, CK => CLK, Q => n23874
                           , QN => n20412);
   REGISTERS_reg_9_8_inst : DFF_X1 port map( D => n6476, CK => CLK, Q => n23872
                           , QN => n20413);
   REGISTERS_reg_9_7_inst : DFF_X1 port map( D => n6475, CK => CLK, Q => n23870
                           , QN => n20414);
   REGISTERS_reg_9_6_inst : DFF_X1 port map( D => n6474, CK => CLK, Q => n23868
                           , QN => n20415);
   REGISTERS_reg_9_5_inst : DFF_X1 port map( D => n6473, CK => CLK, Q => n23866
                           , QN => n20416);
   REGISTERS_reg_9_4_inst : DFF_X1 port map( D => n6472, CK => CLK, Q => n23864
                           , QN => n20417);
   REGISTERS_reg_9_3_inst : DFF_X1 port map( D => n6471, CK => CLK, Q => n23862
                           , QN => n20418);
   REGISTERS_reg_9_2_inst : DFF_X1 port map( D => n6470, CK => CLK, Q => n23860
                           , QN => n20419);
   REGISTERS_reg_9_1_inst : DFF_X1 port map( D => n6469, CK => CLK, Q => n23858
                           , QN => n20420);
   REGISTERS_reg_9_0_inst : DFF_X1 port map( D => n6468, CK => CLK, Q => n23856
                           , QN => n20421);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n7067, CK => CLK, Q => 
                           n17609, QN => n19308);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n7066, CK => CLK, Q => 
                           n17606, QN => n19309);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n7065, CK => CLK, Q => 
                           n17603, QN => n19310);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n7064, CK => CLK, Q => 
                           n17600, QN => n19311);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n7063, CK => CLK, Q => 
                           n17597, QN => n19312);
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n7062, CK => CLK, Q => 
                           n17594, QN => n19313);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n7061, CK => CLK, Q => 
                           n17591, QN => n19314);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n7060, CK => CLK, Q => 
                           n17588, QN => n19315);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n7059, CK => CLK, Q => 
                           n17585, QN => n19316);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n7058, CK => CLK, Q => 
                           n17582, QN => n19317);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n7057, CK => CLK, Q => 
                           n17579, QN => n19318);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n7056, CK => CLK, Q => 
                           n17576, QN => n19319);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n7055, CK => CLK, Q => 
                           n17573, QN => n19320);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n7054, CK => CLK, Q => 
                           n17570, QN => n19321);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n7053, CK => CLK, Q => n17567
                           , QN => n19322);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n7052, CK => CLK, Q => n17564
                           , QN => n19323);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n7051, CK => CLK, Q => n17561
                           , QN => n19324);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n7050, CK => CLK, Q => n17558
                           , QN => n19325);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n7049, CK => CLK, Q => n17555
                           , QN => n19326);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n7048, CK => CLK, Q => n17552
                           , QN => n19327);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n7047, CK => CLK, Q => n17549
                           , QN => n19328);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n7046, CK => CLK, Q => n17546
                           , QN => n19329);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n7045, CK => CLK, Q => n17543
                           , QN => n19330);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n7044, CK => CLK, Q => n17540
                           , QN => n19331);
   REGISTERS_reg_12_59_inst : DFF_X1 port map( D => n6335, CK => CLK, Q => 
                           n8290, QN => n20907);
   REGISTERS_reg_12_58_inst : DFF_X1 port map( D => n6334, CK => CLK, Q => 
                           n8291, QN => n20908);
   REGISTERS_reg_12_57_inst : DFF_X1 port map( D => n6333, CK => CLK, Q => 
                           n8292, QN => n20909);
   REGISTERS_reg_12_56_inst : DFF_X1 port map( D => n6332, CK => CLK, Q => 
                           n8293, QN => n20910);
   REGISTERS_reg_12_55_inst : DFF_X1 port map( D => n6331, CK => CLK, Q => 
                           n8294, QN => n20911);
   REGISTERS_reg_12_54_inst : DFF_X1 port map( D => n6330, CK => CLK, Q => 
                           n8295, QN => n20912);
   REGISTERS_reg_12_53_inst : DFF_X1 port map( D => n6329, CK => CLK, Q => 
                           n8296, QN => n20913);
   REGISTERS_reg_12_52_inst : DFF_X1 port map( D => n6328, CK => CLK, Q => 
                           n8297, QN => n20914);
   REGISTERS_reg_12_51_inst : DFF_X1 port map( D => n6327, CK => CLK, Q => 
                           n8298, QN => n20915);
   REGISTERS_reg_12_50_inst : DFF_X1 port map( D => n6326, CK => CLK, Q => 
                           n8299, QN => n20916);
   REGISTERS_reg_12_49_inst : DFF_X1 port map( D => n6325, CK => CLK, Q => 
                           n8300, QN => n20917);
   REGISTERS_reg_12_48_inst : DFF_X1 port map( D => n6324, CK => CLK, Q => 
                           n8301, QN => n20918);
   REGISTERS_reg_12_47_inst : DFF_X1 port map( D => n6323, CK => CLK, Q => 
                           n8302, QN => n20919);
   REGISTERS_reg_12_46_inst : DFF_X1 port map( D => n6322, CK => CLK, Q => 
                           n8303, QN => n20920);
   REGISTERS_reg_12_45_inst : DFF_X1 port map( D => n6321, CK => CLK, Q => 
                           n8304, QN => n20921);
   REGISTERS_reg_12_44_inst : DFF_X1 port map( D => n6320, CK => CLK, Q => 
                           n8305, QN => n20922);
   REGISTERS_reg_12_43_inst : DFF_X1 port map( D => n6319, CK => CLK, Q => 
                           n8306, QN => n20923);
   REGISTERS_reg_12_42_inst : DFF_X1 port map( D => n6318, CK => CLK, Q => 
                           n8307, QN => n20924);
   REGISTERS_reg_12_41_inst : DFF_X1 port map( D => n6317, CK => CLK, Q => 
                           n8308, QN => n20925);
   REGISTERS_reg_12_40_inst : DFF_X1 port map( D => n6316, CK => CLK, Q => 
                           n8309, QN => n20926);
   REGISTERS_reg_12_39_inst : DFF_X1 port map( D => n6315, CK => CLK, Q => 
                           n8310, QN => n20927);
   REGISTERS_reg_12_38_inst : DFF_X1 port map( D => n6314, CK => CLK, Q => 
                           n8311, QN => n20928);
   REGISTERS_reg_12_37_inst : DFF_X1 port map( D => n6313, CK => CLK, Q => 
                           n8312, QN => n20929);
   REGISTERS_reg_12_36_inst : DFF_X1 port map( D => n6312, CK => CLK, Q => 
                           n8313, QN => n20930);
   REGISTERS_reg_12_35_inst : DFF_X1 port map( D => n6311, CK => CLK, Q => 
                           n8314, QN => n20931);
   REGISTERS_reg_12_34_inst : DFF_X1 port map( D => n6310, CK => CLK, Q => 
                           n8315, QN => n20932);
   REGISTERS_reg_12_33_inst : DFF_X1 port map( D => n6309, CK => CLK, Q => 
                           n8316, QN => n20933);
   REGISTERS_reg_12_32_inst : DFF_X1 port map( D => n6308, CK => CLK, Q => 
                           n8317, QN => n20934);
   REGISTERS_reg_12_31_inst : DFF_X1 port map( D => n6307, CK => CLK, Q => 
                           n8318, QN => n20935);
   REGISTERS_reg_12_30_inst : DFF_X1 port map( D => n6306, CK => CLK, Q => 
                           n8319, QN => n20936);
   REGISTERS_reg_12_29_inst : DFF_X1 port map( D => n6305, CK => CLK, Q => 
                           n8320, QN => n20937);
   REGISTERS_reg_12_28_inst : DFF_X1 port map( D => n6304, CK => CLK, Q => 
                           n8321, QN => n20938);
   REGISTERS_reg_12_27_inst : DFF_X1 port map( D => n6303, CK => CLK, Q => 
                           n8322, QN => n20939);
   REGISTERS_reg_12_26_inst : DFF_X1 port map( D => n6302, CK => CLK, Q => 
                           n8323, QN => n20940);
   REGISTERS_reg_12_25_inst : DFF_X1 port map( D => n6301, CK => CLK, Q => 
                           n8324, QN => n20941);
   REGISTERS_reg_12_24_inst : DFF_X1 port map( D => n6300, CK => CLK, Q => 
                           n8325, QN => n20942);
   REGISTERS_reg_8_59_inst : DFF_X1 port map( D => n6591, CK => CLK, Q => n8034
                           , QN => n20943);
   REGISTERS_reg_8_58_inst : DFF_X1 port map( D => n6590, CK => CLK, Q => n8035
                           , QN => n20944);
   REGISTERS_reg_8_57_inst : DFF_X1 port map( D => n6589, CK => CLK, Q => n8036
                           , QN => n20945);
   REGISTERS_reg_8_56_inst : DFF_X1 port map( D => n6588, CK => CLK, Q => n8037
                           , QN => n20946);
   REGISTERS_reg_8_55_inst : DFF_X1 port map( D => n6587, CK => CLK, Q => n8038
                           , QN => n20947);
   REGISTERS_reg_8_54_inst : DFF_X1 port map( D => n6586, CK => CLK, Q => n8039
                           , QN => n20948);
   REGISTERS_reg_8_53_inst : DFF_X1 port map( D => n6585, CK => CLK, Q => n8040
                           , QN => n20949);
   REGISTERS_reg_8_52_inst : DFF_X1 port map( D => n6584, CK => CLK, Q => n8041
                           , QN => n20950);
   REGISTERS_reg_8_51_inst : DFF_X1 port map( D => n6583, CK => CLK, Q => n8042
                           , QN => n20951);
   REGISTERS_reg_8_50_inst : DFF_X1 port map( D => n6582, CK => CLK, Q => n8043
                           , QN => n20952);
   REGISTERS_reg_8_49_inst : DFF_X1 port map( D => n6581, CK => CLK, Q => n8044
                           , QN => n20953);
   REGISTERS_reg_8_48_inst : DFF_X1 port map( D => n6580, CK => CLK, Q => n8045
                           , QN => n20954);
   REGISTERS_reg_8_47_inst : DFF_X1 port map( D => n6579, CK => CLK, Q => n8046
                           , QN => n20955);
   REGISTERS_reg_8_46_inst : DFF_X1 port map( D => n6578, CK => CLK, Q => n8047
                           , QN => n20956);
   REGISTERS_reg_8_45_inst : DFF_X1 port map( D => n6577, CK => CLK, Q => n8048
                           , QN => n20957);
   REGISTERS_reg_8_44_inst : DFF_X1 port map( D => n6576, CK => CLK, Q => n8049
                           , QN => n20958);
   REGISTERS_reg_8_43_inst : DFF_X1 port map( D => n6575, CK => CLK, Q => n8050
                           , QN => n20959);
   REGISTERS_reg_8_42_inst : DFF_X1 port map( D => n6574, CK => CLK, Q => n8051
                           , QN => n20960);
   REGISTERS_reg_8_41_inst : DFF_X1 port map( D => n6573, CK => CLK, Q => n8052
                           , QN => n20961);
   REGISTERS_reg_8_40_inst : DFF_X1 port map( D => n6572, CK => CLK, Q => n8053
                           , QN => n20962);
   REGISTERS_reg_8_39_inst : DFF_X1 port map( D => n6571, CK => CLK, Q => n8054
                           , QN => n20963);
   REGISTERS_reg_8_38_inst : DFF_X1 port map( D => n6570, CK => CLK, Q => n8055
                           , QN => n20964);
   REGISTERS_reg_8_37_inst : DFF_X1 port map( D => n6569, CK => CLK, Q => n8056
                           , QN => n20965);
   REGISTERS_reg_8_36_inst : DFF_X1 port map( D => n6568, CK => CLK, Q => n8057
                           , QN => n20966);
   REGISTERS_reg_8_35_inst : DFF_X1 port map( D => n6567, CK => CLK, Q => n8058
                           , QN => n20967);
   REGISTERS_reg_8_34_inst : DFF_X1 port map( D => n6566, CK => CLK, Q => n8059
                           , QN => n20968);
   REGISTERS_reg_8_33_inst : DFF_X1 port map( D => n6565, CK => CLK, Q => n8060
                           , QN => n20969);
   REGISTERS_reg_8_32_inst : DFF_X1 port map( D => n6564, CK => CLK, Q => n8061
                           , QN => n20970);
   REGISTERS_reg_8_31_inst : DFF_X1 port map( D => n6563, CK => CLK, Q => n8062
                           , QN => n20971);
   REGISTERS_reg_8_30_inst : DFF_X1 port map( D => n6562, CK => CLK, Q => n8063
                           , QN => n20972);
   REGISTERS_reg_8_29_inst : DFF_X1 port map( D => n6561, CK => CLK, Q => n8064
                           , QN => n20973);
   REGISTERS_reg_8_28_inst : DFF_X1 port map( D => n6560, CK => CLK, Q => n8065
                           , QN => n20974);
   REGISTERS_reg_8_27_inst : DFF_X1 port map( D => n6559, CK => CLK, Q => n8066
                           , QN => n20975);
   REGISTERS_reg_8_26_inst : DFF_X1 port map( D => n6558, CK => CLK, Q => n8067
                           , QN => n20976);
   REGISTERS_reg_8_25_inst : DFF_X1 port map( D => n6557, CK => CLK, Q => n8068
                           , QN => n20977);
   REGISTERS_reg_8_24_inst : DFF_X1 port map( D => n6556, CK => CLK, Q => n8069
                           , QN => n20978);
   REGISTERS_reg_28_59_inst : DFF_X1 port map( D => n5311, CK => CLK, Q => 
                           n24027, QN => n20157);
   REGISTERS_reg_28_58_inst : DFF_X1 port map( D => n5310, CK => CLK, Q => 
                           n24026, QN => n20158);
   REGISTERS_reg_28_57_inst : DFF_X1 port map( D => n5309, CK => CLK, Q => 
                           n24025, QN => n20159);
   REGISTERS_reg_28_56_inst : DFF_X1 port map( D => n5308, CK => CLK, Q => 
                           n24024, QN => n20160);
   REGISTERS_reg_28_55_inst : DFF_X1 port map( D => n5307, CK => CLK, Q => 
                           n24023, QN => n20161);
   REGISTERS_reg_28_54_inst : DFF_X1 port map( D => n5306, CK => CLK, Q => 
                           n24022, QN => n20162);
   REGISTERS_reg_28_53_inst : DFF_X1 port map( D => n5305, CK => CLK, Q => 
                           n24021, QN => n20163);
   REGISTERS_reg_28_52_inst : DFF_X1 port map( D => n5304, CK => CLK, Q => 
                           n24020, QN => n20164);
   REGISTERS_reg_28_51_inst : DFF_X1 port map( D => n5303, CK => CLK, Q => 
                           n24019, QN => n20165);
   REGISTERS_reg_28_50_inst : DFF_X1 port map( D => n5302, CK => CLK, Q => 
                           n24018, QN => n20166);
   REGISTERS_reg_28_49_inst : DFF_X1 port map( D => n5301, CK => CLK, Q => 
                           n24017, QN => n20167);
   REGISTERS_reg_28_48_inst : DFF_X1 port map( D => n5300, CK => CLK, Q => 
                           n24016, QN => n20168);
   REGISTERS_reg_28_47_inst : DFF_X1 port map( D => n5299, CK => CLK, Q => 
                           n24015, QN => n20169);
   REGISTERS_reg_28_46_inst : DFF_X1 port map( D => n5298, CK => CLK, Q => 
                           n24014, QN => n20170);
   REGISTERS_reg_28_45_inst : DFF_X1 port map( D => n5297, CK => CLK, Q => 
                           n24013, QN => n20171);
   REGISTERS_reg_28_44_inst : DFF_X1 port map( D => n5296, CK => CLK, Q => 
                           n24012, QN => n20172);
   REGISTERS_reg_28_43_inst : DFF_X1 port map( D => n5295, CK => CLK, Q => 
                           n24011, QN => n20173);
   REGISTERS_reg_28_42_inst : DFF_X1 port map( D => n5294, CK => CLK, Q => 
                           n24010, QN => n20174);
   REGISTERS_reg_28_41_inst : DFF_X1 port map( D => n5293, CK => CLK, Q => 
                           n24009, QN => n20175);
   REGISTERS_reg_28_40_inst : DFF_X1 port map( D => n5292, CK => CLK, Q => 
                           n24008, QN => n20176);
   REGISTERS_reg_28_39_inst : DFF_X1 port map( D => n5291, CK => CLK, Q => 
                           n24007, QN => n20177);
   REGISTERS_reg_28_38_inst : DFF_X1 port map( D => n5290, CK => CLK, Q => 
                           n24006, QN => n20178);
   REGISTERS_reg_28_37_inst : DFF_X1 port map( D => n5289, CK => CLK, Q => 
                           n24005, QN => n20179);
   REGISTERS_reg_28_36_inst : DFF_X1 port map( D => n5288, CK => CLK, Q => 
                           n24004, QN => n20180);
   REGISTERS_reg_28_35_inst : DFF_X1 port map( D => n5287, CK => CLK, Q => 
                           n24003, QN => n20181);
   REGISTERS_reg_28_34_inst : DFF_X1 port map( D => n5286, CK => CLK, Q => 
                           n24002, QN => n20182);
   REGISTERS_reg_28_33_inst : DFF_X1 port map( D => n5285, CK => CLK, Q => 
                           n24001, QN => n20183);
   REGISTERS_reg_28_32_inst : DFF_X1 port map( D => n5284, CK => CLK, Q => 
                           n24000, QN => n20184);
   REGISTERS_reg_28_31_inst : DFF_X1 port map( D => n5283, CK => CLK, Q => 
                           n23999, QN => n20185);
   REGISTERS_reg_28_30_inst : DFF_X1 port map( D => n5282, CK => CLK, Q => 
                           n23998, QN => n20186);
   REGISTERS_reg_28_29_inst : DFF_X1 port map( D => n5281, CK => CLK, Q => 
                           n23997, QN => n19708);
   REGISTERS_reg_28_28_inst : DFF_X1 port map( D => n5280, CK => CLK, Q => 
                           n23996, QN => n19709);
   REGISTERS_reg_28_27_inst : DFF_X1 port map( D => n5279, CK => CLK, Q => 
                           n23995, QN => n19710);
   REGISTERS_reg_28_26_inst : DFF_X1 port map( D => n5278, CK => CLK, Q => 
                           n23994, QN => n19711);
   REGISTERS_reg_28_25_inst : DFF_X1 port map( D => n5277, CK => CLK, Q => 
                           n23993, QN => n19712);
   REGISTERS_reg_28_24_inst : DFF_X1 port map( D => n5276, CK => CLK, Q => 
                           n23992, QN => n19713);
   REGISTERS_reg_12_23_inst : DFF_X1 port map( D => n6299, CK => CLK, Q => 
                           n8326, QN => n21051);
   REGISTERS_reg_12_22_inst : DFF_X1 port map( D => n6298, CK => CLK, Q => 
                           n8327, QN => n21052);
   REGISTERS_reg_12_21_inst : DFF_X1 port map( D => n6297, CK => CLK, Q => 
                           n8328, QN => n21053);
   REGISTERS_reg_12_20_inst : DFF_X1 port map( D => n6296, CK => CLK, Q => 
                           n8329, QN => n21054);
   REGISTERS_reg_12_19_inst : DFF_X1 port map( D => n6295, CK => CLK, Q => 
                           n8330, QN => n21055);
   REGISTERS_reg_12_18_inst : DFF_X1 port map( D => n6294, CK => CLK, Q => 
                           n8331, QN => n21056);
   REGISTERS_reg_12_17_inst : DFF_X1 port map( D => n6293, CK => CLK, Q => 
                           n8332, QN => n21057);
   REGISTERS_reg_12_16_inst : DFF_X1 port map( D => n6292, CK => CLK, Q => 
                           n8333, QN => n21058);
   REGISTERS_reg_12_15_inst : DFF_X1 port map( D => n6291, CK => CLK, Q => 
                           n8334, QN => n21059);
   REGISTERS_reg_12_14_inst : DFF_X1 port map( D => n6290, CK => CLK, Q => 
                           n8335, QN => n21060);
   REGISTERS_reg_12_13_inst : DFF_X1 port map( D => n6289, CK => CLK, Q => 
                           n8336, QN => n21061);
   REGISTERS_reg_12_12_inst : DFF_X1 port map( D => n6288, CK => CLK, Q => 
                           n8337, QN => n21062);
   REGISTERS_reg_12_11_inst : DFF_X1 port map( D => n6287, CK => CLK, Q => 
                           n8338, QN => n21063);
   REGISTERS_reg_12_10_inst : DFF_X1 port map( D => n6286, CK => CLK, Q => 
                           n8339, QN => n21064);
   REGISTERS_reg_12_9_inst : DFF_X1 port map( D => n6285, CK => CLK, Q => n8340
                           , QN => n21065);
   REGISTERS_reg_12_8_inst : DFF_X1 port map( D => n6284, CK => CLK, Q => n8341
                           , QN => n21066);
   REGISTERS_reg_12_7_inst : DFF_X1 port map( D => n6283, CK => CLK, Q => n8342
                           , QN => n21067);
   REGISTERS_reg_12_6_inst : DFF_X1 port map( D => n6282, CK => CLK, Q => n8343
                           , QN => n21068);
   REGISTERS_reg_12_5_inst : DFF_X1 port map( D => n6281, CK => CLK, Q => n8344
                           , QN => n21069);
   REGISTERS_reg_12_4_inst : DFF_X1 port map( D => n6280, CK => CLK, Q => n8345
                           , QN => n21070);
   REGISTERS_reg_12_3_inst : DFF_X1 port map( D => n6279, CK => CLK, Q => n8346
                           , QN => n21071);
   REGISTERS_reg_12_2_inst : DFF_X1 port map( D => n6278, CK => CLK, Q => n8347
                           , QN => n21072);
   REGISTERS_reg_12_1_inst : DFF_X1 port map( D => n6277, CK => CLK, Q => n8348
                           , QN => n21073);
   REGISTERS_reg_12_0_inst : DFF_X1 port map( D => n6276, CK => CLK, Q => n8349
                           , QN => n21074);
   REGISTERS_reg_8_23_inst : DFF_X1 port map( D => n6555, CK => CLK, Q => n8070
                           , QN => n21075);
   REGISTERS_reg_8_22_inst : DFF_X1 port map( D => n6554, CK => CLK, Q => n8071
                           , QN => n21076);
   REGISTERS_reg_8_21_inst : DFF_X1 port map( D => n6553, CK => CLK, Q => n8072
                           , QN => n21077);
   REGISTERS_reg_8_20_inst : DFF_X1 port map( D => n6552, CK => CLK, Q => n8073
                           , QN => n21078);
   REGISTERS_reg_8_19_inst : DFF_X1 port map( D => n6551, CK => CLK, Q => n8074
                           , QN => n21079);
   REGISTERS_reg_8_18_inst : DFF_X1 port map( D => n6550, CK => CLK, Q => n8075
                           , QN => n21080);
   REGISTERS_reg_8_17_inst : DFF_X1 port map( D => n6549, CK => CLK, Q => n8076
                           , QN => n21081);
   REGISTERS_reg_8_16_inst : DFF_X1 port map( D => n6548, CK => CLK, Q => n8077
                           , QN => n21082);
   REGISTERS_reg_8_15_inst : DFF_X1 port map( D => n6547, CK => CLK, Q => n8078
                           , QN => n21083);
   REGISTERS_reg_8_14_inst : DFF_X1 port map( D => n6546, CK => CLK, Q => n8079
                           , QN => n21084);
   REGISTERS_reg_8_13_inst : DFF_X1 port map( D => n6545, CK => CLK, Q => n8080
                           , QN => n21085);
   REGISTERS_reg_8_12_inst : DFF_X1 port map( D => n6544, CK => CLK, Q => n8081
                           , QN => n21086);
   REGISTERS_reg_8_11_inst : DFF_X1 port map( D => n6543, CK => CLK, Q => n8082
                           , QN => n21087);
   REGISTERS_reg_8_10_inst : DFF_X1 port map( D => n6542, CK => CLK, Q => n8083
                           , QN => n21088);
   REGISTERS_reg_8_9_inst : DFF_X1 port map( D => n6541, CK => CLK, Q => n8084,
                           QN => n21089);
   REGISTERS_reg_8_8_inst : DFF_X1 port map( D => n6540, CK => CLK, Q => n8085,
                           QN => n21090);
   REGISTERS_reg_8_7_inst : DFF_X1 port map( D => n6539, CK => CLK, Q => n8086,
                           QN => n21091);
   REGISTERS_reg_8_6_inst : DFF_X1 port map( D => n6538, CK => CLK, Q => n8087,
                           QN => n21092);
   REGISTERS_reg_8_5_inst : DFF_X1 port map( D => n6537, CK => CLK, Q => n8088,
                           QN => n21093);
   REGISTERS_reg_8_4_inst : DFF_X1 port map( D => n6536, CK => CLK, Q => n8089,
                           QN => n21094);
   REGISTERS_reg_8_3_inst : DFF_X1 port map( D => n6535, CK => CLK, Q => n8090,
                           QN => n21095);
   REGISTERS_reg_8_2_inst : DFF_X1 port map( D => n6534, CK => CLK, Q => n8091,
                           QN => n21096);
   REGISTERS_reg_8_1_inst : DFF_X1 port map( D => n6533, CK => CLK, Q => n8092,
                           QN => n21097);
   REGISTERS_reg_8_0_inst : DFF_X1 port map( D => n6532, CK => CLK, Q => n8093,
                           QN => n21098);
   REGISTERS_reg_30_59_inst : DFF_X1 port map( D => n5183, CK => CLK, Q => 
                           n8674, QN => n20547);
   REGISTERS_reg_30_58_inst : DFF_X1 port map( D => n5182, CK => CLK, Q => 
                           n8675, QN => n20548);
   REGISTERS_reg_30_57_inst : DFF_X1 port map( D => n5181, CK => CLK, Q => 
                           n8676, QN => n20549);
   REGISTERS_reg_30_56_inst : DFF_X1 port map( D => n5180, CK => CLK, Q => 
                           n8677, QN => n20550);
   REGISTERS_reg_30_55_inst : DFF_X1 port map( D => n5179, CK => CLK, Q => 
                           n8678, QN => n20551);
   REGISTERS_reg_30_54_inst : DFF_X1 port map( D => n5178, CK => CLK, Q => 
                           n8679, QN => n20552);
   REGISTERS_reg_30_53_inst : DFF_X1 port map( D => n5177, CK => CLK, Q => 
                           n8680, QN => n20553);
   REGISTERS_reg_30_52_inst : DFF_X1 port map( D => n5176, CK => CLK, Q => 
                           n8681, QN => n20554);
   REGISTERS_reg_30_51_inst : DFF_X1 port map( D => n5175, CK => CLK, Q => 
                           n8682, QN => n20555);
   REGISTERS_reg_30_50_inst : DFF_X1 port map( D => n5174, CK => CLK, Q => 
                           n8683, QN => n20556);
   REGISTERS_reg_30_49_inst : DFF_X1 port map( D => n5173, CK => CLK, Q => 
                           n8684, QN => n20557);
   REGISTERS_reg_30_48_inst : DFF_X1 port map( D => n5172, CK => CLK, Q => 
                           n8685, QN => n20558);
   REGISTERS_reg_30_47_inst : DFF_X1 port map( D => n5171, CK => CLK, Q => 
                           n8686, QN => n20559);
   REGISTERS_reg_30_46_inst : DFF_X1 port map( D => n5170, CK => CLK, Q => 
                           n8687, QN => n20560);
   REGISTERS_reg_30_45_inst : DFF_X1 port map( D => n5169, CK => CLK, Q => 
                           n8688, QN => n20561);
   REGISTERS_reg_30_44_inst : DFF_X1 port map( D => n5168, CK => CLK, Q => 
                           n8689, QN => n20562);
   REGISTERS_reg_30_43_inst : DFF_X1 port map( D => n5167, CK => CLK, Q => 
                           n8690, QN => n20563);
   REGISTERS_reg_30_42_inst : DFF_X1 port map( D => n5166, CK => CLK, Q => 
                           n8691, QN => n20564);
   REGISTERS_reg_30_41_inst : DFF_X1 port map( D => n5165, CK => CLK, Q => 
                           n8692, QN => n20565);
   REGISTERS_reg_30_40_inst : DFF_X1 port map( D => n5164, CK => CLK, Q => 
                           n8693, QN => n20566);
   REGISTERS_reg_30_39_inst : DFF_X1 port map( D => n5163, CK => CLK, Q => 
                           n8694, QN => n20567);
   REGISTERS_reg_30_38_inst : DFF_X1 port map( D => n5162, CK => CLK, Q => 
                           n8695, QN => n20568);
   REGISTERS_reg_30_37_inst : DFF_X1 port map( D => n5161, CK => CLK, Q => 
                           n8696, QN => n20569);
   REGISTERS_reg_30_36_inst : DFF_X1 port map( D => n5160, CK => CLK, Q => 
                           n8697, QN => n20570);
   REGISTERS_reg_30_35_inst : DFF_X1 port map( D => n5159, CK => CLK, Q => 
                           n8698, QN => n20571);
   REGISTERS_reg_30_34_inst : DFF_X1 port map( D => n5158, CK => CLK, Q => 
                           n8699, QN => n20572);
   REGISTERS_reg_30_33_inst : DFF_X1 port map( D => n5157, CK => CLK, Q => 
                           n8700, QN => n20573);
   REGISTERS_reg_30_32_inst : DFF_X1 port map( D => n5156, CK => CLK, Q => 
                           n8701, QN => n20574);
   REGISTERS_reg_30_31_inst : DFF_X1 port map( D => n5155, CK => CLK, Q => 
                           n8702, QN => n20575);
   REGISTERS_reg_30_30_inst : DFF_X1 port map( D => n5154, CK => CLK, Q => 
                           n8703, QN => n20576);
   REGISTERS_reg_30_29_inst : DFF_X1 port map( D => n5153, CK => CLK, Q => 
                           n8704, QN => n20577);
   REGISTERS_reg_30_28_inst : DFF_X1 port map( D => n5152, CK => CLK, Q => 
                           n8705, QN => n20578);
   REGISTERS_reg_30_27_inst : DFF_X1 port map( D => n5151, CK => CLK, Q => 
                           n8706, QN => n20579);
   REGISTERS_reg_30_26_inst : DFF_X1 port map( D => n5150, CK => CLK, Q => 
                           n8707, QN => n20580);
   REGISTERS_reg_30_25_inst : DFF_X1 port map( D => n5149, CK => CLK, Q => 
                           n8708, QN => n20581);
   REGISTERS_reg_30_24_inst : DFF_X1 port map( D => n5148, CK => CLK, Q => 
                           n8709, QN => n20582);
   REGISTERS_reg_26_59_inst : DFF_X1 port map( D => n5439, CK => CLK, Q => 
                           n8354, QN => n20583);
   REGISTERS_reg_26_58_inst : DFF_X1 port map( D => n5438, CK => CLK, Q => 
                           n8355, QN => n20584);
   REGISTERS_reg_26_57_inst : DFF_X1 port map( D => n5437, CK => CLK, Q => 
                           n8356, QN => n20585);
   REGISTERS_reg_26_56_inst : DFF_X1 port map( D => n5436, CK => CLK, Q => 
                           n8357, QN => n20586);
   REGISTERS_reg_26_55_inst : DFF_X1 port map( D => n5435, CK => CLK, Q => 
                           n8358, QN => n20587);
   REGISTERS_reg_26_54_inst : DFF_X1 port map( D => n5434, CK => CLK, Q => 
                           n8359, QN => n20588);
   REGISTERS_reg_26_53_inst : DFF_X1 port map( D => n5433, CK => CLK, Q => 
                           n8360, QN => n20589);
   REGISTERS_reg_26_52_inst : DFF_X1 port map( D => n5432, CK => CLK, Q => 
                           n8361, QN => n20590);
   REGISTERS_reg_26_51_inst : DFF_X1 port map( D => n5431, CK => CLK, Q => 
                           n8362, QN => n20591);
   REGISTERS_reg_26_50_inst : DFF_X1 port map( D => n5430, CK => CLK, Q => 
                           n8363, QN => n20592);
   REGISTERS_reg_26_49_inst : DFF_X1 port map( D => n5429, CK => CLK, Q => 
                           n8364, QN => n20593);
   REGISTERS_reg_26_48_inst : DFF_X1 port map( D => n5428, CK => CLK, Q => 
                           n8365, QN => n20594);
   REGISTERS_reg_26_47_inst : DFF_X1 port map( D => n5427, CK => CLK, Q => 
                           n8366, QN => n20595);
   REGISTERS_reg_26_46_inst : DFF_X1 port map( D => n5426, CK => CLK, Q => 
                           n8367, QN => n20596);
   REGISTERS_reg_26_45_inst : DFF_X1 port map( D => n5425, CK => CLK, Q => 
                           n8368, QN => n20597);
   REGISTERS_reg_26_44_inst : DFF_X1 port map( D => n5424, CK => CLK, Q => 
                           n8369, QN => n20598);
   REGISTERS_reg_26_43_inst : DFF_X1 port map( D => n5423, CK => CLK, Q => 
                           n8370, QN => n20599);
   REGISTERS_reg_26_42_inst : DFF_X1 port map( D => n5422, CK => CLK, Q => 
                           n8371, QN => n20600);
   REGISTERS_reg_26_41_inst : DFF_X1 port map( D => n5421, CK => CLK, Q => 
                           n8372, QN => n20601);
   REGISTERS_reg_26_40_inst : DFF_X1 port map( D => n5420, CK => CLK, Q => 
                           n8373, QN => n20602);
   REGISTERS_reg_26_39_inst : DFF_X1 port map( D => n5419, CK => CLK, Q => 
                           n8374, QN => n20603);
   REGISTERS_reg_26_38_inst : DFF_X1 port map( D => n5418, CK => CLK, Q => 
                           n8375, QN => n20604);
   REGISTERS_reg_26_37_inst : DFF_X1 port map( D => n5417, CK => CLK, Q => 
                           n8376, QN => n20605);
   REGISTERS_reg_26_36_inst : DFF_X1 port map( D => n5416, CK => CLK, Q => 
                           n8377, QN => n20606);
   REGISTERS_reg_26_35_inst : DFF_X1 port map( D => n5415, CK => CLK, Q => 
                           n8378, QN => n20607);
   REGISTERS_reg_26_34_inst : DFF_X1 port map( D => n5414, CK => CLK, Q => 
                           n8379, QN => n20608);
   REGISTERS_reg_26_33_inst : DFF_X1 port map( D => n5413, CK => CLK, Q => 
                           n8380, QN => n20609);
   REGISTERS_reg_26_32_inst : DFF_X1 port map( D => n5412, CK => CLK, Q => 
                           n8381, QN => n20610);
   REGISTERS_reg_26_31_inst : DFF_X1 port map( D => n5411, CK => CLK, Q => 
                           n8382, QN => n20611);
   REGISTERS_reg_26_30_inst : DFF_X1 port map( D => n5410, CK => CLK, Q => 
                           n8383, QN => n20612);
   REGISTERS_reg_26_29_inst : DFF_X1 port map( D => n5409, CK => CLK, Q => 
                           n8384, QN => n20613);
   REGISTERS_reg_26_28_inst : DFF_X1 port map( D => n5408, CK => CLK, Q => 
                           n8385, QN => n20614);
   REGISTERS_reg_26_27_inst : DFF_X1 port map( D => n5407, CK => CLK, Q => 
                           n8386, QN => n20615);
   REGISTERS_reg_26_26_inst : DFF_X1 port map( D => n5406, CK => CLK, Q => 
                           n8387, QN => n20616);
   REGISTERS_reg_26_25_inst : DFF_X1 port map( D => n5405, CK => CLK, Q => 
                           n8388, QN => n20617);
   REGISTERS_reg_26_24_inst : DFF_X1 port map( D => n5404, CK => CLK, Q => 
                           n8389, QN => n20618);
   REGISTERS_reg_28_23_inst : DFF_X1 port map( D => n5275, CK => CLK, Q => 
                           n23991, QN => n19714);
   REGISTERS_reg_28_22_inst : DFF_X1 port map( D => n5274, CK => CLK, Q => 
                           n23990, QN => n19715);
   REGISTERS_reg_28_21_inst : DFF_X1 port map( D => n5273, CK => CLK, Q => 
                           n23989, QN => n19716);
   REGISTERS_reg_28_20_inst : DFF_X1 port map( D => n5272, CK => CLK, Q => 
                           n23988, QN => n19717);
   REGISTERS_reg_28_19_inst : DFF_X1 port map( D => n5271, CK => CLK, Q => 
                           n23987, QN => n19718);
   REGISTERS_reg_28_18_inst : DFF_X1 port map( D => n5270, CK => CLK, Q => 
                           n23986, QN => n19719);
   REGISTERS_reg_28_17_inst : DFF_X1 port map( D => n5269, CK => CLK, Q => 
                           n23985, QN => n19720);
   REGISTERS_reg_28_16_inst : DFF_X1 port map( D => n5268, CK => CLK, Q => 
                           n23984, QN => n19721);
   REGISTERS_reg_28_15_inst : DFF_X1 port map( D => n5267, CK => CLK, Q => 
                           n23983, QN => n19722);
   REGISTERS_reg_28_14_inst : DFF_X1 port map( D => n5266, CK => CLK, Q => 
                           n23982, QN => n19723);
   REGISTERS_reg_28_13_inst : DFF_X1 port map( D => n5265, CK => CLK, Q => 
                           n23981, QN => n19724);
   REGISTERS_reg_28_12_inst : DFF_X1 port map( D => n5264, CK => CLK, Q => 
                           n23980, QN => n19725);
   REGISTERS_reg_28_11_inst : DFF_X1 port map( D => n5263, CK => CLK, Q => 
                           n23979, QN => n19726);
   REGISTERS_reg_28_10_inst : DFF_X1 port map( D => n5262, CK => CLK, Q => 
                           n23978, QN => n19727);
   REGISTERS_reg_28_9_inst : DFF_X1 port map( D => n5261, CK => CLK, Q => 
                           n23977, QN => n19728);
   REGISTERS_reg_28_8_inst : DFF_X1 port map( D => n5260, CK => CLK, Q => 
                           n23976, QN => n19729);
   REGISTERS_reg_28_7_inst : DFF_X1 port map( D => n5259, CK => CLK, Q => 
                           n23975, QN => n19730);
   REGISTERS_reg_28_6_inst : DFF_X1 port map( D => n5258, CK => CLK, Q => 
                           n23974, QN => n19731);
   REGISTERS_reg_28_5_inst : DFF_X1 port map( D => n5257, CK => CLK, Q => 
                           n23973, QN => n19732);
   REGISTERS_reg_28_4_inst : DFF_X1 port map( D => n5256, CK => CLK, Q => 
                           n23972, QN => n19733);
   REGISTERS_reg_28_3_inst : DFF_X1 port map( D => n5255, CK => CLK, Q => 
                           n23971, QN => n19734);
   REGISTERS_reg_28_2_inst : DFF_X1 port map( D => n5254, CK => CLK, Q => 
                           n23970, QN => n19735);
   REGISTERS_reg_28_1_inst : DFF_X1 port map( D => n5253, CK => CLK, Q => 
                           n23969, QN => n19736);
   REGISTERS_reg_28_0_inst : DFF_X1 port map( D => n5252, CK => CLK, Q => 
                           n23968, QN => n19737);
   REGISTERS_reg_30_23_inst : DFF_X1 port map( D => n5147, CK => CLK, Q => 
                           n8710, QN => n20727);
   REGISTERS_reg_30_22_inst : DFF_X1 port map( D => n5146, CK => CLK, Q => 
                           n8711, QN => n20728);
   REGISTERS_reg_30_21_inst : DFF_X1 port map( D => n5145, CK => CLK, Q => 
                           n8712, QN => n20729);
   REGISTERS_reg_30_20_inst : DFF_X1 port map( D => n5144, CK => CLK, Q => 
                           n8713, QN => n20730);
   REGISTERS_reg_30_19_inst : DFF_X1 port map( D => n5143, CK => CLK, Q => 
                           n8714, QN => n20731);
   REGISTERS_reg_30_18_inst : DFF_X1 port map( D => n5142, CK => CLK, Q => 
                           n8715, QN => n20732);
   REGISTERS_reg_30_17_inst : DFF_X1 port map( D => n5141, CK => CLK, Q => 
                           n8716, QN => n20733);
   REGISTERS_reg_30_16_inst : DFF_X1 port map( D => n5140, CK => CLK, Q => 
                           n8717, QN => n20734);
   REGISTERS_reg_30_15_inst : DFF_X1 port map( D => n5139, CK => CLK, Q => 
                           n8718, QN => n20735);
   REGISTERS_reg_30_14_inst : DFF_X1 port map( D => n5138, CK => CLK, Q => 
                           n8719, QN => n20736);
   REGISTERS_reg_30_13_inst : DFF_X1 port map( D => n5137, CK => CLK, Q => 
                           n8720, QN => n20737);
   REGISTERS_reg_30_12_inst : DFF_X1 port map( D => n5136, CK => CLK, Q => 
                           n8721, QN => n20738);
   REGISTERS_reg_30_11_inst : DFF_X1 port map( D => n5135, CK => CLK, Q => 
                           n8722, QN => n20739);
   REGISTERS_reg_30_10_inst : DFF_X1 port map( D => n5134, CK => CLK, Q => 
                           n8723, QN => n20740);
   REGISTERS_reg_30_9_inst : DFF_X1 port map( D => n5133, CK => CLK, Q => n8724
                           , QN => n20741);
   REGISTERS_reg_30_8_inst : DFF_X1 port map( D => n5132, CK => CLK, Q => n8725
                           , QN => n20742);
   REGISTERS_reg_30_7_inst : DFF_X1 port map( D => n5131, CK => CLK, Q => n8726
                           , QN => n20743);
   REGISTERS_reg_30_6_inst : DFF_X1 port map( D => n5130, CK => CLK, Q => n8727
                           , QN => n20744);
   REGISTERS_reg_30_5_inst : DFF_X1 port map( D => n5129, CK => CLK, Q => n8728
                           , QN => n20745);
   REGISTERS_reg_30_4_inst : DFF_X1 port map( D => n5128, CK => CLK, Q => n8729
                           , QN => n20746);
   REGISTERS_reg_30_3_inst : DFF_X1 port map( D => n5127, CK => CLK, Q => n8730
                           , QN => n20747);
   REGISTERS_reg_30_2_inst : DFF_X1 port map( D => n5126, CK => CLK, Q => n8731
                           , QN => n20748);
   REGISTERS_reg_30_1_inst : DFF_X1 port map( D => n5125, CK => CLK, Q => n8732
                           , QN => n20749);
   REGISTERS_reg_30_0_inst : DFF_X1 port map( D => n5124, CK => CLK, Q => n8733
                           , QN => n20750);
   REGISTERS_reg_26_23_inst : DFF_X1 port map( D => n5403, CK => CLK, Q => 
                           n8390, QN => n20751);
   REGISTERS_reg_26_22_inst : DFF_X1 port map( D => n5402, CK => CLK, Q => 
                           n8391, QN => n20752);
   REGISTERS_reg_26_21_inst : DFF_X1 port map( D => n5401, CK => CLK, Q => 
                           n8392, QN => n20753);
   REGISTERS_reg_26_20_inst : DFF_X1 port map( D => n5400, CK => CLK, Q => 
                           n8393, QN => n20754);
   REGISTERS_reg_26_19_inst : DFF_X1 port map( D => n5399, CK => CLK, Q => 
                           n8394, QN => n20755);
   REGISTERS_reg_26_18_inst : DFF_X1 port map( D => n5398, CK => CLK, Q => 
                           n8395, QN => n20756);
   REGISTERS_reg_26_17_inst : DFF_X1 port map( D => n5397, CK => CLK, Q => 
                           n8396, QN => n20757);
   REGISTERS_reg_26_16_inst : DFF_X1 port map( D => n5396, CK => CLK, Q => 
                           n8397, QN => n20758);
   REGISTERS_reg_26_15_inst : DFF_X1 port map( D => n5395, CK => CLK, Q => 
                           n8398, QN => n20759);
   REGISTERS_reg_26_14_inst : DFF_X1 port map( D => n5394, CK => CLK, Q => 
                           n8399, QN => n20760);
   REGISTERS_reg_26_13_inst : DFF_X1 port map( D => n5393, CK => CLK, Q => 
                           n8400, QN => n20761);
   REGISTERS_reg_26_12_inst : DFF_X1 port map( D => n5392, CK => CLK, Q => 
                           n8401, QN => n20762);
   REGISTERS_reg_26_11_inst : DFF_X1 port map( D => n5391, CK => CLK, Q => 
                           n8402, QN => n20763);
   REGISTERS_reg_26_10_inst : DFF_X1 port map( D => n5390, CK => CLK, Q => 
                           n8403, QN => n20764);
   REGISTERS_reg_26_9_inst : DFF_X1 port map( D => n5389, CK => CLK, Q => n8404
                           , QN => n20765);
   REGISTERS_reg_26_8_inst : DFF_X1 port map( D => n5388, CK => CLK, Q => n8405
                           , QN => n20766);
   REGISTERS_reg_26_7_inst : DFF_X1 port map( D => n5387, CK => CLK, Q => n8406
                           , QN => n20767);
   REGISTERS_reg_26_6_inst : DFF_X1 port map( D => n5386, CK => CLK, Q => n8407
                           , QN => n20768);
   REGISTERS_reg_26_5_inst : DFF_X1 port map( D => n5385, CK => CLK, Q => n8408
                           , QN => n20769);
   REGISTERS_reg_26_4_inst : DFF_X1 port map( D => n5384, CK => CLK, Q => n8409
                           , QN => n20770);
   REGISTERS_reg_26_3_inst : DFF_X1 port map( D => n5383, CK => CLK, Q => n8410
                           , QN => n20771);
   REGISTERS_reg_26_2_inst : DFF_X1 port map( D => n5382, CK => CLK, Q => n8411
                           , QN => n20772);
   REGISTERS_reg_26_1_inst : DFF_X1 port map( D => n5381, CK => CLK, Q => n8412
                           , QN => n20773);
   REGISTERS_reg_26_0_inst : DFF_X1 port map( D => n5380, CK => CLK, Q => n8413
                           , QN => n20774);
   REGISTERS_reg_1_62_inst : DFF_X1 port map( D => n7042, CK => CLK, Q => n7647
                           , QN => n21148);
   REGISTERS_reg_1_63_inst : DFF_X1 port map( D => n7043, CK => CLK, Q => n7646
                           , QN => n21149);
   REGISTERS_reg_1_61_inst : DFF_X1 port map( D => n7041, CK => CLK, Q => n7648
                           , QN => n21150);
   REGISTERS_reg_1_60_inst : DFF_X1 port map( D => n7040, CK => CLK, Q => n7649
                           , QN => n21151);
   REGISTERS_reg_1_59_inst : DFF_X1 port map( D => n7039, CK => CLK, Q => n7650
                           , QN => n21152);
   REGISTERS_reg_1_58_inst : DFF_X1 port map( D => n7038, CK => CLK, Q => n7651
                           , QN => n21153);
   REGISTERS_reg_1_57_inst : DFF_X1 port map( D => n7037, CK => CLK, Q => n7652
                           , QN => n21154);
   REGISTERS_reg_1_56_inst : DFF_X1 port map( D => n7036, CK => CLK, Q => n7653
                           , QN => n21155);
   REGISTERS_reg_1_55_inst : DFF_X1 port map( D => n7035, CK => CLK, Q => n7654
                           , QN => n21156);
   REGISTERS_reg_1_54_inst : DFF_X1 port map( D => n7034, CK => CLK, Q => n7655
                           , QN => n21157);
   REGISTERS_reg_1_53_inst : DFF_X1 port map( D => n7033, CK => CLK, Q => n7656
                           , QN => n21158);
   REGISTERS_reg_1_52_inst : DFF_X1 port map( D => n7032, CK => CLK, Q => n7657
                           , QN => n21159);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n7008, CK => CLK, Q => n7681
                           , QN => n21160);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n7007, CK => CLK, Q => n7682
                           , QN => n21161);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n7006, CK => CLK, Q => n7683
                           , QN => n21162);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n7005, CK => CLK, Q => n7684
                           , QN => n21163);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n7004, CK => CLK, Q => n7685
                           , QN => n21164);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n7003, CK => CLK, Q => n7686
                           , QN => n21165);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n7002, CK => CLK, Q => n7687
                           , QN => n21166);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n7001, CK => CLK, Q => n7688
                           , QN => n21167);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n7000, CK => CLK, Q => n7689
                           , QN => n21168);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n6999, CK => CLK, Q => n7690
                           , QN => n21169);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n6998, CK => CLK, Q => n7691
                           , QN => n21170);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n6997, CK => CLK, Q => n7692
                           , QN => n21171);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n6996, CK => CLK, Q => n7693
                           , QN => n21172);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n6995, CK => CLK, Q => n7694
                           , QN => n21173);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n6994, CK => CLK, Q => n7695
                           , QN => n21174);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n6993, CK => CLK, Q => n7696
                           , QN => n21175);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n6992, CK => CLK, Q => n7697
                           , QN => n21176);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n6991, CK => CLK, Q => n7698
                           , QN => n21177);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n6990, CK => CLK, Q => n7699
                           , QN => n21178);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n6989, CK => CLK, Q => n7700,
                           QN => n21179);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n6988, CK => CLK, Q => n7701,
                           QN => n21180);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n6987, CK => CLK, Q => n7702,
                           QN => n21181);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n6986, CK => CLK, Q => n7703,
                           QN => n21182);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n6985, CK => CLK, Q => n7704,
                           QN => n21183);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n6984, CK => CLK, Q => n7705,
                           QN => n21184);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n6983, CK => CLK, Q => n7706,
                           QN => n21185);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n6982, CK => CLK, Q => n7707,
                           QN => n21186);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n6980, CK => CLK, Q => n7709,
                           QN => n21187);
   REGISTERS_reg_27_63_inst : DFF_X1 port map( D => n5379, CK => CLK, Q => 
                           n7966, QN => n20527);
   REGISTERS_reg_27_62_inst : DFF_X1 port map( D => n5378, CK => CLK, Q => 
                           n7967, QN => n20528);
   REGISTERS_reg_27_61_inst : DFF_X1 port map( D => n5377, CK => CLK, Q => 
                           n7968, QN => n20529);
   REGISTERS_reg_27_60_inst : DFF_X1 port map( D => n5376, CK => CLK, Q => 
                           n7969, QN => n20530);
   REGISTERS_reg_27_59_inst : DFF_X1 port map( D => n5375, CK => CLK, Q => 
                           n7970, QN => n20847);
   REGISTERS_reg_27_58_inst : DFF_X1 port map( D => n5374, CK => CLK, Q => 
                           n7971, QN => n20848);
   REGISTERS_reg_27_57_inst : DFF_X1 port map( D => n5373, CK => CLK, Q => 
                           n7972, QN => n20849);
   REGISTERS_reg_27_56_inst : DFF_X1 port map( D => n5372, CK => CLK, Q => 
                           n7973, QN => n20850);
   REGISTERS_reg_27_55_inst : DFF_X1 port map( D => n5371, CK => CLK, Q => 
                           n7974, QN => n20851);
   REGISTERS_reg_27_54_inst : DFF_X1 port map( D => n5370, CK => CLK, Q => 
                           n7975, QN => n20852);
   REGISTERS_reg_27_53_inst : DFF_X1 port map( D => n5369, CK => CLK, Q => 
                           n7976, QN => n20853);
   REGISTERS_reg_27_52_inst : DFF_X1 port map( D => n5368, CK => CLK, Q => 
                           n7977, QN => n20854);
   REGISTERS_reg_27_51_inst : DFF_X1 port map( D => n5367, CK => CLK, Q => 
                           n7978, QN => n20855);
   REGISTERS_reg_27_50_inst : DFF_X1 port map( D => n5366, CK => CLK, Q => 
                           n7979, QN => n20856);
   REGISTERS_reg_27_49_inst : DFF_X1 port map( D => n5365, CK => CLK, Q => 
                           n7980, QN => n20857);
   REGISTERS_reg_27_48_inst : DFF_X1 port map( D => n5364, CK => CLK, Q => 
                           n7981, QN => n20858);
   REGISTERS_reg_27_47_inst : DFF_X1 port map( D => n5363, CK => CLK, Q => 
                           n7982, QN => n20859);
   REGISTERS_reg_27_46_inst : DFF_X1 port map( D => n5362, CK => CLK, Q => 
                           n7983, QN => n20860);
   REGISTERS_reg_27_45_inst : DFF_X1 port map( D => n5361, CK => CLK, Q => 
                           n7984, QN => n20861);
   REGISTERS_reg_27_44_inst : DFF_X1 port map( D => n5360, CK => CLK, Q => 
                           n7985, QN => n20862);
   REGISTERS_reg_27_43_inst : DFF_X1 port map( D => n5359, CK => CLK, Q => 
                           n7986, QN => n20863);
   REGISTERS_reg_27_42_inst : DFF_X1 port map( D => n5358, CK => CLK, Q => 
                           n7987, QN => n20864);
   REGISTERS_reg_27_41_inst : DFF_X1 port map( D => n5357, CK => CLK, Q => 
                           n7988, QN => n20865);
   REGISTERS_reg_27_40_inst : DFF_X1 port map( D => n5356, CK => CLK, Q => 
                           n7989, QN => n20866);
   REGISTERS_reg_27_39_inst : DFF_X1 port map( D => n5355, CK => CLK, Q => 
                           n7990, QN => n20867);
   REGISTERS_reg_27_38_inst : DFF_X1 port map( D => n5354, CK => CLK, Q => 
                           n7991, QN => n20868);
   REGISTERS_reg_27_37_inst : DFF_X1 port map( D => n5353, CK => CLK, Q => 
                           n7992, QN => n20869);
   REGISTERS_reg_27_36_inst : DFF_X1 port map( D => n5352, CK => CLK, Q => 
                           n7993, QN => n20870);
   REGISTERS_reg_27_35_inst : DFF_X1 port map( D => n5351, CK => CLK, Q => 
                           n7994, QN => n20871);
   REGISTERS_reg_27_34_inst : DFF_X1 port map( D => n5350, CK => CLK, Q => 
                           n7995, QN => n20872);
   REGISTERS_reg_27_33_inst : DFF_X1 port map( D => n5349, CK => CLK, Q => 
                           n7996, QN => n20873);
   REGISTERS_reg_27_32_inst : DFF_X1 port map( D => n5348, CK => CLK, Q => 
                           n7997, QN => n20874);
   REGISTERS_reg_27_31_inst : DFF_X1 port map( D => n5347, CK => CLK, Q => 
                           n7998, QN => n20875);
   REGISTERS_reg_27_30_inst : DFF_X1 port map( D => n5346, CK => CLK, Q => 
                           n7999, QN => n20876);
   REGISTERS_reg_27_29_inst : DFF_X1 port map( D => n5345, CK => CLK, Q => 
                           n8000, QN => n20877);
   REGISTERS_reg_27_28_inst : DFF_X1 port map( D => n5344, CK => CLK, Q => 
                           n8001, QN => n20878);
   REGISTERS_reg_27_27_inst : DFF_X1 port map( D => n5343, CK => CLK, Q => 
                           n8002, QN => n20879);
   REGISTERS_reg_27_26_inst : DFF_X1 port map( D => n5342, CK => CLK, Q => 
                           n8003, QN => n20880);
   REGISTERS_reg_27_25_inst : DFF_X1 port map( D => n5341, CK => CLK, Q => 
                           n8004, QN => n20881);
   REGISTERS_reg_27_24_inst : DFF_X1 port map( D => n5340, CK => CLK, Q => 
                           n8005, QN => n20882);
   REGISTERS_reg_27_23_inst : DFF_X1 port map( D => n5339, CK => CLK, Q => 
                           n8006, QN => n20883);
   REGISTERS_reg_27_22_inst : DFF_X1 port map( D => n5338, CK => CLK, Q => 
                           n8007, QN => n20884);
   REGISTERS_reg_27_21_inst : DFF_X1 port map( D => n5337, CK => CLK, Q => 
                           n8008, QN => n20885);
   REGISTERS_reg_27_20_inst : DFF_X1 port map( D => n5336, CK => CLK, Q => 
                           n8009, QN => n20886);
   REGISTERS_reg_27_19_inst : DFF_X1 port map( D => n5335, CK => CLK, Q => 
                           n8010, QN => n20887);
   REGISTERS_reg_27_18_inst : DFF_X1 port map( D => n5334, CK => CLK, Q => 
                           n8011, QN => n20888);
   REGISTERS_reg_27_17_inst : DFF_X1 port map( D => n5333, CK => CLK, Q => 
                           n8012, QN => n20889);
   REGISTERS_reg_27_16_inst : DFF_X1 port map( D => n5332, CK => CLK, Q => 
                           n8013, QN => n20890);
   REGISTERS_reg_27_15_inst : DFF_X1 port map( D => n5331, CK => CLK, Q => 
                           n8014, QN => n20891);
   REGISTERS_reg_27_14_inst : DFF_X1 port map( D => n5330, CK => CLK, Q => 
                           n8015, QN => n20892);
   REGISTERS_reg_27_13_inst : DFF_X1 port map( D => n5329, CK => CLK, Q => 
                           n8016, QN => n20893);
   REGISTERS_reg_27_12_inst : DFF_X1 port map( D => n5328, CK => CLK, Q => 
                           n8017, QN => n20894);
   REGISTERS_reg_27_11_inst : DFF_X1 port map( D => n5327, CK => CLK, Q => 
                           n8018, QN => n20895);
   REGISTERS_reg_27_10_inst : DFF_X1 port map( D => n5326, CK => CLK, Q => 
                           n8019, QN => n20896);
   REGISTERS_reg_27_9_inst : DFF_X1 port map( D => n5325, CK => CLK, Q => n8020
                           , QN => n20897);
   REGISTERS_reg_27_8_inst : DFF_X1 port map( D => n5324, CK => CLK, Q => n8021
                           , QN => n20898);
   REGISTERS_reg_27_7_inst : DFF_X1 port map( D => n5323, CK => CLK, Q => n8022
                           , QN => n20899);
   REGISTERS_reg_27_6_inst : DFF_X1 port map( D => n5322, CK => CLK, Q => n8023
                           , QN => n20900);
   REGISTERS_reg_27_5_inst : DFF_X1 port map( D => n5321, CK => CLK, Q => n8024
                           , QN => n20901);
   REGISTERS_reg_27_4_inst : DFF_X1 port map( D => n5320, CK => CLK, Q => n8025
                           , QN => n20902);
   REGISTERS_reg_27_3_inst : DFF_X1 port map( D => n5319, CK => CLK, Q => n8026
                           , QN => n20903);
   REGISTERS_reg_27_2_inst : DFF_X1 port map( D => n5318, CK => CLK, Q => n8027
                           , QN => n20904);
   REGISTERS_reg_27_1_inst : DFF_X1 port map( D => n5317, CK => CLK, Q => n8028
                           , QN => n20905);
   REGISTERS_reg_27_0_inst : DFF_X1 port map( D => n5316, CK => CLK, Q => n8029
                           , QN => n20906);
   OUT2_reg_63_inst : DFF_X1 port map( D => n4995, CK => CLK, Q => OUT2_63_port
                           , QN => n_1616);
   OUT2_reg_62_inst : DFF_X1 port map( D => n4994, CK => CLK, Q => OUT2_62_port
                           , QN => n_1617);
   OUT2_reg_61_inst : DFF_X1 port map( D => n4993, CK => CLK, Q => OUT2_61_port
                           , QN => n_1618);
   OUT2_reg_60_inst : DFF_X1 port map( D => n4992, CK => CLK, Q => OUT2_60_port
                           , QN => n_1619);
   OUT2_reg_59_inst : DFF_X1 port map( D => n4991, CK => CLK, Q => OUT2_59_port
                           , QN => n_1620);
   OUT2_reg_58_inst : DFF_X1 port map( D => n4990, CK => CLK, Q => OUT2_58_port
                           , QN => n_1621);
   OUT2_reg_57_inst : DFF_X1 port map( D => n4989, CK => CLK, Q => OUT2_57_port
                           , QN => n_1622);
   OUT2_reg_56_inst : DFF_X1 port map( D => n4988, CK => CLK, Q => OUT2_56_port
                           , QN => n_1623);
   OUT2_reg_55_inst : DFF_X1 port map( D => n4987, CK => CLK, Q => OUT2_55_port
                           , QN => n_1624);
   OUT2_reg_54_inst : DFF_X1 port map( D => n4986, CK => CLK, Q => OUT2_54_port
                           , QN => n_1625);
   OUT2_reg_53_inst : DFF_X1 port map( D => n4985, CK => CLK, Q => OUT2_53_port
                           , QN => n_1626);
   OUT2_reg_52_inst : DFF_X1 port map( D => n4984, CK => CLK, Q => OUT2_52_port
                           , QN => n_1627);
   OUT2_reg_51_inst : DFF_X1 port map( D => n4983, CK => CLK, Q => OUT2_51_port
                           , QN => n_1628);
   OUT2_reg_50_inst : DFF_X1 port map( D => n4982, CK => CLK, Q => OUT2_50_port
                           , QN => n_1629);
   OUT2_reg_49_inst : DFF_X1 port map( D => n4981, CK => CLK, Q => OUT2_49_port
                           , QN => n_1630);
   OUT2_reg_48_inst : DFF_X1 port map( D => n4980, CK => CLK, Q => OUT2_48_port
                           , QN => n_1631);
   OUT2_reg_47_inst : DFF_X1 port map( D => n4979, CK => CLK, Q => OUT2_47_port
                           , QN => n_1632);
   OUT2_reg_46_inst : DFF_X1 port map( D => n4978, CK => CLK, Q => OUT2_46_port
                           , QN => n_1633);
   OUT2_reg_45_inst : DFF_X1 port map( D => n4977, CK => CLK, Q => OUT2_45_port
                           , QN => n_1634);
   OUT2_reg_44_inst : DFF_X1 port map( D => n4976, CK => CLK, Q => OUT2_44_port
                           , QN => n_1635);
   OUT2_reg_43_inst : DFF_X1 port map( D => n4975, CK => CLK, Q => OUT2_43_port
                           , QN => n_1636);
   OUT2_reg_42_inst : DFF_X1 port map( D => n4974, CK => CLK, Q => OUT2_42_port
                           , QN => n_1637);
   OUT2_reg_41_inst : DFF_X1 port map( D => n4973, CK => CLK, Q => OUT2_41_port
                           , QN => n_1638);
   OUT2_reg_40_inst : DFF_X1 port map( D => n4972, CK => CLK, Q => OUT2_40_port
                           , QN => n_1639);
   U18625 : NOR2_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), ZN => n22542)
                           ;
   U18626 : INV_X1 port map( A => n24832, ZN => n24818);
   U18627 : INV_X1 port map( A => n24832, ZN => n24817);
   U18628 : INV_X1 port map( A => n25549, ZN => n25535);
   U18629 : INV_X1 port map( A => n25549, ZN => n25536);
   U18630 : INV_X1 port map( A => n24833, ZN => n24819);
   U18631 : INV_X1 port map( A => n25343, ZN => n25329);
   U18632 : INV_X1 port map( A => n25343, ZN => n25328);
   U18633 : INV_X1 port map( A => n25274, ZN => n25260);
   U18634 : INV_X1 port map( A => n25274, ZN => n25261);
   U18635 : INV_X1 port map( A => n25189, ZN => n25175);
   U18636 : INV_X1 port map( A => n25189, ZN => n25176);
   U18637 : INV_X1 port map( A => n25104, ZN => n25090);
   U18638 : INV_X1 port map( A => n25104, ZN => n25091);
   U18639 : INV_X1 port map( A => n25053, ZN => n25039);
   U18640 : INV_X1 port map( A => n25053, ZN => n25040);
   U18641 : INV_X1 port map( A => n25036, ZN => n25022);
   U18642 : INV_X1 port map( A => n25036, ZN => n25023);
   U18643 : INV_X1 port map( A => n24866, ZN => n24852);
   U18644 : INV_X1 port map( A => n24866, ZN => n24853);
   U18645 : INV_X1 port map( A => n24934, ZN => n24920);
   U18646 : INV_X1 port map( A => n24934, ZN => n24921);
   U18647 : INV_X1 port map( A => n24968, ZN => n24954);
   U18648 : INV_X1 port map( A => n24968, ZN => n24955);
   U18649 : INV_X1 port map( A => n24985, ZN => n24971);
   U18650 : INV_X1 port map( A => n24985, ZN => n24972);
   U18651 : INV_X1 port map( A => n25121, ZN => n25107);
   U18652 : INV_X1 port map( A => n25121, ZN => n25108);
   U18653 : INV_X1 port map( A => n25138, ZN => n25124);
   U18654 : INV_X1 port map( A => n25138, ZN => n25125);
   U18655 : INV_X1 port map( A => n25172, ZN => n25158);
   U18656 : INV_X1 port map( A => n25172, ZN => n25159);
   U18657 : INV_X1 port map( A => n25002, ZN => n24988);
   U18658 : INV_X1 port map( A => n25002, ZN => n24989);
   U18659 : INV_X1 port map( A => n25240, ZN => n25226);
   U18660 : INV_X1 port map( A => n25240, ZN => n25227);
   U18661 : INV_X1 port map( A => n25223, ZN => n25209);
   U18662 : INV_X1 port map( A => n25223, ZN => n25210);
   U18663 : INV_X1 port map( A => n25155, ZN => n25141);
   U18664 : INV_X1 port map( A => n25155, ZN => n25142);
   U18665 : INV_X1 port map( A => n24900, ZN => n24886);
   U18666 : INV_X1 port map( A => n24900, ZN => n24887);
   U18667 : INV_X1 port map( A => n25257, ZN => n25243);
   U18668 : INV_X1 port map( A => n25257, ZN => n25244);
   U18669 : INV_X1 port map( A => n25087, ZN => n25073);
   U18670 : INV_X1 port map( A => n25087, ZN => n25074);
   U18671 : INV_X1 port map( A => n25019, ZN => n25005);
   U18672 : INV_X1 port map( A => n25019, ZN => n25006);
   U18673 : INV_X1 port map( A => n24917, ZN => n24903);
   U18674 : INV_X1 port map( A => n24917, ZN => n24904);
   U18675 : INV_X1 port map( A => n24849, ZN => n24835);
   U18676 : INV_X1 port map( A => n24849, ZN => n24836);
   U18677 : INV_X1 port map( A => n25070, ZN => n25056);
   U18678 : INV_X1 port map( A => n25070, ZN => n25057);
   U18679 : INV_X1 port map( A => n25325, ZN => n25311);
   U18680 : INV_X1 port map( A => n25325, ZN => n25312);
   U18681 : INV_X1 port map( A => n25206, ZN => n25192);
   U18682 : INV_X1 port map( A => n25206, ZN => n25193);
   U18683 : INV_X1 port map( A => n25308, ZN => n25294);
   U18684 : INV_X1 port map( A => n25308, ZN => n25295);
   U18685 : INV_X1 port map( A => n24883, ZN => n24869);
   U18686 : INV_X1 port map( A => n24883, ZN => n24870);
   U18687 : INV_X1 port map( A => n24951, ZN => n24937);
   U18688 : INV_X1 port map( A => n24951, ZN => n24938);
   U18689 : INV_X1 port map( A => n25291, ZN => n25277);
   U18690 : INV_X1 port map( A => n25291, ZN => n25278);
   U18691 : BUF_X1 port map( A => n24814, Z => n24832);
   U18692 : BUF_X1 port map( A => n25550, Z => n25549);
   U18693 : BUF_X1 port map( A => n24813, Z => n24831);
   U18694 : BUF_X1 port map( A => n24813, Z => n24830);
   U18695 : BUF_X1 port map( A => n24813, Z => n24829);
   U18696 : BUF_X1 port map( A => n24812, Z => n24828);
   U18697 : BUF_X1 port map( A => n24812, Z => n24827);
   U18698 : BUF_X1 port map( A => n24812, Z => n24826);
   U18699 : BUF_X1 port map( A => n24811, Z => n24825);
   U18700 : BUF_X1 port map( A => n24811, Z => n24824);
   U18701 : BUF_X1 port map( A => n24811, Z => n24823);
   U18702 : BUF_X1 port map( A => n24810, Z => n24822);
   U18703 : BUF_X1 port map( A => n24810, Z => n24821);
   U18704 : BUF_X1 port map( A => n24810, Z => n24820);
   U18705 : BUF_X1 port map( A => n25550, Z => n25537);
   U18706 : BUF_X1 port map( A => n25550, Z => n25538);
   U18707 : BUF_X1 port map( A => n25550, Z => n25539);
   U18708 : BUF_X1 port map( A => n25550, Z => n25540);
   U18709 : BUF_X1 port map( A => n25550, Z => n25541);
   U18710 : BUF_X1 port map( A => n25550, Z => n25542);
   U18711 : BUF_X1 port map( A => n25550, Z => n25543);
   U18712 : BUF_X1 port map( A => n25537, Z => n25544);
   U18713 : BUF_X1 port map( A => n25538, Z => n25545);
   U18714 : BUF_X1 port map( A => n25539, Z => n25546);
   U18715 : BUF_X1 port map( A => n25540, Z => n25547);
   U18716 : BUF_X1 port map( A => n25541, Z => n25548);
   U18717 : BUF_X1 port map( A => n24814, Z => n24833);
   U18718 : BUF_X1 port map( A => n22602, Z => n24442);
   U18719 : BUF_X1 port map( A => n22602, Z => n24438);
   U18720 : BUF_X1 port map( A => n22602, Z => n24439);
   U18721 : BUF_X1 port map( A => n22602, Z => n24440);
   U18722 : BUF_X1 port map( A => n22602, Z => n24441);
   U18723 : BUF_X1 port map( A => n22571, Z => n24586);
   U18724 : BUF_X1 port map( A => n22571, Z => n24582);
   U18725 : BUF_X1 port map( A => n22571, Z => n24583);
   U18726 : BUF_X1 port map( A => n22571, Z => n24584);
   U18727 : BUF_X1 port map( A => n22571, Z => n24585);
   U18728 : BUF_X1 port map( A => n22577, Z => n24556);
   U18729 : BUF_X1 port map( A => n22577, Z => n24552);
   U18730 : BUF_X1 port map( A => n22577, Z => n24553);
   U18731 : BUF_X1 port map( A => n22577, Z => n24554);
   U18732 : BUF_X1 port map( A => n22577, Z => n24555);
   U18733 : BUF_X1 port map( A => n22594, Z => n24490);
   U18734 : BUF_X1 port map( A => n22594, Z => n24486);
   U18735 : BUF_X1 port map( A => n22594, Z => n24487);
   U18736 : BUF_X1 port map( A => n22594, Z => n24488);
   U18737 : BUF_X1 port map( A => n22594, Z => n24489);
   U18738 : BUF_X1 port map( A => n22574, Z => n24568);
   U18739 : BUF_X1 port map( A => n22574, Z => n24564);
   U18740 : BUF_X1 port map( A => n22574, Z => n24565);
   U18741 : BUF_X1 port map( A => n22574, Z => n24566);
   U18742 : BUF_X1 port map( A => n22574, Z => n24567);
   U18743 : BUF_X1 port map( A => n25003, Z => n25002);
   U18744 : BUF_X1 port map( A => n25241, Z => n25240);
   U18745 : BUF_X1 port map( A => n25224, Z => n25223);
   U18746 : BUF_X1 port map( A => n25156, Z => n25155);
   U18747 : BUF_X1 port map( A => n24901, Z => n24900);
   U18748 : BUF_X1 port map( A => n25258, Z => n25257);
   U18749 : BUF_X1 port map( A => n25088, Z => n25087);
   U18750 : BUF_X1 port map( A => n25020, Z => n25019);
   U18751 : BUF_X1 port map( A => n24918, Z => n24917);
   U18752 : BUF_X1 port map( A => n24850, Z => n24849);
   U18753 : BUF_X1 port map( A => n25071, Z => n25070);
   U18754 : BUF_X1 port map( A => n25326, Z => n25325);
   U18755 : BUF_X1 port map( A => n25207, Z => n25206);
   U18756 : BUF_X1 port map( A => n25309, Z => n25308);
   U18757 : BUF_X1 port map( A => n25344, Z => n25342);
   U18758 : BUF_X1 port map( A => n25275, Z => n25274);
   U18759 : BUF_X1 port map( A => n25190, Z => n25189);
   U18760 : BUF_X1 port map( A => n25105, Z => n25104);
   U18761 : BUF_X1 port map( A => n25054, Z => n25053);
   U18762 : BUF_X1 port map( A => n25037, Z => n25036);
   U18763 : BUF_X1 port map( A => n24867, Z => n24866);
   U18764 : BUF_X1 port map( A => n24884, Z => n24883);
   U18765 : BUF_X1 port map( A => n24935, Z => n24934);
   U18766 : BUF_X1 port map( A => n24952, Z => n24951);
   U18767 : BUF_X1 port map( A => n24969, Z => n24968);
   U18768 : BUF_X1 port map( A => n24986, Z => n24985);
   U18769 : BUF_X1 port map( A => n25122, Z => n25121);
   U18770 : BUF_X1 port map( A => n25139, Z => n25138);
   U18771 : BUF_X1 port map( A => n25173, Z => n25172);
   U18772 : BUF_X1 port map( A => n25292, Z => n25291);
   U18773 : BUF_X1 port map( A => n25344, Z => n25331);
   U18774 : BUF_X1 port map( A => n25344, Z => n25332);
   U18775 : BUF_X1 port map( A => n25344, Z => n25333);
   U18776 : BUF_X1 port map( A => n25344, Z => n25334);
   U18777 : BUF_X1 port map( A => n25331, Z => n25341);
   U18778 : BUF_X1 port map( A => n25344, Z => n25330);
   U18779 : BUF_X1 port map( A => n25003, Z => n24990);
   U18780 : BUF_X1 port map( A => n25003, Z => n24991);
   U18781 : BUF_X1 port map( A => n25003, Z => n24992);
   U18782 : BUF_X1 port map( A => n25003, Z => n24993);
   U18783 : BUF_X1 port map( A => n25241, Z => n25228);
   U18784 : BUF_X1 port map( A => n25241, Z => n25229);
   U18785 : BUF_X1 port map( A => n25241, Z => n25230);
   U18786 : BUF_X1 port map( A => n25241, Z => n25231);
   U18787 : BUF_X1 port map( A => n25224, Z => n25211);
   U18788 : BUF_X1 port map( A => n25224, Z => n25212);
   U18789 : BUF_X1 port map( A => n25224, Z => n25213);
   U18790 : BUF_X1 port map( A => n25224, Z => n25214);
   U18791 : BUF_X1 port map( A => n25156, Z => n25143);
   U18792 : BUF_X1 port map( A => n25156, Z => n25144);
   U18793 : BUF_X1 port map( A => n25156, Z => n25145);
   U18794 : BUF_X1 port map( A => n25156, Z => n25146);
   U18795 : BUF_X1 port map( A => n25003, Z => n24994);
   U18796 : BUF_X1 port map( A => n25003, Z => n24995);
   U18797 : BUF_X1 port map( A => n25003, Z => n24996);
   U18798 : BUF_X1 port map( A => n24990, Z => n24997);
   U18799 : BUF_X1 port map( A => n24991, Z => n24998);
   U18800 : BUF_X1 port map( A => n24992, Z => n24999);
   U18801 : BUF_X1 port map( A => n24993, Z => n25000);
   U18802 : BUF_X1 port map( A => n24994, Z => n25001);
   U18803 : BUF_X1 port map( A => n25241, Z => n25232);
   U18804 : BUF_X1 port map( A => n25241, Z => n25233);
   U18805 : BUF_X1 port map( A => n25241, Z => n25234);
   U18806 : BUF_X1 port map( A => n25228, Z => n25235);
   U18807 : BUF_X1 port map( A => n25229, Z => n25236);
   U18808 : BUF_X1 port map( A => n25230, Z => n25237);
   U18809 : BUF_X1 port map( A => n25231, Z => n25238);
   U18810 : BUF_X1 port map( A => n25232, Z => n25239);
   U18811 : BUF_X1 port map( A => n25224, Z => n25215);
   U18812 : BUF_X1 port map( A => n25224, Z => n25216);
   U18813 : BUF_X1 port map( A => n25224, Z => n25217);
   U18814 : BUF_X1 port map( A => n25211, Z => n25218);
   U18815 : BUF_X1 port map( A => n25212, Z => n25219);
   U18816 : BUF_X1 port map( A => n25213, Z => n25220);
   U18817 : BUF_X1 port map( A => n25214, Z => n25221);
   U18818 : BUF_X1 port map( A => n25215, Z => n25222);
   U18819 : BUF_X1 port map( A => n25156, Z => n25147);
   U18820 : BUF_X1 port map( A => n25156, Z => n25148);
   U18821 : BUF_X1 port map( A => n25156, Z => n25149);
   U18822 : BUF_X1 port map( A => n25143, Z => n25150);
   U18823 : BUF_X1 port map( A => n25144, Z => n25151);
   U18824 : BUF_X1 port map( A => n25145, Z => n25152);
   U18825 : BUF_X1 port map( A => n25146, Z => n25153);
   U18826 : BUF_X1 port map( A => n25147, Z => n25154);
   U18827 : BUF_X1 port map( A => n24901, Z => n24888);
   U18828 : BUF_X1 port map( A => n24901, Z => n24889);
   U18829 : BUF_X1 port map( A => n24901, Z => n24890);
   U18830 : BUF_X1 port map( A => n24901, Z => n24891);
   U18831 : BUF_X1 port map( A => n24901, Z => n24892);
   U18832 : BUF_X1 port map( A => n24901, Z => n24893);
   U18833 : BUF_X1 port map( A => n24901, Z => n24894);
   U18834 : BUF_X1 port map( A => n24888, Z => n24895);
   U18835 : BUF_X1 port map( A => n24889, Z => n24896);
   U18836 : BUF_X1 port map( A => n24890, Z => n24897);
   U18837 : BUF_X1 port map( A => n24891, Z => n24898);
   U18838 : BUF_X1 port map( A => n24892, Z => n24899);
   U18839 : BUF_X1 port map( A => n25258, Z => n25245);
   U18840 : BUF_X1 port map( A => n25258, Z => n25246);
   U18841 : BUF_X1 port map( A => n25258, Z => n25247);
   U18842 : BUF_X1 port map( A => n25258, Z => n25248);
   U18843 : BUF_X1 port map( A => n25088, Z => n25075);
   U18844 : BUF_X1 port map( A => n25088, Z => n25076);
   U18845 : BUF_X1 port map( A => n25088, Z => n25077);
   U18846 : BUF_X1 port map( A => n25088, Z => n25078);
   U18847 : BUF_X1 port map( A => n25020, Z => n25007);
   U18848 : BUF_X1 port map( A => n25020, Z => n25008);
   U18849 : BUF_X1 port map( A => n25020, Z => n25009);
   U18850 : BUF_X1 port map( A => n25020, Z => n25010);
   U18851 : BUF_X1 port map( A => n24918, Z => n24905);
   U18852 : BUF_X1 port map( A => n24918, Z => n24906);
   U18853 : BUF_X1 port map( A => n24918, Z => n24907);
   U18854 : BUF_X1 port map( A => n24918, Z => n24908);
   U18855 : BUF_X1 port map( A => n24850, Z => n24837);
   U18856 : BUF_X1 port map( A => n24850, Z => n24838);
   U18857 : BUF_X1 port map( A => n24850, Z => n24839);
   U18858 : BUF_X1 port map( A => n24850, Z => n24840);
   U18859 : BUF_X1 port map( A => n25258, Z => n25249);
   U18860 : BUF_X1 port map( A => n25258, Z => n25250);
   U18861 : BUF_X1 port map( A => n25258, Z => n25251);
   U18862 : BUF_X1 port map( A => n25245, Z => n25252);
   U18863 : BUF_X1 port map( A => n25246, Z => n25253);
   U18864 : BUF_X1 port map( A => n25247, Z => n25254);
   U18865 : BUF_X1 port map( A => n25248, Z => n25255);
   U18866 : BUF_X1 port map( A => n25249, Z => n25256);
   U18867 : BUF_X1 port map( A => n25088, Z => n25079);
   U18868 : BUF_X1 port map( A => n25088, Z => n25080);
   U18869 : BUF_X1 port map( A => n25088, Z => n25081);
   U18870 : BUF_X1 port map( A => n25075, Z => n25082);
   U18871 : BUF_X1 port map( A => n25076, Z => n25083);
   U18872 : BUF_X1 port map( A => n25077, Z => n25084);
   U18873 : BUF_X1 port map( A => n25078, Z => n25085);
   U18874 : BUF_X1 port map( A => n25079, Z => n25086);
   U18875 : BUF_X1 port map( A => n25020, Z => n25011);
   U18876 : BUF_X1 port map( A => n25020, Z => n25012);
   U18877 : BUF_X1 port map( A => n25020, Z => n25013);
   U18878 : BUF_X1 port map( A => n25007, Z => n25014);
   U18879 : BUF_X1 port map( A => n25008, Z => n25015);
   U18880 : BUF_X1 port map( A => n25009, Z => n25016);
   U18881 : BUF_X1 port map( A => n25010, Z => n25017);
   U18882 : BUF_X1 port map( A => n25011, Z => n25018);
   U18883 : BUF_X1 port map( A => n24918, Z => n24909);
   U18884 : BUF_X1 port map( A => n24918, Z => n24910);
   U18885 : BUF_X1 port map( A => n24918, Z => n24911);
   U18886 : BUF_X1 port map( A => n24905, Z => n24912);
   U18887 : BUF_X1 port map( A => n24906, Z => n24913);
   U18888 : BUF_X1 port map( A => n24907, Z => n24914);
   U18889 : BUF_X1 port map( A => n24908, Z => n24915);
   U18890 : BUF_X1 port map( A => n24909, Z => n24916);
   U18891 : BUF_X1 port map( A => n24850, Z => n24841);
   U18892 : BUF_X1 port map( A => n24850, Z => n24842);
   U18893 : BUF_X1 port map( A => n24850, Z => n24843);
   U18894 : BUF_X1 port map( A => n24837, Z => n24844);
   U18895 : BUF_X1 port map( A => n24838, Z => n24845);
   U18896 : BUF_X1 port map( A => n24839, Z => n24846);
   U18897 : BUF_X1 port map( A => n24840, Z => n24847);
   U18898 : BUF_X1 port map( A => n24841, Z => n24848);
   U18899 : BUF_X1 port map( A => n25071, Z => n25058);
   U18900 : BUF_X1 port map( A => n25071, Z => n25059);
   U18901 : BUF_X1 port map( A => n25071, Z => n25060);
   U18902 : BUF_X1 port map( A => n25071, Z => n25061);
   U18903 : BUF_X1 port map( A => n25071, Z => n25062);
   U18904 : BUF_X1 port map( A => n25071, Z => n25063);
   U18905 : BUF_X1 port map( A => n25071, Z => n25064);
   U18906 : BUF_X1 port map( A => n25058, Z => n25065);
   U18907 : BUF_X1 port map( A => n25059, Z => n25066);
   U18908 : BUF_X1 port map( A => n25060, Z => n25067);
   U18909 : BUF_X1 port map( A => n25061, Z => n25068);
   U18910 : BUF_X1 port map( A => n25062, Z => n25069);
   U18911 : BUF_X1 port map( A => n25326, Z => n25313);
   U18912 : BUF_X1 port map( A => n25326, Z => n25314);
   U18913 : BUF_X1 port map( A => n25326, Z => n25315);
   U18914 : BUF_X1 port map( A => n25326, Z => n25316);
   U18915 : BUF_X1 port map( A => n25207, Z => n25194);
   U18916 : BUF_X1 port map( A => n25207, Z => n25195);
   U18917 : BUF_X1 port map( A => n25207, Z => n25196);
   U18918 : BUF_X1 port map( A => n25207, Z => n25197);
   U18919 : BUF_X1 port map( A => n25309, Z => n25296);
   U18920 : BUF_X1 port map( A => n25309, Z => n25297);
   U18921 : BUF_X1 port map( A => n25309, Z => n25298);
   U18922 : BUF_X1 port map( A => n25309, Z => n25299);
   U18923 : BUF_X1 port map( A => n25326, Z => n25317);
   U18924 : BUF_X1 port map( A => n25326, Z => n25318);
   U18925 : BUF_X1 port map( A => n25326, Z => n25319);
   U18926 : BUF_X1 port map( A => n25313, Z => n25320);
   U18927 : BUF_X1 port map( A => n25314, Z => n25321);
   U18928 : BUF_X1 port map( A => n25315, Z => n25322);
   U18929 : BUF_X1 port map( A => n25316, Z => n25323);
   U18930 : BUF_X1 port map( A => n25317, Z => n25324);
   U18931 : BUF_X1 port map( A => n25207, Z => n25198);
   U18932 : BUF_X1 port map( A => n25207, Z => n25199);
   U18933 : BUF_X1 port map( A => n25207, Z => n25200);
   U18934 : BUF_X1 port map( A => n25194, Z => n25201);
   U18935 : BUF_X1 port map( A => n25195, Z => n25202);
   U18936 : BUF_X1 port map( A => n25196, Z => n25203);
   U18937 : BUF_X1 port map( A => n25197, Z => n25204);
   U18938 : BUF_X1 port map( A => n25198, Z => n25205);
   U18939 : BUF_X1 port map( A => n25309, Z => n25300);
   U18940 : BUF_X1 port map( A => n25309, Z => n25301);
   U18941 : BUF_X1 port map( A => n25309, Z => n25302);
   U18942 : BUF_X1 port map( A => n25296, Z => n25303);
   U18943 : BUF_X1 port map( A => n25297, Z => n25304);
   U18944 : BUF_X1 port map( A => n25298, Z => n25305);
   U18945 : BUF_X1 port map( A => n25299, Z => n25306);
   U18946 : BUF_X1 port map( A => n25300, Z => n25307);
   U18947 : BUF_X1 port map( A => n24884, Z => n24877);
   U18948 : BUF_X1 port map( A => n24877, Z => n24878);
   U18949 : BUF_X1 port map( A => n24871, Z => n24879);
   U18950 : BUF_X1 port map( A => n24872, Z => n24880);
   U18951 : BUF_X1 port map( A => n24873, Z => n24881);
   U18952 : BUF_X1 port map( A => n24874, Z => n24882);
   U18953 : BUF_X1 port map( A => n25344, Z => n25335);
   U18954 : BUF_X1 port map( A => n25344, Z => n25336);
   U18955 : BUF_X1 port map( A => n25332, Z => n25337);
   U18956 : BUF_X1 port map( A => n25333, Z => n25338);
   U18957 : BUF_X1 port map( A => n25334, Z => n25339);
   U18958 : BUF_X1 port map( A => n25330, Z => n25340);
   U18959 : BUF_X1 port map( A => n25275, Z => n25262);
   U18960 : BUF_X1 port map( A => n25275, Z => n25263);
   U18961 : BUF_X1 port map( A => n25275, Z => n25264);
   U18962 : BUF_X1 port map( A => n25275, Z => n25265);
   U18963 : BUF_X1 port map( A => n25190, Z => n25177);
   U18964 : BUF_X1 port map( A => n25190, Z => n25178);
   U18965 : BUF_X1 port map( A => n25190, Z => n25179);
   U18966 : BUF_X1 port map( A => n25190, Z => n25180);
   U18967 : BUF_X1 port map( A => n25105, Z => n25092);
   U18968 : BUF_X1 port map( A => n25105, Z => n25093);
   U18969 : BUF_X1 port map( A => n25105, Z => n25094);
   U18970 : BUF_X1 port map( A => n25105, Z => n25095);
   U18971 : BUF_X1 port map( A => n25054, Z => n25041);
   U18972 : BUF_X1 port map( A => n25054, Z => n25042);
   U18973 : BUF_X1 port map( A => n25054, Z => n25043);
   U18974 : BUF_X1 port map( A => n25054, Z => n25044);
   U18975 : BUF_X1 port map( A => n25037, Z => n25024);
   U18976 : BUF_X1 port map( A => n25037, Z => n25025);
   U18977 : BUF_X1 port map( A => n25037, Z => n25026);
   U18978 : BUF_X1 port map( A => n25037, Z => n25027);
   U18979 : BUF_X1 port map( A => n25275, Z => n25266);
   U18980 : BUF_X1 port map( A => n25275, Z => n25267);
   U18981 : BUF_X1 port map( A => n25275, Z => n25268);
   U18982 : BUF_X1 port map( A => n25262, Z => n25269);
   U18983 : BUF_X1 port map( A => n25263, Z => n25270);
   U18984 : BUF_X1 port map( A => n25264, Z => n25271);
   U18985 : BUF_X1 port map( A => n25265, Z => n25272);
   U18986 : BUF_X1 port map( A => n25266, Z => n25273);
   U18987 : BUF_X1 port map( A => n25190, Z => n25181);
   U18988 : BUF_X1 port map( A => n25190, Z => n25182);
   U18989 : BUF_X1 port map( A => n25190, Z => n25183);
   U18990 : BUF_X1 port map( A => n25177, Z => n25184);
   U18991 : BUF_X1 port map( A => n25178, Z => n25185);
   U18992 : BUF_X1 port map( A => n25179, Z => n25186);
   U18993 : BUF_X1 port map( A => n25180, Z => n25187);
   U18994 : BUF_X1 port map( A => n25181, Z => n25188);
   U18995 : BUF_X1 port map( A => n25105, Z => n25096);
   U18996 : BUF_X1 port map( A => n25105, Z => n25097);
   U18997 : BUF_X1 port map( A => n25105, Z => n25098);
   U18998 : BUF_X1 port map( A => n25092, Z => n25099);
   U18999 : BUF_X1 port map( A => n25093, Z => n25100);
   U19000 : BUF_X1 port map( A => n25094, Z => n25101);
   U19001 : BUF_X1 port map( A => n25095, Z => n25102);
   U19002 : BUF_X1 port map( A => n25096, Z => n25103);
   U19003 : BUF_X1 port map( A => n25054, Z => n25045);
   U19004 : BUF_X1 port map( A => n25054, Z => n25046);
   U19005 : BUF_X1 port map( A => n25054, Z => n25047);
   U19006 : BUF_X1 port map( A => n25041, Z => n25048);
   U19007 : BUF_X1 port map( A => n25042, Z => n25049);
   U19008 : BUF_X1 port map( A => n25043, Z => n25050);
   U19009 : BUF_X1 port map( A => n25044, Z => n25051);
   U19010 : BUF_X1 port map( A => n25045, Z => n25052);
   U19011 : BUF_X1 port map( A => n25037, Z => n25028);
   U19012 : BUF_X1 port map( A => n25037, Z => n25029);
   U19013 : BUF_X1 port map( A => n25037, Z => n25030);
   U19014 : BUF_X1 port map( A => n25024, Z => n25031);
   U19015 : BUF_X1 port map( A => n25025, Z => n25032);
   U19016 : BUF_X1 port map( A => n25026, Z => n25033);
   U19017 : BUF_X1 port map( A => n25027, Z => n25034);
   U19018 : BUF_X1 port map( A => n25028, Z => n25035);
   U19019 : BUF_X1 port map( A => n24867, Z => n24854);
   U19020 : BUF_X1 port map( A => n24867, Z => n24855);
   U19021 : BUF_X1 port map( A => n24867, Z => n24856);
   U19022 : BUF_X1 port map( A => n24867, Z => n24857);
   U19023 : BUF_X1 port map( A => n24867, Z => n24858);
   U19024 : BUF_X1 port map( A => n24867, Z => n24859);
   U19025 : BUF_X1 port map( A => n24867, Z => n24860);
   U19026 : BUF_X1 port map( A => n24854, Z => n24861);
   U19027 : BUF_X1 port map( A => n24855, Z => n24862);
   U19028 : BUF_X1 port map( A => n24856, Z => n24863);
   U19029 : BUF_X1 port map( A => n24857, Z => n24864);
   U19030 : BUF_X1 port map( A => n24858, Z => n24865);
   U19031 : BUF_X1 port map( A => n24884, Z => n24871);
   U19032 : BUF_X1 port map( A => n24884, Z => n24872);
   U19033 : BUF_X1 port map( A => n24884, Z => n24873);
   U19034 : BUF_X1 port map( A => n24884, Z => n24874);
   U19035 : BUF_X1 port map( A => n24884, Z => n24875);
   U19036 : BUF_X1 port map( A => n24884, Z => n24876);
   U19037 : BUF_X1 port map( A => n24935, Z => n24922);
   U19038 : BUF_X1 port map( A => n24935, Z => n24923);
   U19039 : BUF_X1 port map( A => n24935, Z => n24924);
   U19040 : BUF_X1 port map( A => n24935, Z => n24925);
   U19041 : BUF_X1 port map( A => n24935, Z => n24926);
   U19042 : BUF_X1 port map( A => n24935, Z => n24927);
   U19043 : BUF_X1 port map( A => n24935, Z => n24928);
   U19044 : BUF_X1 port map( A => n24922, Z => n24929);
   U19045 : BUF_X1 port map( A => n24923, Z => n24930);
   U19046 : BUF_X1 port map( A => n24924, Z => n24931);
   U19047 : BUF_X1 port map( A => n24925, Z => n24932);
   U19048 : BUF_X1 port map( A => n24926, Z => n24933);
   U19049 : BUF_X1 port map( A => n24952, Z => n24939);
   U19050 : BUF_X1 port map( A => n24952, Z => n24940);
   U19051 : BUF_X1 port map( A => n24952, Z => n24941);
   U19052 : BUF_X1 port map( A => n24952, Z => n24942);
   U19053 : BUF_X1 port map( A => n24952, Z => n24943);
   U19054 : BUF_X1 port map( A => n24952, Z => n24944);
   U19055 : BUF_X1 port map( A => n24952, Z => n24945);
   U19056 : BUF_X1 port map( A => n24939, Z => n24946);
   U19057 : BUF_X1 port map( A => n24940, Z => n24947);
   U19058 : BUF_X1 port map( A => n24941, Z => n24948);
   U19059 : BUF_X1 port map( A => n24942, Z => n24949);
   U19060 : BUF_X1 port map( A => n24943, Z => n24950);
   U19061 : BUF_X1 port map( A => n24969, Z => n24956);
   U19062 : BUF_X1 port map( A => n24969, Z => n24957);
   U19063 : BUF_X1 port map( A => n24969, Z => n24958);
   U19064 : BUF_X1 port map( A => n24969, Z => n24959);
   U19065 : BUF_X1 port map( A => n24969, Z => n24960);
   U19066 : BUF_X1 port map( A => n24969, Z => n24961);
   U19067 : BUF_X1 port map( A => n24969, Z => n24962);
   U19068 : BUF_X1 port map( A => n24956, Z => n24963);
   U19069 : BUF_X1 port map( A => n24957, Z => n24964);
   U19070 : BUF_X1 port map( A => n24958, Z => n24965);
   U19071 : BUF_X1 port map( A => n24959, Z => n24966);
   U19072 : BUF_X1 port map( A => n24960, Z => n24967);
   U19073 : BUF_X1 port map( A => n24986, Z => n24973);
   U19074 : BUF_X1 port map( A => n24986, Z => n24974);
   U19075 : BUF_X1 port map( A => n24986, Z => n24975);
   U19076 : BUF_X1 port map( A => n24986, Z => n24976);
   U19077 : BUF_X1 port map( A => n24986, Z => n24977);
   U19078 : BUF_X1 port map( A => n24986, Z => n24978);
   U19079 : BUF_X1 port map( A => n24986, Z => n24979);
   U19080 : BUF_X1 port map( A => n24973, Z => n24980);
   U19081 : BUF_X1 port map( A => n24974, Z => n24981);
   U19082 : BUF_X1 port map( A => n24975, Z => n24982);
   U19083 : BUF_X1 port map( A => n24976, Z => n24983);
   U19084 : BUF_X1 port map( A => n24977, Z => n24984);
   U19085 : BUF_X1 port map( A => n25122, Z => n25109);
   U19086 : BUF_X1 port map( A => n25122, Z => n25110);
   U19087 : BUF_X1 port map( A => n25122, Z => n25111);
   U19088 : BUF_X1 port map( A => n25122, Z => n25112);
   U19089 : BUF_X1 port map( A => n25122, Z => n25113);
   U19090 : BUF_X1 port map( A => n25122, Z => n25114);
   U19091 : BUF_X1 port map( A => n25122, Z => n25115);
   U19092 : BUF_X1 port map( A => n25109, Z => n25116);
   U19093 : BUF_X1 port map( A => n25110, Z => n25117);
   U19094 : BUF_X1 port map( A => n25111, Z => n25118);
   U19095 : BUF_X1 port map( A => n25112, Z => n25119);
   U19096 : BUF_X1 port map( A => n25113, Z => n25120);
   U19097 : BUF_X1 port map( A => n25139, Z => n25126);
   U19098 : BUF_X1 port map( A => n25139, Z => n25127);
   U19099 : BUF_X1 port map( A => n25139, Z => n25128);
   U19100 : BUF_X1 port map( A => n25139, Z => n25129);
   U19101 : BUF_X1 port map( A => n25139, Z => n25130);
   U19102 : BUF_X1 port map( A => n25139, Z => n25131);
   U19103 : BUF_X1 port map( A => n25139, Z => n25132);
   U19104 : BUF_X1 port map( A => n25126, Z => n25133);
   U19105 : BUF_X1 port map( A => n25127, Z => n25134);
   U19106 : BUF_X1 port map( A => n25128, Z => n25135);
   U19107 : BUF_X1 port map( A => n25129, Z => n25136);
   U19108 : BUF_X1 port map( A => n25130, Z => n25137);
   U19109 : BUF_X1 port map( A => n25173, Z => n25160);
   U19110 : BUF_X1 port map( A => n25173, Z => n25161);
   U19111 : BUF_X1 port map( A => n25173, Z => n25162);
   U19112 : BUF_X1 port map( A => n25173, Z => n25163);
   U19113 : BUF_X1 port map( A => n25173, Z => n25164);
   U19114 : BUF_X1 port map( A => n25173, Z => n25165);
   U19115 : BUF_X1 port map( A => n25173, Z => n25166);
   U19116 : BUF_X1 port map( A => n25160, Z => n25167);
   U19117 : BUF_X1 port map( A => n25161, Z => n25168);
   U19118 : BUF_X1 port map( A => n25162, Z => n25169);
   U19119 : BUF_X1 port map( A => n25163, Z => n25170);
   U19120 : BUF_X1 port map( A => n25164, Z => n25171);
   U19121 : BUF_X1 port map( A => n25292, Z => n25279);
   U19122 : BUF_X1 port map( A => n25292, Z => n25280);
   U19123 : BUF_X1 port map( A => n25292, Z => n25281);
   U19124 : BUF_X1 port map( A => n25292, Z => n25282);
   U19125 : BUF_X1 port map( A => n25292, Z => n25283);
   U19126 : BUF_X1 port map( A => n25292, Z => n25284);
   U19127 : BUF_X1 port map( A => n25292, Z => n25285);
   U19128 : BUF_X1 port map( A => n25279, Z => n25286);
   U19129 : BUF_X1 port map( A => n25280, Z => n25287);
   U19130 : BUF_X1 port map( A => n25281, Z => n25288);
   U19131 : BUF_X1 port map( A => n25282, Z => n25289);
   U19132 : BUF_X1 port map( A => n25283, Z => n25290);
   U19133 : BUF_X1 port map( A => n25335, Z => n25343);
   U19134 : BUF_X1 port map( A => n24815, Z => n24813);
   U19135 : BUF_X1 port map( A => n24815, Z => n24812);
   U19136 : BUF_X1 port map( A => n24816, Z => n24811);
   U19137 : BUF_X1 port map( A => n24816, Z => n24810);
   U19138 : BUF_X1 port map( A => n24815, Z => n24814);
   U19139 : INV_X1 port map( A => n25534, ZN => n25550);
   U19140 : BUF_X1 port map( A => n22598, Z => n24466);
   U19141 : BUF_X1 port map( A => n22598, Z => n24462);
   U19142 : BUF_X1 port map( A => n22598, Z => n24463);
   U19143 : BUF_X1 port map( A => n22598, Z => n24464);
   U19144 : BUF_X1 port map( A => n22598, Z => n24465);
   U19145 : BUF_X1 port map( A => n21307, Z => n24786);
   U19146 : BUF_X1 port map( A => n21312, Z => n24762);
   U19147 : BUF_X1 port map( A => n21317, Z => n24738);
   U19148 : BUF_X1 port map( A => n21322, Z => n24714);
   U19149 : BUF_X1 port map( A => n21331, Z => n24690);
   U19150 : BUF_X1 port map( A => n21336, Z => n24666);
   U19151 : BUF_X1 port map( A => n21341, Z => n24642);
   U19152 : BUF_X1 port map( A => n21346, Z => n24618);
   U19153 : BUF_X1 port map( A => n21307, Z => n24787);
   U19154 : BUF_X1 port map( A => n21312, Z => n24763);
   U19155 : BUF_X1 port map( A => n21317, Z => n24739);
   U19156 : BUF_X1 port map( A => n21322, Z => n24715);
   U19157 : BUF_X1 port map( A => n21331, Z => n24691);
   U19158 : BUF_X1 port map( A => n21336, Z => n24667);
   U19159 : BUF_X1 port map( A => n21341, Z => n24643);
   U19160 : BUF_X1 port map( A => n21346, Z => n24619);
   U19161 : BUF_X1 port map( A => n21307, Z => n24788);
   U19162 : BUF_X1 port map( A => n21312, Z => n24764);
   U19163 : BUF_X1 port map( A => n21317, Z => n24740);
   U19164 : BUF_X1 port map( A => n21322, Z => n24716);
   U19165 : BUF_X1 port map( A => n21331, Z => n24692);
   U19166 : BUF_X1 port map( A => n21336, Z => n24668);
   U19167 : BUF_X1 port map( A => n21341, Z => n24644);
   U19168 : BUF_X1 port map( A => n21346, Z => n24620);
   U19169 : BUF_X1 port map( A => n21307, Z => n24789);
   U19170 : BUF_X1 port map( A => n21312, Z => n24765);
   U19171 : BUF_X1 port map( A => n21317, Z => n24741);
   U19172 : BUF_X1 port map( A => n21322, Z => n24717);
   U19173 : BUF_X1 port map( A => n21331, Z => n24693);
   U19174 : BUF_X1 port map( A => n21336, Z => n24669);
   U19175 : BUF_X1 port map( A => n21341, Z => n24645);
   U19176 : BUF_X1 port map( A => n21346, Z => n24621);
   U19177 : BUF_X1 port map( A => n21307, Z => n24790);
   U19178 : BUF_X1 port map( A => n21312, Z => n24766);
   U19179 : BUF_X1 port map( A => n21317, Z => n24742);
   U19180 : BUF_X1 port map( A => n21322, Z => n24718);
   U19181 : BUF_X1 port map( A => n21331, Z => n24694);
   U19182 : BUF_X1 port map( A => n21336, Z => n24670);
   U19183 : BUF_X1 port map( A => n21341, Z => n24646);
   U19184 : BUF_X1 port map( A => n21346, Z => n24622);
   U19185 : BUF_X1 port map( A => n22607, Z => n24418);
   U19186 : BUF_X1 port map( A => n22607, Z => n24414);
   U19187 : BUF_X1 port map( A => n22607, Z => n24415);
   U19188 : BUF_X1 port map( A => n22607, Z => n24416);
   U19189 : BUF_X1 port map( A => n22607, Z => n24417);
   U19190 : BUF_X1 port map( A => n21302, Z => n24792);
   U19191 : BUF_X1 port map( A => n21302, Z => n24793);
   U19192 : BUF_X1 port map( A => n21302, Z => n24794);
   U19193 : BUF_X1 port map( A => n21302, Z => n24795);
   U19194 : BUF_X1 port map( A => n21302, Z => n24796);
   U19195 : BUF_X1 port map( A => n22586, Z => n24514);
   U19196 : BUF_X1 port map( A => n22586, Z => n24510);
   U19197 : BUF_X1 port map( A => n22586, Z => n24511);
   U19198 : BUF_X1 port map( A => n22586, Z => n24512);
   U19199 : BUF_X1 port map( A => n22586, Z => n24513);
   U19200 : BUF_X1 port map( A => n22576, Z => n24562);
   U19201 : BUF_X1 port map( A => n22581, Z => n24538);
   U19202 : BUF_X1 port map( A => n22576, Z => n24558);
   U19203 : BUF_X1 port map( A => n22581, Z => n24534);
   U19204 : BUF_X1 port map( A => n22576, Z => n24559);
   U19205 : BUF_X1 port map( A => n22581, Z => n24535);
   U19206 : BUF_X1 port map( A => n22576, Z => n24560);
   U19207 : BUF_X1 port map( A => n22581, Z => n24536);
   U19208 : BUF_X1 port map( A => n22576, Z => n24561);
   U19209 : BUF_X1 port map( A => n22581, Z => n24537);
   U19210 : BUF_X1 port map( A => n21308, Z => n24780);
   U19211 : BUF_X1 port map( A => n21313, Z => n24756);
   U19212 : BUF_X1 port map( A => n21318, Z => n24732);
   U19213 : BUF_X1 port map( A => n21323, Z => n24708);
   U19214 : BUF_X1 port map( A => n21332, Z => n24684);
   U19215 : BUF_X1 port map( A => n21337, Z => n24660);
   U19216 : BUF_X1 port map( A => n21342, Z => n24636);
   U19217 : BUF_X1 port map( A => n21347, Z => n24612);
   U19218 : BUF_X1 port map( A => n21308, Z => n24781);
   U19219 : BUF_X1 port map( A => n21313, Z => n24757);
   U19220 : BUF_X1 port map( A => n21318, Z => n24733);
   U19221 : BUF_X1 port map( A => n21323, Z => n24709);
   U19222 : BUF_X1 port map( A => n21332, Z => n24685);
   U19223 : BUF_X1 port map( A => n21337, Z => n24661);
   U19224 : BUF_X1 port map( A => n21342, Z => n24637);
   U19225 : BUF_X1 port map( A => n21347, Z => n24613);
   U19226 : BUF_X1 port map( A => n21308, Z => n24782);
   U19227 : BUF_X1 port map( A => n21313, Z => n24758);
   U19228 : BUF_X1 port map( A => n21318, Z => n24734);
   U19229 : BUF_X1 port map( A => n21323, Z => n24710);
   U19230 : BUF_X1 port map( A => n21332, Z => n24686);
   U19231 : BUF_X1 port map( A => n21337, Z => n24662);
   U19232 : BUF_X1 port map( A => n21342, Z => n24638);
   U19233 : BUF_X1 port map( A => n21347, Z => n24614);
   U19234 : BUF_X1 port map( A => n21308, Z => n24783);
   U19235 : BUF_X1 port map( A => n21313, Z => n24759);
   U19236 : BUF_X1 port map( A => n21318, Z => n24735);
   U19237 : BUF_X1 port map( A => n21323, Z => n24711);
   U19238 : BUF_X1 port map( A => n21332, Z => n24687);
   U19239 : BUF_X1 port map( A => n21337, Z => n24663);
   U19240 : BUF_X1 port map( A => n21342, Z => n24639);
   U19241 : BUF_X1 port map( A => n21347, Z => n24615);
   U19242 : BUF_X1 port map( A => n21308, Z => n24784);
   U19243 : BUF_X1 port map( A => n21313, Z => n24760);
   U19244 : BUF_X1 port map( A => n21318, Z => n24736);
   U19245 : BUF_X1 port map( A => n21323, Z => n24712);
   U19246 : BUF_X1 port map( A => n21332, Z => n24688);
   U19247 : BUF_X1 port map( A => n21337, Z => n24664);
   U19248 : BUF_X1 port map( A => n21342, Z => n24640);
   U19249 : BUF_X1 port map( A => n21347, Z => n24616);
   U19250 : BUF_X1 port map( A => n22603, Z => n24436);
   U19251 : BUF_X1 port map( A => n22603, Z => n24432);
   U19252 : BUF_X1 port map( A => n22603, Z => n24433);
   U19253 : BUF_X1 port map( A => n22603, Z => n24434);
   U19254 : BUF_X1 port map( A => n22603, Z => n24435);
   U19255 : BUF_X1 port map( A => n22568, Z => n24598);
   U19256 : BUF_X1 port map( A => n22583, Z => n24526);
   U19257 : BUF_X1 port map( A => n22573, Z => n24574);
   U19258 : BUF_X1 port map( A => n22578, Z => n24550);
   U19259 : BUF_X1 port map( A => n22568, Z => n24595);
   U19260 : BUF_X1 port map( A => n22583, Z => n24523);
   U19261 : BUF_X1 port map( A => n22573, Z => n24571);
   U19262 : BUF_X1 port map( A => n22578, Z => n24547);
   U19263 : BUF_X1 port map( A => n22568, Z => n24596);
   U19264 : BUF_X1 port map( A => n22583, Z => n24524);
   U19265 : BUF_X1 port map( A => n22573, Z => n24572);
   U19266 : BUF_X1 port map( A => n22578, Z => n24548);
   U19267 : BUF_X1 port map( A => n22568, Z => n24597);
   U19268 : BUF_X1 port map( A => n22583, Z => n24525);
   U19269 : BUF_X1 port map( A => n22573, Z => n24573);
   U19270 : BUF_X1 port map( A => n22578, Z => n24549);
   U19271 : BUF_X1 port map( A => n22601, Z => n24448);
   U19272 : BUF_X1 port map( A => n22601, Z => n24444);
   U19273 : BUF_X1 port map( A => n22601, Z => n24445);
   U19274 : BUF_X1 port map( A => n22601, Z => n24446);
   U19275 : BUF_X1 port map( A => n22601, Z => n24447);
   U19276 : BUF_X1 port map( A => n22587, Z => n24508);
   U19277 : BUF_X1 port map( A => n22587, Z => n24504);
   U19278 : BUF_X1 port map( A => n22587, Z => n24505);
   U19279 : BUF_X1 port map( A => n22587, Z => n24506);
   U19280 : BUF_X1 port map( A => n22587, Z => n24507);
   U19281 : BUF_X1 port map( A => n22599, Z => n24460);
   U19282 : BUF_X1 port map( A => n22599, Z => n24456);
   U19283 : BUF_X1 port map( A => n22599, Z => n24457);
   U19284 : BUF_X1 port map( A => n22599, Z => n24458);
   U19285 : BUF_X1 port map( A => n22599, Z => n24459);
   U19286 : BUF_X1 port map( A => n22600, Z => n24454);
   U19287 : BUF_X1 port map( A => n22600, Z => n24450);
   U19288 : BUF_X1 port map( A => n22600, Z => n24451);
   U19289 : BUF_X1 port map( A => n22600, Z => n24452);
   U19290 : BUF_X1 port map( A => n22600, Z => n24453);
   U19291 : BUF_X1 port map( A => n22572, Z => n24580);
   U19292 : BUF_X1 port map( A => n22582, Z => n24532);
   U19293 : BUF_X1 port map( A => n22572, Z => n24576);
   U19294 : BUF_X1 port map( A => n22582, Z => n24528);
   U19295 : BUF_X1 port map( A => n22572, Z => n24577);
   U19296 : BUF_X1 port map( A => n22582, Z => n24529);
   U19297 : BUF_X1 port map( A => n22572, Z => n24578);
   U19298 : BUF_X1 port map( A => n22582, Z => n24530);
   U19299 : BUF_X1 port map( A => n22572, Z => n24579);
   U19300 : BUF_X1 port map( A => n22582, Z => n24531);
   U19301 : BUF_X1 port map( A => n22588, Z => n24502);
   U19302 : BUF_X1 port map( A => n22588, Z => n24498);
   U19303 : BUF_X1 port map( A => n22588, Z => n24499);
   U19304 : BUF_X1 port map( A => n22588, Z => n24500);
   U19305 : BUF_X1 port map( A => n22588, Z => n24501);
   U19306 : BUF_X1 port map( A => n25555, Z => n25562);
   U19307 : BUF_X1 port map( A => n25556, Z => n25563);
   U19308 : BUF_X1 port map( A => n25555, Z => n25561);
   U19309 : BUF_X1 port map( A => n25555, Z => n25560);
   U19310 : BUF_X1 port map( A => n25554, Z => n25559);
   U19311 : BUF_X1 port map( A => n25554, Z => n25558);
   U19312 : BUF_X1 port map( A => n25554, Z => n25557);
   U19313 : BUF_X1 port map( A => n21310, Z => n24774);
   U19314 : BUF_X1 port map( A => n21315, Z => n24750);
   U19315 : BUF_X1 port map( A => n21320, Z => n24726);
   U19316 : BUF_X1 port map( A => n21325, Z => n24702);
   U19317 : BUF_X1 port map( A => n21334, Z => n24678);
   U19318 : BUF_X1 port map( A => n21339, Z => n24654);
   U19319 : BUF_X1 port map( A => n21344, Z => n24630);
   U19320 : BUF_X1 port map( A => n21349, Z => n24606);
   U19321 : BUF_X1 port map( A => n21310, Z => n24775);
   U19322 : BUF_X1 port map( A => n21315, Z => n24751);
   U19323 : BUF_X1 port map( A => n21320, Z => n24727);
   U19324 : BUF_X1 port map( A => n21325, Z => n24703);
   U19325 : BUF_X1 port map( A => n21334, Z => n24679);
   U19326 : BUF_X1 port map( A => n21339, Z => n24655);
   U19327 : BUF_X1 port map( A => n21344, Z => n24631);
   U19328 : BUF_X1 port map( A => n21349, Z => n24607);
   U19329 : BUF_X1 port map( A => n21310, Z => n24776);
   U19330 : BUF_X1 port map( A => n21315, Z => n24752);
   U19331 : BUF_X1 port map( A => n21320, Z => n24728);
   U19332 : BUF_X1 port map( A => n21325, Z => n24704);
   U19333 : BUF_X1 port map( A => n21334, Z => n24680);
   U19334 : BUF_X1 port map( A => n21339, Z => n24656);
   U19335 : BUF_X1 port map( A => n21344, Z => n24632);
   U19336 : BUF_X1 port map( A => n21349, Z => n24608);
   U19337 : BUF_X1 port map( A => n21310, Z => n24777);
   U19338 : BUF_X1 port map( A => n21315, Z => n24753);
   U19339 : BUF_X1 port map( A => n21320, Z => n24729);
   U19340 : BUF_X1 port map( A => n21325, Z => n24705);
   U19341 : BUF_X1 port map( A => n21334, Z => n24681);
   U19342 : BUF_X1 port map( A => n21339, Z => n24657);
   U19343 : BUF_X1 port map( A => n21344, Z => n24633);
   U19344 : BUF_X1 port map( A => n21349, Z => n24609);
   U19345 : BUF_X1 port map( A => n21310, Z => n24778);
   U19346 : BUF_X1 port map( A => n21315, Z => n24754);
   U19347 : BUF_X1 port map( A => n21320, Z => n24730);
   U19348 : BUF_X1 port map( A => n21325, Z => n24706);
   U19349 : BUF_X1 port map( A => n21334, Z => n24682);
   U19350 : BUF_X1 port map( A => n21339, Z => n24658);
   U19351 : BUF_X1 port map( A => n21344, Z => n24634);
   U19352 : BUF_X1 port map( A => n21349, Z => n24610);
   U19353 : BUF_X1 port map( A => n22593, Z => n24496);
   U19354 : BUF_X1 port map( A => n22595, Z => n24484);
   U19355 : BUF_X1 port map( A => n22597, Z => n24472);
   U19356 : BUF_X1 port map( A => n22610, Z => n24406);
   U19357 : BUF_X1 port map( A => n22605, Z => n24430);
   U19358 : BUF_X1 port map( A => n22593, Z => n24492);
   U19359 : BUF_X1 port map( A => n22595, Z => n24480);
   U19360 : BUF_X1 port map( A => n22597, Z => n24468);
   U19361 : BUF_X1 port map( A => n22610, Z => n24402);
   U19362 : BUF_X1 port map( A => n22605, Z => n24426);
   U19363 : BUF_X1 port map( A => n22593, Z => n24493);
   U19364 : BUF_X1 port map( A => n22595, Z => n24481);
   U19365 : BUF_X1 port map( A => n22597, Z => n24469);
   U19366 : BUF_X1 port map( A => n22610, Z => n24403);
   U19367 : BUF_X1 port map( A => n22605, Z => n24427);
   U19368 : BUF_X1 port map( A => n22593, Z => n24494);
   U19369 : BUF_X1 port map( A => n22595, Z => n24482);
   U19370 : BUF_X1 port map( A => n22597, Z => n24470);
   U19371 : BUF_X1 port map( A => n22610, Z => n24404);
   U19372 : BUF_X1 port map( A => n22605, Z => n24428);
   U19373 : BUF_X1 port map( A => n22593, Z => n24495);
   U19374 : BUF_X1 port map( A => n22595, Z => n24483);
   U19375 : BUF_X1 port map( A => n22597, Z => n24471);
   U19376 : BUF_X1 port map( A => n22610, Z => n24405);
   U19377 : BUF_X1 port map( A => n22605, Z => n24429);
   U19378 : BUF_X1 port map( A => n21311, Z => n24768);
   U19379 : BUF_X1 port map( A => n21316, Z => n24744);
   U19380 : BUF_X1 port map( A => n21321, Z => n24720);
   U19381 : BUF_X1 port map( A => n21326, Z => n24696);
   U19382 : BUF_X1 port map( A => n21335, Z => n24672);
   U19383 : BUF_X1 port map( A => n21340, Z => n24648);
   U19384 : BUF_X1 port map( A => n21345, Z => n24624);
   U19385 : BUF_X1 port map( A => n21350, Z => n24600);
   U19386 : BUF_X1 port map( A => n21311, Z => n24769);
   U19387 : BUF_X1 port map( A => n21316, Z => n24745);
   U19388 : BUF_X1 port map( A => n21321, Z => n24721);
   U19389 : BUF_X1 port map( A => n21326, Z => n24697);
   U19390 : BUF_X1 port map( A => n21335, Z => n24673);
   U19391 : BUF_X1 port map( A => n21340, Z => n24649);
   U19392 : BUF_X1 port map( A => n21345, Z => n24625);
   U19393 : BUF_X1 port map( A => n21350, Z => n24601);
   U19394 : BUF_X1 port map( A => n21311, Z => n24770);
   U19395 : BUF_X1 port map( A => n21316, Z => n24746);
   U19396 : BUF_X1 port map( A => n21321, Z => n24722);
   U19397 : BUF_X1 port map( A => n21326, Z => n24698);
   U19398 : BUF_X1 port map( A => n21335, Z => n24674);
   U19399 : BUF_X1 port map( A => n21340, Z => n24650);
   U19400 : BUF_X1 port map( A => n21345, Z => n24626);
   U19401 : BUF_X1 port map( A => n21350, Z => n24602);
   U19402 : BUF_X1 port map( A => n21311, Z => n24771);
   U19403 : BUF_X1 port map( A => n21316, Z => n24747);
   U19404 : BUF_X1 port map( A => n21321, Z => n24723);
   U19405 : BUF_X1 port map( A => n21326, Z => n24699);
   U19406 : BUF_X1 port map( A => n21335, Z => n24675);
   U19407 : BUF_X1 port map( A => n21340, Z => n24651);
   U19408 : BUF_X1 port map( A => n21345, Z => n24627);
   U19409 : BUF_X1 port map( A => n21350, Z => n24603);
   U19410 : BUF_X1 port map( A => n21311, Z => n24772);
   U19411 : BUF_X1 port map( A => n21316, Z => n24748);
   U19412 : BUF_X1 port map( A => n21321, Z => n24724);
   U19413 : BUF_X1 port map( A => n21326, Z => n24700);
   U19414 : BUF_X1 port map( A => n21335, Z => n24676);
   U19415 : BUF_X1 port map( A => n21340, Z => n24652);
   U19416 : BUF_X1 port map( A => n21345, Z => n24628);
   U19417 : BUF_X1 port map( A => n21350, Z => n24604);
   U19418 : BUF_X1 port map( A => n22596, Z => n24478);
   U19419 : BUF_X1 port map( A => n22611, Z => n24400);
   U19420 : BUF_X1 port map( A => n22606, Z => n24424);
   U19421 : BUF_X1 port map( A => n22596, Z => n24474);
   U19422 : BUF_X1 port map( A => n22611, Z => n24396);
   U19423 : BUF_X1 port map( A => n22606, Z => n24420);
   U19424 : BUF_X1 port map( A => n22596, Z => n24475);
   U19425 : BUF_X1 port map( A => n22611, Z => n24397);
   U19426 : BUF_X1 port map( A => n22606, Z => n24421);
   U19427 : BUF_X1 port map( A => n22596, Z => n24476);
   U19428 : BUF_X1 port map( A => n22611, Z => n24398);
   U19429 : BUF_X1 port map( A => n22606, Z => n24422);
   U19430 : BUF_X1 port map( A => n22596, Z => n24477);
   U19431 : BUF_X1 port map( A => n22611, Z => n24399);
   U19432 : BUF_X1 port map( A => n22606, Z => n24423);
   U19433 : NAND2_X1 port map( A1 => n23754, A2 => n23755, ZN => n22594);
   U19434 : NAND2_X1 port map( A1 => n23739, A2 => n23744, ZN => n22574);
   U19435 : BUF_X1 port map( A => n22569, Z => n24592);
   U19436 : BUF_X1 port map( A => n22584, Z => n24520);
   U19437 : BUF_X1 port map( A => n22579, Z => n24544);
   U19438 : BUF_X1 port map( A => n22569, Z => n24588);
   U19439 : BUF_X1 port map( A => n22584, Z => n24516);
   U19440 : BUF_X1 port map( A => n22579, Z => n24540);
   U19441 : BUF_X1 port map( A => n22569, Z => n24589);
   U19442 : BUF_X1 port map( A => n22584, Z => n24517);
   U19443 : BUF_X1 port map( A => n22579, Z => n24541);
   U19444 : BUF_X1 port map( A => n22569, Z => n24590);
   U19445 : BUF_X1 port map( A => n22584, Z => n24518);
   U19446 : BUF_X1 port map( A => n22579, Z => n24542);
   U19447 : BUF_X1 port map( A => n22569, Z => n24591);
   U19448 : BUF_X1 port map( A => n22584, Z => n24519);
   U19449 : BUF_X1 port map( A => n22579, Z => n24543);
   U19450 : BUF_X1 port map( A => n22568, Z => n24594);
   U19451 : BUF_X1 port map( A => n22583, Z => n24522);
   U19452 : BUF_X1 port map( A => n22573, Z => n24570);
   U19453 : BUF_X1 port map( A => n22578, Z => n24546);
   U19454 : BUF_X1 port map( A => n25556, Z => n25564);
   U19455 : AND2_X1 port map( A1 => n23739, A2 => n23740, ZN => n22571);
   U19456 : AND2_X1 port map( A1 => n23739, A2 => n23737, ZN => n22577);
   U19457 : AND2_X1 port map( A1 => n23739, A2 => n23747, ZN => n22602);
   U19458 : BUF_X1 port map( A => n21189, Z => n25534);
   U19459 : OAI21_X1 port map( B1 => n21253, B2 => n21254, A => n25562, ZN => 
                           n21189);
   U19460 : BUF_X1 port map( A => n21296, Z => n24815);
   U19461 : BUF_X1 port map( A => n21296, Z => n24816);
   U19462 : INV_X1 port map( A => n24987, ZN => n25003);
   U19463 : INV_X1 port map( A => n25208, ZN => n25224);
   U19464 : INV_X1 port map( A => n25140, ZN => n25156);
   U19465 : INV_X1 port map( A => n24885, ZN => n24901);
   U19466 : INV_X1 port map( A => n25072, ZN => n25088);
   U19467 : INV_X1 port map( A => n25004, ZN => n25020);
   U19468 : INV_X1 port map( A => n24902, ZN => n24918);
   U19469 : INV_X1 port map( A => n24834, ZN => n24850);
   U19470 : INV_X1 port map( A => n25055, ZN => n25071);
   U19471 : INV_X1 port map( A => n25191, ZN => n25207);
   U19472 : INV_X1 port map( A => n25174, ZN => n25190);
   U19473 : INV_X1 port map( A => n25089, ZN => n25105);
   U19474 : INV_X1 port map( A => n25038, ZN => n25054);
   U19475 : INV_X1 port map( A => n25021, ZN => n25037);
   U19476 : INV_X1 port map( A => n24851, ZN => n24867);
   U19477 : INV_X1 port map( A => n24868, ZN => n24884);
   U19478 : INV_X1 port map( A => n24919, ZN => n24935);
   U19479 : INV_X1 port map( A => n24936, ZN => n24952);
   U19480 : INV_X1 port map( A => n24953, ZN => n24969);
   U19481 : INV_X1 port map( A => n24970, ZN => n24986);
   U19482 : INV_X1 port map( A => n25106, ZN => n25122);
   U19483 : INV_X1 port map( A => n25123, ZN => n25139);
   U19484 : INV_X1 port map( A => n25157, ZN => n25173);
   U19485 : INV_X1 port map( A => n25225, ZN => n25241);
   U19486 : INV_X1 port map( A => n25242, ZN => n25258);
   U19487 : INV_X1 port map( A => n25310, ZN => n25326);
   U19488 : INV_X1 port map( A => n25293, ZN => n25309);
   U19489 : INV_X1 port map( A => n25327, ZN => n25344);
   U19490 : INV_X1 port map( A => n25259, ZN => n25275);
   U19491 : INV_X1 port map( A => n25276, ZN => n25292);
   U19492 : OAI22_X1 port map( A1 => n21151, A2 => n24497, B1 => n20525, B2 => 
                           n24491, ZN => n22663);
   U19493 : OAI22_X1 port map( A1 => n21150, A2 => n24497, B1 => n20524, B2 => 
                           n24491, ZN => n22645);
   U19494 : OAI22_X1 port map( A1 => n21148, A2 => n24497, B1 => n20523, B2 => 
                           n24491, ZN => n22627);
   U19495 : OAI22_X1 port map( A1 => n21149, A2 => n24497, B1 => n20522, B2 => 
                           n24491, ZN => n22592);
   U19496 : OAI22_X1 port map( A1 => n19271, A2 => n24485, B1 => n20261, B2 => 
                           n24479, ZN => n22662);
   U19497 : OAI22_X1 port map( A1 => n19270, A2 => n24485, B1 => n20260, B2 => 
                           n24479, ZN => n22644);
   U19498 : OAI22_X1 port map( A1 => n19269, A2 => n24485, B1 => n20259, B2 => 
                           n24479, ZN => n22626);
   U19499 : OAI22_X1 port map( A1 => n19268, A2 => n24485, B1 => n20258, B2 => 
                           n24479, ZN => n22591);
   U19500 : OAI22_X1 port map( A1 => n20542, A2 => n24473, B1 => n19207, B2 => 
                           n24467, ZN => n22661);
   U19501 : OAI22_X1 port map( A1 => n20541, A2 => n24473, B1 => n19206, B2 => 
                           n24467, ZN => n22643);
   U19502 : OAI22_X1 port map( A1 => n20540, A2 => n24473, B1 => n19205, B2 => 
                           n24467, ZN => n22625);
   U19503 : OAI22_X1 port map( A1 => n20539, A2 => n24473, B1 => n19204, B2 => 
                           n24467, ZN => n22590);
   U19504 : OAI22_X1 port map( A1 => n21159, A2 => n24496, B1 => n20698, B2 => 
                           n24490, ZN => n22807);
   U19505 : OAI22_X1 port map( A1 => n21158, A2 => n24496, B1 => n20697, B2 => 
                           n24490, ZN => n22789);
   U19506 : OAI22_X1 port map( A1 => n21157, A2 => n24496, B1 => n20696, B2 => 
                           n24490, ZN => n22771);
   U19507 : OAI22_X1 port map( A1 => n21156, A2 => n24496, B1 => n20695, B2 => 
                           n24490, ZN => n22753);
   U19508 : OAI22_X1 port map( A1 => n21155, A2 => n24496, B1 => n20694, B2 => 
                           n24490, ZN => n22735);
   U19509 : OAI22_X1 port map( A1 => n21154, A2 => n24496, B1 => n20693, B2 => 
                           n24490, ZN => n22717);
   U19510 : OAI22_X1 port map( A1 => n21153, A2 => n24496, B1 => n20692, B2 => 
                           n24490, ZN => n22699);
   U19511 : OAI22_X1 port map( A1 => n21152, A2 => n24496, B1 => n20691, B2 => 
                           n24490, ZN => n22681);
   U19512 : OAI22_X1 port map( A1 => n21187, A2 => n24492, B1 => n20846, B2 => 
                           n24486, ZN => n23753);
   U19513 : OAI22_X1 port map( A1 => n21147, A2 => n24492, B1 => n20845, B2 => 
                           n24486, ZN => n23725);
   U19514 : OAI22_X1 port map( A1 => n21186, A2 => n24492, B1 => n20844, B2 => 
                           n24486, ZN => n23707);
   U19515 : OAI22_X1 port map( A1 => n21185, A2 => n24492, B1 => n20843, B2 => 
                           n24486, ZN => n23689);
   U19516 : OAI22_X1 port map( A1 => n21184, A2 => n24492, B1 => n20842, B2 => 
                           n24486, ZN => n23671);
   U19517 : OAI22_X1 port map( A1 => n21183, A2 => n24492, B1 => n20841, B2 => 
                           n24486, ZN => n23653);
   U19518 : OAI22_X1 port map( A1 => n21182, A2 => n24492, B1 => n20840, B2 => 
                           n24486, ZN => n23635);
   U19519 : OAI22_X1 port map( A1 => n21181, A2 => n24492, B1 => n20839, B2 => 
                           n24486, ZN => n23617);
   U19520 : OAI22_X1 port map( A1 => n21180, A2 => n24492, B1 => n20838, B2 => 
                           n24486, ZN => n23599);
   U19521 : OAI22_X1 port map( A1 => n21179, A2 => n24492, B1 => n20837, B2 => 
                           n24486, ZN => n23581);
   U19522 : OAI22_X1 port map( A1 => n21178, A2 => n24492, B1 => n20836, B2 => 
                           n24486, ZN => n23563);
   U19523 : OAI22_X1 port map( A1 => n21177, A2 => n24492, B1 => n20835, B2 => 
                           n24486, ZN => n23545);
   U19524 : OAI22_X1 port map( A1 => n21176, A2 => n24493, B1 => n20834, B2 => 
                           n24487, ZN => n23527);
   U19525 : OAI22_X1 port map( A1 => n21175, A2 => n24493, B1 => n20833, B2 => 
                           n24487, ZN => n23509);
   U19526 : OAI22_X1 port map( A1 => n21174, A2 => n24493, B1 => n20832, B2 => 
                           n24487, ZN => n23491);
   U19527 : OAI22_X1 port map( A1 => n21173, A2 => n24493, B1 => n20831, B2 => 
                           n24487, ZN => n23473);
   U19528 : OAI22_X1 port map( A1 => n21172, A2 => n24493, B1 => n20830, B2 => 
                           n24487, ZN => n23455);
   U19529 : OAI22_X1 port map( A1 => n21171, A2 => n24493, B1 => n20829, B2 => 
                           n24487, ZN => n23437);
   U19530 : OAI22_X1 port map( A1 => n21170, A2 => n24493, B1 => n20828, B2 => 
                           n24487, ZN => n23419);
   U19531 : OAI22_X1 port map( A1 => n21169, A2 => n24493, B1 => n20827, B2 => 
                           n24487, ZN => n23401);
   U19532 : OAI22_X1 port map( A1 => n21168, A2 => n24493, B1 => n20826, B2 => 
                           n24487, ZN => n23383);
   U19533 : OAI22_X1 port map( A1 => n21167, A2 => n24493, B1 => n20825, B2 => 
                           n24487, ZN => n23365);
   U19534 : OAI22_X1 port map( A1 => n21166, A2 => n24493, B1 => n20824, B2 => 
                           n24487, ZN => n23347);
   U19535 : OAI22_X1 port map( A1 => n21165, A2 => n24493, B1 => n20823, B2 => 
                           n24487, ZN => n23329);
   U19536 : OAI22_X1 port map( A1 => n21164, A2 => n24494, B1 => n20726, B2 => 
                           n24488, ZN => n23311);
   U19537 : OAI22_X1 port map( A1 => n21163, A2 => n24494, B1 => n20725, B2 => 
                           n24488, ZN => n23293);
   U19538 : OAI22_X1 port map( A1 => n21162, A2 => n24494, B1 => n20724, B2 => 
                           n24488, ZN => n23275);
   U19539 : OAI22_X1 port map( A1 => n21161, A2 => n24494, B1 => n20723, B2 => 
                           n24488, ZN => n23257);
   U19540 : OAI22_X1 port map( A1 => n21160, A2 => n24494, B1 => n20722, B2 => 
                           n24488, ZN => n23239);
   U19541 : OAI22_X1 port map( A1 => n20998, A2 => n24471, B1 => n19227, B2 => 
                           n24465, ZN => n23021);
   U19542 : OAI22_X1 port map( A1 => n20997, A2 => n24471, B1 => n19226, B2 => 
                           n24465, ZN => n23003);
   U19543 : OAI22_X1 port map( A1 => n20996, A2 => n24471, B1 => n19225, B2 => 
                           n24465, ZN => n22985);
   U19544 : OAI22_X1 port map( A1 => n20995, A2 => n24471, B1 => n19224, B2 => 
                           n24465, ZN => n22967);
   U19545 : OAI22_X1 port map( A1 => n20994, A2 => n24471, B1 => n19223, B2 => 
                           n24465, ZN => n22949);
   U19546 : OAI22_X1 port map( A1 => n20993, A2 => n24471, B1 => n19222, B2 => 
                           n24465, ZN => n22931);
   U19547 : OAI22_X1 port map( A1 => n20992, A2 => n24471, B1 => n19221, B2 => 
                           n24465, ZN => n22913);
   U19548 : OAI22_X1 port map( A1 => n20991, A2 => n24471, B1 => n19220, B2 => 
                           n24465, ZN => n22895);
   U19549 : OAI22_X1 port map( A1 => n20990, A2 => n24472, B1 => n19219, B2 => 
                           n24466, ZN => n22877);
   U19550 : OAI22_X1 port map( A1 => n20989, A2 => n24472, B1 => n19218, B2 => 
                           n24466, ZN => n22859);
   U19551 : OAI22_X1 port map( A1 => n20988, A2 => n24472, B1 => n19217, B2 => 
                           n24466, ZN => n22841);
   U19552 : OAI22_X1 port map( A1 => n20987, A2 => n24472, B1 => n19216, B2 => 
                           n24466, ZN => n22823);
   U19553 : OAI22_X1 port map( A1 => n20986, A2 => n24472, B1 => n19215, B2 => 
                           n24466, ZN => n22805);
   U19554 : OAI22_X1 port map( A1 => n20985, A2 => n24472, B1 => n19214, B2 => 
                           n24466, ZN => n22787);
   U19555 : OAI22_X1 port map( A1 => n20984, A2 => n24472, B1 => n19213, B2 => 
                           n24466, ZN => n22769);
   U19556 : OAI22_X1 port map( A1 => n20983, A2 => n24472, B1 => n19212, B2 => 
                           n24466, ZN => n22751);
   U19557 : OAI22_X1 port map( A1 => n20982, A2 => n24472, B1 => n19211, B2 => 
                           n24466, ZN => n22733);
   U19558 : OAI22_X1 port map( A1 => n20981, A2 => n24472, B1 => n19210, B2 => 
                           n24466, ZN => n22715);
   U19559 : OAI22_X1 port map( A1 => n20980, A2 => n24472, B1 => n19209, B2 => 
                           n24466, ZN => n22697);
   U19560 : OAI22_X1 port map( A1 => n20979, A2 => n24472, B1 => n19208, B2 => 
                           n24466, ZN => n22679);
   U19561 : OAI22_X1 port map( A1 => n21122, A2 => n24468, B1 => n19267, B2 => 
                           n24462, ZN => n23751);
   U19562 : OAI22_X1 port map( A1 => n21121, A2 => n24468, B1 => n19266, B2 => 
                           n24462, ZN => n23723);
   U19563 : OAI22_X1 port map( A1 => n21120, A2 => n24468, B1 => n19265, B2 => 
                           n24462, ZN => n23705);
   U19564 : OAI22_X1 port map( A1 => n21119, A2 => n24468, B1 => n19264, B2 => 
                           n24462, ZN => n23687);
   U19565 : OAI22_X1 port map( A1 => n21118, A2 => n24468, B1 => n19263, B2 => 
                           n24462, ZN => n23669);
   U19566 : OAI22_X1 port map( A1 => n21117, A2 => n24468, B1 => n19262, B2 => 
                           n24462, ZN => n23651);
   U19567 : OAI22_X1 port map( A1 => n21116, A2 => n24468, B1 => n19261, B2 => 
                           n24462, ZN => n23633);
   U19568 : OAI22_X1 port map( A1 => n21115, A2 => n24468, B1 => n19260, B2 => 
                           n24462, ZN => n23615);
   U19569 : OAI22_X1 port map( A1 => n21114, A2 => n24468, B1 => n19259, B2 => 
                           n24462, ZN => n23597);
   U19570 : OAI22_X1 port map( A1 => n21113, A2 => n24468, B1 => n19258, B2 => 
                           n24462, ZN => n23579);
   U19571 : OAI22_X1 port map( A1 => n21112, A2 => n24468, B1 => n19257, B2 => 
                           n24462, ZN => n23561);
   U19572 : OAI22_X1 port map( A1 => n21111, A2 => n24468, B1 => n19256, B2 => 
                           n24462, ZN => n23543);
   U19573 : OAI22_X1 port map( A1 => n21110, A2 => n24469, B1 => n19255, B2 => 
                           n24463, ZN => n23525);
   U19574 : OAI22_X1 port map( A1 => n21109, A2 => n24469, B1 => n19254, B2 => 
                           n24463, ZN => n23507);
   U19575 : OAI22_X1 port map( A1 => n21108, A2 => n24469, B1 => n19253, B2 => 
                           n24463, ZN => n23489);
   U19576 : OAI22_X1 port map( A1 => n21107, A2 => n24469, B1 => n19252, B2 => 
                           n24463, ZN => n23471);
   U19577 : OAI22_X1 port map( A1 => n21106, A2 => n24469, B1 => n19251, B2 => 
                           n24463, ZN => n23453);
   U19578 : OAI22_X1 port map( A1 => n21105, A2 => n24469, B1 => n19250, B2 => 
                           n24463, ZN => n23435);
   U19579 : OAI22_X1 port map( A1 => n21104, A2 => n24469, B1 => n19249, B2 => 
                           n24463, ZN => n23417);
   U19580 : OAI22_X1 port map( A1 => n21103, A2 => n24469, B1 => n19248, B2 => 
                           n24463, ZN => n23399);
   U19581 : OAI22_X1 port map( A1 => n21102, A2 => n24469, B1 => n19247, B2 => 
                           n24463, ZN => n23381);
   U19582 : OAI22_X1 port map( A1 => n21101, A2 => n24469, B1 => n19246, B2 => 
                           n24463, ZN => n23363);
   U19583 : OAI22_X1 port map( A1 => n21100, A2 => n24469, B1 => n19245, B2 => 
                           n24463, ZN => n23345);
   U19584 : OAI22_X1 port map( A1 => n21099, A2 => n24469, B1 => n19244, B2 => 
                           n24463, ZN => n23327);
   U19585 : OAI22_X1 port map( A1 => n21014, A2 => n24470, B1 => n19243, B2 => 
                           n24464, ZN => n23309);
   U19586 : OAI22_X1 port map( A1 => n21013, A2 => n24470, B1 => n19242, B2 => 
                           n24464, ZN => n23291);
   U19587 : OAI22_X1 port map( A1 => n21012, A2 => n24470, B1 => n19241, B2 => 
                           n24464, ZN => n23273);
   U19588 : OAI22_X1 port map( A1 => n21011, A2 => n24470, B1 => n19240, B2 => 
                           n24464, ZN => n23255);
   U19589 : OAI22_X1 port map( A1 => n21010, A2 => n24470, B1 => n19239, B2 => 
                           n24464, ZN => n23237);
   U19590 : OAI22_X1 port map( A1 => n21009, A2 => n24470, B1 => n19238, B2 => 
                           n24464, ZN => n23219);
   U19591 : OAI22_X1 port map( A1 => n21008, A2 => n24470, B1 => n19237, B2 => 
                           n24464, ZN => n23201);
   U19592 : OAI22_X1 port map( A1 => n21007, A2 => n24470, B1 => n19236, B2 => 
                           n24464, ZN => n23183);
   U19593 : OAI22_X1 port map( A1 => n21006, A2 => n24470, B1 => n19235, B2 => 
                           n24464, ZN => n23165);
   U19594 : OAI22_X1 port map( A1 => n21005, A2 => n24470, B1 => n19234, B2 => 
                           n24464, ZN => n23147);
   U19595 : OAI22_X1 port map( A1 => n21004, A2 => n24470, B1 => n19233, B2 => 
                           n24464, ZN => n23129);
   U19596 : OAI22_X1 port map( A1 => n21003, A2 => n24470, B1 => n19232, B2 => 
                           n24464, ZN => n23111);
   U19597 : OAI22_X1 port map( A1 => n21002, A2 => n24471, B1 => n19231, B2 => 
                           n24465, ZN => n23093);
   U19598 : OAI22_X1 port map( A1 => n21001, A2 => n24471, B1 => n19230, B2 => 
                           n24465, ZN => n23075);
   U19599 : OAI22_X1 port map( A1 => n21000, A2 => n24471, B1 => n19229, B2 => 
                           n24465, ZN => n23057);
   U19600 : OAI22_X1 port map( A1 => n20999, A2 => n24471, B1 => n19228, B2 => 
                           n24465, ZN => n23039);
   U19601 : OAI22_X1 port map( A1 => n19291, A2 => n24483, B1 => n20357, B2 => 
                           n24477, ZN => n23022);
   U19602 : OAI22_X1 port map( A1 => n19290, A2 => n24483, B1 => n20356, B2 => 
                           n24477, ZN => n23004);
   U19603 : OAI22_X1 port map( A1 => n19289, A2 => n24483, B1 => n20355, B2 => 
                           n24477, ZN => n22986);
   U19604 : OAI22_X1 port map( A1 => n19288, A2 => n24483, B1 => n20354, B2 => 
                           n24477, ZN => n22968);
   U19605 : OAI22_X1 port map( A1 => n19287, A2 => n24483, B1 => n20353, B2 => 
                           n24477, ZN => n22950);
   U19606 : OAI22_X1 port map( A1 => n19286, A2 => n24483, B1 => n20352, B2 => 
                           n24477, ZN => n22932);
   U19607 : OAI22_X1 port map( A1 => n19285, A2 => n24483, B1 => n20351, B2 => 
                           n24477, ZN => n22914);
   U19608 : OAI22_X1 port map( A1 => n19284, A2 => n24483, B1 => n20350, B2 => 
                           n24477, ZN => n22896);
   U19609 : OAI22_X1 port map( A1 => n19283, A2 => n24484, B1 => n20349, B2 => 
                           n24478, ZN => n22878);
   U19610 : OAI22_X1 port map( A1 => n19282, A2 => n24484, B1 => n20348, B2 => 
                           n24478, ZN => n22860);
   U19611 : OAI22_X1 port map( A1 => n19281, A2 => n24484, B1 => n20347, B2 => 
                           n24478, ZN => n22842);
   U19612 : OAI22_X1 port map( A1 => n19280, A2 => n24484, B1 => n20346, B2 => 
                           n24478, ZN => n22824);
   U19613 : OAI22_X1 port map( A1 => n19279, A2 => n24484, B1 => n20345, B2 => 
                           n24478, ZN => n22806);
   U19614 : OAI22_X1 port map( A1 => n19278, A2 => n24484, B1 => n20344, B2 => 
                           n24478, ZN => n22788);
   U19615 : OAI22_X1 port map( A1 => n19277, A2 => n24484, B1 => n20343, B2 => 
                           n24478, ZN => n22770);
   U19616 : OAI22_X1 port map( A1 => n19276, A2 => n24484, B1 => n20342, B2 => 
                           n24478, ZN => n22752);
   U19617 : OAI22_X1 port map( A1 => n19275, A2 => n24484, B1 => n20341, B2 => 
                           n24478, ZN => n22734);
   U19618 : OAI22_X1 port map( A1 => n19274, A2 => n24484, B1 => n20340, B2 => 
                           n24478, ZN => n22716);
   U19619 : OAI22_X1 port map( A1 => n19273, A2 => n24484, B1 => n20339, B2 => 
                           n24478, ZN => n22698);
   U19620 : OAI22_X1 port map( A1 => n19272, A2 => n24484, B1 => n20338, B2 => 
                           n24478, ZN => n22680);
   U19621 : OAI22_X1 port map( A1 => n19331, A2 => n24480, B1 => n20445, B2 => 
                           n24474, ZN => n23752);
   U19622 : OAI22_X1 port map( A1 => n19330, A2 => n24480, B1 => n20444, B2 => 
                           n24474, ZN => n23724);
   U19623 : OAI22_X1 port map( A1 => n19329, A2 => n24480, B1 => n20443, B2 => 
                           n24474, ZN => n23706);
   U19624 : OAI22_X1 port map( A1 => n19328, A2 => n24480, B1 => n20442, B2 => 
                           n24474, ZN => n23688);
   U19625 : OAI22_X1 port map( A1 => n19327, A2 => n24480, B1 => n20441, B2 => 
                           n24474, ZN => n23670);
   U19626 : OAI22_X1 port map( A1 => n19326, A2 => n24480, B1 => n20440, B2 => 
                           n24474, ZN => n23652);
   U19627 : OAI22_X1 port map( A1 => n19325, A2 => n24480, B1 => n20439, B2 => 
                           n24474, ZN => n23634);
   U19628 : OAI22_X1 port map( A1 => n19324, A2 => n24480, B1 => n20438, B2 => 
                           n24474, ZN => n23616);
   U19629 : OAI22_X1 port map( A1 => n19323, A2 => n24480, B1 => n20437, B2 => 
                           n24474, ZN => n23598);
   U19630 : OAI22_X1 port map( A1 => n19322, A2 => n24480, B1 => n20436, B2 => 
                           n24474, ZN => n23580);
   U19631 : OAI22_X1 port map( A1 => n19321, A2 => n24480, B1 => n20435, B2 => 
                           n24474, ZN => n23562);
   U19632 : OAI22_X1 port map( A1 => n19320, A2 => n24480, B1 => n20434, B2 => 
                           n24474, ZN => n23544);
   U19633 : OAI22_X1 port map( A1 => n19319, A2 => n24481, B1 => n20433, B2 => 
                           n24475, ZN => n23526);
   U19634 : OAI22_X1 port map( A1 => n19318, A2 => n24481, B1 => n20432, B2 => 
                           n24475, ZN => n23508);
   U19635 : OAI22_X1 port map( A1 => n19317, A2 => n24481, B1 => n20431, B2 => 
                           n24475, ZN => n23490);
   U19636 : OAI22_X1 port map( A1 => n19316, A2 => n24481, B1 => n20430, B2 => 
                           n24475, ZN => n23472);
   U19637 : OAI22_X1 port map( A1 => n19315, A2 => n24481, B1 => n20429, B2 => 
                           n24475, ZN => n23454);
   U19638 : OAI22_X1 port map( A1 => n19314, A2 => n24481, B1 => n20428, B2 => 
                           n24475, ZN => n23436);
   U19639 : OAI22_X1 port map( A1 => n19313, A2 => n24481, B1 => n20427, B2 => 
                           n24475, ZN => n23418);
   U19640 : OAI22_X1 port map( A1 => n19312, A2 => n24481, B1 => n20426, B2 => 
                           n24475, ZN => n23400);
   U19641 : OAI22_X1 port map( A1 => n19311, A2 => n24481, B1 => n20425, B2 => 
                           n24475, ZN => n23382);
   U19642 : OAI22_X1 port map( A1 => n19310, A2 => n24481, B1 => n20424, B2 => 
                           n24475, ZN => n23364);
   U19643 : OAI22_X1 port map( A1 => n19309, A2 => n24481, B1 => n20423, B2 => 
                           n24475, ZN => n23346);
   U19644 : OAI22_X1 port map( A1 => n19308, A2 => n24481, B1 => n20422, B2 => 
                           n24475, ZN => n23328);
   U19645 : OAI22_X1 port map( A1 => n19307, A2 => n24482, B1 => n20373, B2 => 
                           n24476, ZN => n23310);
   U19646 : OAI22_X1 port map( A1 => n19306, A2 => n24482, B1 => n20372, B2 => 
                           n24476, ZN => n23292);
   U19647 : OAI22_X1 port map( A1 => n19305, A2 => n24482, B1 => n20371, B2 => 
                           n24476, ZN => n23274);
   U19648 : OAI22_X1 port map( A1 => n19304, A2 => n24482, B1 => n20370, B2 => 
                           n24476, ZN => n23256);
   U19649 : OAI22_X1 port map( A1 => n19303, A2 => n24482, B1 => n20369, B2 => 
                           n24476, ZN => n23238);
   U19650 : OAI22_X1 port map( A1 => n19302, A2 => n24482, B1 => n20368, B2 => 
                           n24476, ZN => n23220);
   U19651 : OAI22_X1 port map( A1 => n19301, A2 => n24482, B1 => n20367, B2 => 
                           n24476, ZN => n23202);
   U19652 : OAI22_X1 port map( A1 => n19300, A2 => n24482, B1 => n20366, B2 => 
                           n24476, ZN => n23184);
   U19653 : OAI22_X1 port map( A1 => n19299, A2 => n24482, B1 => n20365, B2 => 
                           n24476, ZN => n23166);
   U19654 : OAI22_X1 port map( A1 => n19298, A2 => n24482, B1 => n20364, B2 => 
                           n24476, ZN => n23148);
   U19655 : OAI22_X1 port map( A1 => n19297, A2 => n24482, B1 => n20363, B2 => 
                           n24476, ZN => n23130);
   U19656 : OAI22_X1 port map( A1 => n19296, A2 => n24482, B1 => n20362, B2 => 
                           n24476, ZN => n23112);
   U19657 : OAI22_X1 port map( A1 => n19295, A2 => n24483, B1 => n20361, B2 => 
                           n24477, ZN => n23094);
   U19658 : OAI22_X1 port map( A1 => n19294, A2 => n24483, B1 => n20360, B2 => 
                           n24477, ZN => n23076);
   U19659 : OAI22_X1 port map( A1 => n19293, A2 => n24483, B1 => n20359, B2 => 
                           n24477, ZN => n23058);
   U19660 : OAI22_X1 port map( A1 => n19292, A2 => n24483, B1 => n20358, B2 => 
                           n24477, ZN => n23040);
   U19661 : OAI22_X1 port map( A1 => n25330, A2 => n25345, B1 => n25328, B2 => 
                           n21187, ZN => n6980);
   U19662 : OAI22_X1 port map( A1 => n25330, A2 => n25351, B1 => n25329, B2 => 
                           n21186, ZN => n6982);
   U19663 : OAI22_X1 port map( A1 => n25330, A2 => n25354, B1 => n25329, B2 => 
                           n21185, ZN => n6983);
   U19664 : OAI22_X1 port map( A1 => n25330, A2 => n25357, B1 => n25329, B2 => 
                           n21184, ZN => n6984);
   U19665 : OAI22_X1 port map( A1 => n25331, A2 => n25360, B1 => n25329, B2 => 
                           n21183, ZN => n6985);
   U19666 : OAI22_X1 port map( A1 => n25331, A2 => n25363, B1 => n25329, B2 => 
                           n21182, ZN => n6986);
   U19667 : OAI22_X1 port map( A1 => n25331, A2 => n25366, B1 => n25329, B2 => 
                           n21181, ZN => n6987);
   U19668 : OAI22_X1 port map( A1 => n25331, A2 => n25369, B1 => n25329, B2 => 
                           n21180, ZN => n6988);
   U19669 : OAI22_X1 port map( A1 => n25331, A2 => n25372, B1 => n25329, B2 => 
                           n21179, ZN => n6989);
   U19670 : OAI22_X1 port map( A1 => n25332, A2 => n25375, B1 => n25329, B2 => 
                           n21178, ZN => n6990);
   U19671 : OAI22_X1 port map( A1 => n25332, A2 => n25378, B1 => n25329, B2 => 
                           n21177, ZN => n6991);
   U19672 : OAI22_X1 port map( A1 => n25332, A2 => n25381, B1 => n25329, B2 => 
                           n21176, ZN => n6992);
   U19673 : OAI22_X1 port map( A1 => n25332, A2 => n25384, B1 => n25329, B2 => 
                           n21175, ZN => n6993);
   U19674 : OAI22_X1 port map( A1 => n25332, A2 => n25387, B1 => n25329, B2 => 
                           n21174, ZN => n6994);
   U19675 : OAI22_X1 port map( A1 => n25333, A2 => n25390, B1 => n25328, B2 => 
                           n21173, ZN => n6995);
   U19676 : OAI22_X1 port map( A1 => n25333, A2 => n25393, B1 => n25328, B2 => 
                           n21172, ZN => n6996);
   U19677 : OAI22_X1 port map( A1 => n25333, A2 => n25396, B1 => n25328, B2 => 
                           n21171, ZN => n6997);
   U19678 : OAI22_X1 port map( A1 => n25333, A2 => n25399, B1 => n25328, B2 => 
                           n21170, ZN => n6998);
   U19679 : OAI22_X1 port map( A1 => n25333, A2 => n25402, B1 => n25328, B2 => 
                           n21169, ZN => n6999);
   U19680 : OAI22_X1 port map( A1 => n25334, A2 => n25405, B1 => n25328, B2 => 
                           n21168, ZN => n7000);
   U19681 : OAI22_X1 port map( A1 => n25334, A2 => n25408, B1 => n25328, B2 => 
                           n21167, ZN => n7001);
   U19682 : OAI22_X1 port map( A1 => n25334, A2 => n25411, B1 => n25328, B2 => 
                           n21166, ZN => n7002);
   U19683 : OAI22_X1 port map( A1 => n25334, A2 => n25414, B1 => n25328, B2 => 
                           n21165, ZN => n7003);
   U19684 : OAI22_X1 port map( A1 => n25334, A2 => n25417, B1 => n25328, B2 => 
                           n21164, ZN => n7004);
   U19685 : OAI22_X1 port map( A1 => n25335, A2 => n25420, B1 => n25328, B2 => 
                           n21163, ZN => n7005);
   U19686 : OAI22_X1 port map( A1 => n25335, A2 => n25423, B1 => n25328, B2 => 
                           n21162, ZN => n7006);
   U19687 : OAI22_X1 port map( A1 => n25335, A2 => n25426, B1 => n25328, B2 => 
                           n21161, ZN => n7007);
   U19688 : OAI22_X1 port map( A1 => n25335, A2 => n25429, B1 => n25327, B2 => 
                           n21160, ZN => n7008);
   U19689 : OAI22_X1 port map( A1 => n25340, A2 => n25501, B1 => n25329, B2 => 
                           n21159, ZN => n7032);
   U19690 : OAI22_X1 port map( A1 => n25340, A2 => n25504, B1 => n25328, B2 => 
                           n21158, ZN => n7033);
   U19691 : OAI22_X1 port map( A1 => n25340, A2 => n25507, B1 => n25327, B2 => 
                           n21157, ZN => n7034);
   U19692 : OAI22_X1 port map( A1 => n25341, A2 => n25510, B1 => n25329, B2 => 
                           n21156, ZN => n7035);
   U19693 : OAI22_X1 port map( A1 => n25341, A2 => n25513, B1 => n25328, B2 => 
                           n21155, ZN => n7036);
   U19694 : OAI22_X1 port map( A1 => n25341, A2 => n25516, B1 => n25327, B2 => 
                           n21154, ZN => n7037);
   U19695 : OAI22_X1 port map( A1 => n25341, A2 => n25519, B1 => n25329, B2 => 
                           n21153, ZN => n7038);
   U19696 : OAI22_X1 port map( A1 => n25341, A2 => n25522, B1 => n25328, B2 => 
                           n21152, ZN => n7039);
   U19697 : OAI22_X1 port map( A1 => n25342, A2 => n25525, B1 => n25327, B2 => 
                           n21151, ZN => n7040);
   U19698 : OAI22_X1 port map( A1 => n25342, A2 => n25528, B1 => n25329, B2 => 
                           n21150, ZN => n7041);
   U19699 : OAI22_X1 port map( A1 => n25342, A2 => n25551, B1 => n25328, B2 => 
                           n21149, ZN => n7043);
   U19700 : OAI22_X1 port map( A1 => n25342, A2 => n25531, B1 => n25327, B2 => 
                           n21148, ZN => n7042);
   U19701 : OAI22_X1 port map( A1 => n24990, A2 => n25346, B1 => n24988, B2 => 
                           n21146, ZN => n5700);
   U19702 : OAI22_X1 port map( A1 => n24990, A2 => n25349, B1 => n24988, B2 => 
                           n21145, ZN => n5701);
   U19703 : OAI22_X1 port map( A1 => n24990, A2 => n25352, B1 => n24988, B2 => 
                           n21144, ZN => n5702);
   U19704 : OAI22_X1 port map( A1 => n24990, A2 => n25355, B1 => n24988, B2 => 
                           n21143, ZN => n5703);
   U19705 : OAI22_X1 port map( A1 => n24990, A2 => n25358, B1 => n24988, B2 => 
                           n21142, ZN => n5704);
   U19706 : OAI22_X1 port map( A1 => n24991, A2 => n25361, B1 => n24988, B2 => 
                           n21141, ZN => n5705);
   U19707 : OAI22_X1 port map( A1 => n24991, A2 => n25364, B1 => n24988, B2 => 
                           n21140, ZN => n5706);
   U19708 : OAI22_X1 port map( A1 => n24991, A2 => n25367, B1 => n24988, B2 => 
                           n21139, ZN => n5707);
   U19709 : OAI22_X1 port map( A1 => n24991, A2 => n25370, B1 => n24988, B2 => 
                           n21138, ZN => n5708);
   U19710 : OAI22_X1 port map( A1 => n24991, A2 => n25373, B1 => n24988, B2 => 
                           n21137, ZN => n5709);
   U19711 : OAI22_X1 port map( A1 => n24992, A2 => n25376, B1 => n24988, B2 => 
                           n21136, ZN => n5710);
   U19712 : OAI22_X1 port map( A1 => n24992, A2 => n25379, B1 => n24988, B2 => 
                           n21135, ZN => n5711);
   U19713 : OAI22_X1 port map( A1 => n24992, A2 => n25382, B1 => n24989, B2 => 
                           n21134, ZN => n5712);
   U19714 : OAI22_X1 port map( A1 => n24992, A2 => n25385, B1 => n24989, B2 => 
                           n21133, ZN => n5713);
   U19715 : OAI22_X1 port map( A1 => n24992, A2 => n25388, B1 => n24989, B2 => 
                           n21132, ZN => n5714);
   U19716 : OAI22_X1 port map( A1 => n24993, A2 => n25391, B1 => n24989, B2 => 
                           n21131, ZN => n5715);
   U19717 : OAI22_X1 port map( A1 => n24993, A2 => n25394, B1 => n24989, B2 => 
                           n21130, ZN => n5716);
   U19718 : OAI22_X1 port map( A1 => n24993, A2 => n25397, B1 => n24989, B2 => 
                           n21129, ZN => n5717);
   U19719 : OAI22_X1 port map( A1 => n24993, A2 => n25400, B1 => n24989, B2 => 
                           n21128, ZN => n5718);
   U19720 : OAI22_X1 port map( A1 => n24993, A2 => n25403, B1 => n24989, B2 => 
                           n21127, ZN => n5719);
   U19721 : OAI22_X1 port map( A1 => n24994, A2 => n25406, B1 => n24989, B2 => 
                           n21126, ZN => n5720);
   U19722 : OAI22_X1 port map( A1 => n24994, A2 => n25409, B1 => n24989, B2 => 
                           n21125, ZN => n5721);
   U19723 : OAI22_X1 port map( A1 => n24994, A2 => n25412, B1 => n24989, B2 => 
                           n21124, ZN => n5722);
   U19724 : OAI22_X1 port map( A1 => n24994, A2 => n25415, B1 => n24989, B2 => 
                           n21123, ZN => n5723);
   U19725 : OAI22_X1 port map( A1 => n25228, A2 => n25345, B1 => n25226, B2 => 
                           n21122, ZN => n6596);
   U19726 : OAI22_X1 port map( A1 => n25228, A2 => n25348, B1 => n25226, B2 => 
                           n21121, ZN => n6597);
   U19727 : OAI22_X1 port map( A1 => n25228, A2 => n25351, B1 => n25226, B2 => 
                           n21120, ZN => n6598);
   U19728 : OAI22_X1 port map( A1 => n25228, A2 => n25354, B1 => n25226, B2 => 
                           n21119, ZN => n6599);
   U19729 : OAI22_X1 port map( A1 => n25228, A2 => n25357, B1 => n25226, B2 => 
                           n21118, ZN => n6600);
   U19730 : OAI22_X1 port map( A1 => n25229, A2 => n25360, B1 => n25226, B2 => 
                           n21117, ZN => n6601);
   U19731 : OAI22_X1 port map( A1 => n25229, A2 => n25363, B1 => n25226, B2 => 
                           n21116, ZN => n6602);
   U19732 : OAI22_X1 port map( A1 => n25229, A2 => n25366, B1 => n25226, B2 => 
                           n21115, ZN => n6603);
   U19733 : OAI22_X1 port map( A1 => n25229, A2 => n25369, B1 => n25226, B2 => 
                           n21114, ZN => n6604);
   U19734 : OAI22_X1 port map( A1 => n25229, A2 => n25372, B1 => n25226, B2 => 
                           n21113, ZN => n6605);
   U19735 : OAI22_X1 port map( A1 => n25230, A2 => n25375, B1 => n25226, B2 => 
                           n21112, ZN => n6606);
   U19736 : OAI22_X1 port map( A1 => n25230, A2 => n25378, B1 => n25226, B2 => 
                           n21111, ZN => n6607);
   U19737 : OAI22_X1 port map( A1 => n25230, A2 => n25381, B1 => n25227, B2 => 
                           n21110, ZN => n6608);
   U19738 : OAI22_X1 port map( A1 => n25230, A2 => n25384, B1 => n25227, B2 => 
                           n21109, ZN => n6609);
   U19739 : OAI22_X1 port map( A1 => n25230, A2 => n25387, B1 => n25227, B2 => 
                           n21108, ZN => n6610);
   U19740 : OAI22_X1 port map( A1 => n25231, A2 => n25390, B1 => n25227, B2 => 
                           n21107, ZN => n6611);
   U19741 : OAI22_X1 port map( A1 => n25231, A2 => n25393, B1 => n25227, B2 => 
                           n21106, ZN => n6612);
   U19742 : OAI22_X1 port map( A1 => n25231, A2 => n25396, B1 => n25227, B2 => 
                           n21105, ZN => n6613);
   U19743 : OAI22_X1 port map( A1 => n25231, A2 => n25399, B1 => n25227, B2 => 
                           n21104, ZN => n6614);
   U19744 : OAI22_X1 port map( A1 => n25231, A2 => n25402, B1 => n25227, B2 => 
                           n21103, ZN => n6615);
   U19745 : OAI22_X1 port map( A1 => n25232, A2 => n25405, B1 => n25227, B2 => 
                           n21102, ZN => n6616);
   U19746 : OAI22_X1 port map( A1 => n25232, A2 => n25408, B1 => n25227, B2 => 
                           n21101, ZN => n6617);
   U19747 : OAI22_X1 port map( A1 => n25232, A2 => n25411, B1 => n25227, B2 => 
                           n21100, ZN => n6618);
   U19748 : OAI22_X1 port map( A1 => n25232, A2 => n25414, B1 => n25227, B2 => 
                           n21099, ZN => n6619);
   U19749 : OAI22_X1 port map( A1 => n25211, A2 => n25345, B1 => n25209, B2 => 
                           n21098, ZN => n6532);
   U19750 : OAI22_X1 port map( A1 => n25211, A2 => n25348, B1 => n25209, B2 => 
                           n21097, ZN => n6533);
   U19751 : OAI22_X1 port map( A1 => n25211, A2 => n25351, B1 => n25209, B2 => 
                           n21096, ZN => n6534);
   U19752 : OAI22_X1 port map( A1 => n25211, A2 => n25354, B1 => n25209, B2 => 
                           n21095, ZN => n6535);
   U19753 : OAI22_X1 port map( A1 => n25211, A2 => n25357, B1 => n25209, B2 => 
                           n21094, ZN => n6536);
   U19754 : OAI22_X1 port map( A1 => n25212, A2 => n25360, B1 => n25209, B2 => 
                           n21093, ZN => n6537);
   U19755 : OAI22_X1 port map( A1 => n25212, A2 => n25363, B1 => n25209, B2 => 
                           n21092, ZN => n6538);
   U19756 : OAI22_X1 port map( A1 => n25212, A2 => n25366, B1 => n25209, B2 => 
                           n21091, ZN => n6539);
   U19757 : OAI22_X1 port map( A1 => n25212, A2 => n25369, B1 => n25209, B2 => 
                           n21090, ZN => n6540);
   U19758 : OAI22_X1 port map( A1 => n25212, A2 => n25372, B1 => n25209, B2 => 
                           n21089, ZN => n6541);
   U19759 : OAI22_X1 port map( A1 => n25213, A2 => n25375, B1 => n25209, B2 => 
                           n21088, ZN => n6542);
   U19760 : OAI22_X1 port map( A1 => n25213, A2 => n25378, B1 => n25209, B2 => 
                           n21087, ZN => n6543);
   U19761 : OAI22_X1 port map( A1 => n25213, A2 => n25381, B1 => n25210, B2 => 
                           n21086, ZN => n6544);
   U19762 : OAI22_X1 port map( A1 => n25213, A2 => n25384, B1 => n25210, B2 => 
                           n21085, ZN => n6545);
   U19763 : OAI22_X1 port map( A1 => n25213, A2 => n25387, B1 => n25210, B2 => 
                           n21084, ZN => n6546);
   U19764 : OAI22_X1 port map( A1 => n25214, A2 => n25390, B1 => n25210, B2 => 
                           n21083, ZN => n6547);
   U19765 : OAI22_X1 port map( A1 => n25214, A2 => n25393, B1 => n25210, B2 => 
                           n21082, ZN => n6548);
   U19766 : OAI22_X1 port map( A1 => n25214, A2 => n25396, B1 => n25210, B2 => 
                           n21081, ZN => n6549);
   U19767 : OAI22_X1 port map( A1 => n25214, A2 => n25399, B1 => n25210, B2 => 
                           n21080, ZN => n6550);
   U19768 : OAI22_X1 port map( A1 => n25214, A2 => n25402, B1 => n25210, B2 => 
                           n21079, ZN => n6551);
   U19769 : OAI22_X1 port map( A1 => n25215, A2 => n25405, B1 => n25210, B2 => 
                           n21078, ZN => n6552);
   U19770 : OAI22_X1 port map( A1 => n25215, A2 => n25408, B1 => n25210, B2 => 
                           n21077, ZN => n6553);
   U19771 : OAI22_X1 port map( A1 => n25215, A2 => n25411, B1 => n25210, B2 => 
                           n21076, ZN => n6554);
   U19772 : OAI22_X1 port map( A1 => n25215, A2 => n25414, B1 => n25210, B2 => 
                           n21075, ZN => n6555);
   U19773 : OAI22_X1 port map( A1 => n25143, A2 => n25346, B1 => n25141, B2 => 
                           n21074, ZN => n6276);
   U19774 : OAI22_X1 port map( A1 => n25143, A2 => n25349, B1 => n25141, B2 => 
                           n21073, ZN => n6277);
   U19775 : OAI22_X1 port map( A1 => n25143, A2 => n25352, B1 => n25141, B2 => 
                           n21072, ZN => n6278);
   U19776 : OAI22_X1 port map( A1 => n25143, A2 => n25355, B1 => n25141, B2 => 
                           n21071, ZN => n6279);
   U19777 : OAI22_X1 port map( A1 => n25143, A2 => n25358, B1 => n25141, B2 => 
                           n21070, ZN => n6280);
   U19778 : OAI22_X1 port map( A1 => n25144, A2 => n25361, B1 => n25141, B2 => 
                           n21069, ZN => n6281);
   U19779 : OAI22_X1 port map( A1 => n25144, A2 => n25364, B1 => n25141, B2 => 
                           n21068, ZN => n6282);
   U19780 : OAI22_X1 port map( A1 => n25144, A2 => n25367, B1 => n25141, B2 => 
                           n21067, ZN => n6283);
   U19781 : OAI22_X1 port map( A1 => n25144, A2 => n25370, B1 => n25141, B2 => 
                           n21066, ZN => n6284);
   U19782 : OAI22_X1 port map( A1 => n25144, A2 => n25373, B1 => n25141, B2 => 
                           n21065, ZN => n6285);
   U19783 : OAI22_X1 port map( A1 => n25145, A2 => n25376, B1 => n25141, B2 => 
                           n21064, ZN => n6286);
   U19784 : OAI22_X1 port map( A1 => n25145, A2 => n25379, B1 => n25141, B2 => 
                           n21063, ZN => n6287);
   U19785 : OAI22_X1 port map( A1 => n25145, A2 => n25382, B1 => n25142, B2 => 
                           n21062, ZN => n6288);
   U19786 : OAI22_X1 port map( A1 => n25145, A2 => n25385, B1 => n25142, B2 => 
                           n21061, ZN => n6289);
   U19787 : OAI22_X1 port map( A1 => n25145, A2 => n25388, B1 => n25142, B2 => 
                           n21060, ZN => n6290);
   U19788 : OAI22_X1 port map( A1 => n25146, A2 => n25391, B1 => n25142, B2 => 
                           n21059, ZN => n6291);
   U19789 : OAI22_X1 port map( A1 => n25146, A2 => n25394, B1 => n25142, B2 => 
                           n21058, ZN => n6292);
   U19790 : OAI22_X1 port map( A1 => n25146, A2 => n25397, B1 => n25142, B2 => 
                           n21057, ZN => n6293);
   U19791 : OAI22_X1 port map( A1 => n25146, A2 => n25400, B1 => n25142, B2 => 
                           n21056, ZN => n6294);
   U19792 : OAI22_X1 port map( A1 => n25146, A2 => n25403, B1 => n25142, B2 => 
                           n21055, ZN => n6295);
   U19793 : OAI22_X1 port map( A1 => n25147, A2 => n25406, B1 => n25142, B2 => 
                           n21054, ZN => n6296);
   U19794 : OAI22_X1 port map( A1 => n25147, A2 => n25409, B1 => n25142, B2 => 
                           n21053, ZN => n6297);
   U19795 : OAI22_X1 port map( A1 => n25147, A2 => n25412, B1 => n25142, B2 => 
                           n21052, ZN => n6298);
   U19796 : OAI22_X1 port map( A1 => n25147, A2 => n25415, B1 => n25142, B2 => 
                           n21051, ZN => n6299);
   U19797 : OAI22_X1 port map( A1 => n25245, A2 => n25345, B1 => n25243, B2 => 
                           n20846, ZN => n6660);
   U19798 : OAI22_X1 port map( A1 => n25245, A2 => n25348, B1 => n25243, B2 => 
                           n20845, ZN => n6661);
   U19799 : OAI22_X1 port map( A1 => n25245, A2 => n25351, B1 => n25243, B2 => 
                           n20844, ZN => n6662);
   U19800 : OAI22_X1 port map( A1 => n25245, A2 => n25354, B1 => n25243, B2 => 
                           n20843, ZN => n6663);
   U19801 : OAI22_X1 port map( A1 => n25245, A2 => n25357, B1 => n25243, B2 => 
                           n20842, ZN => n6664);
   U19802 : OAI22_X1 port map( A1 => n25246, A2 => n25360, B1 => n25243, B2 => 
                           n20841, ZN => n6665);
   U19803 : OAI22_X1 port map( A1 => n25246, A2 => n25363, B1 => n25243, B2 => 
                           n20840, ZN => n6666);
   U19804 : OAI22_X1 port map( A1 => n25246, A2 => n25366, B1 => n25243, B2 => 
                           n20839, ZN => n6667);
   U19805 : OAI22_X1 port map( A1 => n25246, A2 => n25369, B1 => n25243, B2 => 
                           n20838, ZN => n6668);
   U19806 : OAI22_X1 port map( A1 => n25246, A2 => n25372, B1 => n25243, B2 => 
                           n20837, ZN => n6669);
   U19807 : OAI22_X1 port map( A1 => n25247, A2 => n25375, B1 => n25243, B2 => 
                           n20836, ZN => n6670);
   U19808 : OAI22_X1 port map( A1 => n25247, A2 => n25378, B1 => n25243, B2 => 
                           n20835, ZN => n6671);
   U19809 : OAI22_X1 port map( A1 => n25247, A2 => n25381, B1 => n25244, B2 => 
                           n20834, ZN => n6672);
   U19810 : OAI22_X1 port map( A1 => n25247, A2 => n25384, B1 => n25244, B2 => 
                           n20833, ZN => n6673);
   U19811 : OAI22_X1 port map( A1 => n25247, A2 => n25387, B1 => n25244, B2 => 
                           n20832, ZN => n6674);
   U19812 : OAI22_X1 port map( A1 => n25248, A2 => n25390, B1 => n25244, B2 => 
                           n20831, ZN => n6675);
   U19813 : OAI22_X1 port map( A1 => n25248, A2 => n25393, B1 => n25244, B2 => 
                           n20830, ZN => n6676);
   U19814 : OAI22_X1 port map( A1 => n25248, A2 => n25396, B1 => n25244, B2 => 
                           n20829, ZN => n6677);
   U19815 : OAI22_X1 port map( A1 => n25248, A2 => n25399, B1 => n25244, B2 => 
                           n20828, ZN => n6678);
   U19816 : OAI22_X1 port map( A1 => n25248, A2 => n25402, B1 => n25244, B2 => 
                           n20827, ZN => n6679);
   U19817 : OAI22_X1 port map( A1 => n25249, A2 => n25405, B1 => n25244, B2 => 
                           n20826, ZN => n6680);
   U19818 : OAI22_X1 port map( A1 => n25249, A2 => n25408, B1 => n25244, B2 => 
                           n20825, ZN => n6681);
   U19819 : OAI22_X1 port map( A1 => n25249, A2 => n25411, B1 => n25244, B2 => 
                           n20824, ZN => n6682);
   U19820 : OAI22_X1 port map( A1 => n25249, A2 => n25414, B1 => n25244, B2 => 
                           n20823, ZN => n6683);
   U19821 : OAI22_X1 port map( A1 => n25075, A2 => n25346, B1 => n25073, B2 => 
                           n20822, ZN => n6020);
   U19822 : OAI22_X1 port map( A1 => n25075, A2 => n25349, B1 => n25073, B2 => 
                           n20821, ZN => n6021);
   U19823 : OAI22_X1 port map( A1 => n25075, A2 => n25352, B1 => n25073, B2 => 
                           n20820, ZN => n6022);
   U19824 : OAI22_X1 port map( A1 => n25075, A2 => n25355, B1 => n25073, B2 => 
                           n20819, ZN => n6023);
   U19825 : OAI22_X1 port map( A1 => n25075, A2 => n25358, B1 => n25073, B2 => 
                           n20818, ZN => n6024);
   U19826 : OAI22_X1 port map( A1 => n25076, A2 => n25361, B1 => n25073, B2 => 
                           n20817, ZN => n6025);
   U19827 : OAI22_X1 port map( A1 => n25076, A2 => n25364, B1 => n25073, B2 => 
                           n20816, ZN => n6026);
   U19828 : OAI22_X1 port map( A1 => n25076, A2 => n25367, B1 => n25073, B2 => 
                           n20815, ZN => n6027);
   U19829 : OAI22_X1 port map( A1 => n25076, A2 => n25370, B1 => n25073, B2 => 
                           n20814, ZN => n6028);
   U19830 : OAI22_X1 port map( A1 => n25076, A2 => n25373, B1 => n25073, B2 => 
                           n20813, ZN => n6029);
   U19831 : OAI22_X1 port map( A1 => n25077, A2 => n25376, B1 => n25073, B2 => 
                           n20812, ZN => n6030);
   U19832 : OAI22_X1 port map( A1 => n25077, A2 => n25379, B1 => n25073, B2 => 
                           n20811, ZN => n6031);
   U19833 : OAI22_X1 port map( A1 => n25077, A2 => n25382, B1 => n25074, B2 => 
                           n20810, ZN => n6032);
   U19834 : OAI22_X1 port map( A1 => n25077, A2 => n25385, B1 => n25074, B2 => 
                           n20809, ZN => n6033);
   U19835 : OAI22_X1 port map( A1 => n25077, A2 => n25388, B1 => n25074, B2 => 
                           n20808, ZN => n6034);
   U19836 : OAI22_X1 port map( A1 => n25078, A2 => n25391, B1 => n25074, B2 => 
                           n20807, ZN => n6035);
   U19837 : OAI22_X1 port map( A1 => n25078, A2 => n25394, B1 => n25074, B2 => 
                           n20806, ZN => n6036);
   U19838 : OAI22_X1 port map( A1 => n25078, A2 => n25397, B1 => n25074, B2 => 
                           n20805, ZN => n6037);
   U19839 : OAI22_X1 port map( A1 => n25078, A2 => n25400, B1 => n25074, B2 => 
                           n20804, ZN => n6038);
   U19840 : OAI22_X1 port map( A1 => n25078, A2 => n25403, B1 => n25074, B2 => 
                           n20803, ZN => n6039);
   U19841 : OAI22_X1 port map( A1 => n25079, A2 => n25406, B1 => n25074, B2 => 
                           n20802, ZN => n6040);
   U19842 : OAI22_X1 port map( A1 => n25079, A2 => n25409, B1 => n25074, B2 => 
                           n20801, ZN => n6041);
   U19843 : OAI22_X1 port map( A1 => n25079, A2 => n25412, B1 => n25074, B2 => 
                           n20800, ZN => n6042);
   U19844 : OAI22_X1 port map( A1 => n25079, A2 => n25415, B1 => n25074, B2 => 
                           n20799, ZN => n6043);
   U19845 : OAI22_X1 port map( A1 => n25007, A2 => n25346, B1 => n25005, B2 => 
                           n20798, ZN => n5764);
   U19846 : OAI22_X1 port map( A1 => n25007, A2 => n25349, B1 => n25005, B2 => 
                           n20797, ZN => n5765);
   U19847 : OAI22_X1 port map( A1 => n25007, A2 => n25352, B1 => n25005, B2 => 
                           n20796, ZN => n5766);
   U19848 : OAI22_X1 port map( A1 => n25007, A2 => n25355, B1 => n25005, B2 => 
                           n20795, ZN => n5767);
   U19849 : OAI22_X1 port map( A1 => n25007, A2 => n25358, B1 => n25005, B2 => 
                           n20794, ZN => n5768);
   U19850 : OAI22_X1 port map( A1 => n25008, A2 => n25361, B1 => n25005, B2 => 
                           n20793, ZN => n5769);
   U19851 : OAI22_X1 port map( A1 => n25008, A2 => n25364, B1 => n25005, B2 => 
                           n20792, ZN => n5770);
   U19852 : OAI22_X1 port map( A1 => n25008, A2 => n25367, B1 => n25005, B2 => 
                           n20791, ZN => n5771);
   U19853 : OAI22_X1 port map( A1 => n25008, A2 => n25370, B1 => n25005, B2 => 
                           n20790, ZN => n5772);
   U19854 : OAI22_X1 port map( A1 => n25008, A2 => n25373, B1 => n25005, B2 => 
                           n20789, ZN => n5773);
   U19855 : OAI22_X1 port map( A1 => n25009, A2 => n25376, B1 => n25005, B2 => 
                           n20788, ZN => n5774);
   U19856 : OAI22_X1 port map( A1 => n25009, A2 => n25379, B1 => n25005, B2 => 
                           n20787, ZN => n5775);
   U19857 : OAI22_X1 port map( A1 => n25009, A2 => n25382, B1 => n25006, B2 => 
                           n20786, ZN => n5776);
   U19858 : OAI22_X1 port map( A1 => n25009, A2 => n25385, B1 => n25006, B2 => 
                           n20785, ZN => n5777);
   U19859 : OAI22_X1 port map( A1 => n25009, A2 => n25388, B1 => n25006, B2 => 
                           n20784, ZN => n5778);
   U19860 : OAI22_X1 port map( A1 => n25010, A2 => n25391, B1 => n25006, B2 => 
                           n20783, ZN => n5779);
   U19861 : OAI22_X1 port map( A1 => n25010, A2 => n25394, B1 => n25006, B2 => 
                           n20782, ZN => n5780);
   U19862 : OAI22_X1 port map( A1 => n25010, A2 => n25397, B1 => n25006, B2 => 
                           n20781, ZN => n5781);
   U19863 : OAI22_X1 port map( A1 => n25010, A2 => n25400, B1 => n25006, B2 => 
                           n20780, ZN => n5782);
   U19864 : OAI22_X1 port map( A1 => n25010, A2 => n25403, B1 => n25006, B2 => 
                           n20779, ZN => n5783);
   U19865 : OAI22_X1 port map( A1 => n25011, A2 => n25406, B1 => n25006, B2 => 
                           n20778, ZN => n5784);
   U19866 : OAI22_X1 port map( A1 => n25011, A2 => n25409, B1 => n25006, B2 => 
                           n20777, ZN => n5785);
   U19867 : OAI22_X1 port map( A1 => n25011, A2 => n25412, B1 => n25006, B2 => 
                           n20776, ZN => n5786);
   U19868 : OAI22_X1 port map( A1 => n25011, A2 => n25415, B1 => n25006, B2 => 
                           n20775, ZN => n5787);
   U19869 : OAI22_X1 port map( A1 => n24905, A2 => n25347, B1 => n24903, B2 => 
                           n20774, ZN => n5380);
   U19870 : OAI22_X1 port map( A1 => n24905, A2 => n25350, B1 => n24903, B2 => 
                           n20773, ZN => n5381);
   U19871 : OAI22_X1 port map( A1 => n24905, A2 => n25353, B1 => n24903, B2 => 
                           n20772, ZN => n5382);
   U19872 : OAI22_X1 port map( A1 => n24905, A2 => n25356, B1 => n24903, B2 => 
                           n20771, ZN => n5383);
   U19873 : OAI22_X1 port map( A1 => n24905, A2 => n25359, B1 => n24903, B2 => 
                           n20770, ZN => n5384);
   U19874 : OAI22_X1 port map( A1 => n24906, A2 => n25362, B1 => n24903, B2 => 
                           n20769, ZN => n5385);
   U19875 : OAI22_X1 port map( A1 => n24906, A2 => n25365, B1 => n24903, B2 => 
                           n20768, ZN => n5386);
   U19876 : OAI22_X1 port map( A1 => n24906, A2 => n25368, B1 => n24903, B2 => 
                           n20767, ZN => n5387);
   U19877 : OAI22_X1 port map( A1 => n24906, A2 => n25371, B1 => n24903, B2 => 
                           n20766, ZN => n5388);
   U19878 : OAI22_X1 port map( A1 => n24906, A2 => n25374, B1 => n24903, B2 => 
                           n20765, ZN => n5389);
   U19879 : OAI22_X1 port map( A1 => n24907, A2 => n25377, B1 => n24903, B2 => 
                           n20764, ZN => n5390);
   U19880 : OAI22_X1 port map( A1 => n24907, A2 => n25380, B1 => n24903, B2 => 
                           n20763, ZN => n5391);
   U19881 : OAI22_X1 port map( A1 => n24907, A2 => n25383, B1 => n24904, B2 => 
                           n20762, ZN => n5392);
   U19882 : OAI22_X1 port map( A1 => n24907, A2 => n25386, B1 => n24904, B2 => 
                           n20761, ZN => n5393);
   U19883 : OAI22_X1 port map( A1 => n24907, A2 => n25389, B1 => n24904, B2 => 
                           n20760, ZN => n5394);
   U19884 : OAI22_X1 port map( A1 => n24908, A2 => n25392, B1 => n24904, B2 => 
                           n20759, ZN => n5395);
   U19885 : OAI22_X1 port map( A1 => n24908, A2 => n25395, B1 => n24904, B2 => 
                           n20758, ZN => n5396);
   U19886 : OAI22_X1 port map( A1 => n24908, A2 => n25398, B1 => n24904, B2 => 
                           n20757, ZN => n5397);
   U19887 : OAI22_X1 port map( A1 => n24908, A2 => n25401, B1 => n24904, B2 => 
                           n20756, ZN => n5398);
   U19888 : OAI22_X1 port map( A1 => n24908, A2 => n25404, B1 => n24904, B2 => 
                           n20755, ZN => n5399);
   U19889 : OAI22_X1 port map( A1 => n24909, A2 => n25407, B1 => n24904, B2 => 
                           n20754, ZN => n5400);
   U19890 : OAI22_X1 port map( A1 => n24909, A2 => n25410, B1 => n24904, B2 => 
                           n20753, ZN => n5401);
   U19891 : OAI22_X1 port map( A1 => n24909, A2 => n25413, B1 => n24904, B2 => 
                           n20752, ZN => n5402);
   U19892 : OAI22_X1 port map( A1 => n24909, A2 => n25416, B1 => n24904, B2 => 
                           n20751, ZN => n5403);
   U19893 : OAI22_X1 port map( A1 => n24837, A2 => n25347, B1 => n24835, B2 => 
                           n20750, ZN => n5124);
   U19894 : OAI22_X1 port map( A1 => n24837, A2 => n25350, B1 => n24835, B2 => 
                           n20749, ZN => n5125);
   U19895 : OAI22_X1 port map( A1 => n24837, A2 => n25353, B1 => n24835, B2 => 
                           n20748, ZN => n5126);
   U19896 : OAI22_X1 port map( A1 => n24837, A2 => n25356, B1 => n24835, B2 => 
                           n20747, ZN => n5127);
   U19897 : OAI22_X1 port map( A1 => n24837, A2 => n25359, B1 => n24835, B2 => 
                           n20746, ZN => n5128);
   U19898 : OAI22_X1 port map( A1 => n24838, A2 => n25362, B1 => n24835, B2 => 
                           n20745, ZN => n5129);
   U19899 : OAI22_X1 port map( A1 => n24838, A2 => n25365, B1 => n24835, B2 => 
                           n20744, ZN => n5130);
   U19900 : OAI22_X1 port map( A1 => n24838, A2 => n25368, B1 => n24835, B2 => 
                           n20743, ZN => n5131);
   U19901 : OAI22_X1 port map( A1 => n24838, A2 => n25371, B1 => n24835, B2 => 
                           n20742, ZN => n5132);
   U19902 : OAI22_X1 port map( A1 => n24838, A2 => n25374, B1 => n24835, B2 => 
                           n20741, ZN => n5133);
   U19903 : OAI22_X1 port map( A1 => n24839, A2 => n25377, B1 => n24835, B2 => 
                           n20740, ZN => n5134);
   U19904 : OAI22_X1 port map( A1 => n24839, A2 => n25380, B1 => n24835, B2 => 
                           n20739, ZN => n5135);
   U19905 : OAI22_X1 port map( A1 => n24839, A2 => n25383, B1 => n24836, B2 => 
                           n20738, ZN => n5136);
   U19906 : OAI22_X1 port map( A1 => n24839, A2 => n25386, B1 => n24836, B2 => 
                           n20737, ZN => n5137);
   U19907 : OAI22_X1 port map( A1 => n24839, A2 => n25389, B1 => n24836, B2 => 
                           n20736, ZN => n5138);
   U19908 : OAI22_X1 port map( A1 => n24840, A2 => n25392, B1 => n24836, B2 => 
                           n20735, ZN => n5139);
   U19909 : OAI22_X1 port map( A1 => n24840, A2 => n25395, B1 => n24836, B2 => 
                           n20734, ZN => n5140);
   U19910 : OAI22_X1 port map( A1 => n24840, A2 => n25398, B1 => n24836, B2 => 
                           n20733, ZN => n5141);
   U19911 : OAI22_X1 port map( A1 => n24840, A2 => n25401, B1 => n24836, B2 => 
                           n20732, ZN => n5142);
   U19912 : OAI22_X1 port map( A1 => n24840, A2 => n25404, B1 => n24836, B2 => 
                           n20731, ZN => n5143);
   U19913 : OAI22_X1 port map( A1 => n24841, A2 => n25407, B1 => n24836, B2 => 
                           n20730, ZN => n5144);
   U19914 : OAI22_X1 port map( A1 => n24841, A2 => n25410, B1 => n24836, B2 => 
                           n20729, ZN => n5145);
   U19915 : OAI22_X1 port map( A1 => n24841, A2 => n25413, B1 => n24836, B2 => 
                           n20728, ZN => n5146);
   U19916 : OAI22_X1 port map( A1 => n24841, A2 => n25416, B1 => n24836, B2 => 
                           n20727, ZN => n5147);
   U19917 : OAI22_X1 port map( A1 => n25058, A2 => n25346, B1 => n25056, B2 => 
                           n20505, ZN => n5956);
   U19918 : OAI22_X1 port map( A1 => n25058, A2 => n25349, B1 => n25056, B2 => 
                           n20504, ZN => n5957);
   U19919 : OAI22_X1 port map( A1 => n25058, A2 => n25352, B1 => n25056, B2 => 
                           n20503, ZN => n5958);
   U19920 : OAI22_X1 port map( A1 => n25058, A2 => n25355, B1 => n25056, B2 => 
                           n20502, ZN => n5959);
   U19921 : OAI22_X1 port map( A1 => n25058, A2 => n25358, B1 => n25056, B2 => 
                           n20501, ZN => n5960);
   U19922 : OAI22_X1 port map( A1 => n25059, A2 => n25361, B1 => n25056, B2 => 
                           n20500, ZN => n5961);
   U19923 : OAI22_X1 port map( A1 => n25059, A2 => n25364, B1 => n25056, B2 => 
                           n20499, ZN => n5962);
   U19924 : OAI22_X1 port map( A1 => n25059, A2 => n25367, B1 => n25056, B2 => 
                           n20498, ZN => n5963);
   U19925 : OAI22_X1 port map( A1 => n25059, A2 => n25370, B1 => n25056, B2 => 
                           n20497, ZN => n5964);
   U19926 : OAI22_X1 port map( A1 => n25059, A2 => n25373, B1 => n25056, B2 => 
                           n20496, ZN => n5965);
   U19927 : OAI22_X1 port map( A1 => n25060, A2 => n25376, B1 => n25056, B2 => 
                           n20495, ZN => n5966);
   U19928 : OAI22_X1 port map( A1 => n25060, A2 => n25379, B1 => n25056, B2 => 
                           n20494, ZN => n5967);
   U19929 : OAI22_X1 port map( A1 => n25060, A2 => n25382, B1 => n25057, B2 => 
                           n20493, ZN => n5968);
   U19930 : OAI22_X1 port map( A1 => n25060, A2 => n25385, B1 => n25057, B2 => 
                           n20492, ZN => n5969);
   U19931 : OAI22_X1 port map( A1 => n25060, A2 => n25388, B1 => n25057, B2 => 
                           n20491, ZN => n5970);
   U19932 : OAI22_X1 port map( A1 => n25061, A2 => n25391, B1 => n25057, B2 => 
                           n20490, ZN => n5971);
   U19933 : OAI22_X1 port map( A1 => n25061, A2 => n25394, B1 => n25057, B2 => 
                           n20489, ZN => n5972);
   U19934 : OAI22_X1 port map( A1 => n25061, A2 => n25397, B1 => n25057, B2 => 
                           n20488, ZN => n5973);
   U19935 : OAI22_X1 port map( A1 => n25061, A2 => n25400, B1 => n25057, B2 => 
                           n20487, ZN => n5974);
   U19936 : OAI22_X1 port map( A1 => n25061, A2 => n25403, B1 => n25057, B2 => 
                           n20486, ZN => n5975);
   U19937 : OAI22_X1 port map( A1 => n25062, A2 => n25406, B1 => n25057, B2 => 
                           n20485, ZN => n5976);
   U19938 : OAI22_X1 port map( A1 => n25062, A2 => n25409, B1 => n25057, B2 => 
                           n20484, ZN => n5977);
   U19939 : OAI22_X1 port map( A1 => n25062, A2 => n25412, B1 => n25057, B2 => 
                           n20483, ZN => n5978);
   U19940 : OAI22_X1 port map( A1 => n25062, A2 => n25415, B1 => n25057, B2 => 
                           n20482, ZN => n5979);
   U19941 : OAI22_X1 port map( A1 => n25313, A2 => n25345, B1 => n25311, B2 => 
                           n20445, ZN => n6916);
   U19942 : OAI22_X1 port map( A1 => n25313, A2 => n25348, B1 => n25311, B2 => 
                           n20444, ZN => n6917);
   U19943 : OAI22_X1 port map( A1 => n25313, A2 => n25351, B1 => n25311, B2 => 
                           n20443, ZN => n6918);
   U19944 : OAI22_X1 port map( A1 => n25313, A2 => n25354, B1 => n25311, B2 => 
                           n20442, ZN => n6919);
   U19945 : OAI22_X1 port map( A1 => n25313, A2 => n25357, B1 => n25311, B2 => 
                           n20441, ZN => n6920);
   U19946 : OAI22_X1 port map( A1 => n25314, A2 => n25360, B1 => n25311, B2 => 
                           n20440, ZN => n6921);
   U19947 : OAI22_X1 port map( A1 => n25314, A2 => n25363, B1 => n25311, B2 => 
                           n20439, ZN => n6922);
   U19948 : OAI22_X1 port map( A1 => n25314, A2 => n25366, B1 => n25311, B2 => 
                           n20438, ZN => n6923);
   U19949 : OAI22_X1 port map( A1 => n25314, A2 => n25369, B1 => n25311, B2 => 
                           n20437, ZN => n6924);
   U19950 : OAI22_X1 port map( A1 => n25314, A2 => n25372, B1 => n25311, B2 => 
                           n20436, ZN => n6925);
   U19951 : OAI22_X1 port map( A1 => n25315, A2 => n25375, B1 => n25311, B2 => 
                           n20435, ZN => n6926);
   U19952 : OAI22_X1 port map( A1 => n25315, A2 => n25378, B1 => n25311, B2 => 
                           n20434, ZN => n6927);
   U19953 : OAI22_X1 port map( A1 => n25315, A2 => n25381, B1 => n25312, B2 => 
                           n20433, ZN => n6928);
   U19954 : OAI22_X1 port map( A1 => n25315, A2 => n25384, B1 => n25312, B2 => 
                           n20432, ZN => n6929);
   U19955 : OAI22_X1 port map( A1 => n25315, A2 => n25387, B1 => n25312, B2 => 
                           n20431, ZN => n6930);
   U19956 : OAI22_X1 port map( A1 => n25316, A2 => n25390, B1 => n25312, B2 => 
                           n20430, ZN => n6931);
   U19957 : OAI22_X1 port map( A1 => n25316, A2 => n25393, B1 => n25312, B2 => 
                           n20429, ZN => n6932);
   U19958 : OAI22_X1 port map( A1 => n25316, A2 => n25396, B1 => n25312, B2 => 
                           n20428, ZN => n6933);
   U19959 : OAI22_X1 port map( A1 => n25316, A2 => n25399, B1 => n25312, B2 => 
                           n20427, ZN => n6934);
   U19960 : OAI22_X1 port map( A1 => n25316, A2 => n25402, B1 => n25312, B2 => 
                           n20426, ZN => n6935);
   U19961 : OAI22_X1 port map( A1 => n25317, A2 => n25405, B1 => n25312, B2 => 
                           n20425, ZN => n6936);
   U19962 : OAI22_X1 port map( A1 => n25317, A2 => n25408, B1 => n25312, B2 => 
                           n20424, ZN => n6937);
   U19963 : OAI22_X1 port map( A1 => n25317, A2 => n25411, B1 => n25312, B2 => 
                           n20423, ZN => n6938);
   U19964 : OAI22_X1 port map( A1 => n25317, A2 => n25414, B1 => n25312, B2 => 
                           n20422, ZN => n6939);
   U19965 : OAI22_X1 port map( A1 => n25194, A2 => n25345, B1 => n25192, B2 => 
                           n20421, ZN => n6468);
   U19966 : OAI22_X1 port map( A1 => n25194, A2 => n25348, B1 => n25192, B2 => 
                           n20420, ZN => n6469);
   U19967 : OAI22_X1 port map( A1 => n25194, A2 => n25351, B1 => n25192, B2 => 
                           n20419, ZN => n6470);
   U19968 : OAI22_X1 port map( A1 => n25194, A2 => n25354, B1 => n25192, B2 => 
                           n20418, ZN => n6471);
   U19969 : OAI22_X1 port map( A1 => n25194, A2 => n25357, B1 => n25192, B2 => 
                           n20417, ZN => n6472);
   U19970 : OAI22_X1 port map( A1 => n25195, A2 => n25360, B1 => n25192, B2 => 
                           n20416, ZN => n6473);
   U19971 : OAI22_X1 port map( A1 => n25195, A2 => n25363, B1 => n25192, B2 => 
                           n20415, ZN => n6474);
   U19972 : OAI22_X1 port map( A1 => n25195, A2 => n25366, B1 => n25192, B2 => 
                           n20414, ZN => n6475);
   U19973 : OAI22_X1 port map( A1 => n25195, A2 => n25369, B1 => n25192, B2 => 
                           n20413, ZN => n6476);
   U19974 : OAI22_X1 port map( A1 => n25195, A2 => n25372, B1 => n25192, B2 => 
                           n20412, ZN => n6477);
   U19975 : OAI22_X1 port map( A1 => n25196, A2 => n25375, B1 => n25192, B2 => 
                           n20411, ZN => n6478);
   U19976 : OAI22_X1 port map( A1 => n25196, A2 => n25378, B1 => n25192, B2 => 
                           n20410, ZN => n6479);
   U19977 : OAI22_X1 port map( A1 => n25196, A2 => n25381, B1 => n25193, B2 => 
                           n20409, ZN => n6480);
   U19978 : OAI22_X1 port map( A1 => n25196, A2 => n25384, B1 => n25193, B2 => 
                           n20408, ZN => n6481);
   U19979 : OAI22_X1 port map( A1 => n25196, A2 => n25387, B1 => n25193, B2 => 
                           n20407, ZN => n6482);
   U19980 : OAI22_X1 port map( A1 => n25197, A2 => n25390, B1 => n25193, B2 => 
                           n20406, ZN => n6483);
   U19981 : OAI22_X1 port map( A1 => n25197, A2 => n25393, B1 => n25193, B2 => 
                           n20405, ZN => n6484);
   U19982 : OAI22_X1 port map( A1 => n25197, A2 => n25396, B1 => n25193, B2 => 
                           n20404, ZN => n6485);
   U19983 : OAI22_X1 port map( A1 => n25197, A2 => n25399, B1 => n25193, B2 => 
                           n20403, ZN => n6486);
   U19984 : OAI22_X1 port map( A1 => n25197, A2 => n25402, B1 => n25193, B2 => 
                           n20402, ZN => n6487);
   U19985 : OAI22_X1 port map( A1 => n25198, A2 => n25405, B1 => n25193, B2 => 
                           n20401, ZN => n6488);
   U19986 : OAI22_X1 port map( A1 => n25198, A2 => n25408, B1 => n25193, B2 => 
                           n20400, ZN => n6489);
   U19987 : OAI22_X1 port map( A1 => n25198, A2 => n25411, B1 => n25193, B2 => 
                           n20399, ZN => n6490);
   U19988 : OAI22_X1 port map( A1 => n25198, A2 => n25414, B1 => n25193, B2 => 
                           n20398, ZN => n6491);
   U19989 : OAI22_X1 port map( A1 => n25296, A2 => n25345, B1 => n25294, B2 => 
                           n20397, ZN => n6852);
   U19990 : OAI22_X1 port map( A1 => n25296, A2 => n25348, B1 => n25294, B2 => 
                           n20396, ZN => n6853);
   U19991 : OAI22_X1 port map( A1 => n25296, A2 => n25351, B1 => n25294, B2 => 
                           n20395, ZN => n6854);
   U19992 : OAI22_X1 port map( A1 => n25296, A2 => n25354, B1 => n25294, B2 => 
                           n20394, ZN => n6855);
   U19993 : OAI22_X1 port map( A1 => n25296, A2 => n25357, B1 => n25294, B2 => 
                           n20393, ZN => n6856);
   U19994 : OAI22_X1 port map( A1 => n25297, A2 => n25360, B1 => n25294, B2 => 
                           n20392, ZN => n6857);
   U19995 : OAI22_X1 port map( A1 => n25297, A2 => n25363, B1 => n25294, B2 => 
                           n20391, ZN => n6858);
   U19996 : OAI22_X1 port map( A1 => n25297, A2 => n25366, B1 => n25294, B2 => 
                           n20390, ZN => n6859);
   U19997 : OAI22_X1 port map( A1 => n25297, A2 => n25369, B1 => n25294, B2 => 
                           n20389, ZN => n6860);
   U19998 : OAI22_X1 port map( A1 => n25297, A2 => n25372, B1 => n25294, B2 => 
                           n20388, ZN => n6861);
   U19999 : OAI22_X1 port map( A1 => n25298, A2 => n25375, B1 => n25294, B2 => 
                           n20387, ZN => n6862);
   U20000 : OAI22_X1 port map( A1 => n25298, A2 => n25378, B1 => n25294, B2 => 
                           n20386, ZN => n6863);
   U20001 : OAI22_X1 port map( A1 => n25298, A2 => n25381, B1 => n25295, B2 => 
                           n20385, ZN => n6864);
   U20002 : OAI22_X1 port map( A1 => n25298, A2 => n25384, B1 => n25295, B2 => 
                           n20384, ZN => n6865);
   U20003 : OAI22_X1 port map( A1 => n25298, A2 => n25387, B1 => n25295, B2 => 
                           n20383, ZN => n6866);
   U20004 : OAI22_X1 port map( A1 => n25299, A2 => n25390, B1 => n25295, B2 => 
                           n20382, ZN => n6867);
   U20005 : OAI22_X1 port map( A1 => n25299, A2 => n25393, B1 => n25295, B2 => 
                           n20381, ZN => n6868);
   U20006 : OAI22_X1 port map( A1 => n25299, A2 => n25396, B1 => n25295, B2 => 
                           n20380, ZN => n6869);
   U20007 : OAI22_X1 port map( A1 => n25299, A2 => n25399, B1 => n25295, B2 => 
                           n20379, ZN => n6870);
   U20008 : OAI22_X1 port map( A1 => n25299, A2 => n25402, B1 => n25295, B2 => 
                           n20378, ZN => n6871);
   U20009 : OAI22_X1 port map( A1 => n25300, A2 => n25405, B1 => n25295, B2 => 
                           n20377, ZN => n6872);
   U20010 : OAI22_X1 port map( A1 => n25300, A2 => n25408, B1 => n25295, B2 => 
                           n20376, ZN => n6873);
   U20011 : OAI22_X1 port map( A1 => n25300, A2 => n25411, B1 => n25295, B2 => 
                           n20375, ZN => n6874);
   U20012 : OAI22_X1 port map( A1 => n25300, A2 => n25414, B1 => n25295, B2 => 
                           n20374, ZN => n6875);
   U20013 : OAI22_X1 port map( A1 => n24871, A2 => n25347, B1 => n24869, B2 => 
                           n19737, ZN => n5252);
   U20014 : OAI22_X1 port map( A1 => n24871, A2 => n25350, B1 => n24869, B2 => 
                           n19736, ZN => n5253);
   U20015 : OAI22_X1 port map( A1 => n24871, A2 => n25353, B1 => n24869, B2 => 
                           n19735, ZN => n5254);
   U20016 : OAI22_X1 port map( A1 => n24871, A2 => n25356, B1 => n24869, B2 => 
                           n19734, ZN => n5255);
   U20017 : OAI22_X1 port map( A1 => n24871, A2 => n25359, B1 => n24869, B2 => 
                           n19733, ZN => n5256);
   U20018 : OAI22_X1 port map( A1 => n24872, A2 => n25362, B1 => n24869, B2 => 
                           n19732, ZN => n5257);
   U20019 : OAI22_X1 port map( A1 => n24872, A2 => n25365, B1 => n24869, B2 => 
                           n19731, ZN => n5258);
   U20020 : OAI22_X1 port map( A1 => n24872, A2 => n25368, B1 => n24869, B2 => 
                           n19730, ZN => n5259);
   U20021 : OAI22_X1 port map( A1 => n24872, A2 => n25371, B1 => n24869, B2 => 
                           n19729, ZN => n5260);
   U20022 : OAI22_X1 port map( A1 => n24872, A2 => n25374, B1 => n24869, B2 => 
                           n19728, ZN => n5261);
   U20023 : OAI22_X1 port map( A1 => n24873, A2 => n25377, B1 => n24869, B2 => 
                           n19727, ZN => n5262);
   U20024 : OAI22_X1 port map( A1 => n24873, A2 => n25380, B1 => n24869, B2 => 
                           n19726, ZN => n5263);
   U20025 : OAI22_X1 port map( A1 => n24873, A2 => n25383, B1 => n24870, B2 => 
                           n19725, ZN => n5264);
   U20026 : OAI22_X1 port map( A1 => n24873, A2 => n25386, B1 => n24870, B2 => 
                           n19724, ZN => n5265);
   U20027 : OAI22_X1 port map( A1 => n24873, A2 => n25389, B1 => n24870, B2 => 
                           n19723, ZN => n5266);
   U20028 : OAI22_X1 port map( A1 => n24874, A2 => n25392, B1 => n24870, B2 => 
                           n19722, ZN => n5267);
   U20029 : OAI22_X1 port map( A1 => n24874, A2 => n25395, B1 => n24870, B2 => 
                           n19721, ZN => n5268);
   U20030 : OAI22_X1 port map( A1 => n24874, A2 => n25398, B1 => n24870, B2 => 
                           n19720, ZN => n5269);
   U20031 : OAI22_X1 port map( A1 => n24874, A2 => n25401, B1 => n24870, B2 => 
                           n19719, ZN => n5270);
   U20032 : OAI22_X1 port map( A1 => n24874, A2 => n25404, B1 => n24870, B2 => 
                           n19718, ZN => n5271);
   U20033 : OAI22_X1 port map( A1 => n24875, A2 => n25407, B1 => n24870, B2 => 
                           n19717, ZN => n5272);
   U20034 : OAI22_X1 port map( A1 => n24875, A2 => n25410, B1 => n24870, B2 => 
                           n19716, ZN => n5273);
   U20035 : OAI22_X1 port map( A1 => n24875, A2 => n25413, B1 => n24870, B2 => 
                           n19715, ZN => n5274);
   U20036 : OAI22_X1 port map( A1 => n24875, A2 => n25416, B1 => n24870, B2 => 
                           n19714, ZN => n5275);
   U20037 : OAI22_X1 port map( A1 => n24939, A2 => n25347, B1 => n24937, B2 => 
                           n19707, ZN => n5508);
   U20038 : OAI22_X1 port map( A1 => n24939, A2 => n25350, B1 => n24937, B2 => 
                           n19706, ZN => n5509);
   U20039 : OAI22_X1 port map( A1 => n24939, A2 => n25353, B1 => n24937, B2 => 
                           n19705, ZN => n5510);
   U20040 : OAI22_X1 port map( A1 => n24939, A2 => n25356, B1 => n24937, B2 => 
                           n19704, ZN => n5511);
   U20041 : OAI22_X1 port map( A1 => n24939, A2 => n25359, B1 => n24937, B2 => 
                           n19703, ZN => n5512);
   U20042 : OAI22_X1 port map( A1 => n24940, A2 => n25362, B1 => n24937, B2 => 
                           n19702, ZN => n5513);
   U20043 : OAI22_X1 port map( A1 => n24940, A2 => n25365, B1 => n24937, B2 => 
                           n19701, ZN => n5514);
   U20044 : OAI22_X1 port map( A1 => n24940, A2 => n25368, B1 => n24937, B2 => 
                           n19700, ZN => n5515);
   U20045 : OAI22_X1 port map( A1 => n24940, A2 => n25371, B1 => n24937, B2 => 
                           n19699, ZN => n5516);
   U20046 : OAI22_X1 port map( A1 => n24940, A2 => n25374, B1 => n24937, B2 => 
                           n19698, ZN => n5517);
   U20047 : OAI22_X1 port map( A1 => n24941, A2 => n25377, B1 => n24937, B2 => 
                           n19697, ZN => n5518);
   U20048 : OAI22_X1 port map( A1 => n24941, A2 => n25380, B1 => n24937, B2 => 
                           n19696, ZN => n5519);
   U20049 : OAI22_X1 port map( A1 => n24941, A2 => n25383, B1 => n24938, B2 => 
                           n19695, ZN => n5520);
   U20050 : OAI22_X1 port map( A1 => n24941, A2 => n25386, B1 => n24938, B2 => 
                           n19694, ZN => n5521);
   U20051 : OAI22_X1 port map( A1 => n24941, A2 => n25389, B1 => n24938, B2 => 
                           n19693, ZN => n5522);
   U20052 : OAI22_X1 port map( A1 => n24942, A2 => n25392, B1 => n24938, B2 => 
                           n19692, ZN => n5523);
   U20053 : OAI22_X1 port map( A1 => n24942, A2 => n25395, B1 => n24938, B2 => 
                           n19691, ZN => n5524);
   U20054 : OAI22_X1 port map( A1 => n24942, A2 => n25398, B1 => n24938, B2 => 
                           n19690, ZN => n5525);
   U20055 : OAI22_X1 port map( A1 => n24942, A2 => n25401, B1 => n24938, B2 => 
                           n19689, ZN => n5526);
   U20056 : OAI22_X1 port map( A1 => n24942, A2 => n25404, B1 => n24938, B2 => 
                           n19688, ZN => n5527);
   U20057 : OAI22_X1 port map( A1 => n24943, A2 => n25407, B1 => n24938, B2 => 
                           n19687, ZN => n5528);
   U20058 : OAI22_X1 port map( A1 => n24943, A2 => n25410, B1 => n24938, B2 => 
                           n19686, ZN => n5529);
   U20059 : OAI22_X1 port map( A1 => n24943, A2 => n25413, B1 => n24938, B2 => 
                           n19685, ZN => n5530);
   U20060 : OAI22_X1 port map( A1 => n24943, A2 => n25416, B1 => n24938, B2 => 
                           n19684, ZN => n5531);
   U20061 : OAI22_X1 port map( A1 => n25279, A2 => n25345, B1 => n25277, B2 => 
                           n19395, ZN => n6788);
   U20062 : OAI22_X1 port map( A1 => n25279, A2 => n25348, B1 => n25277, B2 => 
                           n19394, ZN => n6789);
   U20063 : OAI22_X1 port map( A1 => n25279, A2 => n25351, B1 => n25277, B2 => 
                           n19393, ZN => n6790);
   U20064 : OAI22_X1 port map( A1 => n25279, A2 => n25354, B1 => n25277, B2 => 
                           n19392, ZN => n6791);
   U20065 : OAI22_X1 port map( A1 => n25279, A2 => n25357, B1 => n25277, B2 => 
                           n19391, ZN => n6792);
   U20066 : OAI22_X1 port map( A1 => n25280, A2 => n25360, B1 => n25277, B2 => 
                           n19390, ZN => n6793);
   U20067 : OAI22_X1 port map( A1 => n25280, A2 => n25363, B1 => n25277, B2 => 
                           n19389, ZN => n6794);
   U20068 : OAI22_X1 port map( A1 => n25280, A2 => n25366, B1 => n25277, B2 => 
                           n19388, ZN => n6795);
   U20069 : OAI22_X1 port map( A1 => n25280, A2 => n25369, B1 => n25277, B2 => 
                           n19387, ZN => n6796);
   U20070 : OAI22_X1 port map( A1 => n25280, A2 => n25372, B1 => n25277, B2 => 
                           n19386, ZN => n6797);
   U20071 : OAI22_X1 port map( A1 => n25281, A2 => n25375, B1 => n25277, B2 => 
                           n19385, ZN => n6798);
   U20072 : OAI22_X1 port map( A1 => n25281, A2 => n25378, B1 => n25277, B2 => 
                           n19384, ZN => n6799);
   U20073 : OAI22_X1 port map( A1 => n25281, A2 => n25381, B1 => n25278, B2 => 
                           n19383, ZN => n6800);
   U20074 : OAI22_X1 port map( A1 => n25281, A2 => n25384, B1 => n25278, B2 => 
                           n19382, ZN => n6801);
   U20075 : OAI22_X1 port map( A1 => n25281, A2 => n25387, B1 => n25278, B2 => 
                           n19381, ZN => n6802);
   U20076 : OAI22_X1 port map( A1 => n25282, A2 => n25390, B1 => n25278, B2 => 
                           n19380, ZN => n6803);
   U20077 : OAI22_X1 port map( A1 => n25282, A2 => n25393, B1 => n25278, B2 => 
                           n19379, ZN => n6804);
   U20078 : OAI22_X1 port map( A1 => n25282, A2 => n25396, B1 => n25278, B2 => 
                           n19378, ZN => n6805);
   U20079 : OAI22_X1 port map( A1 => n25282, A2 => n25399, B1 => n25278, B2 => 
                           n19377, ZN => n6806);
   U20080 : OAI22_X1 port map( A1 => n25282, A2 => n25402, B1 => n25278, B2 => 
                           n19376, ZN => n6807);
   U20081 : OAI22_X1 port map( A1 => n25283, A2 => n25405, B1 => n25278, B2 => 
                           n19375, ZN => n6808);
   U20082 : OAI22_X1 port map( A1 => n25283, A2 => n25408, B1 => n25278, B2 => 
                           n19374, ZN => n6809);
   U20083 : OAI22_X1 port map( A1 => n25283, A2 => n25411, B1 => n25278, B2 => 
                           n19373, ZN => n6810);
   U20084 : OAI22_X1 port map( A1 => n25283, A2 => n25414, B1 => n25278, B2 => 
                           n19372, ZN => n6811);
   U20085 : OAI22_X1 port map( A1 => n25537, A2 => n25345, B1 => n25535, B2 => 
                           n19331, ZN => n7044);
   U20086 : OAI22_X1 port map( A1 => n25537, A2 => n25348, B1 => n25535, B2 => 
                           n19330, ZN => n7045);
   U20087 : OAI22_X1 port map( A1 => n25537, A2 => n25351, B1 => n25535, B2 => 
                           n19329, ZN => n7046);
   U20088 : OAI22_X1 port map( A1 => n25537, A2 => n25354, B1 => n25535, B2 => 
                           n19328, ZN => n7047);
   U20089 : OAI22_X1 port map( A1 => n25537, A2 => n25357, B1 => n25535, B2 => 
                           n19327, ZN => n7048);
   U20090 : OAI22_X1 port map( A1 => n25538, A2 => n25360, B1 => n25535, B2 => 
                           n19326, ZN => n7049);
   U20091 : OAI22_X1 port map( A1 => n25538, A2 => n25363, B1 => n25535, B2 => 
                           n19325, ZN => n7050);
   U20092 : OAI22_X1 port map( A1 => n25538, A2 => n25366, B1 => n25535, B2 => 
                           n19324, ZN => n7051);
   U20093 : OAI22_X1 port map( A1 => n25538, A2 => n25369, B1 => n25535, B2 => 
                           n19323, ZN => n7052);
   U20094 : OAI22_X1 port map( A1 => n25538, A2 => n25372, B1 => n25535, B2 => 
                           n19322, ZN => n7053);
   U20095 : OAI22_X1 port map( A1 => n25539, A2 => n25375, B1 => n25535, B2 => 
                           n19321, ZN => n7054);
   U20096 : OAI22_X1 port map( A1 => n25539, A2 => n25378, B1 => n25535, B2 => 
                           n19320, ZN => n7055);
   U20097 : OAI22_X1 port map( A1 => n25539, A2 => n25381, B1 => n25536, B2 => 
                           n19319, ZN => n7056);
   U20098 : OAI22_X1 port map( A1 => n25539, A2 => n25384, B1 => n25536, B2 => 
                           n19318, ZN => n7057);
   U20099 : OAI22_X1 port map( A1 => n25539, A2 => n25387, B1 => n25536, B2 => 
                           n19317, ZN => n7058);
   U20100 : OAI22_X1 port map( A1 => n25540, A2 => n25390, B1 => n25536, B2 => 
                           n19316, ZN => n7059);
   U20101 : OAI22_X1 port map( A1 => n25540, A2 => n25393, B1 => n25536, B2 => 
                           n19315, ZN => n7060);
   U20102 : OAI22_X1 port map( A1 => n25540, A2 => n25396, B1 => n25536, B2 => 
                           n19314, ZN => n7061);
   U20103 : OAI22_X1 port map( A1 => n25540, A2 => n25399, B1 => n25536, B2 => 
                           n19313, ZN => n7062);
   U20104 : OAI22_X1 port map( A1 => n25540, A2 => n25402, B1 => n25536, B2 => 
                           n19312, ZN => n7063);
   U20105 : OAI22_X1 port map( A1 => n25541, A2 => n25405, B1 => n25536, B2 => 
                           n19311, ZN => n7064);
   U20106 : OAI22_X1 port map( A1 => n25541, A2 => n25408, B1 => n25536, B2 => 
                           n19310, ZN => n7065);
   U20107 : OAI22_X1 port map( A1 => n25541, A2 => n25411, B1 => n25536, B2 => 
                           n19309, ZN => n7066);
   U20108 : OAI22_X1 port map( A1 => n25541, A2 => n25414, B1 => n25536, B2 => 
                           n19308, ZN => n7067);
   U20109 : OAI22_X1 port map( A1 => n24994, A2 => n25418, B1 => n24988, B2 => 
                           n21050, ZN => n5724);
   U20110 : OAI22_X1 port map( A1 => n24995, A2 => n25421, B1 => n24989, B2 => 
                           n21049, ZN => n5725);
   U20111 : OAI22_X1 port map( A1 => n24995, A2 => n25424, B1 => n24987, B2 => 
                           n21048, ZN => n5726);
   U20112 : OAI22_X1 port map( A1 => n24995, A2 => n25427, B1 => n24988, B2 => 
                           n21047, ZN => n5727);
   U20113 : OAI22_X1 port map( A1 => n24995, A2 => n25430, B1 => n24989, B2 => 
                           n21046, ZN => n5728);
   U20114 : OAI22_X1 port map( A1 => n24995, A2 => n25433, B1 => n24987, B2 => 
                           n21045, ZN => n5729);
   U20115 : OAI22_X1 port map( A1 => n24996, A2 => n25436, B1 => n24988, B2 => 
                           n21044, ZN => n5730);
   U20116 : OAI22_X1 port map( A1 => n24996, A2 => n25439, B1 => n24989, B2 => 
                           n21043, ZN => n5731);
   U20117 : OAI22_X1 port map( A1 => n24996, A2 => n25442, B1 => n24987, B2 => 
                           n21042, ZN => n5732);
   U20118 : OAI22_X1 port map( A1 => n24996, A2 => n25445, B1 => n24988, B2 => 
                           n21041, ZN => n5733);
   U20119 : OAI22_X1 port map( A1 => n24996, A2 => n25448, B1 => n24989, B2 => 
                           n21040, ZN => n5734);
   U20120 : OAI22_X1 port map( A1 => n24997, A2 => n25451, B1 => n24987, B2 => 
                           n21039, ZN => n5735);
   U20121 : OAI22_X1 port map( A1 => n24997, A2 => n25454, B1 => n21285, B2 => 
                           n21038, ZN => n5736);
   U20122 : OAI22_X1 port map( A1 => n24997, A2 => n25457, B1 => n24987, B2 => 
                           n21037, ZN => n5737);
   U20123 : OAI22_X1 port map( A1 => n24997, A2 => n25460, B1 => n21285, B2 => 
                           n21036, ZN => n5738);
   U20124 : OAI22_X1 port map( A1 => n24997, A2 => n25463, B1 => n24987, B2 => 
                           n21035, ZN => n5739);
   U20125 : OAI22_X1 port map( A1 => n24998, A2 => n25466, B1 => n21285, B2 => 
                           n21034, ZN => n5740);
   U20126 : OAI22_X1 port map( A1 => n24998, A2 => n25469, B1 => n24987, B2 => 
                           n21033, ZN => n5741);
   U20127 : OAI22_X1 port map( A1 => n24998, A2 => n25472, B1 => n24988, B2 => 
                           n21032, ZN => n5742);
   U20128 : OAI22_X1 port map( A1 => n24998, A2 => n25475, B1 => n24989, B2 => 
                           n21031, ZN => n5743);
   U20129 : OAI22_X1 port map( A1 => n24998, A2 => n25478, B1 => n24987, B2 => 
                           n21030, ZN => n5744);
   U20130 : OAI22_X1 port map( A1 => n24999, A2 => n25481, B1 => n24987, B2 => 
                           n21029, ZN => n5745);
   U20131 : OAI22_X1 port map( A1 => n24999, A2 => n25484, B1 => n24988, B2 => 
                           n21028, ZN => n5746);
   U20132 : OAI22_X1 port map( A1 => n24999, A2 => n25487, B1 => n24989, B2 => 
                           n21027, ZN => n5747);
   U20133 : OAI22_X1 port map( A1 => n24999, A2 => n25490, B1 => n24987, B2 => 
                           n21026, ZN => n5748);
   U20134 : OAI22_X1 port map( A1 => n24999, A2 => n25493, B1 => n24987, B2 => 
                           n21025, ZN => n5749);
   U20135 : OAI22_X1 port map( A1 => n25000, A2 => n25496, B1 => n21285, B2 => 
                           n21024, ZN => n5750);
   U20136 : OAI22_X1 port map( A1 => n25000, A2 => n25499, B1 => n24987, B2 => 
                           n21023, ZN => n5751);
   U20137 : OAI22_X1 port map( A1 => n25000, A2 => n25502, B1 => n21285, B2 => 
                           n21022, ZN => n5752);
   U20138 : OAI22_X1 port map( A1 => n25000, A2 => n25505, B1 => n24987, B2 => 
                           n21021, ZN => n5753);
   U20139 : OAI22_X1 port map( A1 => n25000, A2 => n25508, B1 => n21285, B2 => 
                           n21020, ZN => n5754);
   U20140 : OAI22_X1 port map( A1 => n25001, A2 => n25511, B1 => n24987, B2 => 
                           n21019, ZN => n5755);
   U20141 : OAI22_X1 port map( A1 => n25001, A2 => n25514, B1 => n21285, B2 => 
                           n21018, ZN => n5756);
   U20142 : OAI22_X1 port map( A1 => n25001, A2 => n25517, B1 => n24987, B2 => 
                           n21017, ZN => n5757);
   U20143 : OAI22_X1 port map( A1 => n25001, A2 => n25520, B1 => n21285, B2 => 
                           n21016, ZN => n5758);
   U20144 : OAI22_X1 port map( A1 => n25001, A2 => n25523, B1 => n24987, B2 => 
                           n21015, ZN => n5759);
   U20145 : OAI22_X1 port map( A1 => n25232, A2 => n25417, B1 => n25226, B2 => 
                           n21014, ZN => n6620);
   U20146 : OAI22_X1 port map( A1 => n25233, A2 => n25420, B1 => n25227, B2 => 
                           n21013, ZN => n6621);
   U20147 : OAI22_X1 port map( A1 => n25233, A2 => n25423, B1 => n25225, B2 => 
                           n21012, ZN => n6622);
   U20148 : OAI22_X1 port map( A1 => n25233, A2 => n25426, B1 => n25226, B2 => 
                           n21011, ZN => n6623);
   U20149 : OAI22_X1 port map( A1 => n25233, A2 => n25429, B1 => n25227, B2 => 
                           n21010, ZN => n6624);
   U20150 : OAI22_X1 port map( A1 => n25233, A2 => n25432, B1 => n25225, B2 => 
                           n21009, ZN => n6625);
   U20151 : OAI22_X1 port map( A1 => n25234, A2 => n25435, B1 => n25226, B2 => 
                           n21008, ZN => n6626);
   U20152 : OAI22_X1 port map( A1 => n25234, A2 => n25438, B1 => n25227, B2 => 
                           n21007, ZN => n6627);
   U20153 : OAI22_X1 port map( A1 => n25234, A2 => n25441, B1 => n25225, B2 => 
                           n21006, ZN => n6628);
   U20154 : OAI22_X1 port map( A1 => n25234, A2 => n25444, B1 => n25226, B2 => 
                           n21005, ZN => n6629);
   U20155 : OAI22_X1 port map( A1 => n25234, A2 => n25447, B1 => n25227, B2 => 
                           n21004, ZN => n6630);
   U20156 : OAI22_X1 port map( A1 => n25235, A2 => n25450, B1 => n25225, B2 => 
                           n21003, ZN => n6631);
   U20157 : OAI22_X1 port map( A1 => n25235, A2 => n25453, B1 => n21267, B2 => 
                           n21002, ZN => n6632);
   U20158 : OAI22_X1 port map( A1 => n25235, A2 => n25456, B1 => n25225, B2 => 
                           n21001, ZN => n6633);
   U20159 : OAI22_X1 port map( A1 => n25235, A2 => n25459, B1 => n21267, B2 => 
                           n21000, ZN => n6634);
   U20160 : OAI22_X1 port map( A1 => n25235, A2 => n25462, B1 => n25225, B2 => 
                           n20999, ZN => n6635);
   U20161 : OAI22_X1 port map( A1 => n25236, A2 => n25465, B1 => n21267, B2 => 
                           n20998, ZN => n6636);
   U20162 : OAI22_X1 port map( A1 => n25236, A2 => n25468, B1 => n25225, B2 => 
                           n20997, ZN => n6637);
   U20163 : OAI22_X1 port map( A1 => n25236, A2 => n25471, B1 => n25226, B2 => 
                           n20996, ZN => n6638);
   U20164 : OAI22_X1 port map( A1 => n25236, A2 => n25474, B1 => n25227, B2 => 
                           n20995, ZN => n6639);
   U20165 : OAI22_X1 port map( A1 => n25236, A2 => n25477, B1 => n25225, B2 => 
                           n20994, ZN => n6640);
   U20166 : OAI22_X1 port map( A1 => n25237, A2 => n25480, B1 => n25225, B2 => 
                           n20993, ZN => n6641);
   U20167 : OAI22_X1 port map( A1 => n25237, A2 => n25483, B1 => n25226, B2 => 
                           n20992, ZN => n6642);
   U20168 : OAI22_X1 port map( A1 => n25237, A2 => n25486, B1 => n25227, B2 => 
                           n20991, ZN => n6643);
   U20169 : OAI22_X1 port map( A1 => n25237, A2 => n25489, B1 => n25225, B2 => 
                           n20990, ZN => n6644);
   U20170 : OAI22_X1 port map( A1 => n25237, A2 => n25492, B1 => n25225, B2 => 
                           n20989, ZN => n6645);
   U20171 : OAI22_X1 port map( A1 => n25238, A2 => n25495, B1 => n21267, B2 => 
                           n20988, ZN => n6646);
   U20172 : OAI22_X1 port map( A1 => n25238, A2 => n25498, B1 => n25225, B2 => 
                           n20987, ZN => n6647);
   U20173 : OAI22_X1 port map( A1 => n25238, A2 => n25501, B1 => n21267, B2 => 
                           n20986, ZN => n6648);
   U20174 : OAI22_X1 port map( A1 => n25238, A2 => n25504, B1 => n25225, B2 => 
                           n20985, ZN => n6649);
   U20175 : OAI22_X1 port map( A1 => n25238, A2 => n25507, B1 => n21267, B2 => 
                           n20984, ZN => n6650);
   U20176 : OAI22_X1 port map( A1 => n25239, A2 => n25510, B1 => n25225, B2 => 
                           n20983, ZN => n6651);
   U20177 : OAI22_X1 port map( A1 => n25239, A2 => n25513, B1 => n21267, B2 => 
                           n20982, ZN => n6652);
   U20178 : OAI22_X1 port map( A1 => n25239, A2 => n25516, B1 => n25225, B2 => 
                           n20981, ZN => n6653);
   U20179 : OAI22_X1 port map( A1 => n25239, A2 => n25519, B1 => n21267, B2 => 
                           n20980, ZN => n6654);
   U20180 : OAI22_X1 port map( A1 => n25239, A2 => n25522, B1 => n25225, B2 => 
                           n20979, ZN => n6655);
   U20181 : OAI22_X1 port map( A1 => n25215, A2 => n25417, B1 => n25209, B2 => 
                           n20978, ZN => n6556);
   U20182 : OAI22_X1 port map( A1 => n25216, A2 => n25420, B1 => n25210, B2 => 
                           n20977, ZN => n6557);
   U20183 : OAI22_X1 port map( A1 => n25216, A2 => n25423, B1 => n25208, B2 => 
                           n20976, ZN => n6558);
   U20184 : OAI22_X1 port map( A1 => n25216, A2 => n25426, B1 => n25209, B2 => 
                           n20975, ZN => n6559);
   U20185 : OAI22_X1 port map( A1 => n25216, A2 => n25429, B1 => n25210, B2 => 
                           n20974, ZN => n6560);
   U20186 : OAI22_X1 port map( A1 => n25216, A2 => n25432, B1 => n25208, B2 => 
                           n20973, ZN => n6561);
   U20187 : OAI22_X1 port map( A1 => n25217, A2 => n25435, B1 => n25209, B2 => 
                           n20972, ZN => n6562);
   U20188 : OAI22_X1 port map( A1 => n25217, A2 => n25438, B1 => n25210, B2 => 
                           n20971, ZN => n6563);
   U20189 : OAI22_X1 port map( A1 => n25217, A2 => n25441, B1 => n25208, B2 => 
                           n20970, ZN => n6564);
   U20190 : OAI22_X1 port map( A1 => n25217, A2 => n25444, B1 => n25209, B2 => 
                           n20969, ZN => n6565);
   U20191 : OAI22_X1 port map( A1 => n25217, A2 => n25447, B1 => n25210, B2 => 
                           n20968, ZN => n6566);
   U20192 : OAI22_X1 port map( A1 => n25218, A2 => n25450, B1 => n25208, B2 => 
                           n20967, ZN => n6567);
   U20193 : OAI22_X1 port map( A1 => n25218, A2 => n25453, B1 => n21270, B2 => 
                           n20966, ZN => n6568);
   U20194 : OAI22_X1 port map( A1 => n25218, A2 => n25456, B1 => n25208, B2 => 
                           n20965, ZN => n6569);
   U20195 : OAI22_X1 port map( A1 => n25218, A2 => n25459, B1 => n21270, B2 => 
                           n20964, ZN => n6570);
   U20196 : OAI22_X1 port map( A1 => n25218, A2 => n25462, B1 => n25208, B2 => 
                           n20963, ZN => n6571);
   U20197 : OAI22_X1 port map( A1 => n25219, A2 => n25465, B1 => n21270, B2 => 
                           n20962, ZN => n6572);
   U20198 : OAI22_X1 port map( A1 => n25219, A2 => n25468, B1 => n25208, B2 => 
                           n20961, ZN => n6573);
   U20199 : OAI22_X1 port map( A1 => n25219, A2 => n25471, B1 => n25209, B2 => 
                           n20960, ZN => n6574);
   U20200 : OAI22_X1 port map( A1 => n25219, A2 => n25474, B1 => n25210, B2 => 
                           n20959, ZN => n6575);
   U20201 : OAI22_X1 port map( A1 => n25219, A2 => n25477, B1 => n25208, B2 => 
                           n20958, ZN => n6576);
   U20202 : OAI22_X1 port map( A1 => n25220, A2 => n25480, B1 => n25208, B2 => 
                           n20957, ZN => n6577);
   U20203 : OAI22_X1 port map( A1 => n25220, A2 => n25483, B1 => n25209, B2 => 
                           n20956, ZN => n6578);
   U20204 : OAI22_X1 port map( A1 => n25220, A2 => n25486, B1 => n25210, B2 => 
                           n20955, ZN => n6579);
   U20205 : OAI22_X1 port map( A1 => n25220, A2 => n25489, B1 => n25208, B2 => 
                           n20954, ZN => n6580);
   U20206 : OAI22_X1 port map( A1 => n25220, A2 => n25492, B1 => n25208, B2 => 
                           n20953, ZN => n6581);
   U20207 : OAI22_X1 port map( A1 => n25221, A2 => n25495, B1 => n21270, B2 => 
                           n20952, ZN => n6582);
   U20208 : OAI22_X1 port map( A1 => n25221, A2 => n25498, B1 => n25208, B2 => 
                           n20951, ZN => n6583);
   U20209 : OAI22_X1 port map( A1 => n25221, A2 => n25501, B1 => n21270, B2 => 
                           n20950, ZN => n6584);
   U20210 : OAI22_X1 port map( A1 => n25221, A2 => n25504, B1 => n25208, B2 => 
                           n20949, ZN => n6585);
   U20211 : OAI22_X1 port map( A1 => n25221, A2 => n25507, B1 => n21270, B2 => 
                           n20948, ZN => n6586);
   U20212 : OAI22_X1 port map( A1 => n25222, A2 => n25510, B1 => n25208, B2 => 
                           n20947, ZN => n6587);
   U20213 : OAI22_X1 port map( A1 => n25222, A2 => n25513, B1 => n21270, B2 => 
                           n20946, ZN => n6588);
   U20214 : OAI22_X1 port map( A1 => n25222, A2 => n25516, B1 => n25208, B2 => 
                           n20945, ZN => n6589);
   U20215 : OAI22_X1 port map( A1 => n25222, A2 => n25519, B1 => n21270, B2 => 
                           n20944, ZN => n6590);
   U20216 : OAI22_X1 port map( A1 => n25222, A2 => n25522, B1 => n25208, B2 => 
                           n20943, ZN => n6591);
   U20217 : OAI22_X1 port map( A1 => n25147, A2 => n25418, B1 => n25141, B2 => 
                           n20942, ZN => n6300);
   U20218 : OAI22_X1 port map( A1 => n25148, A2 => n25421, B1 => n25142, B2 => 
                           n20941, ZN => n6301);
   U20219 : OAI22_X1 port map( A1 => n25148, A2 => n25424, B1 => n25140, B2 => 
                           n20940, ZN => n6302);
   U20220 : OAI22_X1 port map( A1 => n25148, A2 => n25427, B1 => n25141, B2 => 
                           n20939, ZN => n6303);
   U20221 : OAI22_X1 port map( A1 => n25148, A2 => n25430, B1 => n25142, B2 => 
                           n20938, ZN => n6304);
   U20222 : OAI22_X1 port map( A1 => n25148, A2 => n25433, B1 => n25140, B2 => 
                           n20937, ZN => n6305);
   U20223 : OAI22_X1 port map( A1 => n25149, A2 => n25436, B1 => n25141, B2 => 
                           n20936, ZN => n6306);
   U20224 : OAI22_X1 port map( A1 => n25149, A2 => n25439, B1 => n25142, B2 => 
                           n20935, ZN => n6307);
   U20225 : OAI22_X1 port map( A1 => n25149, A2 => n25442, B1 => n25140, B2 => 
                           n20934, ZN => n6308);
   U20226 : OAI22_X1 port map( A1 => n25149, A2 => n25445, B1 => n25141, B2 => 
                           n20933, ZN => n6309);
   U20227 : OAI22_X1 port map( A1 => n25149, A2 => n25448, B1 => n25142, B2 => 
                           n20932, ZN => n6310);
   U20228 : OAI22_X1 port map( A1 => n25150, A2 => n25451, B1 => n25140, B2 => 
                           n20931, ZN => n6311);
   U20229 : OAI22_X1 port map( A1 => n25150, A2 => n25454, B1 => n21275, B2 => 
                           n20930, ZN => n6312);
   U20230 : OAI22_X1 port map( A1 => n25150, A2 => n25457, B1 => n25140, B2 => 
                           n20929, ZN => n6313);
   U20231 : OAI22_X1 port map( A1 => n25150, A2 => n25460, B1 => n21275, B2 => 
                           n20928, ZN => n6314);
   U20232 : OAI22_X1 port map( A1 => n25150, A2 => n25463, B1 => n25140, B2 => 
                           n20927, ZN => n6315);
   U20233 : OAI22_X1 port map( A1 => n25151, A2 => n25466, B1 => n21275, B2 => 
                           n20926, ZN => n6316);
   U20234 : OAI22_X1 port map( A1 => n25151, A2 => n25469, B1 => n25140, B2 => 
                           n20925, ZN => n6317);
   U20235 : OAI22_X1 port map( A1 => n25151, A2 => n25472, B1 => n25141, B2 => 
                           n20924, ZN => n6318);
   U20236 : OAI22_X1 port map( A1 => n25151, A2 => n25475, B1 => n25142, B2 => 
                           n20923, ZN => n6319);
   U20237 : OAI22_X1 port map( A1 => n25151, A2 => n25478, B1 => n25140, B2 => 
                           n20922, ZN => n6320);
   U20238 : OAI22_X1 port map( A1 => n25152, A2 => n25481, B1 => n25140, B2 => 
                           n20921, ZN => n6321);
   U20239 : OAI22_X1 port map( A1 => n25152, A2 => n25484, B1 => n25141, B2 => 
                           n20920, ZN => n6322);
   U20240 : OAI22_X1 port map( A1 => n25152, A2 => n25487, B1 => n25142, B2 => 
                           n20919, ZN => n6323);
   U20241 : OAI22_X1 port map( A1 => n25152, A2 => n25490, B1 => n25140, B2 => 
                           n20918, ZN => n6324);
   U20242 : OAI22_X1 port map( A1 => n25152, A2 => n25493, B1 => n25140, B2 => 
                           n20917, ZN => n6325);
   U20243 : OAI22_X1 port map( A1 => n25153, A2 => n25496, B1 => n21275, B2 => 
                           n20916, ZN => n6326);
   U20244 : OAI22_X1 port map( A1 => n25153, A2 => n25499, B1 => n25140, B2 => 
                           n20915, ZN => n6327);
   U20245 : OAI22_X1 port map( A1 => n25153, A2 => n25502, B1 => n21275, B2 => 
                           n20914, ZN => n6328);
   U20246 : OAI22_X1 port map( A1 => n25153, A2 => n25505, B1 => n25140, B2 => 
                           n20913, ZN => n6329);
   U20247 : OAI22_X1 port map( A1 => n25153, A2 => n25508, B1 => n21275, B2 => 
                           n20912, ZN => n6330);
   U20248 : OAI22_X1 port map( A1 => n25154, A2 => n25511, B1 => n25140, B2 => 
                           n20911, ZN => n6331);
   U20249 : OAI22_X1 port map( A1 => n25154, A2 => n25514, B1 => n21275, B2 => 
                           n20910, ZN => n6332);
   U20250 : OAI22_X1 port map( A1 => n25154, A2 => n25517, B1 => n25140, B2 => 
                           n20909, ZN => n6333);
   U20251 : OAI22_X1 port map( A1 => n25154, A2 => n25520, B1 => n21275, B2 => 
                           n20908, ZN => n6334);
   U20252 : OAI22_X1 port map( A1 => n25154, A2 => n25523, B1 => n25140, B2 => 
                           n20907, ZN => n6335);
   U20253 : OAI22_X1 port map( A1 => n25249, A2 => n25417, B1 => n25243, B2 => 
                           n20726, ZN => n6684);
   U20254 : OAI22_X1 port map( A1 => n25250, A2 => n25420, B1 => n25244, B2 => 
                           n20725, ZN => n6685);
   U20255 : OAI22_X1 port map( A1 => n25250, A2 => n25423, B1 => n25242, B2 => 
                           n20724, ZN => n6686);
   U20256 : OAI22_X1 port map( A1 => n25250, A2 => n25426, B1 => n25243, B2 => 
                           n20723, ZN => n6687);
   U20257 : OAI22_X1 port map( A1 => n25250, A2 => n25429, B1 => n25244, B2 => 
                           n20722, ZN => n6688);
   U20258 : OAI22_X1 port map( A1 => n25250, A2 => n25432, B1 => n25242, B2 => 
                           n20721, ZN => n6689);
   U20259 : OAI22_X1 port map( A1 => n25251, A2 => n25435, B1 => n25243, B2 => 
                           n20720, ZN => n6690);
   U20260 : OAI22_X1 port map( A1 => n25251, A2 => n25438, B1 => n25244, B2 => 
                           n20719, ZN => n6691);
   U20261 : OAI22_X1 port map( A1 => n25251, A2 => n25441, B1 => n25242, B2 => 
                           n20718, ZN => n6692);
   U20262 : OAI22_X1 port map( A1 => n25251, A2 => n25444, B1 => n25243, B2 => 
                           n20717, ZN => n6693);
   U20263 : OAI22_X1 port map( A1 => n25251, A2 => n25447, B1 => n25244, B2 => 
                           n20716, ZN => n6694);
   U20264 : OAI22_X1 port map( A1 => n25252, A2 => n25450, B1 => n25242, B2 => 
                           n20715, ZN => n6695);
   U20265 : OAI22_X1 port map( A1 => n25252, A2 => n25453, B1 => n21265, B2 => 
                           n20714, ZN => n6696);
   U20266 : OAI22_X1 port map( A1 => n25252, A2 => n25456, B1 => n25242, B2 => 
                           n20713, ZN => n6697);
   U20267 : OAI22_X1 port map( A1 => n25252, A2 => n25459, B1 => n21265, B2 => 
                           n20712, ZN => n6698);
   U20268 : OAI22_X1 port map( A1 => n25252, A2 => n25462, B1 => n25242, B2 => 
                           n20711, ZN => n6699);
   U20269 : OAI22_X1 port map( A1 => n25253, A2 => n25465, B1 => n21265, B2 => 
                           n20710, ZN => n6700);
   U20270 : OAI22_X1 port map( A1 => n25253, A2 => n25468, B1 => n25242, B2 => 
                           n20709, ZN => n6701);
   U20271 : OAI22_X1 port map( A1 => n25253, A2 => n25471, B1 => n25243, B2 => 
                           n20708, ZN => n6702);
   U20272 : OAI22_X1 port map( A1 => n25253, A2 => n25474, B1 => n25244, B2 => 
                           n20707, ZN => n6703);
   U20273 : OAI22_X1 port map( A1 => n25253, A2 => n25477, B1 => n25242, B2 => 
                           n20706, ZN => n6704);
   U20274 : OAI22_X1 port map( A1 => n25254, A2 => n25480, B1 => n25242, B2 => 
                           n20705, ZN => n6705);
   U20275 : OAI22_X1 port map( A1 => n25254, A2 => n25483, B1 => n25243, B2 => 
                           n20704, ZN => n6706);
   U20276 : OAI22_X1 port map( A1 => n25254, A2 => n25486, B1 => n25244, B2 => 
                           n20703, ZN => n6707);
   U20277 : OAI22_X1 port map( A1 => n25254, A2 => n25489, B1 => n25242, B2 => 
                           n20702, ZN => n6708);
   U20278 : OAI22_X1 port map( A1 => n25254, A2 => n25492, B1 => n25242, B2 => 
                           n20701, ZN => n6709);
   U20279 : OAI22_X1 port map( A1 => n25255, A2 => n25495, B1 => n21265, B2 => 
                           n20700, ZN => n6710);
   U20280 : OAI22_X1 port map( A1 => n25255, A2 => n25498, B1 => n25242, B2 => 
                           n20699, ZN => n6711);
   U20281 : OAI22_X1 port map( A1 => n25255, A2 => n25501, B1 => n21265, B2 => 
                           n20698, ZN => n6712);
   U20282 : OAI22_X1 port map( A1 => n25255, A2 => n25504, B1 => n25242, B2 => 
                           n20697, ZN => n6713);
   U20283 : OAI22_X1 port map( A1 => n25255, A2 => n25507, B1 => n21265, B2 => 
                           n20696, ZN => n6714);
   U20284 : OAI22_X1 port map( A1 => n25256, A2 => n25510, B1 => n25242, B2 => 
                           n20695, ZN => n6715);
   U20285 : OAI22_X1 port map( A1 => n25256, A2 => n25513, B1 => n21265, B2 => 
                           n20694, ZN => n6716);
   U20286 : OAI22_X1 port map( A1 => n25256, A2 => n25516, B1 => n25242, B2 => 
                           n20693, ZN => n6717);
   U20287 : OAI22_X1 port map( A1 => n25256, A2 => n25519, B1 => n21265, B2 => 
                           n20692, ZN => n6718);
   U20288 : OAI22_X1 port map( A1 => n25256, A2 => n25522, B1 => n25242, B2 => 
                           n20691, ZN => n6719);
   U20289 : OAI22_X1 port map( A1 => n25079, A2 => n25418, B1 => n25073, B2 => 
                           n20690, ZN => n6044);
   U20290 : OAI22_X1 port map( A1 => n25080, A2 => n25421, B1 => n25074, B2 => 
                           n20689, ZN => n6045);
   U20291 : OAI22_X1 port map( A1 => n25080, A2 => n25424, B1 => n25072, B2 => 
                           n20688, ZN => n6046);
   U20292 : OAI22_X1 port map( A1 => n25080, A2 => n25427, B1 => n25073, B2 => 
                           n20687, ZN => n6047);
   U20293 : OAI22_X1 port map( A1 => n25080, A2 => n25430, B1 => n25074, B2 => 
                           n20686, ZN => n6048);
   U20294 : OAI22_X1 port map( A1 => n25080, A2 => n25433, B1 => n25072, B2 => 
                           n20685, ZN => n6049);
   U20295 : OAI22_X1 port map( A1 => n25081, A2 => n25436, B1 => n25073, B2 => 
                           n20684, ZN => n6050);
   U20296 : OAI22_X1 port map( A1 => n25081, A2 => n25439, B1 => n25074, B2 => 
                           n20683, ZN => n6051);
   U20297 : OAI22_X1 port map( A1 => n25081, A2 => n25442, B1 => n25072, B2 => 
                           n20682, ZN => n6052);
   U20298 : OAI22_X1 port map( A1 => n25081, A2 => n25445, B1 => n25073, B2 => 
                           n20681, ZN => n6053);
   U20299 : OAI22_X1 port map( A1 => n25081, A2 => n25448, B1 => n25074, B2 => 
                           n20680, ZN => n6054);
   U20300 : OAI22_X1 port map( A1 => n25082, A2 => n25451, B1 => n25072, B2 => 
                           n20679, ZN => n6055);
   U20301 : OAI22_X1 port map( A1 => n25082, A2 => n25454, B1 => n21279, B2 => 
                           n20678, ZN => n6056);
   U20302 : OAI22_X1 port map( A1 => n25082, A2 => n25457, B1 => n25072, B2 => 
                           n20677, ZN => n6057);
   U20303 : OAI22_X1 port map( A1 => n25082, A2 => n25460, B1 => n21279, B2 => 
                           n20676, ZN => n6058);
   U20304 : OAI22_X1 port map( A1 => n25082, A2 => n25463, B1 => n25072, B2 => 
                           n20675, ZN => n6059);
   U20305 : OAI22_X1 port map( A1 => n25083, A2 => n25466, B1 => n21279, B2 => 
                           n20674, ZN => n6060);
   U20306 : OAI22_X1 port map( A1 => n25083, A2 => n25469, B1 => n25072, B2 => 
                           n20673, ZN => n6061);
   U20307 : OAI22_X1 port map( A1 => n25083, A2 => n25472, B1 => n25073, B2 => 
                           n20672, ZN => n6062);
   U20308 : OAI22_X1 port map( A1 => n25083, A2 => n25475, B1 => n25074, B2 => 
                           n20671, ZN => n6063);
   U20309 : OAI22_X1 port map( A1 => n25083, A2 => n25478, B1 => n25072, B2 => 
                           n20670, ZN => n6064);
   U20310 : OAI22_X1 port map( A1 => n25084, A2 => n25481, B1 => n25072, B2 => 
                           n20669, ZN => n6065);
   U20311 : OAI22_X1 port map( A1 => n25084, A2 => n25484, B1 => n25073, B2 => 
                           n20668, ZN => n6066);
   U20312 : OAI22_X1 port map( A1 => n25084, A2 => n25487, B1 => n25074, B2 => 
                           n20667, ZN => n6067);
   U20313 : OAI22_X1 port map( A1 => n25084, A2 => n25490, B1 => n25072, B2 => 
                           n20666, ZN => n6068);
   U20314 : OAI22_X1 port map( A1 => n25084, A2 => n25493, B1 => n25072, B2 => 
                           n20665, ZN => n6069);
   U20315 : OAI22_X1 port map( A1 => n25085, A2 => n25496, B1 => n21279, B2 => 
                           n20664, ZN => n6070);
   U20316 : OAI22_X1 port map( A1 => n25085, A2 => n25499, B1 => n25072, B2 => 
                           n20663, ZN => n6071);
   U20317 : OAI22_X1 port map( A1 => n25085, A2 => n25502, B1 => n21279, B2 => 
                           n20662, ZN => n6072);
   U20318 : OAI22_X1 port map( A1 => n25085, A2 => n25505, B1 => n25072, B2 => 
                           n20661, ZN => n6073);
   U20319 : OAI22_X1 port map( A1 => n25085, A2 => n25508, B1 => n21279, B2 => 
                           n20660, ZN => n6074);
   U20320 : OAI22_X1 port map( A1 => n25086, A2 => n25511, B1 => n25072, B2 => 
                           n20659, ZN => n6075);
   U20321 : OAI22_X1 port map( A1 => n25086, A2 => n25514, B1 => n21279, B2 => 
                           n20658, ZN => n6076);
   U20322 : OAI22_X1 port map( A1 => n25086, A2 => n25517, B1 => n25072, B2 => 
                           n20657, ZN => n6077);
   U20323 : OAI22_X1 port map( A1 => n25086, A2 => n25520, B1 => n21279, B2 => 
                           n20656, ZN => n6078);
   U20324 : OAI22_X1 port map( A1 => n25086, A2 => n25523, B1 => n25072, B2 => 
                           n20655, ZN => n6079);
   U20325 : OAI22_X1 port map( A1 => n25011, A2 => n25418, B1 => n25005, B2 => 
                           n20654, ZN => n5788);
   U20326 : OAI22_X1 port map( A1 => n25012, A2 => n25421, B1 => n25006, B2 => 
                           n20653, ZN => n5789);
   U20327 : OAI22_X1 port map( A1 => n25012, A2 => n25424, B1 => n25004, B2 => 
                           n20652, ZN => n5790);
   U20328 : OAI22_X1 port map( A1 => n25012, A2 => n25427, B1 => n25005, B2 => 
                           n20651, ZN => n5791);
   U20329 : OAI22_X1 port map( A1 => n25012, A2 => n25430, B1 => n25006, B2 => 
                           n20650, ZN => n5792);
   U20330 : OAI22_X1 port map( A1 => n25012, A2 => n25433, B1 => n25004, B2 => 
                           n20649, ZN => n5793);
   U20331 : OAI22_X1 port map( A1 => n25013, A2 => n25436, B1 => n25005, B2 => 
                           n20648, ZN => n5794);
   U20332 : OAI22_X1 port map( A1 => n25013, A2 => n25439, B1 => n25006, B2 => 
                           n20647, ZN => n5795);
   U20333 : OAI22_X1 port map( A1 => n25013, A2 => n25442, B1 => n25004, B2 => 
                           n20646, ZN => n5796);
   U20334 : OAI22_X1 port map( A1 => n25013, A2 => n25445, B1 => n25005, B2 => 
                           n20645, ZN => n5797);
   U20335 : OAI22_X1 port map( A1 => n25013, A2 => n25448, B1 => n25006, B2 => 
                           n20644, ZN => n5798);
   U20336 : OAI22_X1 port map( A1 => n25014, A2 => n25451, B1 => n25004, B2 => 
                           n20643, ZN => n5799);
   U20337 : OAI22_X1 port map( A1 => n25014, A2 => n25454, B1 => n21284, B2 => 
                           n20642, ZN => n5800);
   U20338 : OAI22_X1 port map( A1 => n25014, A2 => n25457, B1 => n25004, B2 => 
                           n20641, ZN => n5801);
   U20339 : OAI22_X1 port map( A1 => n25014, A2 => n25460, B1 => n21284, B2 => 
                           n20640, ZN => n5802);
   U20340 : OAI22_X1 port map( A1 => n25014, A2 => n25463, B1 => n25004, B2 => 
                           n20639, ZN => n5803);
   U20341 : OAI22_X1 port map( A1 => n25015, A2 => n25466, B1 => n21284, B2 => 
                           n20638, ZN => n5804);
   U20342 : OAI22_X1 port map( A1 => n25015, A2 => n25469, B1 => n25004, B2 => 
                           n20637, ZN => n5805);
   U20343 : OAI22_X1 port map( A1 => n25015, A2 => n25472, B1 => n25005, B2 => 
                           n20636, ZN => n5806);
   U20344 : OAI22_X1 port map( A1 => n25015, A2 => n25475, B1 => n25006, B2 => 
                           n20635, ZN => n5807);
   U20345 : OAI22_X1 port map( A1 => n25015, A2 => n25478, B1 => n25004, B2 => 
                           n20634, ZN => n5808);
   U20346 : OAI22_X1 port map( A1 => n25016, A2 => n25481, B1 => n25004, B2 => 
                           n20633, ZN => n5809);
   U20347 : OAI22_X1 port map( A1 => n25016, A2 => n25484, B1 => n25005, B2 => 
                           n20632, ZN => n5810);
   U20348 : OAI22_X1 port map( A1 => n25016, A2 => n25487, B1 => n25006, B2 => 
                           n20631, ZN => n5811);
   U20349 : OAI22_X1 port map( A1 => n25016, A2 => n25490, B1 => n25004, B2 => 
                           n20630, ZN => n5812);
   U20350 : OAI22_X1 port map( A1 => n25016, A2 => n25493, B1 => n25004, B2 => 
                           n20629, ZN => n5813);
   U20351 : OAI22_X1 port map( A1 => n25017, A2 => n25496, B1 => n21284, B2 => 
                           n20628, ZN => n5814);
   U20352 : OAI22_X1 port map( A1 => n25017, A2 => n25499, B1 => n25004, B2 => 
                           n20627, ZN => n5815);
   U20353 : OAI22_X1 port map( A1 => n25017, A2 => n25502, B1 => n21284, B2 => 
                           n20626, ZN => n5816);
   U20354 : OAI22_X1 port map( A1 => n25017, A2 => n25505, B1 => n25004, B2 => 
                           n20625, ZN => n5817);
   U20355 : OAI22_X1 port map( A1 => n25017, A2 => n25508, B1 => n21284, B2 => 
                           n20624, ZN => n5818);
   U20356 : OAI22_X1 port map( A1 => n25018, A2 => n25511, B1 => n25004, B2 => 
                           n20623, ZN => n5819);
   U20357 : OAI22_X1 port map( A1 => n25018, A2 => n25514, B1 => n21284, B2 => 
                           n20622, ZN => n5820);
   U20358 : OAI22_X1 port map( A1 => n25018, A2 => n25517, B1 => n25004, B2 => 
                           n20621, ZN => n5821);
   U20359 : OAI22_X1 port map( A1 => n25018, A2 => n25520, B1 => n21284, B2 => 
                           n20620, ZN => n5822);
   U20360 : OAI22_X1 port map( A1 => n25018, A2 => n25523, B1 => n25004, B2 => 
                           n20619, ZN => n5823);
   U20361 : OAI22_X1 port map( A1 => n24909, A2 => n25419, B1 => n24903, B2 => 
                           n20618, ZN => n5404);
   U20362 : OAI22_X1 port map( A1 => n24910, A2 => n25422, B1 => n24904, B2 => 
                           n20617, ZN => n5405);
   U20363 : OAI22_X1 port map( A1 => n24910, A2 => n25425, B1 => n24902, B2 => 
                           n20616, ZN => n5406);
   U20364 : OAI22_X1 port map( A1 => n24910, A2 => n25428, B1 => n24903, B2 => 
                           n20615, ZN => n5407);
   U20365 : OAI22_X1 port map( A1 => n24910, A2 => n25431, B1 => n24904, B2 => 
                           n20614, ZN => n5408);
   U20366 : OAI22_X1 port map( A1 => n24910, A2 => n25434, B1 => n24902, B2 => 
                           n20613, ZN => n5409);
   U20367 : OAI22_X1 port map( A1 => n24911, A2 => n25437, B1 => n24903, B2 => 
                           n20612, ZN => n5410);
   U20368 : OAI22_X1 port map( A1 => n24911, A2 => n25440, B1 => n24904, B2 => 
                           n20611, ZN => n5411);
   U20369 : OAI22_X1 port map( A1 => n24911, A2 => n25443, B1 => n24902, B2 => 
                           n20610, ZN => n5412);
   U20370 : OAI22_X1 port map( A1 => n24911, A2 => n25446, B1 => n24903, B2 => 
                           n20609, ZN => n5413);
   U20371 : OAI22_X1 port map( A1 => n24911, A2 => n25449, B1 => n24904, B2 => 
                           n20608, ZN => n5414);
   U20372 : OAI22_X1 port map( A1 => n24912, A2 => n25452, B1 => n24902, B2 => 
                           n20607, ZN => n5415);
   U20373 : OAI22_X1 port map( A1 => n24912, A2 => n25455, B1 => n21291, B2 => 
                           n20606, ZN => n5416);
   U20374 : OAI22_X1 port map( A1 => n24912, A2 => n25458, B1 => n24902, B2 => 
                           n20605, ZN => n5417);
   U20375 : OAI22_X1 port map( A1 => n24912, A2 => n25461, B1 => n21291, B2 => 
                           n20604, ZN => n5418);
   U20376 : OAI22_X1 port map( A1 => n24912, A2 => n25464, B1 => n24902, B2 => 
                           n20603, ZN => n5419);
   U20377 : OAI22_X1 port map( A1 => n24913, A2 => n25467, B1 => n21291, B2 => 
                           n20602, ZN => n5420);
   U20378 : OAI22_X1 port map( A1 => n24913, A2 => n25470, B1 => n24902, B2 => 
                           n20601, ZN => n5421);
   U20379 : OAI22_X1 port map( A1 => n24913, A2 => n25473, B1 => n24903, B2 => 
                           n20600, ZN => n5422);
   U20380 : OAI22_X1 port map( A1 => n24913, A2 => n25476, B1 => n24904, B2 => 
                           n20599, ZN => n5423);
   U20381 : OAI22_X1 port map( A1 => n24913, A2 => n25479, B1 => n24902, B2 => 
                           n20598, ZN => n5424);
   U20382 : OAI22_X1 port map( A1 => n24914, A2 => n25482, B1 => n24902, B2 => 
                           n20597, ZN => n5425);
   U20383 : OAI22_X1 port map( A1 => n24914, A2 => n25485, B1 => n24903, B2 => 
                           n20596, ZN => n5426);
   U20384 : OAI22_X1 port map( A1 => n24914, A2 => n25488, B1 => n24904, B2 => 
                           n20595, ZN => n5427);
   U20385 : OAI22_X1 port map( A1 => n24914, A2 => n25491, B1 => n24902, B2 => 
                           n20594, ZN => n5428);
   U20386 : OAI22_X1 port map( A1 => n24914, A2 => n25494, B1 => n24902, B2 => 
                           n20593, ZN => n5429);
   U20387 : OAI22_X1 port map( A1 => n24915, A2 => n25497, B1 => n21291, B2 => 
                           n20592, ZN => n5430);
   U20388 : OAI22_X1 port map( A1 => n24915, A2 => n25500, B1 => n24902, B2 => 
                           n20591, ZN => n5431);
   U20389 : OAI22_X1 port map( A1 => n24915, A2 => n25503, B1 => n21291, B2 => 
                           n20590, ZN => n5432);
   U20390 : OAI22_X1 port map( A1 => n24915, A2 => n25506, B1 => n24902, B2 => 
                           n20589, ZN => n5433);
   U20391 : OAI22_X1 port map( A1 => n24915, A2 => n25509, B1 => n21291, B2 => 
                           n20588, ZN => n5434);
   U20392 : OAI22_X1 port map( A1 => n24916, A2 => n25512, B1 => n24902, B2 => 
                           n20587, ZN => n5435);
   U20393 : OAI22_X1 port map( A1 => n24916, A2 => n25515, B1 => n21291, B2 => 
                           n20586, ZN => n5436);
   U20394 : OAI22_X1 port map( A1 => n24916, A2 => n25518, B1 => n24902, B2 => 
                           n20585, ZN => n5437);
   U20395 : OAI22_X1 port map( A1 => n24916, A2 => n25521, B1 => n21291, B2 => 
                           n20584, ZN => n5438);
   U20396 : OAI22_X1 port map( A1 => n24916, A2 => n25524, B1 => n24902, B2 => 
                           n20583, ZN => n5439);
   U20397 : OAI22_X1 port map( A1 => n24841, A2 => n25419, B1 => n24835, B2 => 
                           n20582, ZN => n5148);
   U20398 : OAI22_X1 port map( A1 => n24842, A2 => n25422, B1 => n24836, B2 => 
                           n20581, ZN => n5149);
   U20399 : OAI22_X1 port map( A1 => n24842, A2 => n25425, B1 => n24834, B2 => 
                           n20580, ZN => n5150);
   U20400 : OAI22_X1 port map( A1 => n24842, A2 => n25428, B1 => n24835, B2 => 
                           n20579, ZN => n5151);
   U20401 : OAI22_X1 port map( A1 => n24842, A2 => n25431, B1 => n24836, B2 => 
                           n20578, ZN => n5152);
   U20402 : OAI22_X1 port map( A1 => n24842, A2 => n25434, B1 => n24834, B2 => 
                           n20577, ZN => n5153);
   U20403 : OAI22_X1 port map( A1 => n24843, A2 => n25437, B1 => n24835, B2 => 
                           n20576, ZN => n5154);
   U20404 : OAI22_X1 port map( A1 => n24843, A2 => n25440, B1 => n24836, B2 => 
                           n20575, ZN => n5155);
   U20405 : OAI22_X1 port map( A1 => n24843, A2 => n25443, B1 => n24834, B2 => 
                           n20574, ZN => n5156);
   U20406 : OAI22_X1 port map( A1 => n24843, A2 => n25446, B1 => n24835, B2 => 
                           n20573, ZN => n5157);
   U20407 : OAI22_X1 port map( A1 => n24843, A2 => n25449, B1 => n24836, B2 => 
                           n20572, ZN => n5158);
   U20408 : OAI22_X1 port map( A1 => n24844, A2 => n25452, B1 => n24834, B2 => 
                           n20571, ZN => n5159);
   U20409 : OAI22_X1 port map( A1 => n24844, A2 => n25455, B1 => n21295, B2 => 
                           n20570, ZN => n5160);
   U20410 : OAI22_X1 port map( A1 => n24844, A2 => n25458, B1 => n24834, B2 => 
                           n20569, ZN => n5161);
   U20411 : OAI22_X1 port map( A1 => n24844, A2 => n25461, B1 => n21295, B2 => 
                           n20568, ZN => n5162);
   U20412 : OAI22_X1 port map( A1 => n24844, A2 => n25464, B1 => n24834, B2 => 
                           n20567, ZN => n5163);
   U20413 : OAI22_X1 port map( A1 => n24845, A2 => n25467, B1 => n21295, B2 => 
                           n20566, ZN => n5164);
   U20414 : OAI22_X1 port map( A1 => n24845, A2 => n25470, B1 => n24834, B2 => 
                           n20565, ZN => n5165);
   U20415 : OAI22_X1 port map( A1 => n24845, A2 => n25473, B1 => n24835, B2 => 
                           n20564, ZN => n5166);
   U20416 : OAI22_X1 port map( A1 => n24845, A2 => n25476, B1 => n24836, B2 => 
                           n20563, ZN => n5167);
   U20417 : OAI22_X1 port map( A1 => n24845, A2 => n25479, B1 => n24834, B2 => 
                           n20562, ZN => n5168);
   U20418 : OAI22_X1 port map( A1 => n24846, A2 => n25482, B1 => n24834, B2 => 
                           n20561, ZN => n5169);
   U20419 : OAI22_X1 port map( A1 => n24846, A2 => n25485, B1 => n24835, B2 => 
                           n20560, ZN => n5170);
   U20420 : OAI22_X1 port map( A1 => n24846, A2 => n25488, B1 => n24836, B2 => 
                           n20559, ZN => n5171);
   U20421 : OAI22_X1 port map( A1 => n24846, A2 => n25491, B1 => n24834, B2 => 
                           n20558, ZN => n5172);
   U20422 : OAI22_X1 port map( A1 => n24846, A2 => n25494, B1 => n24834, B2 => 
                           n20557, ZN => n5173);
   U20423 : OAI22_X1 port map( A1 => n24847, A2 => n25497, B1 => n21295, B2 => 
                           n20556, ZN => n5174);
   U20424 : OAI22_X1 port map( A1 => n24847, A2 => n25500, B1 => n24834, B2 => 
                           n20555, ZN => n5175);
   U20425 : OAI22_X1 port map( A1 => n24847, A2 => n25503, B1 => n21295, B2 => 
                           n20554, ZN => n5176);
   U20426 : OAI22_X1 port map( A1 => n24847, A2 => n25506, B1 => n24834, B2 => 
                           n20553, ZN => n5177);
   U20427 : OAI22_X1 port map( A1 => n24847, A2 => n25509, B1 => n21295, B2 => 
                           n20552, ZN => n5178);
   U20428 : OAI22_X1 port map( A1 => n24848, A2 => n25512, B1 => n24834, B2 => 
                           n20551, ZN => n5179);
   U20429 : OAI22_X1 port map( A1 => n24848, A2 => n25515, B1 => n21295, B2 => 
                           n20550, ZN => n5180);
   U20430 : OAI22_X1 port map( A1 => n24848, A2 => n25518, B1 => n24834, B2 => 
                           n20549, ZN => n5181);
   U20431 : OAI22_X1 port map( A1 => n24848, A2 => n25521, B1 => n21295, B2 => 
                           n20548, ZN => n5182);
   U20432 : OAI22_X1 port map( A1 => n24848, A2 => n25524, B1 => n24834, B2 => 
                           n20547, ZN => n5183);
   U20433 : OAI22_X1 port map( A1 => n25062, A2 => n25418, B1 => n25056, B2 => 
                           n20481, ZN => n5980);
   U20434 : OAI22_X1 port map( A1 => n25063, A2 => n25421, B1 => n25057, B2 => 
                           n20480, ZN => n5981);
   U20435 : OAI22_X1 port map( A1 => n25063, A2 => n25424, B1 => n25055, B2 => 
                           n20479, ZN => n5982);
   U20436 : OAI22_X1 port map( A1 => n25063, A2 => n25427, B1 => n25056, B2 => 
                           n20478, ZN => n5983);
   U20437 : OAI22_X1 port map( A1 => n25063, A2 => n25430, B1 => n25057, B2 => 
                           n20477, ZN => n5984);
   U20438 : OAI22_X1 port map( A1 => n25063, A2 => n25433, B1 => n25055, B2 => 
                           n20476, ZN => n5985);
   U20439 : OAI22_X1 port map( A1 => n25064, A2 => n25436, B1 => n25056, B2 => 
                           n20475, ZN => n5986);
   U20440 : OAI22_X1 port map( A1 => n25064, A2 => n25439, B1 => n25057, B2 => 
                           n20474, ZN => n5987);
   U20441 : OAI22_X1 port map( A1 => n25064, A2 => n25442, B1 => n25055, B2 => 
                           n20473, ZN => n5988);
   U20442 : OAI22_X1 port map( A1 => n25064, A2 => n25445, B1 => n25056, B2 => 
                           n20472, ZN => n5989);
   U20443 : OAI22_X1 port map( A1 => n25064, A2 => n25448, B1 => n25057, B2 => 
                           n20471, ZN => n5990);
   U20444 : OAI22_X1 port map( A1 => n25065, A2 => n25451, B1 => n25055, B2 => 
                           n20470, ZN => n5991);
   U20445 : OAI22_X1 port map( A1 => n25065, A2 => n25454, B1 => n21281, B2 => 
                           n20469, ZN => n5992);
   U20446 : OAI22_X1 port map( A1 => n25065, A2 => n25457, B1 => n25055, B2 => 
                           n20468, ZN => n5993);
   U20447 : OAI22_X1 port map( A1 => n25065, A2 => n25460, B1 => n21281, B2 => 
                           n20467, ZN => n5994);
   U20448 : OAI22_X1 port map( A1 => n25065, A2 => n25463, B1 => n25055, B2 => 
                           n20466, ZN => n5995);
   U20449 : OAI22_X1 port map( A1 => n25066, A2 => n25466, B1 => n21281, B2 => 
                           n20465, ZN => n5996);
   U20450 : OAI22_X1 port map( A1 => n25066, A2 => n25469, B1 => n25055, B2 => 
                           n20464, ZN => n5997);
   U20451 : OAI22_X1 port map( A1 => n25066, A2 => n25472, B1 => n25056, B2 => 
                           n20463, ZN => n5998);
   U20452 : OAI22_X1 port map( A1 => n25066, A2 => n25475, B1 => n25057, B2 => 
                           n20462, ZN => n5999);
   U20453 : OAI22_X1 port map( A1 => n25066, A2 => n25478, B1 => n25055, B2 => 
                           n20461, ZN => n6000);
   U20454 : OAI22_X1 port map( A1 => n25067, A2 => n25481, B1 => n25055, B2 => 
                           n20460, ZN => n6001);
   U20455 : OAI22_X1 port map( A1 => n25067, A2 => n25484, B1 => n25056, B2 => 
                           n20459, ZN => n6002);
   U20456 : OAI22_X1 port map( A1 => n25067, A2 => n25487, B1 => n25057, B2 => 
                           n20458, ZN => n6003);
   U20457 : OAI22_X1 port map( A1 => n25067, A2 => n25490, B1 => n25055, B2 => 
                           n20457, ZN => n6004);
   U20458 : OAI22_X1 port map( A1 => n25067, A2 => n25493, B1 => n25055, B2 => 
                           n20456, ZN => n6005);
   U20459 : OAI22_X1 port map( A1 => n25068, A2 => n25496, B1 => n21281, B2 => 
                           n20455, ZN => n6006);
   U20460 : OAI22_X1 port map( A1 => n25068, A2 => n25499, B1 => n25055, B2 => 
                           n20454, ZN => n6007);
   U20461 : OAI22_X1 port map( A1 => n25068, A2 => n25502, B1 => n21281, B2 => 
                           n20453, ZN => n6008);
   U20462 : OAI22_X1 port map( A1 => n25068, A2 => n25505, B1 => n25055, B2 => 
                           n20452, ZN => n6009);
   U20463 : OAI22_X1 port map( A1 => n25068, A2 => n25508, B1 => n21281, B2 => 
                           n20451, ZN => n6010);
   U20464 : OAI22_X1 port map( A1 => n25069, A2 => n25511, B1 => n25055, B2 => 
                           n20450, ZN => n6011);
   U20465 : OAI22_X1 port map( A1 => n25069, A2 => n25514, B1 => n21281, B2 => 
                           n20449, ZN => n6012);
   U20466 : OAI22_X1 port map( A1 => n25069, A2 => n25517, B1 => n25055, B2 => 
                           n20448, ZN => n6013);
   U20467 : OAI22_X1 port map( A1 => n25069, A2 => n25520, B1 => n21281, B2 => 
                           n20447, ZN => n6014);
   U20468 : OAI22_X1 port map( A1 => n25069, A2 => n25523, B1 => n25055, B2 => 
                           n20446, ZN => n6015);
   U20469 : OAI22_X1 port map( A1 => n25317, A2 => n25417, B1 => n25311, B2 => 
                           n20373, ZN => n6940);
   U20470 : OAI22_X1 port map( A1 => n25318, A2 => n25420, B1 => n25312, B2 => 
                           n20372, ZN => n6941);
   U20471 : OAI22_X1 port map( A1 => n25318, A2 => n25423, B1 => n25310, B2 => 
                           n20371, ZN => n6942);
   U20472 : OAI22_X1 port map( A1 => n25318, A2 => n25426, B1 => n25311, B2 => 
                           n20370, ZN => n6943);
   U20473 : OAI22_X1 port map( A1 => n25318, A2 => n25429, B1 => n25312, B2 => 
                           n20369, ZN => n6944);
   U20474 : OAI22_X1 port map( A1 => n25318, A2 => n25432, B1 => n25310, B2 => 
                           n20368, ZN => n6945);
   U20475 : OAI22_X1 port map( A1 => n25319, A2 => n25435, B1 => n25311, B2 => 
                           n20367, ZN => n6946);
   U20476 : OAI22_X1 port map( A1 => n25319, A2 => n25438, B1 => n25312, B2 => 
                           n20366, ZN => n6947);
   U20477 : OAI22_X1 port map( A1 => n25319, A2 => n25441, B1 => n25310, B2 => 
                           n20365, ZN => n6948);
   U20478 : OAI22_X1 port map( A1 => n25319, A2 => n25444, B1 => n25311, B2 => 
                           n20364, ZN => n6949);
   U20479 : OAI22_X1 port map( A1 => n25319, A2 => n25447, B1 => n25312, B2 => 
                           n20363, ZN => n6950);
   U20480 : OAI22_X1 port map( A1 => n25320, A2 => n25450, B1 => n25310, B2 => 
                           n20362, ZN => n6951);
   U20481 : OAI22_X1 port map( A1 => n25320, A2 => n25453, B1 => n21257, B2 => 
                           n20361, ZN => n6952);
   U20482 : OAI22_X1 port map( A1 => n25320, A2 => n25456, B1 => n25310, B2 => 
                           n20360, ZN => n6953);
   U20483 : OAI22_X1 port map( A1 => n25320, A2 => n25459, B1 => n21257, B2 => 
                           n20359, ZN => n6954);
   U20484 : OAI22_X1 port map( A1 => n25320, A2 => n25462, B1 => n25310, B2 => 
                           n20358, ZN => n6955);
   U20485 : OAI22_X1 port map( A1 => n25321, A2 => n25465, B1 => n21257, B2 => 
                           n20357, ZN => n6956);
   U20486 : OAI22_X1 port map( A1 => n25321, A2 => n25468, B1 => n25310, B2 => 
                           n20356, ZN => n6957);
   U20487 : OAI22_X1 port map( A1 => n25321, A2 => n25471, B1 => n25311, B2 => 
                           n20355, ZN => n6958);
   U20488 : OAI22_X1 port map( A1 => n25321, A2 => n25474, B1 => n25312, B2 => 
                           n20354, ZN => n6959);
   U20489 : OAI22_X1 port map( A1 => n25321, A2 => n25477, B1 => n25310, B2 => 
                           n20353, ZN => n6960);
   U20490 : OAI22_X1 port map( A1 => n25322, A2 => n25480, B1 => n25310, B2 => 
                           n20352, ZN => n6961);
   U20491 : OAI22_X1 port map( A1 => n25322, A2 => n25483, B1 => n25311, B2 => 
                           n20351, ZN => n6962);
   U20492 : OAI22_X1 port map( A1 => n25322, A2 => n25486, B1 => n25312, B2 => 
                           n20350, ZN => n6963);
   U20493 : OAI22_X1 port map( A1 => n25322, A2 => n25489, B1 => n25310, B2 => 
                           n20349, ZN => n6964);
   U20494 : OAI22_X1 port map( A1 => n25322, A2 => n25492, B1 => n25310, B2 => 
                           n20348, ZN => n6965);
   U20495 : OAI22_X1 port map( A1 => n25323, A2 => n25495, B1 => n21257, B2 => 
                           n20347, ZN => n6966);
   U20496 : OAI22_X1 port map( A1 => n25323, A2 => n25498, B1 => n25310, B2 => 
                           n20346, ZN => n6967);
   U20497 : OAI22_X1 port map( A1 => n25323, A2 => n25501, B1 => n21257, B2 => 
                           n20345, ZN => n6968);
   U20498 : OAI22_X1 port map( A1 => n25323, A2 => n25504, B1 => n25310, B2 => 
                           n20344, ZN => n6969);
   U20499 : OAI22_X1 port map( A1 => n25323, A2 => n25507, B1 => n21257, B2 => 
                           n20343, ZN => n6970);
   U20500 : OAI22_X1 port map( A1 => n25324, A2 => n25510, B1 => n25310, B2 => 
                           n20342, ZN => n6971);
   U20501 : OAI22_X1 port map( A1 => n25324, A2 => n25513, B1 => n21257, B2 => 
                           n20341, ZN => n6972);
   U20502 : OAI22_X1 port map( A1 => n25324, A2 => n25516, B1 => n25310, B2 => 
                           n20340, ZN => n6973);
   U20503 : OAI22_X1 port map( A1 => n25324, A2 => n25519, B1 => n21257, B2 => 
                           n20339, ZN => n6974);
   U20504 : OAI22_X1 port map( A1 => n25324, A2 => n25522, B1 => n25310, B2 => 
                           n20338, ZN => n6975);
   U20505 : OAI22_X1 port map( A1 => n25198, A2 => n25417, B1 => n25192, B2 => 
                           n20337, ZN => n6492);
   U20506 : OAI22_X1 port map( A1 => n25199, A2 => n25420, B1 => n25193, B2 => 
                           n20336, ZN => n6493);
   U20507 : OAI22_X1 port map( A1 => n25199, A2 => n25423, B1 => n25191, B2 => 
                           n20335, ZN => n6494);
   U20508 : OAI22_X1 port map( A1 => n25199, A2 => n25426, B1 => n25192, B2 => 
                           n20334, ZN => n6495);
   U20509 : OAI22_X1 port map( A1 => n25199, A2 => n25429, B1 => n25193, B2 => 
                           n20333, ZN => n6496);
   U20510 : OAI22_X1 port map( A1 => n25199, A2 => n25432, B1 => n25191, B2 => 
                           n20332, ZN => n6497);
   U20511 : OAI22_X1 port map( A1 => n25200, A2 => n25435, B1 => n25192, B2 => 
                           n20331, ZN => n6498);
   U20512 : OAI22_X1 port map( A1 => n25200, A2 => n25438, B1 => n25193, B2 => 
                           n20330, ZN => n6499);
   U20513 : OAI22_X1 port map( A1 => n25200, A2 => n25441, B1 => n25191, B2 => 
                           n20329, ZN => n6500);
   U20514 : OAI22_X1 port map( A1 => n25200, A2 => n25444, B1 => n25192, B2 => 
                           n20328, ZN => n6501);
   U20515 : OAI22_X1 port map( A1 => n25200, A2 => n25447, B1 => n25193, B2 => 
                           n20327, ZN => n6502);
   U20516 : OAI22_X1 port map( A1 => n25201, A2 => n25450, B1 => n25191, B2 => 
                           n20326, ZN => n6503);
   U20517 : OAI22_X1 port map( A1 => n25201, A2 => n25453, B1 => n21272, B2 => 
                           n20325, ZN => n6504);
   U20518 : OAI22_X1 port map( A1 => n25201, A2 => n25456, B1 => n25191, B2 => 
                           n20324, ZN => n6505);
   U20519 : OAI22_X1 port map( A1 => n25201, A2 => n25459, B1 => n21272, B2 => 
                           n20323, ZN => n6506);
   U20520 : OAI22_X1 port map( A1 => n25201, A2 => n25462, B1 => n25191, B2 => 
                           n20322, ZN => n6507);
   U20521 : OAI22_X1 port map( A1 => n25202, A2 => n25465, B1 => n21272, B2 => 
                           n20321, ZN => n6508);
   U20522 : OAI22_X1 port map( A1 => n25202, A2 => n25468, B1 => n25191, B2 => 
                           n20320, ZN => n6509);
   U20523 : OAI22_X1 port map( A1 => n25202, A2 => n25471, B1 => n25192, B2 => 
                           n20319, ZN => n6510);
   U20524 : OAI22_X1 port map( A1 => n25202, A2 => n25474, B1 => n25193, B2 => 
                           n20318, ZN => n6511);
   U20525 : OAI22_X1 port map( A1 => n25202, A2 => n25477, B1 => n25191, B2 => 
                           n20317, ZN => n6512);
   U20526 : OAI22_X1 port map( A1 => n25203, A2 => n25480, B1 => n25191, B2 => 
                           n20316, ZN => n6513);
   U20527 : OAI22_X1 port map( A1 => n25203, A2 => n25483, B1 => n25192, B2 => 
                           n20315, ZN => n6514);
   U20528 : OAI22_X1 port map( A1 => n25203, A2 => n25486, B1 => n25193, B2 => 
                           n20314, ZN => n6515);
   U20529 : OAI22_X1 port map( A1 => n25203, A2 => n25489, B1 => n25191, B2 => 
                           n20313, ZN => n6516);
   U20530 : OAI22_X1 port map( A1 => n25203, A2 => n25492, B1 => n25191, B2 => 
                           n20312, ZN => n6517);
   U20531 : OAI22_X1 port map( A1 => n25204, A2 => n25495, B1 => n21272, B2 => 
                           n20311, ZN => n6518);
   U20532 : OAI22_X1 port map( A1 => n25204, A2 => n25498, B1 => n25191, B2 => 
                           n20310, ZN => n6519);
   U20533 : OAI22_X1 port map( A1 => n25204, A2 => n25501, B1 => n21272, B2 => 
                           n20309, ZN => n6520);
   U20534 : OAI22_X1 port map( A1 => n25204, A2 => n25504, B1 => n25191, B2 => 
                           n20308, ZN => n6521);
   U20535 : OAI22_X1 port map( A1 => n25204, A2 => n25507, B1 => n21272, B2 => 
                           n20307, ZN => n6522);
   U20536 : OAI22_X1 port map( A1 => n25205, A2 => n25510, B1 => n25191, B2 => 
                           n20306, ZN => n6523);
   U20537 : OAI22_X1 port map( A1 => n25205, A2 => n25513, B1 => n21272, B2 => 
                           n20305, ZN => n6524);
   U20538 : OAI22_X1 port map( A1 => n25205, A2 => n25516, B1 => n25191, B2 => 
                           n20304, ZN => n6525);
   U20539 : OAI22_X1 port map( A1 => n25205, A2 => n25519, B1 => n21272, B2 => 
                           n20303, ZN => n6526);
   U20540 : OAI22_X1 port map( A1 => n25205, A2 => n25522, B1 => n25191, B2 => 
                           n20302, ZN => n6527);
   U20541 : OAI22_X1 port map( A1 => n25300, A2 => n25417, B1 => n25294, B2 => 
                           n20301, ZN => n6876);
   U20542 : OAI22_X1 port map( A1 => n25301, A2 => n25420, B1 => n25295, B2 => 
                           n20300, ZN => n6877);
   U20543 : OAI22_X1 port map( A1 => n25301, A2 => n25423, B1 => n25293, B2 => 
                           n20299, ZN => n6878);
   U20544 : OAI22_X1 port map( A1 => n25301, A2 => n25426, B1 => n25294, B2 => 
                           n20298, ZN => n6879);
   U20545 : OAI22_X1 port map( A1 => n25301, A2 => n25429, B1 => n25295, B2 => 
                           n20297, ZN => n6880);
   U20546 : OAI22_X1 port map( A1 => n25301, A2 => n25432, B1 => n25293, B2 => 
                           n20296, ZN => n6881);
   U20547 : OAI22_X1 port map( A1 => n25302, A2 => n25435, B1 => n25294, B2 => 
                           n20295, ZN => n6882);
   U20548 : OAI22_X1 port map( A1 => n25302, A2 => n25438, B1 => n25295, B2 => 
                           n20294, ZN => n6883);
   U20549 : OAI22_X1 port map( A1 => n25302, A2 => n25441, B1 => n25293, B2 => 
                           n20293, ZN => n6884);
   U20550 : OAI22_X1 port map( A1 => n25302, A2 => n25444, B1 => n25294, B2 => 
                           n20292, ZN => n6885);
   U20551 : OAI22_X1 port map( A1 => n25302, A2 => n25447, B1 => n25295, B2 => 
                           n20291, ZN => n6886);
   U20552 : OAI22_X1 port map( A1 => n25303, A2 => n25450, B1 => n25293, B2 => 
                           n20290, ZN => n6887);
   U20553 : OAI22_X1 port map( A1 => n25303, A2 => n25453, B1 => n21259, B2 => 
                           n20289, ZN => n6888);
   U20554 : OAI22_X1 port map( A1 => n25303, A2 => n25456, B1 => n25293, B2 => 
                           n20288, ZN => n6889);
   U20555 : OAI22_X1 port map( A1 => n25303, A2 => n25459, B1 => n21259, B2 => 
                           n20287, ZN => n6890);
   U20556 : OAI22_X1 port map( A1 => n25303, A2 => n25462, B1 => n25293, B2 => 
                           n20286, ZN => n6891);
   U20557 : OAI22_X1 port map( A1 => n25304, A2 => n25465, B1 => n21259, B2 => 
                           n20285, ZN => n6892);
   U20558 : OAI22_X1 port map( A1 => n25304, A2 => n25468, B1 => n25293, B2 => 
                           n20284, ZN => n6893);
   U20559 : OAI22_X1 port map( A1 => n25304, A2 => n25471, B1 => n25294, B2 => 
                           n20283, ZN => n6894);
   U20560 : OAI22_X1 port map( A1 => n25304, A2 => n25474, B1 => n25295, B2 => 
                           n20282, ZN => n6895);
   U20561 : OAI22_X1 port map( A1 => n25304, A2 => n25477, B1 => n25293, B2 => 
                           n20281, ZN => n6896);
   U20562 : OAI22_X1 port map( A1 => n25305, A2 => n25480, B1 => n25293, B2 => 
                           n20280, ZN => n6897);
   U20563 : OAI22_X1 port map( A1 => n25305, A2 => n25483, B1 => n25294, B2 => 
                           n20279, ZN => n6898);
   U20564 : OAI22_X1 port map( A1 => n25305, A2 => n25486, B1 => n25295, B2 => 
                           n20278, ZN => n6899);
   U20565 : OAI22_X1 port map( A1 => n25305, A2 => n25489, B1 => n25293, B2 => 
                           n20277, ZN => n6900);
   U20566 : OAI22_X1 port map( A1 => n25305, A2 => n25492, B1 => n25293, B2 => 
                           n20276, ZN => n6901);
   U20567 : OAI22_X1 port map( A1 => n25306, A2 => n25495, B1 => n21259, B2 => 
                           n20275, ZN => n6902);
   U20568 : OAI22_X1 port map( A1 => n25306, A2 => n25498, B1 => n25293, B2 => 
                           n20274, ZN => n6903);
   U20569 : OAI22_X1 port map( A1 => n25306, A2 => n25501, B1 => n21259, B2 => 
                           n20273, ZN => n6904);
   U20570 : OAI22_X1 port map( A1 => n25306, A2 => n25504, B1 => n25293, B2 => 
                           n20272, ZN => n6905);
   U20571 : OAI22_X1 port map( A1 => n25306, A2 => n25507, B1 => n21259, B2 => 
                           n20271, ZN => n6906);
   U20572 : OAI22_X1 port map( A1 => n25307, A2 => n25510, B1 => n25293, B2 => 
                           n20270, ZN => n6907);
   U20573 : OAI22_X1 port map( A1 => n25307, A2 => n25513, B1 => n21259, B2 => 
                           n20269, ZN => n6908);
   U20574 : OAI22_X1 port map( A1 => n25307, A2 => n25516, B1 => n25293, B2 => 
                           n20268, ZN => n6909);
   U20575 : OAI22_X1 port map( A1 => n25307, A2 => n25519, B1 => n21259, B2 => 
                           n20267, ZN => n6910);
   U20576 : OAI22_X1 port map( A1 => n25307, A2 => n25522, B1 => n25293, B2 => 
                           n20266, ZN => n6911);
   U20577 : OAI22_X1 port map( A1 => n24877, A2 => n25437, B1 => n24868, B2 => 
                           n20186, ZN => n5282);
   U20578 : OAI22_X1 port map( A1 => n24877, A2 => n25440, B1 => n24868, B2 => 
                           n20185, ZN => n5283);
   U20579 : OAI22_X1 port map( A1 => n24877, A2 => n25443, B1 => n21293, B2 => 
                           n20184, ZN => n5284);
   U20580 : OAI22_X1 port map( A1 => n24877, A2 => n25446, B1 => n24868, B2 => 
                           n20183, ZN => n5285);
   U20581 : OAI22_X1 port map( A1 => n24877, A2 => n25449, B1 => n21293, B2 => 
                           n20182, ZN => n5286);
   U20582 : OAI22_X1 port map( A1 => n24878, A2 => n25452, B1 => n24868, B2 => 
                           n20181, ZN => n5287);
   U20583 : OAI22_X1 port map( A1 => n24878, A2 => n25455, B1 => n24869, B2 => 
                           n20180, ZN => n5288);
   U20584 : OAI22_X1 port map( A1 => n24878, A2 => n25458, B1 => n24870, B2 => 
                           n20179, ZN => n5289);
   U20585 : OAI22_X1 port map( A1 => n24878, A2 => n25461, B1 => n24868, B2 => 
                           n20178, ZN => n5290);
   U20586 : OAI22_X1 port map( A1 => n24878, A2 => n25464, B1 => n24869, B2 => 
                           n20177, ZN => n5291);
   U20587 : OAI22_X1 port map( A1 => n24879, A2 => n25467, B1 => n24870, B2 => 
                           n20176, ZN => n5292);
   U20588 : OAI22_X1 port map( A1 => n24879, A2 => n25470, B1 => n24868, B2 => 
                           n20175, ZN => n5293);
   U20589 : OAI22_X1 port map( A1 => n24879, A2 => n25473, B1 => n24869, B2 => 
                           n20174, ZN => n5294);
   U20590 : OAI22_X1 port map( A1 => n24879, A2 => n25476, B1 => n24870, B2 => 
                           n20173, ZN => n5295);
   U20591 : OAI22_X1 port map( A1 => n24879, A2 => n25479, B1 => n24868, B2 => 
                           n20172, ZN => n5296);
   U20592 : OAI22_X1 port map( A1 => n24880, A2 => n25482, B1 => n24869, B2 => 
                           n20171, ZN => n5297);
   U20593 : OAI22_X1 port map( A1 => n24880, A2 => n25485, B1 => n24870, B2 => 
                           n20170, ZN => n5298);
   U20594 : OAI22_X1 port map( A1 => n24880, A2 => n25488, B1 => n24868, B2 => 
                           n20169, ZN => n5299);
   U20595 : OAI22_X1 port map( A1 => n24880, A2 => n25491, B1 => n21293, B2 => 
                           n20168, ZN => n5300);
   U20596 : OAI22_X1 port map( A1 => n24880, A2 => n25494, B1 => n24868, B2 => 
                           n20167, ZN => n5301);
   U20597 : OAI22_X1 port map( A1 => n24881, A2 => n25497, B1 => n21293, B2 => 
                           n20166, ZN => n5302);
   U20598 : OAI22_X1 port map( A1 => n24881, A2 => n25500, B1 => n24868, B2 => 
                           n20165, ZN => n5303);
   U20599 : OAI22_X1 port map( A1 => n24881, A2 => n25503, B1 => n21293, B2 => 
                           n20164, ZN => n5304);
   U20600 : OAI22_X1 port map( A1 => n24881, A2 => n25506, B1 => n24868, B2 => 
                           n20163, ZN => n5305);
   U20601 : OAI22_X1 port map( A1 => n24881, A2 => n25509, B1 => n24869, B2 => 
                           n20162, ZN => n5306);
   U20602 : OAI22_X1 port map( A1 => n24882, A2 => n25512, B1 => n24870, B2 => 
                           n20161, ZN => n5307);
   U20603 : OAI22_X1 port map( A1 => n24882, A2 => n25515, B1 => n24868, B2 => 
                           n20160, ZN => n5308);
   U20604 : OAI22_X1 port map( A1 => n24882, A2 => n25518, B1 => n24868, B2 => 
                           n20159, ZN => n5309);
   U20605 : OAI22_X1 port map( A1 => n24882, A2 => n25521, B1 => n24869, B2 => 
                           n20158, ZN => n5310);
   U20606 : OAI22_X1 port map( A1 => n24882, A2 => n25524, B1 => n24870, B2 => 
                           n20157, ZN => n5311);
   U20607 : OAI22_X1 port map( A1 => n24875, A2 => n25419, B1 => n21293, B2 => 
                           n19713, ZN => n5276);
   U20608 : OAI22_X1 port map( A1 => n24876, A2 => n25422, B1 => n24868, B2 => 
                           n19712, ZN => n5277);
   U20609 : OAI22_X1 port map( A1 => n24876, A2 => n25425, B1 => n21293, B2 => 
                           n19711, ZN => n5278);
   U20610 : OAI22_X1 port map( A1 => n24876, A2 => n25428, B1 => n24868, B2 => 
                           n19710, ZN => n5279);
   U20611 : OAI22_X1 port map( A1 => n24876, A2 => n25431, B1 => n21293, B2 => 
                           n19709, ZN => n5280);
   U20612 : OAI22_X1 port map( A1 => n24876, A2 => n25434, B1 => n24868, B2 => 
                           n19708, ZN => n5281);
   U20613 : OAI22_X1 port map( A1 => n24943, A2 => n25419, B1 => n24937, B2 => 
                           n19683, ZN => n5532);
   U20614 : OAI22_X1 port map( A1 => n24944, A2 => n25422, B1 => n24938, B2 => 
                           n19682, ZN => n5533);
   U20615 : OAI22_X1 port map( A1 => n24944, A2 => n25425, B1 => n24936, B2 => 
                           n19681, ZN => n5534);
   U20616 : OAI22_X1 port map( A1 => n24944, A2 => n25428, B1 => n24937, B2 => 
                           n19680, ZN => n5535);
   U20617 : OAI22_X1 port map( A1 => n24944, A2 => n25431, B1 => n24938, B2 => 
                           n19679, ZN => n5536);
   U20618 : OAI22_X1 port map( A1 => n24944, A2 => n25434, B1 => n24936, B2 => 
                           n19678, ZN => n5537);
   U20619 : OAI22_X1 port map( A1 => n24945, A2 => n25437, B1 => n24937, B2 => 
                           n19677, ZN => n5538);
   U20620 : OAI22_X1 port map( A1 => n24945, A2 => n25440, B1 => n24938, B2 => 
                           n19676, ZN => n5539);
   U20621 : OAI22_X1 port map( A1 => n24945, A2 => n25443, B1 => n24936, B2 => 
                           n19675, ZN => n5540);
   U20622 : OAI22_X1 port map( A1 => n24945, A2 => n25446, B1 => n24937, B2 => 
                           n19674, ZN => n5541);
   U20623 : OAI22_X1 port map( A1 => n24945, A2 => n25449, B1 => n24938, B2 => 
                           n19673, ZN => n5542);
   U20624 : OAI22_X1 port map( A1 => n24946, A2 => n25452, B1 => n24936, B2 => 
                           n19672, ZN => n5543);
   U20625 : OAI22_X1 port map( A1 => n24946, A2 => n25455, B1 => n21288, B2 => 
                           n19671, ZN => n5544);
   U20626 : OAI22_X1 port map( A1 => n24946, A2 => n25458, B1 => n24936, B2 => 
                           n19670, ZN => n5545);
   U20627 : OAI22_X1 port map( A1 => n24946, A2 => n25461, B1 => n21288, B2 => 
                           n19669, ZN => n5546);
   U20628 : OAI22_X1 port map( A1 => n24946, A2 => n25464, B1 => n24936, B2 => 
                           n19668, ZN => n5547);
   U20629 : OAI22_X1 port map( A1 => n24947, A2 => n25467, B1 => n21288, B2 => 
                           n19667, ZN => n5548);
   U20630 : OAI22_X1 port map( A1 => n24947, A2 => n25470, B1 => n24936, B2 => 
                           n19666, ZN => n5549);
   U20631 : OAI22_X1 port map( A1 => n24947, A2 => n25473, B1 => n24937, B2 => 
                           n19665, ZN => n5550);
   U20632 : OAI22_X1 port map( A1 => n24947, A2 => n25476, B1 => n24938, B2 => 
                           n19664, ZN => n5551);
   U20633 : OAI22_X1 port map( A1 => n24947, A2 => n25479, B1 => n24936, B2 => 
                           n19663, ZN => n5552);
   U20634 : OAI22_X1 port map( A1 => n24948, A2 => n25482, B1 => n24936, B2 => 
                           n19662, ZN => n5553);
   U20635 : OAI22_X1 port map( A1 => n24948, A2 => n25485, B1 => n24937, B2 => 
                           n19661, ZN => n5554);
   U20636 : OAI22_X1 port map( A1 => n24948, A2 => n25488, B1 => n24938, B2 => 
                           n19660, ZN => n5555);
   U20637 : OAI22_X1 port map( A1 => n24948, A2 => n25491, B1 => n24936, B2 => 
                           n19659, ZN => n5556);
   U20638 : OAI22_X1 port map( A1 => n24948, A2 => n25494, B1 => n24936, B2 => 
                           n19658, ZN => n5557);
   U20639 : OAI22_X1 port map( A1 => n24949, A2 => n25497, B1 => n21288, B2 => 
                           n19657, ZN => n5558);
   U20640 : OAI22_X1 port map( A1 => n24949, A2 => n25500, B1 => n24936, B2 => 
                           n19656, ZN => n5559);
   U20641 : OAI22_X1 port map( A1 => n24949, A2 => n25503, B1 => n21288, B2 => 
                           n19655, ZN => n5560);
   U20642 : OAI22_X1 port map( A1 => n24949, A2 => n25506, B1 => n24936, B2 => 
                           n19654, ZN => n5561);
   U20643 : OAI22_X1 port map( A1 => n24949, A2 => n25509, B1 => n21288, B2 => 
                           n19653, ZN => n5562);
   U20644 : OAI22_X1 port map( A1 => n24950, A2 => n25512, B1 => n24936, B2 => 
                           n19652, ZN => n5563);
   U20645 : OAI22_X1 port map( A1 => n24950, A2 => n25515, B1 => n21288, B2 => 
                           n19651, ZN => n5564);
   U20646 : OAI22_X1 port map( A1 => n24950, A2 => n25518, B1 => n24936, B2 => 
                           n19650, ZN => n5565);
   U20647 : OAI22_X1 port map( A1 => n24950, A2 => n25521, B1 => n21288, B2 => 
                           n19649, ZN => n5566);
   U20648 : OAI22_X1 port map( A1 => n24950, A2 => n25524, B1 => n24936, B2 => 
                           n19648, ZN => n5567);
   U20649 : OAI22_X1 port map( A1 => n25283, A2 => n25417, B1 => n25277, B2 => 
                           n19371, ZN => n6812);
   U20650 : OAI22_X1 port map( A1 => n25284, A2 => n25420, B1 => n25278, B2 => 
                           n19370, ZN => n6813);
   U20651 : OAI22_X1 port map( A1 => n25284, A2 => n25423, B1 => n25276, B2 => 
                           n19369, ZN => n6814);
   U20652 : OAI22_X1 port map( A1 => n25284, A2 => n25426, B1 => n25277, B2 => 
                           n19368, ZN => n6815);
   U20653 : OAI22_X1 port map( A1 => n25284, A2 => n25429, B1 => n25278, B2 => 
                           n19367, ZN => n6816);
   U20654 : OAI22_X1 port map( A1 => n25284, A2 => n25432, B1 => n25276, B2 => 
                           n19366, ZN => n6817);
   U20655 : OAI22_X1 port map( A1 => n25285, A2 => n25435, B1 => n25277, B2 => 
                           n19365, ZN => n6818);
   U20656 : OAI22_X1 port map( A1 => n25285, A2 => n25438, B1 => n25278, B2 => 
                           n19364, ZN => n6819);
   U20657 : OAI22_X1 port map( A1 => n25285, A2 => n25441, B1 => n25276, B2 => 
                           n19363, ZN => n6820);
   U20658 : OAI22_X1 port map( A1 => n25285, A2 => n25444, B1 => n25277, B2 => 
                           n19362, ZN => n6821);
   U20659 : OAI22_X1 port map( A1 => n25285, A2 => n25447, B1 => n25278, B2 => 
                           n19361, ZN => n6822);
   U20660 : OAI22_X1 port map( A1 => n25286, A2 => n25450, B1 => n25276, B2 => 
                           n19360, ZN => n6823);
   U20661 : OAI22_X1 port map( A1 => n25286, A2 => n25453, B1 => n21261, B2 => 
                           n19359, ZN => n6824);
   U20662 : OAI22_X1 port map( A1 => n25286, A2 => n25456, B1 => n25276, B2 => 
                           n19358, ZN => n6825);
   U20663 : OAI22_X1 port map( A1 => n25286, A2 => n25459, B1 => n21261, B2 => 
                           n19357, ZN => n6826);
   U20664 : OAI22_X1 port map( A1 => n25286, A2 => n25462, B1 => n25276, B2 => 
                           n19356, ZN => n6827);
   U20665 : OAI22_X1 port map( A1 => n25287, A2 => n25465, B1 => n21261, B2 => 
                           n19355, ZN => n6828);
   U20666 : OAI22_X1 port map( A1 => n25287, A2 => n25468, B1 => n25276, B2 => 
                           n19354, ZN => n6829);
   U20667 : OAI22_X1 port map( A1 => n25287, A2 => n25471, B1 => n25277, B2 => 
                           n19353, ZN => n6830);
   U20668 : OAI22_X1 port map( A1 => n25287, A2 => n25474, B1 => n25278, B2 => 
                           n19352, ZN => n6831);
   U20669 : OAI22_X1 port map( A1 => n25287, A2 => n25477, B1 => n25276, B2 => 
                           n19351, ZN => n6832);
   U20670 : OAI22_X1 port map( A1 => n25288, A2 => n25480, B1 => n25276, B2 => 
                           n19350, ZN => n6833);
   U20671 : OAI22_X1 port map( A1 => n25288, A2 => n25483, B1 => n25277, B2 => 
                           n19349, ZN => n6834);
   U20672 : OAI22_X1 port map( A1 => n25288, A2 => n25486, B1 => n25278, B2 => 
                           n19348, ZN => n6835);
   U20673 : OAI22_X1 port map( A1 => n25288, A2 => n25489, B1 => n25276, B2 => 
                           n19347, ZN => n6836);
   U20674 : OAI22_X1 port map( A1 => n25288, A2 => n25492, B1 => n25276, B2 => 
                           n19346, ZN => n6837);
   U20675 : OAI22_X1 port map( A1 => n25289, A2 => n25495, B1 => n21261, B2 => 
                           n19345, ZN => n6838);
   U20676 : OAI22_X1 port map( A1 => n25289, A2 => n25498, B1 => n25276, B2 => 
                           n19344, ZN => n6839);
   U20677 : OAI22_X1 port map( A1 => n25289, A2 => n25501, B1 => n21261, B2 => 
                           n19343, ZN => n6840);
   U20678 : OAI22_X1 port map( A1 => n25289, A2 => n25504, B1 => n25276, B2 => 
                           n19342, ZN => n6841);
   U20679 : OAI22_X1 port map( A1 => n25289, A2 => n25507, B1 => n21261, B2 => 
                           n19341, ZN => n6842);
   U20680 : OAI22_X1 port map( A1 => n25290, A2 => n25510, B1 => n25276, B2 => 
                           n19340, ZN => n6843);
   U20681 : OAI22_X1 port map( A1 => n25290, A2 => n25513, B1 => n21261, B2 => 
                           n19339, ZN => n6844);
   U20682 : OAI22_X1 port map( A1 => n25290, A2 => n25516, B1 => n25276, B2 => 
                           n19338, ZN => n6845);
   U20683 : OAI22_X1 port map( A1 => n25290, A2 => n25519, B1 => n21261, B2 => 
                           n19337, ZN => n6846);
   U20684 : OAI22_X1 port map( A1 => n25290, A2 => n25522, B1 => n25276, B2 => 
                           n19336, ZN => n6847);
   U20685 : OAI22_X1 port map( A1 => n25541, A2 => n25417, B1 => n25535, B2 => 
                           n19307, ZN => n7068);
   U20686 : OAI22_X1 port map( A1 => n25542, A2 => n25420, B1 => n25536, B2 => 
                           n19306, ZN => n7069);
   U20687 : OAI22_X1 port map( A1 => n25542, A2 => n25423, B1 => n25534, B2 => 
                           n19305, ZN => n7070);
   U20688 : OAI22_X1 port map( A1 => n25542, A2 => n25426, B1 => n25535, B2 => 
                           n19304, ZN => n7071);
   U20689 : OAI22_X1 port map( A1 => n25542, A2 => n25429, B1 => n25536, B2 => 
                           n19303, ZN => n7072);
   U20690 : OAI22_X1 port map( A1 => n25542, A2 => n25432, B1 => n25534, B2 => 
                           n19302, ZN => n7073);
   U20691 : OAI22_X1 port map( A1 => n25543, A2 => n25435, B1 => n25535, B2 => 
                           n19301, ZN => n7074);
   U20692 : OAI22_X1 port map( A1 => n25543, A2 => n25438, B1 => n25536, B2 => 
                           n19300, ZN => n7075);
   U20693 : OAI22_X1 port map( A1 => n25543, A2 => n25441, B1 => n25534, B2 => 
                           n19299, ZN => n7076);
   U20694 : OAI22_X1 port map( A1 => n25543, A2 => n25444, B1 => n25535, B2 => 
                           n19298, ZN => n7077);
   U20695 : OAI22_X1 port map( A1 => n25543, A2 => n25447, B1 => n25536, B2 => 
                           n19297, ZN => n7078);
   U20696 : OAI22_X1 port map( A1 => n25544, A2 => n25450, B1 => n25534, B2 => 
                           n19296, ZN => n7079);
   U20697 : OAI22_X1 port map( A1 => n25544, A2 => n25453, B1 => n21189, B2 => 
                           n19295, ZN => n7080);
   U20698 : OAI22_X1 port map( A1 => n25544, A2 => n25456, B1 => n25534, B2 => 
                           n19294, ZN => n7081);
   U20699 : OAI22_X1 port map( A1 => n25544, A2 => n25459, B1 => n21189, B2 => 
                           n19293, ZN => n7082);
   U20700 : OAI22_X1 port map( A1 => n25544, A2 => n25462, B1 => n25534, B2 => 
                           n19292, ZN => n7083);
   U20701 : OAI22_X1 port map( A1 => n25545, A2 => n25465, B1 => n21189, B2 => 
                           n19291, ZN => n7084);
   U20702 : OAI22_X1 port map( A1 => n25545, A2 => n25468, B1 => n25534, B2 => 
                           n19290, ZN => n7085);
   U20703 : OAI22_X1 port map( A1 => n25545, A2 => n25471, B1 => n25535, B2 => 
                           n19289, ZN => n7086);
   U20704 : OAI22_X1 port map( A1 => n25545, A2 => n25474, B1 => n25536, B2 => 
                           n19288, ZN => n7087);
   U20705 : OAI22_X1 port map( A1 => n25545, A2 => n25477, B1 => n25534, B2 => 
                           n19287, ZN => n7088);
   U20706 : OAI22_X1 port map( A1 => n25546, A2 => n25480, B1 => n25534, B2 => 
                           n19286, ZN => n7089);
   U20707 : OAI22_X1 port map( A1 => n25546, A2 => n25483, B1 => n25535, B2 => 
                           n19285, ZN => n7090);
   U20708 : OAI22_X1 port map( A1 => n25546, A2 => n25486, B1 => n25536, B2 => 
                           n19284, ZN => n7091);
   U20709 : OAI22_X1 port map( A1 => n25546, A2 => n25489, B1 => n25534, B2 => 
                           n19283, ZN => n7092);
   U20710 : OAI22_X1 port map( A1 => n25546, A2 => n25492, B1 => n25534, B2 => 
                           n19282, ZN => n7093);
   U20711 : OAI22_X1 port map( A1 => n25547, A2 => n25495, B1 => n21189, B2 => 
                           n19281, ZN => n7094);
   U20712 : OAI22_X1 port map( A1 => n25547, A2 => n25498, B1 => n25534, B2 => 
                           n19280, ZN => n7095);
   U20713 : OAI22_X1 port map( A1 => n25547, A2 => n25501, B1 => n21189, B2 => 
                           n19279, ZN => n7096);
   U20714 : OAI22_X1 port map( A1 => n25547, A2 => n25504, B1 => n25534, B2 => 
                           n19278, ZN => n7097);
   U20715 : OAI22_X1 port map( A1 => n25547, A2 => n25507, B1 => n21189, B2 => 
                           n19277, ZN => n7098);
   U20716 : OAI22_X1 port map( A1 => n25548, A2 => n25510, B1 => n25534, B2 => 
                           n19276, ZN => n7099);
   U20717 : OAI22_X1 port map( A1 => n25548, A2 => n25513, B1 => n21189, B2 => 
                           n19275, ZN => n7100);
   U20718 : OAI22_X1 port map( A1 => n25548, A2 => n25516, B1 => n25534, B2 => 
                           n19274, ZN => n7101);
   U20719 : OAI22_X1 port map( A1 => n25548, A2 => n25519, B1 => n21189, B2 => 
                           n19273, ZN => n7102);
   U20720 : OAI22_X1 port map( A1 => n25548, A2 => n25522, B1 => n25534, B2 => 
                           n19272, ZN => n7103);
   U20721 : OAI22_X1 port map( A1 => n25330, A2 => n25348, B1 => n21255, B2 => 
                           n21147, ZN => n6981);
   U20722 : OAI22_X1 port map( A1 => n25002, A2 => n25526, B1 => n21285, B2 => 
                           n20546, ZN => n5760);
   U20723 : OAI22_X1 port map( A1 => n25002, A2 => n25529, B1 => n21285, B2 => 
                           n20545, ZN => n5761);
   U20724 : OAI22_X1 port map( A1 => n25002, A2 => n25532, B1 => n24987, B2 => 
                           n20544, ZN => n5762);
   U20725 : OAI22_X1 port map( A1 => n25002, A2 => n25552, B1 => n21285, B2 => 
                           n20543, ZN => n5763);
   U20726 : OAI22_X1 port map( A1 => n25240, A2 => n25525, B1 => n21267, B2 => 
                           n20542, ZN => n6656);
   U20727 : OAI22_X1 port map( A1 => n25240, A2 => n25528, B1 => n21267, B2 => 
                           n20541, ZN => n6657);
   U20728 : OAI22_X1 port map( A1 => n25240, A2 => n25531, B1 => n25225, B2 => 
                           n20540, ZN => n6658);
   U20729 : OAI22_X1 port map( A1 => n25240, A2 => n25551, B1 => n21267, B2 => 
                           n20539, ZN => n6659);
   U20730 : OAI22_X1 port map( A1 => n25223, A2 => n25525, B1 => n21270, B2 => 
                           n20538, ZN => n6592);
   U20731 : OAI22_X1 port map( A1 => n25223, A2 => n25528, B1 => n21270, B2 => 
                           n20537, ZN => n6593);
   U20732 : OAI22_X1 port map( A1 => n25223, A2 => n25531, B1 => n25208, B2 => 
                           n20536, ZN => n6594);
   U20733 : OAI22_X1 port map( A1 => n25223, A2 => n25551, B1 => n21270, B2 => 
                           n20535, ZN => n6595);
   U20734 : OAI22_X1 port map( A1 => n25155, A2 => n25526, B1 => n21275, B2 => 
                           n20534, ZN => n6336);
   U20735 : OAI22_X1 port map( A1 => n25155, A2 => n25529, B1 => n21275, B2 => 
                           n20533, ZN => n6337);
   U20736 : OAI22_X1 port map( A1 => n25155, A2 => n25532, B1 => n25140, B2 => 
                           n20532, ZN => n6338);
   U20737 : OAI22_X1 port map( A1 => n25155, A2 => n25552, B1 => n21275, B2 => 
                           n20531, ZN => n6339);
   U20738 : OAI22_X1 port map( A1 => n25257, A2 => n25525, B1 => n21265, B2 => 
                           n20525, ZN => n6720);
   U20739 : OAI22_X1 port map( A1 => n25257, A2 => n25528, B1 => n21265, B2 => 
                           n20524, ZN => n6721);
   U20740 : OAI22_X1 port map( A1 => n25257, A2 => n25531, B1 => n25242, B2 => 
                           n20523, ZN => n6722);
   U20741 : OAI22_X1 port map( A1 => n25257, A2 => n25551, B1 => n21265, B2 => 
                           n20522, ZN => n6723);
   U20742 : OAI22_X1 port map( A1 => n25087, A2 => n25526, B1 => n21279, B2 => 
                           n20521, ZN => n6080);
   U20743 : OAI22_X1 port map( A1 => n25087, A2 => n25529, B1 => n21279, B2 => 
                           n20520, ZN => n6081);
   U20744 : OAI22_X1 port map( A1 => n25087, A2 => n25532, B1 => n25072, B2 => 
                           n20519, ZN => n6082);
   U20745 : OAI22_X1 port map( A1 => n25087, A2 => n25552, B1 => n21279, B2 => 
                           n20518, ZN => n6083);
   U20746 : OAI22_X1 port map( A1 => n25019, A2 => n25526, B1 => n21284, B2 => 
                           n20517, ZN => n5824);
   U20747 : OAI22_X1 port map( A1 => n25019, A2 => n25529, B1 => n21284, B2 => 
                           n20516, ZN => n5825);
   U20748 : OAI22_X1 port map( A1 => n25019, A2 => n25532, B1 => n25004, B2 => 
                           n20515, ZN => n5826);
   U20749 : OAI22_X1 port map( A1 => n25019, A2 => n25552, B1 => n21284, B2 => 
                           n20514, ZN => n5827);
   U20750 : OAI22_X1 port map( A1 => n24917, A2 => n25527, B1 => n21291, B2 => 
                           n20513, ZN => n5440);
   U20751 : OAI22_X1 port map( A1 => n24917, A2 => n25530, B1 => n21291, B2 => 
                           n20512, ZN => n5441);
   U20752 : OAI22_X1 port map( A1 => n24917, A2 => n25533, B1 => n24902, B2 => 
                           n20511, ZN => n5442);
   U20753 : OAI22_X1 port map( A1 => n24917, A2 => n25553, B1 => n21291, B2 => 
                           n20510, ZN => n5443);
   U20754 : OAI22_X1 port map( A1 => n24849, A2 => n25527, B1 => n21295, B2 => 
                           n20509, ZN => n5184);
   U20755 : OAI22_X1 port map( A1 => n24849, A2 => n25530, B1 => n21295, B2 => 
                           n20508, ZN => n5185);
   U20756 : OAI22_X1 port map( A1 => n24849, A2 => n25533, B1 => n24834, B2 => 
                           n20507, ZN => n5186);
   U20757 : OAI22_X1 port map( A1 => n24849, A2 => n25553, B1 => n21295, B2 => 
                           n20506, ZN => n5187);
   U20758 : OAI22_X1 port map( A1 => n25070, A2 => n25526, B1 => n21281, B2 => 
                           n20265, ZN => n6016);
   U20759 : OAI22_X1 port map( A1 => n25070, A2 => n25529, B1 => n21281, B2 => 
                           n20264, ZN => n6017);
   U20760 : OAI22_X1 port map( A1 => n25070, A2 => n25532, B1 => n25055, B2 => 
                           n20263, ZN => n6018);
   U20761 : OAI22_X1 port map( A1 => n25070, A2 => n25552, B1 => n21281, B2 => 
                           n20262, ZN => n6019);
   U20762 : OAI22_X1 port map( A1 => n25325, A2 => n25525, B1 => n21257, B2 => 
                           n20261, ZN => n6976);
   U20763 : OAI22_X1 port map( A1 => n25325, A2 => n25528, B1 => n21257, B2 => 
                           n20260, ZN => n6977);
   U20764 : OAI22_X1 port map( A1 => n25325, A2 => n25531, B1 => n25310, B2 => 
                           n20259, ZN => n6978);
   U20765 : OAI22_X1 port map( A1 => n25325, A2 => n25551, B1 => n21257, B2 => 
                           n20258, ZN => n6979);
   U20766 : OAI22_X1 port map( A1 => n25206, A2 => n25525, B1 => n21272, B2 => 
                           n20257, ZN => n6528);
   U20767 : OAI22_X1 port map( A1 => n25206, A2 => n25528, B1 => n21272, B2 => 
                           n20256, ZN => n6529);
   U20768 : OAI22_X1 port map( A1 => n25206, A2 => n25531, B1 => n25191, B2 => 
                           n20255, ZN => n6530);
   U20769 : OAI22_X1 port map( A1 => n25206, A2 => n25551, B1 => n21272, B2 => 
                           n20254, ZN => n6531);
   U20770 : OAI22_X1 port map( A1 => n25308, A2 => n25525, B1 => n21259, B2 => 
                           n20253, ZN => n6912);
   U20771 : OAI22_X1 port map( A1 => n25308, A2 => n25528, B1 => n21259, B2 => 
                           n20252, ZN => n6913);
   U20772 : OAI22_X1 port map( A1 => n25308, A2 => n25531, B1 => n25293, B2 => 
                           n20251, ZN => n6914);
   U20773 : OAI22_X1 port map( A1 => n25308, A2 => n25551, B1 => n21259, B2 => 
                           n20250, ZN => n6915);
   U20774 : OAI22_X1 port map( A1 => n24951, A2 => n25527, B1 => n21288, B2 => 
                           n20152, ZN => n5568);
   U20775 : OAI22_X1 port map( A1 => n24951, A2 => n25530, B1 => n21288, B2 => 
                           n20151, ZN => n5569);
   U20776 : OAI22_X1 port map( A1 => n24951, A2 => n25533, B1 => n24936, B2 => 
                           n20150, ZN => n5570);
   U20777 : OAI22_X1 port map( A1 => n24951, A2 => n25553, B1 => n21288, B2 => 
                           n20149, ZN => n5571);
   U20778 : OAI22_X1 port map( A1 => n24883, A2 => n25527, B1 => n21293, B2 => 
                           n20148, ZN => n5312);
   U20779 : OAI22_X1 port map( A1 => n24883, A2 => n25530, B1 => n21293, B2 => 
                           n20147, ZN => n5313);
   U20780 : OAI22_X1 port map( A1 => n24883, A2 => n25533, B1 => n24868, B2 => 
                           n20146, ZN => n5314);
   U20781 : OAI22_X1 port map( A1 => n24883, A2 => n25553, B1 => n21293, B2 => 
                           n20145, ZN => n5315);
   U20782 : OAI22_X1 port map( A1 => n25291, A2 => n25525, B1 => n21261, B2 => 
                           n19335, ZN => n6848);
   U20783 : OAI22_X1 port map( A1 => n25291, A2 => n25528, B1 => n21261, B2 => 
                           n19334, ZN => n6849);
   U20784 : OAI22_X1 port map( A1 => n25291, A2 => n25531, B1 => n25276, B2 => 
                           n19333, ZN => n6850);
   U20785 : OAI22_X1 port map( A1 => n25291, A2 => n25551, B1 => n21261, B2 => 
                           n19332, ZN => n6851);
   U20786 : OAI22_X1 port map( A1 => n25549, A2 => n25525, B1 => n21189, B2 => 
                           n19271, ZN => n7104);
   U20787 : OAI22_X1 port map( A1 => n25549, A2 => n25528, B1 => n21189, B2 => 
                           n19270, ZN => n7105);
   U20788 : OAI22_X1 port map( A1 => n25549, A2 => n25531, B1 => n25534, B2 => 
                           n19269, ZN => n7106);
   U20789 : OAI22_X1 port map( A1 => n25549, A2 => n25551, B1 => n21189, B2 => 
                           n19268, ZN => n7107);
   U20790 : NOR3_X1 port map( A1 => n19203, A2 => n19199, A3 => n19200, ZN => 
                           n23739);
   U20791 : BUF_X1 port map( A => n21298, Z => n24802);
   U20792 : BUF_X1 port map( A => n21298, Z => n24801);
   U20793 : BUF_X1 port map( A => n21298, Z => n24799);
   U20794 : BUF_X1 port map( A => n21298, Z => n24798);
   U20795 : BUF_X1 port map( A => n21298, Z => n24800);
   U20796 : BUF_X1 port map( A => n22608, Z => n24409);
   U20797 : BUF_X1 port map( A => n22608, Z => n24412);
   U20798 : BUF_X1 port map( A => n22608, Z => n24411);
   U20799 : BUF_X1 port map( A => n22608, Z => n24410);
   U20800 : BUF_X1 port map( A => n21297, Z => n24805);
   U20801 : BUF_X1 port map( A => n21297, Z => n24806);
   U20802 : BUF_X1 port map( A => n21297, Z => n24807);
   U20803 : BUF_X1 port map( A => n21297, Z => n24808);
   U20804 : NAND2_X1 port map( A1 => n22542, A2 => n22554, ZN => n21339);
   U20805 : NAND2_X1 port map( A1 => n22542, A2 => n22553, ZN => n21340);
   U20806 : NAND2_X1 port map( A1 => n23748, A2 => n23744, ZN => n22610);
   U20807 : NAND2_X1 port map( A1 => n23742, A2 => n23747, ZN => n22584);
   U20808 : NOR2_X1 port map( A1 => n19202, A2 => n19201, ZN => n23755);
   U20809 : BUF_X1 port map( A => n21252, Z => n25346);
   U20810 : BUF_X1 port map( A => n21251, Z => n25349);
   U20811 : BUF_X1 port map( A => n21250, Z => n25352);
   U20812 : BUF_X1 port map( A => n21249, Z => n25355);
   U20813 : BUF_X1 port map( A => n21248, Z => n25358);
   U20814 : BUF_X1 port map( A => n21247, Z => n25361);
   U20815 : BUF_X1 port map( A => n21246, Z => n25364);
   U20816 : BUF_X1 port map( A => n21245, Z => n25367);
   U20817 : BUF_X1 port map( A => n21244, Z => n25370);
   U20818 : BUF_X1 port map( A => n21243, Z => n25373);
   U20819 : BUF_X1 port map( A => n21242, Z => n25376);
   U20820 : BUF_X1 port map( A => n21241, Z => n25379);
   U20821 : BUF_X1 port map( A => n21240, Z => n25382);
   U20822 : BUF_X1 port map( A => n21239, Z => n25385);
   U20823 : BUF_X1 port map( A => n21238, Z => n25388);
   U20824 : BUF_X1 port map( A => n21237, Z => n25391);
   U20825 : BUF_X1 port map( A => n21236, Z => n25394);
   U20826 : BUF_X1 port map( A => n21235, Z => n25397);
   U20827 : BUF_X1 port map( A => n21234, Z => n25400);
   U20828 : BUF_X1 port map( A => n21233, Z => n25403);
   U20829 : BUF_X1 port map( A => n21232, Z => n25406);
   U20830 : BUF_X1 port map( A => n21231, Z => n25409);
   U20831 : BUF_X1 port map( A => n21230, Z => n25412);
   U20832 : BUF_X1 port map( A => n21229, Z => n25415);
   U20833 : BUF_X1 port map( A => n21228, Z => n25418);
   U20834 : BUF_X1 port map( A => n21227, Z => n25421);
   U20835 : BUF_X1 port map( A => n21226, Z => n25424);
   U20836 : BUF_X1 port map( A => n21225, Z => n25427);
   U20837 : BUF_X1 port map( A => n21224, Z => n25430);
   U20838 : BUF_X1 port map( A => n21223, Z => n25433);
   U20839 : BUF_X1 port map( A => n21222, Z => n25436);
   U20840 : BUF_X1 port map( A => n21221, Z => n25439);
   U20841 : BUF_X1 port map( A => n21220, Z => n25442);
   U20842 : BUF_X1 port map( A => n21219, Z => n25445);
   U20843 : BUF_X1 port map( A => n21218, Z => n25448);
   U20844 : BUF_X1 port map( A => n21217, Z => n25451);
   U20845 : BUF_X1 port map( A => n21216, Z => n25454);
   U20846 : BUF_X1 port map( A => n21215, Z => n25457);
   U20847 : BUF_X1 port map( A => n21214, Z => n25460);
   U20848 : BUF_X1 port map( A => n21213, Z => n25463);
   U20849 : BUF_X1 port map( A => n21212, Z => n25466);
   U20850 : BUF_X1 port map( A => n21211, Z => n25469);
   U20851 : BUF_X1 port map( A => n21210, Z => n25472);
   U20852 : BUF_X1 port map( A => n21209, Z => n25475);
   U20853 : BUF_X1 port map( A => n21208, Z => n25478);
   U20854 : BUF_X1 port map( A => n21207, Z => n25481);
   U20855 : BUF_X1 port map( A => n21206, Z => n25484);
   U20856 : BUF_X1 port map( A => n21205, Z => n25487);
   U20857 : BUF_X1 port map( A => n21204, Z => n25490);
   U20858 : BUF_X1 port map( A => n21203, Z => n25493);
   U20859 : BUF_X1 port map( A => n21202, Z => n25496);
   U20860 : BUF_X1 port map( A => n21201, Z => n25499);
   U20861 : BUF_X1 port map( A => n21200, Z => n25502);
   U20862 : BUF_X1 port map( A => n21199, Z => n25505);
   U20863 : BUF_X1 port map( A => n21198, Z => n25508);
   U20864 : BUF_X1 port map( A => n21197, Z => n25511);
   U20865 : BUF_X1 port map( A => n21196, Z => n25514);
   U20866 : BUF_X1 port map( A => n21195, Z => n25517);
   U20867 : BUF_X1 port map( A => n21194, Z => n25520);
   U20868 : BUF_X1 port map( A => n21193, Z => n25523);
   U20869 : BUF_X1 port map( A => n21192, Z => n25526);
   U20870 : BUF_X1 port map( A => n21191, Z => n25529);
   U20871 : BUF_X1 port map( A => n21190, Z => n25532);
   U20872 : BUF_X1 port map( A => n21188, Z => n25552);
   U20873 : BUF_X1 port map( A => n21252, Z => n25345);
   U20874 : BUF_X1 port map( A => n21251, Z => n25348);
   U20875 : BUF_X1 port map( A => n21250, Z => n25351);
   U20876 : BUF_X1 port map( A => n21249, Z => n25354);
   U20877 : BUF_X1 port map( A => n21248, Z => n25357);
   U20878 : BUF_X1 port map( A => n21247, Z => n25360);
   U20879 : BUF_X1 port map( A => n21246, Z => n25363);
   U20880 : BUF_X1 port map( A => n21245, Z => n25366);
   U20881 : BUF_X1 port map( A => n21244, Z => n25369);
   U20882 : BUF_X1 port map( A => n21243, Z => n25372);
   U20883 : BUF_X1 port map( A => n21242, Z => n25375);
   U20884 : BUF_X1 port map( A => n21241, Z => n25378);
   U20885 : BUF_X1 port map( A => n21240, Z => n25381);
   U20886 : BUF_X1 port map( A => n21239, Z => n25384);
   U20887 : BUF_X1 port map( A => n21238, Z => n25387);
   U20888 : BUF_X1 port map( A => n21237, Z => n25390);
   U20889 : BUF_X1 port map( A => n21236, Z => n25393);
   U20890 : BUF_X1 port map( A => n21235, Z => n25396);
   U20891 : BUF_X1 port map( A => n21234, Z => n25399);
   U20892 : BUF_X1 port map( A => n21233, Z => n25402);
   U20893 : BUF_X1 port map( A => n21232, Z => n25405);
   U20894 : BUF_X1 port map( A => n21231, Z => n25408);
   U20895 : BUF_X1 port map( A => n21230, Z => n25411);
   U20896 : BUF_X1 port map( A => n21229, Z => n25414);
   U20897 : BUF_X1 port map( A => n21228, Z => n25417);
   U20898 : BUF_X1 port map( A => n21227, Z => n25420);
   U20899 : BUF_X1 port map( A => n21226, Z => n25423);
   U20900 : BUF_X1 port map( A => n21225, Z => n25426);
   U20901 : BUF_X1 port map( A => n21224, Z => n25429);
   U20902 : BUF_X1 port map( A => n21223, Z => n25432);
   U20903 : BUF_X1 port map( A => n21222, Z => n25435);
   U20904 : BUF_X1 port map( A => n21221, Z => n25438);
   U20905 : BUF_X1 port map( A => n21220, Z => n25441);
   U20906 : BUF_X1 port map( A => n21219, Z => n25444);
   U20907 : BUF_X1 port map( A => n21218, Z => n25447);
   U20908 : BUF_X1 port map( A => n21217, Z => n25450);
   U20909 : BUF_X1 port map( A => n21216, Z => n25453);
   U20910 : BUF_X1 port map( A => n21215, Z => n25456);
   U20911 : BUF_X1 port map( A => n21214, Z => n25459);
   U20912 : BUF_X1 port map( A => n21213, Z => n25462);
   U20913 : BUF_X1 port map( A => n21212, Z => n25465);
   U20914 : BUF_X1 port map( A => n21211, Z => n25468);
   U20915 : BUF_X1 port map( A => n21210, Z => n25471);
   U20916 : BUF_X1 port map( A => n21209, Z => n25474);
   U20917 : BUF_X1 port map( A => n21208, Z => n25477);
   U20918 : BUF_X1 port map( A => n21207, Z => n25480);
   U20919 : BUF_X1 port map( A => n21206, Z => n25483);
   U20920 : BUF_X1 port map( A => n21205, Z => n25486);
   U20921 : BUF_X1 port map( A => n21204, Z => n25489);
   U20922 : BUF_X1 port map( A => n21203, Z => n25492);
   U20923 : BUF_X1 port map( A => n21202, Z => n25495);
   U20924 : BUF_X1 port map( A => n21201, Z => n25498);
   U20925 : BUF_X1 port map( A => n21200, Z => n25501);
   U20926 : BUF_X1 port map( A => n21199, Z => n25504);
   U20927 : BUF_X1 port map( A => n21198, Z => n25507);
   U20928 : BUF_X1 port map( A => n21197, Z => n25510);
   U20929 : BUF_X1 port map( A => n21196, Z => n25513);
   U20930 : BUF_X1 port map( A => n21195, Z => n25516);
   U20931 : BUF_X1 port map( A => n21194, Z => n25519);
   U20932 : BUF_X1 port map( A => n21193, Z => n25522);
   U20933 : BUF_X1 port map( A => n21192, Z => n25525);
   U20934 : BUF_X1 port map( A => n21191, Z => n25528);
   U20935 : BUF_X1 port map( A => n21190, Z => n25531);
   U20936 : BUF_X1 port map( A => n21188, Z => n25551);
   U20937 : NAND2_X1 port map( A1 => n22554, A2 => n22538, ZN => n21334);
   U20938 : NAND2_X1 port map( A1 => n22539, A2 => n22538, ZN => n21310);
   U20939 : NAND2_X1 port map( A1 => n22537, A2 => n22538, ZN => n21311);
   U20940 : NAND2_X1 port map( A1 => n22546, A2 => n22538, ZN => n21320);
   U20941 : NAND2_X1 port map( A1 => n22545, A2 => n22538, ZN => n21321);
   U20942 : NAND2_X1 port map( A1 => n23756, A2 => n23757, ZN => n22593);
   U20943 : NAND2_X1 port map( A1 => n23754, A2 => n23757, ZN => n22595);
   U20944 : NAND2_X1 port map( A1 => n23754, A2 => n23758, ZN => n22596);
   U20945 : NAND2_X1 port map( A1 => n23756, A2 => n23755, ZN => n22597);
   U20946 : NAND2_X1 port map( A1 => n22538, A2 => n22553, ZN => n21335);
   U20947 : NAND2_X1 port map( A1 => n23740, A2 => n23741, ZN => n22569);
   U20948 : NAND2_X1 port map( A1 => n23747, A2 => n23738, ZN => n22579);
   U20949 : NAND2_X1 port map( A1 => n22558, A2 => n22540, ZN => n21344);
   U20950 : NAND2_X1 port map( A1 => n22557, A2 => n22540, ZN => n21345);
   U20951 : NAND2_X1 port map( A1 => n22558, A2 => n22543, ZN => n21349);
   U20952 : NAND2_X1 port map( A1 => n22557, A2 => n22543, ZN => n21350);
   U20953 : NAND2_X1 port map( A1 => n23740, A2 => n23745, ZN => n22611);
   U20954 : NAND2_X1 port map( A1 => n23740, A2 => n23742, ZN => n22605);
   U20955 : NAND2_X1 port map( A1 => n23737, A2 => n23745, ZN => n22606);
   U20956 : NAND2_X1 port map( A1 => n22539, A2 => n22542, ZN => n21315);
   U20957 : NAND2_X1 port map( A1 => n22537, A2 => n22542, ZN => n21316);
   U20958 : NAND2_X1 port map( A1 => n22546, A2 => n22542, ZN => n21325);
   U20959 : NAND2_X1 port map( A1 => n22545, A2 => n22542, ZN => n21326);
   U20960 : BUF_X1 port map( A => n22608, Z => n24408);
   U20961 : BUF_X1 port map( A => n21297, Z => n24804);
   U20962 : BUF_X1 port map( A => n21192, Z => n25527);
   U20963 : BUF_X1 port map( A => n21191, Z => n25530);
   U20964 : BUF_X1 port map( A => n21190, Z => n25533);
   U20965 : BUF_X1 port map( A => n21188, Z => n25553);
   U20966 : BUF_X1 port map( A => n21252, Z => n25347);
   U20967 : BUF_X1 port map( A => n21251, Z => n25350);
   U20968 : BUF_X1 port map( A => n21250, Z => n25353);
   U20969 : BUF_X1 port map( A => n21249, Z => n25356);
   U20970 : BUF_X1 port map( A => n21248, Z => n25359);
   U20971 : BUF_X1 port map( A => n21247, Z => n25362);
   U20972 : BUF_X1 port map( A => n21246, Z => n25365);
   U20973 : BUF_X1 port map( A => n21245, Z => n25368);
   U20974 : BUF_X1 port map( A => n21244, Z => n25371);
   U20975 : BUF_X1 port map( A => n21243, Z => n25374);
   U20976 : BUF_X1 port map( A => n21242, Z => n25377);
   U20977 : BUF_X1 port map( A => n21241, Z => n25380);
   U20978 : BUF_X1 port map( A => n21240, Z => n25383);
   U20979 : BUF_X1 port map( A => n21239, Z => n25386);
   U20980 : BUF_X1 port map( A => n21238, Z => n25389);
   U20981 : BUF_X1 port map( A => n21237, Z => n25392);
   U20982 : BUF_X1 port map( A => n21236, Z => n25395);
   U20983 : BUF_X1 port map( A => n21235, Z => n25398);
   U20984 : BUF_X1 port map( A => n21234, Z => n25401);
   U20985 : BUF_X1 port map( A => n21233, Z => n25404);
   U20986 : BUF_X1 port map( A => n21232, Z => n25407);
   U20987 : BUF_X1 port map( A => n21231, Z => n25410);
   U20988 : BUF_X1 port map( A => n21230, Z => n25413);
   U20989 : BUF_X1 port map( A => n21229, Z => n25416);
   U20990 : BUF_X1 port map( A => n21228, Z => n25419);
   U20991 : BUF_X1 port map( A => n21227, Z => n25422);
   U20992 : BUF_X1 port map( A => n21226, Z => n25425);
   U20993 : BUF_X1 port map( A => n21225, Z => n25428);
   U20994 : BUF_X1 port map( A => n21224, Z => n25431);
   U20995 : BUF_X1 port map( A => n21223, Z => n25434);
   U20996 : BUF_X1 port map( A => n21222, Z => n25437);
   U20997 : BUF_X1 port map( A => n21221, Z => n25440);
   U20998 : BUF_X1 port map( A => n21220, Z => n25443);
   U20999 : BUF_X1 port map( A => n21219, Z => n25446);
   U21000 : BUF_X1 port map( A => n21218, Z => n25449);
   U21001 : BUF_X1 port map( A => n21217, Z => n25452);
   U21002 : BUF_X1 port map( A => n21216, Z => n25455);
   U21003 : BUF_X1 port map( A => n21215, Z => n25458);
   U21004 : BUF_X1 port map( A => n21214, Z => n25461);
   U21005 : BUF_X1 port map( A => n21213, Z => n25464);
   U21006 : BUF_X1 port map( A => n21212, Z => n25467);
   U21007 : BUF_X1 port map( A => n21211, Z => n25470);
   U21008 : BUF_X1 port map( A => n21210, Z => n25473);
   U21009 : BUF_X1 port map( A => n21209, Z => n25476);
   U21010 : BUF_X1 port map( A => n21208, Z => n25479);
   U21011 : BUF_X1 port map( A => n21207, Z => n25482);
   U21012 : BUF_X1 port map( A => n21206, Z => n25485);
   U21013 : BUF_X1 port map( A => n21205, Z => n25488);
   U21014 : BUF_X1 port map( A => n21204, Z => n25491);
   U21015 : BUF_X1 port map( A => n21203, Z => n25494);
   U21016 : BUF_X1 port map( A => n21202, Z => n25497);
   U21017 : BUF_X1 port map( A => n21201, Z => n25500);
   U21018 : BUF_X1 port map( A => n21200, Z => n25503);
   U21019 : BUF_X1 port map( A => n21199, Z => n25506);
   U21020 : BUF_X1 port map( A => n21198, Z => n25509);
   U21021 : BUF_X1 port map( A => n21197, Z => n25512);
   U21022 : BUF_X1 port map( A => n21196, Z => n25515);
   U21023 : BUF_X1 port map( A => n21195, Z => n25518);
   U21024 : BUF_X1 port map( A => n21194, Z => n25521);
   U21025 : BUF_X1 port map( A => n21193, Z => n25524);
   U21026 : OAI21_X1 port map( B1 => n21268, B2 => n21289, A => n25564, ZN => 
                           n21296);
   U21027 : NAND2_X1 port map( A1 => n23745, A2 => n23744, ZN => n22573);
   U21028 : AND2_X1 port map( A1 => n23758, A2 => n23761, ZN => n23740);
   U21029 : NAND2_X1 port map( A1 => n23742, A2 => n23737, ZN => n22568);
   U21030 : AND2_X1 port map( A1 => n23761, A2 => n23757, ZN => n23744);
   U21031 : AND2_X1 port map( A1 => n23755, A2 => n23761, ZN => n23737);
   U21032 : AND2_X1 port map( A1 => n23759, A2 => n23761, ZN => n23747);
   U21033 : NAND2_X1 port map( A1 => n23737, A2 => n23748, ZN => n22583);
   U21034 : NAND2_X1 port map( A1 => n23740, A2 => n23748, ZN => n22578);
   U21035 : AND2_X1 port map( A1 => n23760, A2 => n19203, ZN => n23754);
   U21036 : OR2_X1 port map( A1 => n24413, A2 => n19190, ZN => n22598);
   U21037 : NAND2_X1 port map( A1 => n23754, A2 => n23759, ZN => n22601);
   U21038 : NAND2_X1 port map( A1 => n23756, A2 => n23758, ZN => n22599);
   U21039 : NAND2_X1 port map( A1 => n23756, A2 => n23759, ZN => n22600);
   U21040 : AND2_X1 port map( A1 => n23748, A2 => n23747, ZN => n22586);
   U21041 : AND2_X1 port map( A1 => n23745, A2 => n23747, ZN => n22588);
   U21042 : AND2_X1 port map( A1 => n23742, A2 => n23744, ZN => n22582);
   U21043 : AND2_X1 port map( A1 => n22543, A2 => n22554, ZN => n21336);
   U21044 : AND2_X1 port map( A1 => n22543, A2 => n22553, ZN => n21337);
   U21045 : AND2_X1 port map( A1 => n22558, A2 => n22542, ZN => n21346);
   U21046 : AND2_X1 port map( A1 => n22557, A2 => n22542, ZN => n21347);
   U21047 : AND2_X1 port map( A1 => n22558, A2 => n22538, ZN => n21341);
   U21048 : AND2_X1 port map( A1 => n22557, A2 => n22538, ZN => n21342);
   U21049 : AND2_X1 port map( A1 => n23738, A2 => n23744, ZN => n22587);
   U21050 : AND2_X1 port map( A1 => n23741, A2 => n23744, ZN => n22576);
   U21051 : AND2_X1 port map( A1 => n23741, A2 => n23747, ZN => n22581);
   U21052 : AND2_X1 port map( A1 => n23741, A2 => n23737, ZN => n22607);
   U21053 : AND2_X1 port map( A1 => n24803, A2 => n19190, ZN => n21302);
   U21054 : AND2_X1 port map( A1 => n22540, A2 => n22553, ZN => n21332);
   U21055 : AND2_X1 port map( A1 => n22539, A2 => n22543, ZN => n21312);
   U21056 : AND2_X1 port map( A1 => n22537, A2 => n22543, ZN => n21313);
   U21057 : AND2_X1 port map( A1 => n22546, A2 => n22543, ZN => n21322);
   U21058 : AND2_X1 port map( A1 => n22545, A2 => n22543, ZN => n21323);
   U21059 : AND2_X1 port map( A1 => n22540, A2 => n22554, ZN => n21331);
   U21060 : AND2_X1 port map( A1 => n23737, A2 => n23738, ZN => n22572);
   U21061 : AND2_X1 port map( A1 => n23740, A2 => n23738, ZN => n22603);
   U21062 : AND2_X1 port map( A1 => n22539, A2 => n22540, ZN => n21307);
   U21063 : AND2_X1 port map( A1 => n22537, A2 => n22540, ZN => n21308);
   U21064 : AND2_X1 port map( A1 => n22546, A2 => n22540, ZN => n21317);
   U21065 : AND2_X1 port map( A1 => n22545, A2 => n22540, ZN => n21318);
   U21066 : AND3_X1 port map( A1 => n19200, A2 => n19199, A3 => n23761, ZN => 
                           n23760);
   U21067 : BUF_X1 port map( A => n21267, Z => n25225);
   U21068 : OAI21_X1 port map( B1 => n21253, B2 => n21268, A => n25564, ZN => 
                           n21267);
   U21069 : BUF_X1 port map( A => n21265, Z => n25242);
   U21070 : OAI21_X1 port map( B1 => n21253, B2 => n21266, A => n25564, ZN => 
                           n21265);
   U21071 : BUF_X1 port map( A => n21257, Z => n25310);
   U21072 : OAI21_X1 port map( B1 => n21253, B2 => n21258, A => n25564, ZN => 
                           n21257);
   U21073 : BUF_X1 port map( A => n21259, Z => n25293);
   U21074 : OAI21_X1 port map( B1 => n21253, B2 => n21260, A => n25564, ZN => 
                           n21259);
   U21075 : BUF_X1 port map( A => n21255, Z => n25327);
   U21076 : OAI21_X1 port map( B1 => n21253, B2 => n21256, A => n25564, ZN => 
                           n21255);
   U21077 : BUF_X1 port map( A => n21263, Z => n25259);
   U21078 : OAI21_X1 port map( B1 => n21253, B2 => n21264, A => n25564, ZN => 
                           n21263);
   U21079 : BUF_X1 port map( A => n21261, Z => n25276);
   U21080 : OAI21_X1 port map( B1 => n21253, B2 => n21262, A => n25564, ZN => 
                           n21261);
   U21081 : BUF_X1 port map( A => n21285, Z => n24987);
   U21082 : OAI21_X1 port map( B1 => n21264, B2 => n21280, A => n25563, ZN => 
                           n21285);
   U21083 : BUF_X1 port map( A => n21270, Z => n25208);
   U21084 : OAI21_X1 port map( B1 => n21254, B2 => n21271, A => n25564, ZN => 
                           n21270);
   U21085 : BUF_X1 port map( A => n21275, Z => n25140);
   U21086 : OAI21_X1 port map( B1 => n21262, B2 => n21271, A => n25563, ZN => 
                           n21275);
   U21087 : BUF_X1 port map( A => n21292, Z => n24885);
   U21088 : OAI21_X1 port map( B1 => n21260, B2 => n21289, A => n25562, ZN => 
                           n21292);
   U21089 : BUF_X1 port map( A => n21279, Z => n25072);
   U21090 : OAI21_X1 port map( B1 => n21254, B2 => n21280, A => n25563, ZN => 
                           n21279);
   U21091 : BUF_X1 port map( A => n21284, Z => n25004);
   U21092 : OAI21_X1 port map( B1 => n21262, B2 => n21280, A => n25563, ZN => 
                           n21284);
   U21093 : BUF_X1 port map( A => n21291, Z => n24902);
   U21094 : OAI21_X1 port map( B1 => n21258, B2 => n21289, A => n25562, ZN => 
                           n21291);
   U21095 : BUF_X1 port map( A => n21295, Z => n24834);
   U21096 : OAI21_X1 port map( B1 => n21266, B2 => n21289, A => n25562, ZN => 
                           n21295);
   U21097 : BUF_X1 port map( A => n21281, Z => n25055);
   U21098 : OAI21_X1 port map( B1 => n21256, B2 => n21280, A => n25563, ZN => 
                           n21281);
   U21099 : BUF_X1 port map( A => n21272, Z => n25191);
   U21100 : OAI21_X1 port map( B1 => n21256, B2 => n21271, A => n25564, ZN => 
                           n21272);
   U21101 : BUF_X1 port map( A => n21273, Z => n25174);
   U21102 : OAI21_X1 port map( B1 => n21258, B2 => n21271, A => n25563, ZN => 
                           n21273);
   U21103 : BUF_X1 port map( A => n21278, Z => n25089);
   U21104 : OAI21_X1 port map( B1 => n21268, B2 => n21271, A => n25563, ZN => 
                           n21278);
   U21105 : BUF_X1 port map( A => n21282, Z => n25038);
   U21106 : OAI21_X1 port map( B1 => n21258, B2 => n21280, A => n25563, ZN => 
                           n21282);
   U21107 : BUF_X1 port map( A => n21283, Z => n25021);
   U21108 : OAI21_X1 port map( B1 => n21260, B2 => n21280, A => n25563, ZN => 
                           n21283);
   U21109 : BUF_X1 port map( A => n21294, Z => n24851);
   U21110 : OAI21_X1 port map( B1 => n21264, B2 => n21289, A => n25562, ZN => 
                           n21294);
   U21111 : BUF_X1 port map( A => n21293, Z => n24868);
   U21112 : OAI21_X1 port map( B1 => n21262, B2 => n21289, A => n25562, ZN => 
                           n21293);
   U21113 : BUF_X1 port map( A => n21290, Z => n24919);
   U21114 : OAI21_X1 port map( B1 => n21256, B2 => n21289, A => n25562, ZN => 
                           n21290);
   U21115 : BUF_X1 port map( A => n21288, Z => n24936);
   U21116 : OAI21_X1 port map( B1 => n21254, B2 => n21289, A => n25562, ZN => 
                           n21288);
   U21117 : BUF_X1 port map( A => n21287, Z => n24953);
   U21118 : OAI21_X1 port map( B1 => n21268, B2 => n21280, A => n25562, ZN => 
                           n21287);
   U21119 : BUF_X1 port map( A => n21286, Z => n24970);
   U21120 : OAI21_X1 port map( B1 => n21266, B2 => n21280, A => n25563, ZN => 
                           n21286);
   U21121 : BUF_X1 port map( A => n21277, Z => n25106);
   U21122 : OAI21_X1 port map( B1 => n21266, B2 => n21271, A => n25563, ZN => 
                           n21277);
   U21123 : BUF_X1 port map( A => n21276, Z => n25123);
   U21124 : OAI21_X1 port map( B1 => n21264, B2 => n21271, A => n25563, ZN => 
                           n21276);
   U21125 : BUF_X1 port map( A => n21274, Z => n25157);
   U21126 : OAI21_X1 port map( B1 => n21260, B2 => n21271, A => n25563, ZN => 
                           n21274);
   U21127 : AOI222_X1 port map( A1 => n24513, A2 => n24008, B1 => n24507, B2 =>
                           n8629, C1 => n24501, C2 => n8501, ZN => n23019);
   U21128 : AOI222_X1 port map( A1 => n24513, A2 => n24009, B1 => n24507, B2 =>
                           n8628, C1 => n24501, C2 => n8500, ZN => n23001);
   U21129 : AOI222_X1 port map( A1 => n24513, A2 => n24010, B1 => n24507, B2 =>
                           n8627, C1 => n24501, C2 => n8499, ZN => n22983);
   U21130 : AOI222_X1 port map( A1 => n24513, A2 => n24011, B1 => n24507, B2 =>
                           n8626, C1 => n24501, C2 => n8498, ZN => n22965);
   U21131 : AOI222_X1 port map( A1 => n24513, A2 => n24012, B1 => n24507, B2 =>
                           n8625, C1 => n24501, C2 => n8497, ZN => n22947);
   U21132 : AOI222_X1 port map( A1 => n24513, A2 => n24013, B1 => n24507, B2 =>
                           n8624, C1 => n24501, C2 => n8496, ZN => n22929);
   U21133 : AOI222_X1 port map( A1 => n24513, A2 => n24014, B1 => n24507, B2 =>
                           n8623, C1 => n24501, C2 => n8495, ZN => n22911);
   U21134 : AOI222_X1 port map( A1 => n24513, A2 => n24015, B1 => n24507, B2 =>
                           n8622, C1 => n24501, C2 => n8494, ZN => n22893);
   U21135 : AOI222_X1 port map( A1 => n24514, A2 => n24016, B1 => n24508, B2 =>
                           n8621, C1 => n24502, C2 => n8493, ZN => n22875);
   U21136 : AOI222_X1 port map( A1 => n24514, A2 => n24017, B1 => n24508, B2 =>
                           n8620, C1 => n24502, C2 => n8492, ZN => n22857);
   U21137 : AOI222_X1 port map( A1 => n24514, A2 => n24018, B1 => n24508, B2 =>
                           n8619, C1 => n24502, C2 => n8491, ZN => n22839);
   U21138 : AOI222_X1 port map( A1 => n24514, A2 => n24019, B1 => n24508, B2 =>
                           n8618, C1 => n24502, C2 => n8490, ZN => n22821);
   U21139 : AOI222_X1 port map( A1 => n24514, A2 => n24020, B1 => n24508, B2 =>
                           n8617, C1 => n24502, C2 => n8489, ZN => n22803);
   U21140 : AOI222_X1 port map( A1 => n24514, A2 => n24021, B1 => n24508, B2 =>
                           n8616, C1 => n24502, C2 => n8488, ZN => n22785);
   U21141 : AOI222_X1 port map( A1 => n24514, A2 => n24022, B1 => n24508, B2 =>
                           n8615, C1 => n24502, C2 => n8487, ZN => n22767);
   U21142 : AOI222_X1 port map( A1 => n24514, A2 => n24023, B1 => n24508, B2 =>
                           n8614, C1 => n24502, C2 => n8486, ZN => n22749);
   U21143 : AOI222_X1 port map( A1 => n24514, A2 => n24024, B1 => n24508, B2 =>
                           n8613, C1 => n24502, C2 => n8485, ZN => n22731);
   U21144 : AOI222_X1 port map( A1 => n24514, A2 => n24025, B1 => n24508, B2 =>
                           n8612, C1 => n24502, C2 => n8484, ZN => n22713);
   U21145 : AOI222_X1 port map( A1 => n24514, A2 => n24026, B1 => n24508, B2 =>
                           n8611, C1 => n24502, C2 => n8483, ZN => n22695);
   U21146 : AOI222_X1 port map( A1 => n24514, A2 => n24027, B1 => n24508, B2 =>
                           n8610, C1 => n24502, C2 => n8482, ZN => n22677);
   U21147 : AOI222_X1 port map( A1 => n24515, A2 => n24028, B1 => n24509, B2 =>
                           n8609, C1 => n24503, C2 => n8481, ZN => n22659);
   U21148 : AOI222_X1 port map( A1 => n24515, A2 => n24029, B1 => n24509, B2 =>
                           n8608, C1 => n24503, C2 => n8480, ZN => n22641);
   U21149 : AOI222_X1 port map( A1 => n24515, A2 => n24030, B1 => n24509, B2 =>
                           n8607, C1 => n24503, C2 => n8479, ZN => n22623);
   U21150 : AOI222_X1 port map( A1 => n24515, A2 => n24031, B1 => n24509, B2 =>
                           n8606, C1 => n24503, C2 => n8478, ZN => n22585);
   U21151 : AOI222_X1 port map( A1 => n24510, A2 => n23968, B1 => n24504, B2 =>
                           n8669, C1 => n24498, C2 => n8541, ZN => n23749);
   U21152 : AOI222_X1 port map( A1 => n24510, A2 => n23969, B1 => n24504, B2 =>
                           n8668, C1 => n24498, C2 => n8540, ZN => n23721);
   U21153 : AOI222_X1 port map( A1 => n24510, A2 => n23970, B1 => n24504, B2 =>
                           n8667, C1 => n24498, C2 => n8539, ZN => n23703);
   U21154 : AOI222_X1 port map( A1 => n24510, A2 => n23971, B1 => n24504, B2 =>
                           n8666, C1 => n24498, C2 => n8538, ZN => n23685);
   U21155 : AOI222_X1 port map( A1 => n24510, A2 => n23972, B1 => n24504, B2 =>
                           n8665, C1 => n24498, C2 => n8537, ZN => n23667);
   U21156 : AOI222_X1 port map( A1 => n24510, A2 => n23973, B1 => n24504, B2 =>
                           n8664, C1 => n24498, C2 => n8536, ZN => n23649);
   U21157 : AOI222_X1 port map( A1 => n24510, A2 => n23974, B1 => n24504, B2 =>
                           n8663, C1 => n24498, C2 => n8535, ZN => n23631);
   U21158 : AOI222_X1 port map( A1 => n24510, A2 => n23975, B1 => n24504, B2 =>
                           n8662, C1 => n24498, C2 => n8534, ZN => n23613);
   U21159 : AOI222_X1 port map( A1 => n24510, A2 => n23976, B1 => n24504, B2 =>
                           n8661, C1 => n24498, C2 => n8533, ZN => n23595);
   U21160 : AOI222_X1 port map( A1 => n24510, A2 => n23977, B1 => n24504, B2 =>
                           n8660, C1 => n24498, C2 => n8532, ZN => n23577);
   U21161 : AOI222_X1 port map( A1 => n24510, A2 => n23978, B1 => n24504, B2 =>
                           n8659, C1 => n24498, C2 => n8531, ZN => n23559);
   U21162 : AOI222_X1 port map( A1 => n24510, A2 => n23979, B1 => n24504, B2 =>
                           n8658, C1 => n24498, C2 => n8530, ZN => n23541);
   U21163 : AOI222_X1 port map( A1 => n24511, A2 => n23980, B1 => n24505, B2 =>
                           n8657, C1 => n24499, C2 => n8529, ZN => n23523);
   U21164 : AOI222_X1 port map( A1 => n24511, A2 => n23981, B1 => n24505, B2 =>
                           n8656, C1 => n24499, C2 => n8528, ZN => n23505);
   U21165 : AOI222_X1 port map( A1 => n24511, A2 => n23982, B1 => n24505, B2 =>
                           n8655, C1 => n24499, C2 => n8527, ZN => n23487);
   U21166 : AOI222_X1 port map( A1 => n24511, A2 => n23983, B1 => n24505, B2 =>
                           n8654, C1 => n24499, C2 => n8526, ZN => n23469);
   U21167 : AOI222_X1 port map( A1 => n24511, A2 => n23984, B1 => n24505, B2 =>
                           n8653, C1 => n24499, C2 => n8525, ZN => n23451);
   U21168 : AOI222_X1 port map( A1 => n24511, A2 => n23985, B1 => n24505, B2 =>
                           n8652, C1 => n24499, C2 => n8524, ZN => n23433);
   U21169 : AOI222_X1 port map( A1 => n24511, A2 => n23986, B1 => n24505, B2 =>
                           n8651, C1 => n24499, C2 => n8523, ZN => n23415);
   U21170 : AOI222_X1 port map( A1 => n24511, A2 => n23987, B1 => n24505, B2 =>
                           n8650, C1 => n24499, C2 => n8522, ZN => n23397);
   U21171 : AOI222_X1 port map( A1 => n24511, A2 => n23988, B1 => n24505, B2 =>
                           n8649, C1 => n24499, C2 => n8521, ZN => n23379);
   U21172 : AOI222_X1 port map( A1 => n24511, A2 => n23989, B1 => n24505, B2 =>
                           n8648, C1 => n24499, C2 => n8520, ZN => n23361);
   U21173 : AOI222_X1 port map( A1 => n24511, A2 => n23990, B1 => n24505, B2 =>
                           n8647, C1 => n24499, C2 => n8519, ZN => n23343);
   U21174 : AOI222_X1 port map( A1 => n24511, A2 => n23991, B1 => n24505, B2 =>
                           n8646, C1 => n24499, C2 => n8518, ZN => n23325);
   U21175 : AOI222_X1 port map( A1 => n24512, A2 => n23992, B1 => n24506, B2 =>
                           n8645, C1 => n24500, C2 => n8517, ZN => n23307);
   U21176 : AOI222_X1 port map( A1 => n24512, A2 => n23993, B1 => n24506, B2 =>
                           n8644, C1 => n24500, C2 => n8516, ZN => n23289);
   U21177 : AOI222_X1 port map( A1 => n24512, A2 => n23994, B1 => n24506, B2 =>
                           n8643, C1 => n24500, C2 => n8515, ZN => n23271);
   U21178 : AOI222_X1 port map( A1 => n24512, A2 => n23995, B1 => n24506, B2 =>
                           n8642, C1 => n24500, C2 => n8514, ZN => n23253);
   U21179 : AOI222_X1 port map( A1 => n24512, A2 => n23996, B1 => n24506, B2 =>
                           n8641, C1 => n24500, C2 => n8513, ZN => n23235);
   U21180 : AOI222_X1 port map( A1 => n24512, A2 => n23997, B1 => n24506, B2 =>
                           n8640, C1 => n24500, C2 => n8512, ZN => n23217);
   U21181 : AOI222_X1 port map( A1 => n24512, A2 => n23998, B1 => n24506, B2 =>
                           n8639, C1 => n24500, C2 => n8511, ZN => n23199);
   U21182 : AOI222_X1 port map( A1 => n24512, A2 => n23999, B1 => n24506, B2 =>
                           n8638, C1 => n24500, C2 => n8510, ZN => n23181);
   U21183 : AOI222_X1 port map( A1 => n24512, A2 => n24000, B1 => n24506, B2 =>
                           n8637, C1 => n24500, C2 => n8509, ZN => n23163);
   U21184 : AOI222_X1 port map( A1 => n24512, A2 => n24001, B1 => n24506, B2 =>
                           n8636, C1 => n24500, C2 => n8508, ZN => n23145);
   U21185 : AOI222_X1 port map( A1 => n24512, A2 => n24002, B1 => n24506, B2 =>
                           n8635, C1 => n24500, C2 => n8507, ZN => n23127);
   U21186 : AOI222_X1 port map( A1 => n24512, A2 => n24003, B1 => n24506, B2 =>
                           n8634, C1 => n24500, C2 => n8506, ZN => n23109);
   U21187 : AOI222_X1 port map( A1 => n24513, A2 => n24004, B1 => n24507, B2 =>
                           n8633, C1 => n24501, C2 => n8505, ZN => n23091);
   U21188 : AOI222_X1 port map( A1 => n24513, A2 => n24005, B1 => n24507, B2 =>
                           n8632, C1 => n24501, C2 => n8504, ZN => n23073);
   U21189 : AOI222_X1 port map( A1 => n24513, A2 => n24006, B1 => n24507, B2 =>
                           n8631, C1 => n24501, C2 => n8503, ZN => n23055);
   U21190 : AOI222_X1 port map( A1 => n24513, A2 => n24007, B1 => n24507, B2 =>
                           n8630, C1 => n24501, C2 => n8502, ZN => n23037);
   U21191 : OAI222_X1 port map( A1 => n20285, A2 => n24459, B1 => n17290, B2 =>
                           n24453, C1 => n19355, C2 => n24447, ZN => n23020);
   U21192 : OAI222_X1 port map( A1 => n20284, A2 => n24459, B1 => n17287, B2 =>
                           n24453, C1 => n19354, C2 => n24447, ZN => n23002);
   U21193 : OAI222_X1 port map( A1 => n20283, A2 => n24459, B1 => n17284, B2 =>
                           n24453, C1 => n19353, C2 => n24447, ZN => n22984);
   U21194 : OAI222_X1 port map( A1 => n20282, A2 => n24459, B1 => n17281, B2 =>
                           n24453, C1 => n19352, C2 => n24447, ZN => n22966);
   U21195 : OAI222_X1 port map( A1 => n20281, A2 => n24459, B1 => n17278, B2 =>
                           n24453, C1 => n19351, C2 => n24447, ZN => n22948);
   U21196 : OAI222_X1 port map( A1 => n20280, A2 => n24459, B1 => n17275, B2 =>
                           n24453, C1 => n19350, C2 => n24447, ZN => n22930);
   U21197 : OAI222_X1 port map( A1 => n20279, A2 => n24459, B1 => n17272, B2 =>
                           n24453, C1 => n19349, C2 => n24447, ZN => n22912);
   U21198 : OAI222_X1 port map( A1 => n20278, A2 => n24459, B1 => n17269, B2 =>
                           n24453, C1 => n19348, C2 => n24447, ZN => n22894);
   U21199 : OAI222_X1 port map( A1 => n20277, A2 => n24460, B1 => n17266, B2 =>
                           n24454, C1 => n19347, C2 => n24448, ZN => n22876);
   U21200 : OAI222_X1 port map( A1 => n20276, A2 => n24460, B1 => n17263, B2 =>
                           n24454, C1 => n19346, C2 => n24448, ZN => n22858);
   U21201 : OAI222_X1 port map( A1 => n20275, A2 => n24460, B1 => n17260, B2 =>
                           n24454, C1 => n19345, C2 => n24448, ZN => n22840);
   U21202 : OAI222_X1 port map( A1 => n20274, A2 => n24460, B1 => n17257, B2 =>
                           n24454, C1 => n19344, C2 => n24448, ZN => n22822);
   U21203 : OAI222_X1 port map( A1 => n20273, A2 => n24460, B1 => n17254, B2 =>
                           n24454, C1 => n19343, C2 => n24448, ZN => n22804);
   U21204 : OAI222_X1 port map( A1 => n20272, A2 => n24460, B1 => n17251, B2 =>
                           n24454, C1 => n19342, C2 => n24448, ZN => n22786);
   U21205 : OAI222_X1 port map( A1 => n20271, A2 => n24460, B1 => n17248, B2 =>
                           n24454, C1 => n19341, C2 => n24448, ZN => n22768);
   U21206 : OAI222_X1 port map( A1 => n20270, A2 => n24460, B1 => n17245, B2 =>
                           n24454, C1 => n19340, C2 => n24448, ZN => n22750);
   U21207 : OAI222_X1 port map( A1 => n20269, A2 => n24460, B1 => n17242, B2 =>
                           n24454, C1 => n19339, C2 => n24448, ZN => n22732);
   U21208 : OAI222_X1 port map( A1 => n20268, A2 => n24460, B1 => n17239, B2 =>
                           n24454, C1 => n19338, C2 => n24448, ZN => n22714);
   U21209 : OAI222_X1 port map( A1 => n20267, A2 => n24460, B1 => n17236, B2 =>
                           n24454, C1 => n19337, C2 => n24448, ZN => n22696);
   U21210 : OAI222_X1 port map( A1 => n20266, A2 => n24460, B1 => n17233, B2 =>
                           n24454, C1 => n19336, C2 => n24448, ZN => n22678);
   U21211 : OAI222_X1 port map( A1 => n20397, A2 => n24456, B1 => n17410, B2 =>
                           n24450, C1 => n19395, C2 => n24444, ZN => n23750);
   U21212 : OAI222_X1 port map( A1 => n20396, A2 => n24456, B1 => n17407, B2 =>
                           n24450, C1 => n19394, C2 => n24444, ZN => n23722);
   U21213 : OAI222_X1 port map( A1 => n20395, A2 => n24456, B1 => n17404, B2 =>
                           n24450, C1 => n19393, C2 => n24444, ZN => n23704);
   U21214 : OAI222_X1 port map( A1 => n20394, A2 => n24456, B1 => n17401, B2 =>
                           n24450, C1 => n19392, C2 => n24444, ZN => n23686);
   U21215 : OAI222_X1 port map( A1 => n20393, A2 => n24456, B1 => n17398, B2 =>
                           n24450, C1 => n19391, C2 => n24444, ZN => n23668);
   U21216 : OAI222_X1 port map( A1 => n20392, A2 => n24456, B1 => n17395, B2 =>
                           n24450, C1 => n19390, C2 => n24444, ZN => n23650);
   U21217 : OAI222_X1 port map( A1 => n20391, A2 => n24456, B1 => n17392, B2 =>
                           n24450, C1 => n19389, C2 => n24444, ZN => n23632);
   U21218 : OAI222_X1 port map( A1 => n20390, A2 => n24456, B1 => n17389, B2 =>
                           n24450, C1 => n19388, C2 => n24444, ZN => n23614);
   U21219 : OAI222_X1 port map( A1 => n20389, A2 => n24456, B1 => n17386, B2 =>
                           n24450, C1 => n19387, C2 => n24444, ZN => n23596);
   U21220 : OAI222_X1 port map( A1 => n20388, A2 => n24456, B1 => n17383, B2 =>
                           n24450, C1 => n19386, C2 => n24444, ZN => n23578);
   U21221 : OAI222_X1 port map( A1 => n20387, A2 => n24456, B1 => n17380, B2 =>
                           n24450, C1 => n19385, C2 => n24444, ZN => n23560);
   U21222 : OAI222_X1 port map( A1 => n20386, A2 => n24456, B1 => n17377, B2 =>
                           n24450, C1 => n19384, C2 => n24444, ZN => n23542);
   U21223 : OAI222_X1 port map( A1 => n20385, A2 => n24457, B1 => n17374, B2 =>
                           n24451, C1 => n19383, C2 => n24445, ZN => n23524);
   U21224 : OAI222_X1 port map( A1 => n20384, A2 => n24457, B1 => n17371, B2 =>
                           n24451, C1 => n19382, C2 => n24445, ZN => n23506);
   U21225 : OAI222_X1 port map( A1 => n20383, A2 => n24457, B1 => n17368, B2 =>
                           n24451, C1 => n19381, C2 => n24445, ZN => n23488);
   U21226 : OAI222_X1 port map( A1 => n20382, A2 => n24457, B1 => n17365, B2 =>
                           n24451, C1 => n19380, C2 => n24445, ZN => n23470);
   U21227 : OAI222_X1 port map( A1 => n20381, A2 => n24457, B1 => n17362, B2 =>
                           n24451, C1 => n19379, C2 => n24445, ZN => n23452);
   U21228 : OAI222_X1 port map( A1 => n20380, A2 => n24457, B1 => n17359, B2 =>
                           n24451, C1 => n19378, C2 => n24445, ZN => n23434);
   U21229 : OAI222_X1 port map( A1 => n20379, A2 => n24457, B1 => n17356, B2 =>
                           n24451, C1 => n19377, C2 => n24445, ZN => n23416);
   U21230 : OAI222_X1 port map( A1 => n20378, A2 => n24457, B1 => n17353, B2 =>
                           n24451, C1 => n19376, C2 => n24445, ZN => n23398);
   U21231 : OAI222_X1 port map( A1 => n20377, A2 => n24457, B1 => n17350, B2 =>
                           n24451, C1 => n19375, C2 => n24445, ZN => n23380);
   U21232 : OAI222_X1 port map( A1 => n20376, A2 => n24457, B1 => n17347, B2 =>
                           n24451, C1 => n19374, C2 => n24445, ZN => n23362);
   U21233 : OAI222_X1 port map( A1 => n20375, A2 => n24457, B1 => n17344, B2 =>
                           n24451, C1 => n19373, C2 => n24445, ZN => n23344);
   U21234 : OAI222_X1 port map( A1 => n20374, A2 => n24457, B1 => n17341, B2 =>
                           n24451, C1 => n19372, C2 => n24445, ZN => n23326);
   U21235 : OAI222_X1 port map( A1 => n20301, A2 => n24458, B1 => n17338, B2 =>
                           n24452, C1 => n19371, C2 => n24446, ZN => n23308);
   U21236 : OAI222_X1 port map( A1 => n20300, A2 => n24458, B1 => n17335, B2 =>
                           n24452, C1 => n19370, C2 => n24446, ZN => n23290);
   U21237 : OAI222_X1 port map( A1 => n20299, A2 => n24458, B1 => n17332, B2 =>
                           n24452, C1 => n19369, C2 => n24446, ZN => n23272);
   U21238 : OAI222_X1 port map( A1 => n20298, A2 => n24458, B1 => n17329, B2 =>
                           n24452, C1 => n19368, C2 => n24446, ZN => n23254);
   U21239 : OAI222_X1 port map( A1 => n20297, A2 => n24458, B1 => n17326, B2 =>
                           n24452, C1 => n19367, C2 => n24446, ZN => n23236);
   U21240 : OAI222_X1 port map( A1 => n20296, A2 => n24458, B1 => n17323, B2 =>
                           n24452, C1 => n19366, C2 => n24446, ZN => n23218);
   U21241 : OAI222_X1 port map( A1 => n20295, A2 => n24458, B1 => n17320, B2 =>
                           n24452, C1 => n19365, C2 => n24446, ZN => n23200);
   U21242 : OAI222_X1 port map( A1 => n20294, A2 => n24458, B1 => n17317, B2 =>
                           n24452, C1 => n19364, C2 => n24446, ZN => n23182);
   U21243 : OAI222_X1 port map( A1 => n20293, A2 => n24458, B1 => n17314, B2 =>
                           n24452, C1 => n19363, C2 => n24446, ZN => n23164);
   U21244 : OAI222_X1 port map( A1 => n20292, A2 => n24458, B1 => n17311, B2 =>
                           n24452, C1 => n19362, C2 => n24446, ZN => n23146);
   U21245 : OAI222_X1 port map( A1 => n20291, A2 => n24458, B1 => n17308, B2 =>
                           n24452, C1 => n19361, C2 => n24446, ZN => n23128);
   U21246 : OAI222_X1 port map( A1 => n20290, A2 => n24458, B1 => n17305, B2 =>
                           n24452, C1 => n19360, C2 => n24446, ZN => n23110);
   U21247 : OAI222_X1 port map( A1 => n20289, A2 => n24459, B1 => n17302, B2 =>
                           n24453, C1 => n19359, C2 => n24447, ZN => n23092);
   U21248 : OAI222_X1 port map( A1 => n20288, A2 => n24459, B1 => n17299, B2 =>
                           n24453, C1 => n19358, C2 => n24447, ZN => n23074);
   U21249 : OAI222_X1 port map( A1 => n20287, A2 => n24459, B1 => n17296, B2 =>
                           n24453, C1 => n19357, C2 => n24447, ZN => n23056);
   U21250 : OAI222_X1 port map( A1 => n20286, A2 => n24459, B1 => n17293, B2 =>
                           n24453, C1 => n19356, C2 => n24447, ZN => n23038);
   U21251 : OAI222_X1 port map( A1 => n20253, A2 => n24461, B1 => n17230, B2 =>
                           n24455, C1 => n19335, C2 => n24449, ZN => n22660);
   U21252 : OAI222_X1 port map( A1 => n20252, A2 => n24461, B1 => n17227, B2 =>
                           n24455, C1 => n19334, C2 => n24449, ZN => n22642);
   U21253 : OAI222_X1 port map( A1 => n20251, A2 => n24461, B1 => n17224, B2 =>
                           n24455, C1 => n19333, C2 => n24449, ZN => n22624);
   U21254 : OAI222_X1 port map( A1 => n20250, A2 => n24461, B1 => n17221, B2 =>
                           n24455, C1 => n19332, C2 => n24449, ZN => n22589);
   U21255 : NOR4_X1 port map( A1 => n22652, A2 => n22653, A3 => n22654, A4 => 
                           n22655, ZN => n22651);
   U21256 : OAI221_X1 port map( B1 => n20513, B2 => n24551, C1 => n20517, C2 =>
                           n24545, A => n22658, ZN => n22653);
   U21257 : OAI221_X1 port map( B1 => n20265, B2 => n24575, C1 => n7307, C2 => 
                           n24569, A => n22657, ZN => n22654);
   U21258 : OAI221_X1 port map( B1 => n20509, B2 => n24527, C1 => n836, C2 => 
                           n24521, A => n22659, ZN => n22652);
   U21259 : NOR4_X1 port map( A1 => n22634, A2 => n22635, A3 => n22636, A4 => 
                           n22637, ZN => n22633);
   U21260 : OAI221_X1 port map( B1 => n20512, B2 => n24551, C1 => n20516, C2 =>
                           n24545, A => n22640, ZN => n22635);
   U21261 : OAI221_X1 port map( B1 => n20264, B2 => n24575, C1 => n7305, C2 => 
                           n24569, A => n22639, ZN => n22636);
   U21262 : OAI221_X1 port map( B1 => n20508, B2 => n24527, C1 => n835, C2 => 
                           n24521, A => n22641, ZN => n22634);
   U21263 : NOR4_X1 port map( A1 => n22616, A2 => n22617, A3 => n22618, A4 => 
                           n22619, ZN => n22615);
   U21264 : OAI221_X1 port map( B1 => n20511, B2 => n24551, C1 => n20515, C2 =>
                           n24545, A => n22622, ZN => n22617);
   U21265 : OAI221_X1 port map( B1 => n20263, B2 => n24575, C1 => n7303, C2 => 
                           n24569, A => n22621, ZN => n22618);
   U21266 : OAI221_X1 port map( B1 => n20507, B2 => n24527, C1 => n834, C2 => 
                           n24521, A => n22623, ZN => n22616);
   U21267 : NOR4_X1 port map( A1 => n22564, A2 => n22565, A3 => n22566, A4 => 
                           n22567, ZN => n22563);
   U21268 : OAI221_X1 port map( B1 => n20510, B2 => n24551, C1 => n20514, C2 =>
                           n24545, A => n22580, ZN => n22565);
   U21269 : OAI221_X1 port map( B1 => n20262, B2 => n24575, C1 => n7301, C2 => 
                           n24569, A => n22575, ZN => n22566);
   U21270 : OAI221_X1 port map( B1 => n20506, B2 => n24527, C1 => n833, C2 => 
                           n24521, A => n22585, ZN => n22564);
   U21271 : NOR4_X1 port map( A1 => n23012, A2 => n23013, A3 => n23014, A4 => 
                           n23015, ZN => n23011);
   U21272 : OAI221_X1 port map( B1 => n20602, B2 => n24549, C1 => n20638, C2 =>
                           n24543, A => n23018, ZN => n23013);
   U21273 : OAI221_X1 port map( B1 => n20465, B2 => n24573, C1 => n7347, C2 => 
                           n24567, A => n23017, ZN => n23014);
   U21274 : OAI221_X1 port map( B1 => n20566, B2 => n24525, C1 => n856, C2 => 
                           n24519, A => n23019, ZN => n23012);
   U21275 : NOR4_X1 port map( A1 => n22994, A2 => n22995, A3 => n22996, A4 => 
                           n22997, ZN => n22993);
   U21276 : OAI221_X1 port map( B1 => n20601, B2 => n24549, C1 => n20637, C2 =>
                           n24543, A => n23000, ZN => n22995);
   U21277 : OAI221_X1 port map( B1 => n20464, B2 => n24573, C1 => n7345, C2 => 
                           n24567, A => n22999, ZN => n22996);
   U21278 : OAI221_X1 port map( B1 => n20565, B2 => n24525, C1 => n855, C2 => 
                           n24519, A => n23001, ZN => n22994);
   U21279 : NOR4_X1 port map( A1 => n22976, A2 => n22977, A3 => n22978, A4 => 
                           n22979, ZN => n22975);
   U21280 : OAI221_X1 port map( B1 => n20600, B2 => n24549, C1 => n20636, C2 =>
                           n24543, A => n22982, ZN => n22977);
   U21281 : OAI221_X1 port map( B1 => n20463, B2 => n24573, C1 => n7343, C2 => 
                           n24567, A => n22981, ZN => n22978);
   U21282 : OAI221_X1 port map( B1 => n20564, B2 => n24525, C1 => n854, C2 => 
                           n24519, A => n22983, ZN => n22976);
   U21283 : NOR4_X1 port map( A1 => n22958, A2 => n22959, A3 => n22960, A4 => 
                           n22961, ZN => n22957);
   U21284 : OAI221_X1 port map( B1 => n20599, B2 => n24549, C1 => n20635, C2 =>
                           n24543, A => n22964, ZN => n22959);
   U21285 : OAI221_X1 port map( B1 => n20462, B2 => n24573, C1 => n7341, C2 => 
                           n24567, A => n22963, ZN => n22960);
   U21286 : OAI221_X1 port map( B1 => n20563, B2 => n24525, C1 => n853, C2 => 
                           n24519, A => n22965, ZN => n22958);
   U21287 : NOR4_X1 port map( A1 => n22940, A2 => n22941, A3 => n22942, A4 => 
                           n22943, ZN => n22939);
   U21288 : OAI221_X1 port map( B1 => n20598, B2 => n24549, C1 => n20634, C2 =>
                           n24543, A => n22946, ZN => n22941);
   U21289 : OAI221_X1 port map( B1 => n20461, B2 => n24573, C1 => n7339, C2 => 
                           n24567, A => n22945, ZN => n22942);
   U21290 : OAI221_X1 port map( B1 => n20562, B2 => n24525, C1 => n852, C2 => 
                           n24519, A => n22947, ZN => n22940);
   U21291 : NOR4_X1 port map( A1 => n22922, A2 => n22923, A3 => n22924, A4 => 
                           n22925, ZN => n22921);
   U21292 : OAI221_X1 port map( B1 => n20597, B2 => n24549, C1 => n20633, C2 =>
                           n24543, A => n22928, ZN => n22923);
   U21293 : OAI221_X1 port map( B1 => n20460, B2 => n24573, C1 => n7337, C2 => 
                           n24567, A => n22927, ZN => n22924);
   U21294 : OAI221_X1 port map( B1 => n20561, B2 => n24525, C1 => n851, C2 => 
                           n24519, A => n22929, ZN => n22922);
   U21295 : NOR4_X1 port map( A1 => n22904, A2 => n22905, A3 => n22906, A4 => 
                           n22907, ZN => n22903);
   U21296 : OAI221_X1 port map( B1 => n20596, B2 => n24549, C1 => n20632, C2 =>
                           n24543, A => n22910, ZN => n22905);
   U21297 : OAI221_X1 port map( B1 => n20459, B2 => n24573, C1 => n7335, C2 => 
                           n24567, A => n22909, ZN => n22906);
   U21298 : OAI221_X1 port map( B1 => n20560, B2 => n24525, C1 => n850, C2 => 
                           n24519, A => n22911, ZN => n22904);
   U21299 : NOR4_X1 port map( A1 => n22886, A2 => n22887, A3 => n22888, A4 => 
                           n22889, ZN => n22885);
   U21300 : OAI221_X1 port map( B1 => n20595, B2 => n24549, C1 => n20631, C2 =>
                           n24543, A => n22892, ZN => n22887);
   U21301 : OAI221_X1 port map( B1 => n20458, B2 => n24573, C1 => n7333, C2 => 
                           n24567, A => n22891, ZN => n22888);
   U21302 : OAI221_X1 port map( B1 => n20559, B2 => n24525, C1 => n849, C2 => 
                           n24519, A => n22893, ZN => n22886);
   U21303 : NOR4_X1 port map( A1 => n22868, A2 => n22869, A3 => n22870, A4 => 
                           n22871, ZN => n22867);
   U21304 : OAI221_X1 port map( B1 => n20594, B2 => n24550, C1 => n20630, C2 =>
                           n24544, A => n22874, ZN => n22869);
   U21305 : OAI221_X1 port map( B1 => n20457, B2 => n24574, C1 => n7331, C2 => 
                           n24568, A => n22873, ZN => n22870);
   U21306 : OAI221_X1 port map( B1 => n20558, B2 => n24526, C1 => n848, C2 => 
                           n24520, A => n22875, ZN => n22868);
   U21307 : NOR4_X1 port map( A1 => n22850, A2 => n22851, A3 => n22852, A4 => 
                           n22853, ZN => n22849);
   U21308 : OAI221_X1 port map( B1 => n20593, B2 => n24550, C1 => n20629, C2 =>
                           n24544, A => n22856, ZN => n22851);
   U21309 : OAI221_X1 port map( B1 => n20456, B2 => n24574, C1 => n7329, C2 => 
                           n24568, A => n22855, ZN => n22852);
   U21310 : OAI221_X1 port map( B1 => n20557, B2 => n24526, C1 => n847, C2 => 
                           n24520, A => n22857, ZN => n22850);
   U21311 : NOR4_X1 port map( A1 => n22832, A2 => n22833, A3 => n22834, A4 => 
                           n22835, ZN => n22831);
   U21312 : OAI221_X1 port map( B1 => n20592, B2 => n24550, C1 => n20628, C2 =>
                           n24544, A => n22838, ZN => n22833);
   U21313 : OAI221_X1 port map( B1 => n20455, B2 => n24574, C1 => n7327, C2 => 
                           n24568, A => n22837, ZN => n22834);
   U21314 : OAI221_X1 port map( B1 => n20556, B2 => n24526, C1 => n846, C2 => 
                           n24520, A => n22839, ZN => n22832);
   U21315 : NOR4_X1 port map( A1 => n22814, A2 => n22815, A3 => n22816, A4 => 
                           n22817, ZN => n22813);
   U21316 : OAI221_X1 port map( B1 => n20591, B2 => n24550, C1 => n20627, C2 =>
                           n24544, A => n22820, ZN => n22815);
   U21317 : OAI221_X1 port map( B1 => n20454, B2 => n24574, C1 => n7325, C2 => 
                           n24568, A => n22819, ZN => n22816);
   U21318 : OAI221_X1 port map( B1 => n20555, B2 => n24526, C1 => n845, C2 => 
                           n24520, A => n22821, ZN => n22814);
   U21319 : NOR4_X1 port map( A1 => n22796, A2 => n22797, A3 => n22798, A4 => 
                           n22799, ZN => n22795);
   U21320 : OAI221_X1 port map( B1 => n20590, B2 => n24550, C1 => n20626, C2 =>
                           n24544, A => n22802, ZN => n22797);
   U21321 : OAI221_X1 port map( B1 => n20453, B2 => n24574, C1 => n7323, C2 => 
                           n24568, A => n22801, ZN => n22798);
   U21322 : OAI221_X1 port map( B1 => n20554, B2 => n24526, C1 => n844, C2 => 
                           n24520, A => n22803, ZN => n22796);
   U21323 : NOR4_X1 port map( A1 => n22778, A2 => n22779, A3 => n22780, A4 => 
                           n22781, ZN => n22777);
   U21324 : OAI221_X1 port map( B1 => n20589, B2 => n24550, C1 => n20625, C2 =>
                           n24544, A => n22784, ZN => n22779);
   U21325 : OAI221_X1 port map( B1 => n20452, B2 => n24574, C1 => n7321, C2 => 
                           n24568, A => n22783, ZN => n22780);
   U21326 : OAI221_X1 port map( B1 => n20553, B2 => n24526, C1 => n843, C2 => 
                           n24520, A => n22785, ZN => n22778);
   U21327 : NOR4_X1 port map( A1 => n22760, A2 => n22761, A3 => n22762, A4 => 
                           n22763, ZN => n22759);
   U21328 : OAI221_X1 port map( B1 => n20588, B2 => n24550, C1 => n20624, C2 =>
                           n24544, A => n22766, ZN => n22761);
   U21329 : OAI221_X1 port map( B1 => n20451, B2 => n24574, C1 => n7319, C2 => 
                           n24568, A => n22765, ZN => n22762);
   U21330 : OAI221_X1 port map( B1 => n20552, B2 => n24526, C1 => n842, C2 => 
                           n24520, A => n22767, ZN => n22760);
   U21331 : NOR4_X1 port map( A1 => n22742, A2 => n22743, A3 => n22744, A4 => 
                           n22745, ZN => n22741);
   U21332 : OAI221_X1 port map( B1 => n20587, B2 => n24550, C1 => n20623, C2 =>
                           n24544, A => n22748, ZN => n22743);
   U21333 : OAI221_X1 port map( B1 => n20450, B2 => n24574, C1 => n7317, C2 => 
                           n24568, A => n22747, ZN => n22744);
   U21334 : OAI221_X1 port map( B1 => n20551, B2 => n24526, C1 => n841, C2 => 
                           n24520, A => n22749, ZN => n22742);
   U21335 : NOR4_X1 port map( A1 => n22724, A2 => n22725, A3 => n22726, A4 => 
                           n22727, ZN => n22723);
   U21336 : OAI221_X1 port map( B1 => n20586, B2 => n24550, C1 => n20622, C2 =>
                           n24544, A => n22730, ZN => n22725);
   U21337 : OAI221_X1 port map( B1 => n20449, B2 => n24574, C1 => n7315, C2 => 
                           n24568, A => n22729, ZN => n22726);
   U21338 : OAI221_X1 port map( B1 => n20550, B2 => n24526, C1 => n840, C2 => 
                           n24520, A => n22731, ZN => n22724);
   U21339 : NOR4_X1 port map( A1 => n22706, A2 => n22707, A3 => n22708, A4 => 
                           n22709, ZN => n22705);
   U21340 : OAI221_X1 port map( B1 => n20585, B2 => n24550, C1 => n20621, C2 =>
                           n24544, A => n22712, ZN => n22707);
   U21341 : OAI221_X1 port map( B1 => n20448, B2 => n24574, C1 => n7313, C2 => 
                           n24568, A => n22711, ZN => n22708);
   U21342 : OAI221_X1 port map( B1 => n20549, B2 => n24526, C1 => n839, C2 => 
                           n24520, A => n22713, ZN => n22706);
   U21343 : NOR4_X1 port map( A1 => n22688, A2 => n22689, A3 => n22690, A4 => 
                           n22691, ZN => n22687);
   U21344 : OAI221_X1 port map( B1 => n20584, B2 => n24550, C1 => n20620, C2 =>
                           n24544, A => n22694, ZN => n22689);
   U21345 : OAI221_X1 port map( B1 => n20447, B2 => n24574, C1 => n7311, C2 => 
                           n24568, A => n22693, ZN => n22690);
   U21346 : OAI221_X1 port map( B1 => n20548, B2 => n24526, C1 => n838, C2 => 
                           n24520, A => n22695, ZN => n22688);
   U21347 : NOR4_X1 port map( A1 => n22670, A2 => n22671, A3 => n22672, A4 => 
                           n22673, ZN => n22669);
   U21348 : OAI221_X1 port map( B1 => n20583, B2 => n24550, C1 => n20619, C2 =>
                           n24544, A => n22676, ZN => n22671);
   U21349 : OAI221_X1 port map( B1 => n20446, B2 => n24574, C1 => n7309, C2 => 
                           n24568, A => n22675, ZN => n22672);
   U21350 : OAI221_X1 port map( B1 => n20547, B2 => n24526, C1 => n837, C2 => 
                           n24520, A => n22677, ZN => n22670);
   U21351 : NOR4_X1 port map( A1 => n23732, A2 => n23733, A3 => n23734, A4 => 
                           n23735, ZN => n23731);
   U21352 : OAI221_X1 port map( B1 => n20774, B2 => n24546, C1 => n20798, C2 =>
                           n24540, A => n23746, ZN => n23733);
   U21353 : OAI221_X1 port map( B1 => n20505, B2 => n24570, C1 => n7427, C2 => 
                           n24564, A => n23743, ZN => n23734);
   U21354 : OAI221_X1 port map( B1 => n20750, B2 => n24522, C1 => n896, C2 => 
                           n24516, A => n23749, ZN => n23732);
   U21355 : NOR4_X1 port map( A1 => n23714, A2 => n23715, A3 => n23716, A4 => 
                           n23717, ZN => n23713);
   U21356 : OAI221_X1 port map( B1 => n20773, B2 => n24546, C1 => n20797, C2 =>
                           n24540, A => n23720, ZN => n23715);
   U21357 : OAI221_X1 port map( B1 => n20504, B2 => n24570, C1 => n7425, C2 => 
                           n24564, A => n23719, ZN => n23716);
   U21358 : OAI221_X1 port map( B1 => n20749, B2 => n24522, C1 => n895, C2 => 
                           n24516, A => n23721, ZN => n23714);
   U21359 : NOR4_X1 port map( A1 => n23696, A2 => n23697, A3 => n23698, A4 => 
                           n23699, ZN => n23695);
   U21360 : OAI221_X1 port map( B1 => n20772, B2 => n24546, C1 => n20796, C2 =>
                           n24540, A => n23702, ZN => n23697);
   U21361 : OAI221_X1 port map( B1 => n20503, B2 => n24570, C1 => n7423, C2 => 
                           n24564, A => n23701, ZN => n23698);
   U21362 : OAI221_X1 port map( B1 => n20748, B2 => n24522, C1 => n894, C2 => 
                           n24516, A => n23703, ZN => n23696);
   U21363 : NOR4_X1 port map( A1 => n23678, A2 => n23679, A3 => n23680, A4 => 
                           n23681, ZN => n23677);
   U21364 : OAI221_X1 port map( B1 => n20771, B2 => n24546, C1 => n20795, C2 =>
                           n24540, A => n23684, ZN => n23679);
   U21365 : OAI221_X1 port map( B1 => n20502, B2 => n24570, C1 => n7421, C2 => 
                           n24564, A => n23683, ZN => n23680);
   U21366 : OAI221_X1 port map( B1 => n20747, B2 => n24522, C1 => n893, C2 => 
                           n24516, A => n23685, ZN => n23678);
   U21367 : NOR4_X1 port map( A1 => n23660, A2 => n23661, A3 => n23662, A4 => 
                           n23663, ZN => n23659);
   U21368 : OAI221_X1 port map( B1 => n20770, B2 => n24546, C1 => n20794, C2 =>
                           n24540, A => n23666, ZN => n23661);
   U21369 : OAI221_X1 port map( B1 => n20501, B2 => n24570, C1 => n7419, C2 => 
                           n24564, A => n23665, ZN => n23662);
   U21370 : OAI221_X1 port map( B1 => n20746, B2 => n24522, C1 => n892, C2 => 
                           n24516, A => n23667, ZN => n23660);
   U21371 : NOR4_X1 port map( A1 => n23642, A2 => n23643, A3 => n23644, A4 => 
                           n23645, ZN => n23641);
   U21372 : OAI221_X1 port map( B1 => n20769, B2 => n24546, C1 => n20793, C2 =>
                           n24540, A => n23648, ZN => n23643);
   U21373 : OAI221_X1 port map( B1 => n20500, B2 => n24570, C1 => n7417, C2 => 
                           n24564, A => n23647, ZN => n23644);
   U21374 : OAI221_X1 port map( B1 => n20745, B2 => n24522, C1 => n891, C2 => 
                           n24516, A => n23649, ZN => n23642);
   U21375 : NOR4_X1 port map( A1 => n23624, A2 => n23625, A3 => n23626, A4 => 
                           n23627, ZN => n23623);
   U21376 : OAI221_X1 port map( B1 => n20768, B2 => n24546, C1 => n20792, C2 =>
                           n24540, A => n23630, ZN => n23625);
   U21377 : OAI221_X1 port map( B1 => n20499, B2 => n24570, C1 => n7415, C2 => 
                           n24564, A => n23629, ZN => n23626);
   U21378 : OAI221_X1 port map( B1 => n20744, B2 => n24522, C1 => n890, C2 => 
                           n24516, A => n23631, ZN => n23624);
   U21379 : NOR4_X1 port map( A1 => n23606, A2 => n23607, A3 => n23608, A4 => 
                           n23609, ZN => n23605);
   U21380 : OAI221_X1 port map( B1 => n20767, B2 => n24546, C1 => n20791, C2 =>
                           n24540, A => n23612, ZN => n23607);
   U21381 : OAI221_X1 port map( B1 => n20498, B2 => n24570, C1 => n7413, C2 => 
                           n24564, A => n23611, ZN => n23608);
   U21382 : OAI221_X1 port map( B1 => n20743, B2 => n24522, C1 => n889, C2 => 
                           n24516, A => n23613, ZN => n23606);
   U21383 : NOR4_X1 port map( A1 => n23588, A2 => n23589, A3 => n23590, A4 => 
                           n23591, ZN => n23587);
   U21384 : OAI221_X1 port map( B1 => n20766, B2 => n24546, C1 => n20790, C2 =>
                           n24540, A => n23594, ZN => n23589);
   U21385 : OAI221_X1 port map( B1 => n20497, B2 => n24570, C1 => n7411, C2 => 
                           n24564, A => n23593, ZN => n23590);
   U21386 : OAI221_X1 port map( B1 => n20742, B2 => n24522, C1 => n888, C2 => 
                           n24516, A => n23595, ZN => n23588);
   U21387 : NOR4_X1 port map( A1 => n23570, A2 => n23571, A3 => n23572, A4 => 
                           n23573, ZN => n23569);
   U21388 : OAI221_X1 port map( B1 => n20765, B2 => n24546, C1 => n20789, C2 =>
                           n24540, A => n23576, ZN => n23571);
   U21389 : OAI221_X1 port map( B1 => n20496, B2 => n24570, C1 => n7409, C2 => 
                           n24564, A => n23575, ZN => n23572);
   U21390 : OAI221_X1 port map( B1 => n20741, B2 => n24522, C1 => n887, C2 => 
                           n24516, A => n23577, ZN => n23570);
   U21391 : NOR4_X1 port map( A1 => n23552, A2 => n23553, A3 => n23554, A4 => 
                           n23555, ZN => n23551);
   U21392 : OAI221_X1 port map( B1 => n20764, B2 => n24546, C1 => n20788, C2 =>
                           n24540, A => n23558, ZN => n23553);
   U21393 : OAI221_X1 port map( B1 => n20495, B2 => n24570, C1 => n7407, C2 => 
                           n24564, A => n23557, ZN => n23554);
   U21394 : OAI221_X1 port map( B1 => n20740, B2 => n24522, C1 => n886, C2 => 
                           n24516, A => n23559, ZN => n23552);
   U21395 : NOR4_X1 port map( A1 => n23534, A2 => n23535, A3 => n23536, A4 => 
                           n23537, ZN => n23533);
   U21396 : OAI221_X1 port map( B1 => n20763, B2 => n24546, C1 => n20787, C2 =>
                           n24540, A => n23540, ZN => n23535);
   U21397 : OAI221_X1 port map( B1 => n20494, B2 => n24570, C1 => n7405, C2 => 
                           n24564, A => n23539, ZN => n23536);
   U21398 : OAI221_X1 port map( B1 => n20739, B2 => n24522, C1 => n885, C2 => 
                           n24516, A => n23541, ZN => n23534);
   U21399 : NOR4_X1 port map( A1 => n23516, A2 => n23517, A3 => n23518, A4 => 
                           n23519, ZN => n23515);
   U21400 : OAI221_X1 port map( B1 => n20762, B2 => n24547, C1 => n20786, C2 =>
                           n24541, A => n23522, ZN => n23517);
   U21401 : OAI221_X1 port map( B1 => n20493, B2 => n24571, C1 => n7403, C2 => 
                           n24565, A => n23521, ZN => n23518);
   U21402 : OAI221_X1 port map( B1 => n20738, B2 => n24523, C1 => n884, C2 => 
                           n24517, A => n23523, ZN => n23516);
   U21403 : NOR4_X1 port map( A1 => n23498, A2 => n23499, A3 => n23500, A4 => 
                           n23501, ZN => n23497);
   U21404 : OAI221_X1 port map( B1 => n20761, B2 => n24547, C1 => n20785, C2 =>
                           n24541, A => n23504, ZN => n23499);
   U21405 : OAI221_X1 port map( B1 => n20492, B2 => n24571, C1 => n7401, C2 => 
                           n24565, A => n23503, ZN => n23500);
   U21406 : OAI221_X1 port map( B1 => n20737, B2 => n24523, C1 => n883, C2 => 
                           n24517, A => n23505, ZN => n23498);
   U21407 : NOR4_X1 port map( A1 => n23480, A2 => n23481, A3 => n23482, A4 => 
                           n23483, ZN => n23479);
   U21408 : OAI221_X1 port map( B1 => n20760, B2 => n24547, C1 => n20784, C2 =>
                           n24541, A => n23486, ZN => n23481);
   U21409 : OAI221_X1 port map( B1 => n20491, B2 => n24571, C1 => n7399, C2 => 
                           n24565, A => n23485, ZN => n23482);
   U21410 : OAI221_X1 port map( B1 => n20736, B2 => n24523, C1 => n882, C2 => 
                           n24517, A => n23487, ZN => n23480);
   U21411 : NOR4_X1 port map( A1 => n23462, A2 => n23463, A3 => n23464, A4 => 
                           n23465, ZN => n23461);
   U21412 : OAI221_X1 port map( B1 => n20759, B2 => n24547, C1 => n20783, C2 =>
                           n24541, A => n23468, ZN => n23463);
   U21413 : OAI221_X1 port map( B1 => n20490, B2 => n24571, C1 => n7397, C2 => 
                           n24565, A => n23467, ZN => n23464);
   U21414 : OAI221_X1 port map( B1 => n20735, B2 => n24523, C1 => n881, C2 => 
                           n24517, A => n23469, ZN => n23462);
   U21415 : NOR4_X1 port map( A1 => n23444, A2 => n23445, A3 => n23446, A4 => 
                           n23447, ZN => n23443);
   U21416 : OAI221_X1 port map( B1 => n20758, B2 => n24547, C1 => n20782, C2 =>
                           n24541, A => n23450, ZN => n23445);
   U21417 : OAI221_X1 port map( B1 => n20489, B2 => n24571, C1 => n7395, C2 => 
                           n24565, A => n23449, ZN => n23446);
   U21418 : OAI221_X1 port map( B1 => n20734, B2 => n24523, C1 => n880, C2 => 
                           n24517, A => n23451, ZN => n23444);
   U21419 : NOR4_X1 port map( A1 => n23426, A2 => n23427, A3 => n23428, A4 => 
                           n23429, ZN => n23425);
   U21420 : OAI221_X1 port map( B1 => n20757, B2 => n24547, C1 => n20781, C2 =>
                           n24541, A => n23432, ZN => n23427);
   U21421 : OAI221_X1 port map( B1 => n20488, B2 => n24571, C1 => n7393, C2 => 
                           n24565, A => n23431, ZN => n23428);
   U21422 : OAI221_X1 port map( B1 => n20733, B2 => n24523, C1 => n879, C2 => 
                           n24517, A => n23433, ZN => n23426);
   U21423 : NOR4_X1 port map( A1 => n23408, A2 => n23409, A3 => n23410, A4 => 
                           n23411, ZN => n23407);
   U21424 : OAI221_X1 port map( B1 => n20756, B2 => n24547, C1 => n20780, C2 =>
                           n24541, A => n23414, ZN => n23409);
   U21425 : OAI221_X1 port map( B1 => n20487, B2 => n24571, C1 => n7391, C2 => 
                           n24565, A => n23413, ZN => n23410);
   U21426 : OAI221_X1 port map( B1 => n20732, B2 => n24523, C1 => n878, C2 => 
                           n24517, A => n23415, ZN => n23408);
   U21427 : NOR4_X1 port map( A1 => n23390, A2 => n23391, A3 => n23392, A4 => 
                           n23393, ZN => n23389);
   U21428 : OAI221_X1 port map( B1 => n20755, B2 => n24547, C1 => n20779, C2 =>
                           n24541, A => n23396, ZN => n23391);
   U21429 : OAI221_X1 port map( B1 => n20486, B2 => n24571, C1 => n7389, C2 => 
                           n24565, A => n23395, ZN => n23392);
   U21430 : OAI221_X1 port map( B1 => n20731, B2 => n24523, C1 => n877, C2 => 
                           n24517, A => n23397, ZN => n23390);
   U21431 : NOR4_X1 port map( A1 => n23372, A2 => n23373, A3 => n23374, A4 => 
                           n23375, ZN => n23371);
   U21432 : OAI221_X1 port map( B1 => n20754, B2 => n24547, C1 => n20778, C2 =>
                           n24541, A => n23378, ZN => n23373);
   U21433 : OAI221_X1 port map( B1 => n20485, B2 => n24571, C1 => n7387, C2 => 
                           n24565, A => n23377, ZN => n23374);
   U21434 : OAI221_X1 port map( B1 => n20730, B2 => n24523, C1 => n876, C2 => 
                           n24517, A => n23379, ZN => n23372);
   U21435 : NOR4_X1 port map( A1 => n23354, A2 => n23355, A3 => n23356, A4 => 
                           n23357, ZN => n23353);
   U21436 : OAI221_X1 port map( B1 => n20753, B2 => n24547, C1 => n20777, C2 =>
                           n24541, A => n23360, ZN => n23355);
   U21437 : OAI221_X1 port map( B1 => n20484, B2 => n24571, C1 => n7385, C2 => 
                           n24565, A => n23359, ZN => n23356);
   U21438 : OAI221_X1 port map( B1 => n20729, B2 => n24523, C1 => n875, C2 => 
                           n24517, A => n23361, ZN => n23354);
   U21439 : NOR4_X1 port map( A1 => n23336, A2 => n23337, A3 => n23338, A4 => 
                           n23339, ZN => n23335);
   U21440 : OAI221_X1 port map( B1 => n20752, B2 => n24547, C1 => n20776, C2 =>
                           n24541, A => n23342, ZN => n23337);
   U21441 : OAI221_X1 port map( B1 => n20483, B2 => n24571, C1 => n7383, C2 => 
                           n24565, A => n23341, ZN => n23338);
   U21442 : OAI221_X1 port map( B1 => n20728, B2 => n24523, C1 => n874, C2 => 
                           n24517, A => n23343, ZN => n23336);
   U21443 : NOR4_X1 port map( A1 => n23318, A2 => n23319, A3 => n23320, A4 => 
                           n23321, ZN => n23317);
   U21444 : OAI221_X1 port map( B1 => n20751, B2 => n24547, C1 => n20775, C2 =>
                           n24541, A => n23324, ZN => n23319);
   U21445 : OAI221_X1 port map( B1 => n20482, B2 => n24571, C1 => n7381, C2 => 
                           n24565, A => n23323, ZN => n23320);
   U21446 : OAI221_X1 port map( B1 => n20727, B2 => n24523, C1 => n873, C2 => 
                           n24517, A => n23325, ZN => n23318);
   U21447 : NOR4_X1 port map( A1 => n23300, A2 => n23301, A3 => n23302, A4 => 
                           n23303, ZN => n23299);
   U21448 : OAI221_X1 port map( B1 => n20618, B2 => n24548, C1 => n20654, C2 =>
                           n24542, A => n23306, ZN => n23301);
   U21449 : OAI221_X1 port map( B1 => n20481, B2 => n24572, C1 => n7379, C2 => 
                           n24566, A => n23305, ZN => n23302);
   U21450 : OAI221_X1 port map( B1 => n20582, B2 => n24524, C1 => n872, C2 => 
                           n24518, A => n23307, ZN => n23300);
   U21451 : NOR4_X1 port map( A1 => n23282, A2 => n23283, A3 => n23284, A4 => 
                           n23285, ZN => n23281);
   U21452 : OAI221_X1 port map( B1 => n20617, B2 => n24548, C1 => n20653, C2 =>
                           n24542, A => n23288, ZN => n23283);
   U21453 : OAI221_X1 port map( B1 => n20480, B2 => n24572, C1 => n7377, C2 => 
                           n24566, A => n23287, ZN => n23284);
   U21454 : OAI221_X1 port map( B1 => n20581, B2 => n24524, C1 => n871, C2 => 
                           n24518, A => n23289, ZN => n23282);
   U21455 : NOR4_X1 port map( A1 => n23264, A2 => n23265, A3 => n23266, A4 => 
                           n23267, ZN => n23263);
   U21456 : OAI221_X1 port map( B1 => n20616, B2 => n24548, C1 => n20652, C2 =>
                           n24542, A => n23270, ZN => n23265);
   U21457 : OAI221_X1 port map( B1 => n20479, B2 => n24572, C1 => n7375, C2 => 
                           n24566, A => n23269, ZN => n23266);
   U21458 : OAI221_X1 port map( B1 => n20580, B2 => n24524, C1 => n870, C2 => 
                           n24518, A => n23271, ZN => n23264);
   U21459 : NOR4_X1 port map( A1 => n23246, A2 => n23247, A3 => n23248, A4 => 
                           n23249, ZN => n23245);
   U21460 : OAI221_X1 port map( B1 => n20615, B2 => n24548, C1 => n20651, C2 =>
                           n24542, A => n23252, ZN => n23247);
   U21461 : OAI221_X1 port map( B1 => n20478, B2 => n24572, C1 => n7373, C2 => 
                           n24566, A => n23251, ZN => n23248);
   U21462 : OAI221_X1 port map( B1 => n20579, B2 => n24524, C1 => n869, C2 => 
                           n24518, A => n23253, ZN => n23246);
   U21463 : NOR4_X1 port map( A1 => n23228, A2 => n23229, A3 => n23230, A4 => 
                           n23231, ZN => n23227);
   U21464 : OAI221_X1 port map( B1 => n20614, B2 => n24548, C1 => n20650, C2 =>
                           n24542, A => n23234, ZN => n23229);
   U21465 : OAI221_X1 port map( B1 => n20477, B2 => n24572, C1 => n7371, C2 => 
                           n24566, A => n23233, ZN => n23230);
   U21466 : OAI221_X1 port map( B1 => n20578, B2 => n24524, C1 => n868, C2 => 
                           n24518, A => n23235, ZN => n23228);
   U21467 : NOR4_X1 port map( A1 => n23210, A2 => n23211, A3 => n23212, A4 => 
                           n23213, ZN => n23209);
   U21468 : OAI221_X1 port map( B1 => n20613, B2 => n24548, C1 => n20649, C2 =>
                           n24542, A => n23216, ZN => n23211);
   U21469 : OAI221_X1 port map( B1 => n20476, B2 => n24572, C1 => n7369, C2 => 
                           n24566, A => n23215, ZN => n23212);
   U21470 : OAI221_X1 port map( B1 => n20577, B2 => n24524, C1 => n867, C2 => 
                           n24518, A => n23217, ZN => n23210);
   U21471 : NOR4_X1 port map( A1 => n23192, A2 => n23193, A3 => n23194, A4 => 
                           n23195, ZN => n23191);
   U21472 : OAI221_X1 port map( B1 => n20612, B2 => n24548, C1 => n20648, C2 =>
                           n24542, A => n23198, ZN => n23193);
   U21473 : OAI221_X1 port map( B1 => n20475, B2 => n24572, C1 => n7367, C2 => 
                           n24566, A => n23197, ZN => n23194);
   U21474 : OAI221_X1 port map( B1 => n20576, B2 => n24524, C1 => n866, C2 => 
                           n24518, A => n23199, ZN => n23192);
   U21475 : NOR4_X1 port map( A1 => n23174, A2 => n23175, A3 => n23176, A4 => 
                           n23177, ZN => n23173);
   U21476 : OAI221_X1 port map( B1 => n20611, B2 => n24548, C1 => n20647, C2 =>
                           n24542, A => n23180, ZN => n23175);
   U21477 : OAI221_X1 port map( B1 => n20474, B2 => n24572, C1 => n7365, C2 => 
                           n24566, A => n23179, ZN => n23176);
   U21478 : OAI221_X1 port map( B1 => n20575, B2 => n24524, C1 => n865, C2 => 
                           n24518, A => n23181, ZN => n23174);
   U21479 : NOR4_X1 port map( A1 => n23156, A2 => n23157, A3 => n23158, A4 => 
                           n23159, ZN => n23155);
   U21480 : OAI221_X1 port map( B1 => n20610, B2 => n24548, C1 => n20646, C2 =>
                           n24542, A => n23162, ZN => n23157);
   U21481 : OAI221_X1 port map( B1 => n20473, B2 => n24572, C1 => n7363, C2 => 
                           n24566, A => n23161, ZN => n23158);
   U21482 : OAI221_X1 port map( B1 => n20574, B2 => n24524, C1 => n864, C2 => 
                           n24518, A => n23163, ZN => n23156);
   U21483 : NOR4_X1 port map( A1 => n23138, A2 => n23139, A3 => n23140, A4 => 
                           n23141, ZN => n23137);
   U21484 : OAI221_X1 port map( B1 => n20609, B2 => n24548, C1 => n20645, C2 =>
                           n24542, A => n23144, ZN => n23139);
   U21485 : OAI221_X1 port map( B1 => n20472, B2 => n24572, C1 => n7361, C2 => 
                           n24566, A => n23143, ZN => n23140);
   U21486 : OAI221_X1 port map( B1 => n20573, B2 => n24524, C1 => n863, C2 => 
                           n24518, A => n23145, ZN => n23138);
   U21487 : NOR4_X1 port map( A1 => n23120, A2 => n23121, A3 => n23122, A4 => 
                           n23123, ZN => n23119);
   U21488 : OAI221_X1 port map( B1 => n20608, B2 => n24548, C1 => n20644, C2 =>
                           n24542, A => n23126, ZN => n23121);
   U21489 : OAI221_X1 port map( B1 => n20471, B2 => n24572, C1 => n7359, C2 => 
                           n24566, A => n23125, ZN => n23122);
   U21490 : OAI221_X1 port map( B1 => n20572, B2 => n24524, C1 => n862, C2 => 
                           n24518, A => n23127, ZN => n23120);
   U21491 : NOR4_X1 port map( A1 => n23102, A2 => n23103, A3 => n23104, A4 => 
                           n23105, ZN => n23101);
   U21492 : OAI221_X1 port map( B1 => n20607, B2 => n24548, C1 => n20643, C2 =>
                           n24542, A => n23108, ZN => n23103);
   U21493 : OAI221_X1 port map( B1 => n20470, B2 => n24572, C1 => n7357, C2 => 
                           n24566, A => n23107, ZN => n23104);
   U21494 : OAI221_X1 port map( B1 => n20571, B2 => n24524, C1 => n861, C2 => 
                           n24518, A => n23109, ZN => n23102);
   U21495 : NOR4_X1 port map( A1 => n23084, A2 => n23085, A3 => n23086, A4 => 
                           n23087, ZN => n23083);
   U21496 : OAI221_X1 port map( B1 => n20606, B2 => n24549, C1 => n20642, C2 =>
                           n24543, A => n23090, ZN => n23085);
   U21497 : OAI221_X1 port map( B1 => n20469, B2 => n24573, C1 => n7355, C2 => 
                           n24567, A => n23089, ZN => n23086);
   U21498 : OAI221_X1 port map( B1 => n20570, B2 => n24525, C1 => n860, C2 => 
                           n24519, A => n23091, ZN => n23084);
   U21499 : NOR4_X1 port map( A1 => n23066, A2 => n23067, A3 => n23068, A4 => 
                           n23069, ZN => n23065);
   U21500 : OAI221_X1 port map( B1 => n20605, B2 => n24549, C1 => n20641, C2 =>
                           n24543, A => n23072, ZN => n23067);
   U21501 : OAI221_X1 port map( B1 => n20468, B2 => n24573, C1 => n7353, C2 => 
                           n24567, A => n23071, ZN => n23068);
   U21502 : OAI221_X1 port map( B1 => n20569, B2 => n24525, C1 => n859, C2 => 
                           n24519, A => n23073, ZN => n23066);
   U21503 : NOR4_X1 port map( A1 => n23048, A2 => n23049, A3 => n23050, A4 => 
                           n23051, ZN => n23047);
   U21504 : OAI221_X1 port map( B1 => n20604, B2 => n24549, C1 => n20640, C2 =>
                           n24543, A => n23054, ZN => n23049);
   U21505 : OAI221_X1 port map( B1 => n20467, B2 => n24573, C1 => n7351, C2 => 
                           n24567, A => n23053, ZN => n23050);
   U21506 : OAI221_X1 port map( B1 => n20568, B2 => n24525, C1 => n858, C2 => 
                           n24519, A => n23055, ZN => n23048);
   U21507 : NOR4_X1 port map( A1 => n23030, A2 => n23031, A3 => n23032, A4 => 
                           n23033, ZN => n23029);
   U21508 : OAI221_X1 port map( B1 => n20603, B2 => n24549, C1 => n20639, C2 =>
                           n24543, A => n23036, ZN => n23031);
   U21509 : OAI221_X1 port map( B1 => n20466, B2 => n24573, C1 => n7349, C2 => 
                           n24567, A => n23035, ZN => n23032);
   U21510 : OAI221_X1 port map( B1 => n20567, B2 => n24525, C1 => n857, C2 => 
                           n24519, A => n23037, ZN => n23030);
   U21511 : AOI221_X1 port map( B1 => n24786, B2 => n8285, C1 => n24780, C2 => 
                           n8733, A => n22536, ZN => n22535);
   U21512 : OAI22_X1 port map( A1 => n8988, A2 => n24774, B1 => n19737, B2 => 
                           n24768, ZN => n22536);
   U21513 : AOI221_X1 port map( B1 => n24786, B2 => n8284, C1 => n24780, C2 => 
                           n8732, A => n22517, ZN => n22516);
   U21514 : OAI22_X1 port map( A1 => n8986, A2 => n24774, B1 => n19736, B2 => 
                           n24768, ZN => n22517);
   U21515 : AOI221_X1 port map( B1 => n24786, B2 => n8283, C1 => n24780, C2 => 
                           n8731, A => n22498, ZN => n22497);
   U21516 : OAI22_X1 port map( A1 => n8984, A2 => n24774, B1 => n19735, B2 => 
                           n24768, ZN => n22498);
   U21517 : AOI221_X1 port map( B1 => n24786, B2 => n8282, C1 => n24780, C2 => 
                           n8730, A => n22479, ZN => n22478);
   U21518 : OAI22_X1 port map( A1 => n8982, A2 => n24774, B1 => n19734, B2 => 
                           n24768, ZN => n22479);
   U21519 : AOI221_X1 port map( B1 => n24786, B2 => n8281, C1 => n24780, C2 => 
                           n8729, A => n22460, ZN => n22459);
   U21520 : OAI22_X1 port map( A1 => n8980, A2 => n24774, B1 => n19733, B2 => 
                           n24768, ZN => n22460);
   U21521 : AOI221_X1 port map( B1 => n24786, B2 => n8280, C1 => n24780, C2 => 
                           n8728, A => n22441, ZN => n22440);
   U21522 : OAI22_X1 port map( A1 => n8978, A2 => n24774, B1 => n19732, B2 => 
                           n24768, ZN => n22441);
   U21523 : AOI221_X1 port map( B1 => n24786, B2 => n8279, C1 => n24780, C2 => 
                           n8727, A => n22422, ZN => n22421);
   U21524 : OAI22_X1 port map( A1 => n8976, A2 => n24774, B1 => n19731, B2 => 
                           n24768, ZN => n22422);
   U21525 : AOI221_X1 port map( B1 => n24786, B2 => n8278, C1 => n24780, C2 => 
                           n8726, A => n22403, ZN => n22402);
   U21526 : OAI22_X1 port map( A1 => n8974, A2 => n24774, B1 => n19730, B2 => 
                           n24768, ZN => n22403);
   U21527 : AOI221_X1 port map( B1 => n24786, B2 => n8277, C1 => n24780, C2 => 
                           n8725, A => n22384, ZN => n22383);
   U21528 : OAI22_X1 port map( A1 => n8972, A2 => n24774, B1 => n19729, B2 => 
                           n24768, ZN => n22384);
   U21529 : AOI221_X1 port map( B1 => n24786, B2 => n8276, C1 => n24780, C2 => 
                           n8724, A => n22365, ZN => n22364);
   U21530 : OAI22_X1 port map( A1 => n8970, A2 => n24774, B1 => n19728, B2 => 
                           n24768, ZN => n22365);
   U21531 : AOI221_X1 port map( B1 => n24786, B2 => n8275, C1 => n24780, C2 => 
                           n8723, A => n22346, ZN => n22345);
   U21532 : OAI22_X1 port map( A1 => n8968, A2 => n24774, B1 => n19727, B2 => 
                           n24768, ZN => n22346);
   U21533 : AOI221_X1 port map( B1 => n24786, B2 => n8274, C1 => n24780, C2 => 
                           n8722, A => n22327, ZN => n22326);
   U21534 : OAI22_X1 port map( A1 => n8966, A2 => n24774, B1 => n19726, B2 => 
                           n24768, ZN => n22327);
   U21535 : AOI221_X1 port map( B1 => n24787, B2 => n8273, C1 => n24781, C2 => 
                           n8721, A => n22308, ZN => n22307);
   U21536 : OAI22_X1 port map( A1 => n8964, A2 => n24775, B1 => n19725, B2 => 
                           n24769, ZN => n22308);
   U21537 : AOI221_X1 port map( B1 => n24787, B2 => n8272, C1 => n24781, C2 => 
                           n8720, A => n22289, ZN => n22288);
   U21538 : OAI22_X1 port map( A1 => n8962, A2 => n24775, B1 => n19724, B2 => 
                           n24769, ZN => n22289);
   U21539 : AOI221_X1 port map( B1 => n24787, B2 => n8271, C1 => n24781, C2 => 
                           n8719, A => n22270, ZN => n22269);
   U21540 : OAI22_X1 port map( A1 => n8960, A2 => n24775, B1 => n19723, B2 => 
                           n24769, ZN => n22270);
   U21541 : AOI221_X1 port map( B1 => n24787, B2 => n8270, C1 => n24781, C2 => 
                           n8718, A => n22251, ZN => n22250);
   U21542 : OAI22_X1 port map( A1 => n8958, A2 => n24775, B1 => n19722, B2 => 
                           n24769, ZN => n22251);
   U21543 : AOI221_X1 port map( B1 => n24787, B2 => n8269, C1 => n24781, C2 => 
                           n8717, A => n22232, ZN => n22231);
   U21544 : OAI22_X1 port map( A1 => n8956, A2 => n24775, B1 => n19721, B2 => 
                           n24769, ZN => n22232);
   U21545 : AOI221_X1 port map( B1 => n24787, B2 => n8268, C1 => n24781, C2 => 
                           n8716, A => n22213, ZN => n22212);
   U21546 : OAI22_X1 port map( A1 => n8954, A2 => n24775, B1 => n19720, B2 => 
                           n24769, ZN => n22213);
   U21547 : AOI221_X1 port map( B1 => n24787, B2 => n8267, C1 => n24781, C2 => 
                           n8715, A => n22194, ZN => n22193);
   U21548 : OAI22_X1 port map( A1 => n8952, A2 => n24775, B1 => n19719, B2 => 
                           n24769, ZN => n22194);
   U21549 : AOI221_X1 port map( B1 => n24787, B2 => n8266, C1 => n24781, C2 => 
                           n8714, A => n22175, ZN => n22174);
   U21550 : OAI22_X1 port map( A1 => n8950, A2 => n24775, B1 => n19718, B2 => 
                           n24769, ZN => n22175);
   U21551 : AOI221_X1 port map( B1 => n24787, B2 => n8265, C1 => n24781, C2 => 
                           n8713, A => n22156, ZN => n22155);
   U21552 : OAI22_X1 port map( A1 => n8948, A2 => n24775, B1 => n19717, B2 => 
                           n24769, ZN => n22156);
   U21553 : AOI221_X1 port map( B1 => n24787, B2 => n8264, C1 => n24781, C2 => 
                           n8712, A => n22137, ZN => n22136);
   U21554 : OAI22_X1 port map( A1 => n8946, A2 => n24775, B1 => n19716, B2 => 
                           n24769, ZN => n22137);
   U21555 : AOI221_X1 port map( B1 => n24787, B2 => n8263, C1 => n24781, C2 => 
                           n8711, A => n22118, ZN => n22117);
   U21556 : OAI22_X1 port map( A1 => n8944, A2 => n24775, B1 => n19715, B2 => 
                           n24769, ZN => n22118);
   U21557 : AOI221_X1 port map( B1 => n24787, B2 => n8262, C1 => n24781, C2 => 
                           n8710, A => n22099, ZN => n22098);
   U21558 : OAI22_X1 port map( A1 => n8942, A2 => n24775, B1 => n19714, B2 => 
                           n24769, ZN => n22099);
   U21559 : AOI221_X1 port map( B1 => n24788, B2 => n8261, C1 => n24782, C2 => 
                           n8709, A => n22080, ZN => n22079);
   U21560 : OAI22_X1 port map( A1 => n8940, A2 => n24776, B1 => n19713, B2 => 
                           n24770, ZN => n22080);
   U21561 : AOI221_X1 port map( B1 => n24788, B2 => n8260, C1 => n24782, C2 => 
                           n8708, A => n22061, ZN => n22060);
   U21562 : OAI22_X1 port map( A1 => n8938, A2 => n24776, B1 => n19712, B2 => 
                           n24770, ZN => n22061);
   U21563 : AOI221_X1 port map( B1 => n24788, B2 => n8259, C1 => n24782, C2 => 
                           n8707, A => n22042, ZN => n22041);
   U21564 : OAI22_X1 port map( A1 => n8936, A2 => n24776, B1 => n19711, B2 => 
                           n24770, ZN => n22042);
   U21565 : AOI221_X1 port map( B1 => n24788, B2 => n8258, C1 => n24782, C2 => 
                           n8706, A => n22023, ZN => n22022);
   U21566 : OAI22_X1 port map( A1 => n8934, A2 => n24776, B1 => n19710, B2 => 
                           n24770, ZN => n22023);
   U21567 : AOI221_X1 port map( B1 => n24788, B2 => n8257, C1 => n24782, C2 => 
                           n8705, A => n22004, ZN => n22003);
   U21568 : OAI22_X1 port map( A1 => n8932, A2 => n24776, B1 => n19709, B2 => 
                           n24770, ZN => n22004);
   U21569 : AOI221_X1 port map( B1 => n24788, B2 => n8256, C1 => n24782, C2 => 
                           n8704, A => n21985, ZN => n21984);
   U21570 : OAI22_X1 port map( A1 => n8930, A2 => n24776, B1 => n19708, B2 => 
                           n24770, ZN => n21985);
   U21571 : AOI221_X1 port map( B1 => n24788, B2 => n8255, C1 => n24782, C2 => 
                           n8703, A => n21966, ZN => n21965);
   U21572 : OAI22_X1 port map( A1 => n8928, A2 => n24776, B1 => n20186, B2 => 
                           n24770, ZN => n21966);
   U21573 : AOI221_X1 port map( B1 => n24788, B2 => n8254, C1 => n24782, C2 => 
                           n8702, A => n21947, ZN => n21946);
   U21574 : OAI22_X1 port map( A1 => n8926, A2 => n24776, B1 => n20185, B2 => 
                           n24770, ZN => n21947);
   U21575 : AOI221_X1 port map( B1 => n24788, B2 => n8253, C1 => n24782, C2 => 
                           n8701, A => n21928, ZN => n21927);
   U21576 : OAI22_X1 port map( A1 => n8924, A2 => n24776, B1 => n20184, B2 => 
                           n24770, ZN => n21928);
   U21577 : AOI221_X1 port map( B1 => n24788, B2 => n8252, C1 => n24782, C2 => 
                           n8700, A => n21909, ZN => n21908);
   U21578 : OAI22_X1 port map( A1 => n8922, A2 => n24776, B1 => n20183, B2 => 
                           n24770, ZN => n21909);
   U21579 : AOI221_X1 port map( B1 => n24788, B2 => n8251, C1 => n24782, C2 => 
                           n8699, A => n21890, ZN => n21889);
   U21580 : OAI22_X1 port map( A1 => n8920, A2 => n24776, B1 => n20182, B2 => 
                           n24770, ZN => n21890);
   U21581 : AOI221_X1 port map( B1 => n24788, B2 => n8250, C1 => n24782, C2 => 
                           n8698, A => n21871, ZN => n21870);
   U21582 : OAI22_X1 port map( A1 => n8918, A2 => n24776, B1 => n20181, B2 => 
                           n24770, ZN => n21871);
   U21583 : AOI221_X1 port map( B1 => n24789, B2 => n8249, C1 => n24783, C2 => 
                           n8697, A => n21852, ZN => n21851);
   U21584 : OAI22_X1 port map( A1 => n8916, A2 => n24777, B1 => n20180, B2 => 
                           n24771, ZN => n21852);
   U21585 : AOI221_X1 port map( B1 => n24789, B2 => n8248, C1 => n24783, C2 => 
                           n8696, A => n21833, ZN => n21832);
   U21586 : OAI22_X1 port map( A1 => n8914, A2 => n24777, B1 => n20179, B2 => 
                           n24771, ZN => n21833);
   U21587 : AOI221_X1 port map( B1 => n24789, B2 => n8247, C1 => n24783, C2 => 
                           n8695, A => n21814, ZN => n21813);
   U21588 : OAI22_X1 port map( A1 => n8912, A2 => n24777, B1 => n20178, B2 => 
                           n24771, ZN => n21814);
   U21589 : AOI221_X1 port map( B1 => n24789, B2 => n8246, C1 => n24783, C2 => 
                           n8694, A => n21795, ZN => n21794);
   U21590 : OAI22_X1 port map( A1 => n8910, A2 => n24777, B1 => n20177, B2 => 
                           n24771, ZN => n21795);
   U21591 : AOI221_X1 port map( B1 => n24789, B2 => n8245, C1 => n24783, C2 => 
                           n8693, A => n21776, ZN => n21775);
   U21592 : OAI22_X1 port map( A1 => n8908, A2 => n24777, B1 => n20176, B2 => 
                           n24771, ZN => n21776);
   U21593 : AOI221_X1 port map( B1 => n24789, B2 => n8244, C1 => n24783, C2 => 
                           n8692, A => n21757, ZN => n21756);
   U21594 : OAI22_X1 port map( A1 => n8906, A2 => n24777, B1 => n20175, B2 => 
                           n24771, ZN => n21757);
   U21595 : AOI221_X1 port map( B1 => n24789, B2 => n8243, C1 => n24783, C2 => 
                           n8691, A => n21738, ZN => n21737);
   U21596 : OAI22_X1 port map( A1 => n8904, A2 => n24777, B1 => n20174, B2 => 
                           n24771, ZN => n21738);
   U21597 : AOI221_X1 port map( B1 => n24789, B2 => n8242, C1 => n24783, C2 => 
                           n8690, A => n21719, ZN => n21718);
   U21598 : OAI22_X1 port map( A1 => n8902, A2 => n24777, B1 => n20173, B2 => 
                           n24771, ZN => n21719);
   U21599 : AOI221_X1 port map( B1 => n24789, B2 => n8241, C1 => n24783, C2 => 
                           n8689, A => n21700, ZN => n21699);
   U21600 : OAI22_X1 port map( A1 => n8900, A2 => n24777, B1 => n20172, B2 => 
                           n24771, ZN => n21700);
   U21601 : AOI221_X1 port map( B1 => n24789, B2 => n8240, C1 => n24783, C2 => 
                           n8688, A => n21681, ZN => n21680);
   U21602 : OAI22_X1 port map( A1 => n8898, A2 => n24777, B1 => n20171, B2 => 
                           n24771, ZN => n21681);
   U21603 : AOI221_X1 port map( B1 => n24789, B2 => n8239, C1 => n24783, C2 => 
                           n8687, A => n21662, ZN => n21661);
   U21604 : OAI22_X1 port map( A1 => n8896, A2 => n24777, B1 => n20170, B2 => 
                           n24771, ZN => n21662);
   U21605 : AOI221_X1 port map( B1 => n24789, B2 => n8238, C1 => n24783, C2 => 
                           n8686, A => n21643, ZN => n21642);
   U21606 : OAI22_X1 port map( A1 => n8894, A2 => n24777, B1 => n20169, B2 => 
                           n24771, ZN => n21643);
   U21607 : AOI221_X1 port map( B1 => n24790, B2 => n8237, C1 => n24784, C2 => 
                           n8685, A => n21624, ZN => n21623);
   U21608 : OAI22_X1 port map( A1 => n8892, A2 => n24778, B1 => n20168, B2 => 
                           n24772, ZN => n21624);
   U21609 : AOI221_X1 port map( B1 => n24790, B2 => n8236, C1 => n24784, C2 => 
                           n8684, A => n21605, ZN => n21604);
   U21610 : OAI22_X1 port map( A1 => n8890, A2 => n24778, B1 => n20167, B2 => 
                           n24772, ZN => n21605);
   U21611 : AOI221_X1 port map( B1 => n24790, B2 => n8235, C1 => n24784, C2 => 
                           n8683, A => n21586, ZN => n21585);
   U21612 : OAI22_X1 port map( A1 => n8888, A2 => n24778, B1 => n20166, B2 => 
                           n24772, ZN => n21586);
   U21613 : AOI221_X1 port map( B1 => n24790, B2 => n8234, C1 => n24784, C2 => 
                           n8682, A => n21567, ZN => n21566);
   U21614 : OAI22_X1 port map( A1 => n8886, A2 => n24778, B1 => n20165, B2 => 
                           n24772, ZN => n21567);
   U21615 : AOI221_X1 port map( B1 => n24790, B2 => n8233, C1 => n24784, C2 => 
                           n8681, A => n21548, ZN => n21547);
   U21616 : OAI22_X1 port map( A1 => n8884, A2 => n24778, B1 => n20164, B2 => 
                           n24772, ZN => n21548);
   U21617 : AOI221_X1 port map( B1 => n24790, B2 => n8232, C1 => n24784, C2 => 
                           n8680, A => n21529, ZN => n21528);
   U21618 : OAI22_X1 port map( A1 => n8882, A2 => n24778, B1 => n20163, B2 => 
                           n24772, ZN => n21529);
   U21619 : AOI221_X1 port map( B1 => n24790, B2 => n8231, C1 => n24784, C2 => 
                           n8679, A => n21510, ZN => n21509);
   U21620 : OAI22_X1 port map( A1 => n8880, A2 => n24778, B1 => n20162, B2 => 
                           n24772, ZN => n21510);
   U21621 : AOI221_X1 port map( B1 => n24790, B2 => n8230, C1 => n24784, C2 => 
                           n8678, A => n21491, ZN => n21490);
   U21622 : OAI22_X1 port map( A1 => n8878, A2 => n24778, B1 => n20161, B2 => 
                           n24772, ZN => n21491);
   U21623 : AOI221_X1 port map( B1 => n24790, B2 => n8229, C1 => n24784, C2 => 
                           n8677, A => n21472, ZN => n21471);
   U21624 : OAI22_X1 port map( A1 => n8876, A2 => n24778, B1 => n20160, B2 => 
                           n24772, ZN => n21472);
   U21625 : AOI221_X1 port map( B1 => n24790, B2 => n8228, C1 => n24784, C2 => 
                           n8676, A => n21453, ZN => n21452);
   U21626 : OAI22_X1 port map( A1 => n8874, A2 => n24778, B1 => n20159, B2 => 
                           n24772, ZN => n21453);
   U21627 : AOI221_X1 port map( B1 => n24790, B2 => n8227, C1 => n24784, C2 => 
                           n8675, A => n21434, ZN => n21433);
   U21628 : OAI22_X1 port map( A1 => n8872, A2 => n24778, B1 => n20158, B2 => 
                           n24772, ZN => n21434);
   U21629 : AOI221_X1 port map( B1 => n24790, B2 => n8226, C1 => n24784, C2 => 
                           n8674, A => n21415, ZN => n21414);
   U21630 : OAI22_X1 port map( A1 => n8870, A2 => n24778, B1 => n20157, B2 => 
                           n24772, ZN => n21415);
   U21631 : AOI221_X1 port map( B1 => n24791, B2 => n8225, C1 => n24785, C2 => 
                           n8673, A => n21396, ZN => n21395);
   U21632 : OAI22_X1 port map( A1 => n8868, A2 => n24779, B1 => n20148, B2 => 
                           n24773, ZN => n21396);
   U21633 : AOI221_X1 port map( B1 => n24791, B2 => n8224, C1 => n24785, C2 => 
                           n8672, A => n21377, ZN => n21376);
   U21634 : OAI22_X1 port map( A1 => n8866, A2 => n24779, B1 => n20147, B2 => 
                           n24773, ZN => n21377);
   U21635 : AOI221_X1 port map( B1 => n24791, B2 => n8223, C1 => n24785, C2 => 
                           n8671, A => n21358, ZN => n21357);
   U21636 : OAI22_X1 port map( A1 => n8864, A2 => n24779, B1 => n20146, B2 => 
                           n24773, ZN => n21358);
   U21637 : AOI221_X1 port map( B1 => n24791, B2 => n8222, C1 => n24785, C2 => 
                           n8670, A => n21309, ZN => n21306);
   U21638 : OAI22_X1 port map( A1 => n8862, A2 => n24779, B1 => n20145, B2 => 
                           n24773, ZN => n21309);
   U21639 : AOI221_X1 port map( B1 => n24690, B2 => n20073, C1 => n24684, C2 =>
                           n19523, A => n22552, ZN => n22551);
   U21640 : OAI22_X1 port map( A1 => n896, A2 => n24678, B1 => n21074, B2 => 
                           n24672, ZN => n22552);
   U21641 : AOI221_X1 port map( B1 => n24690, B2 => n20072, C1 => n24684, C2 =>
                           n19522, A => n22525, ZN => n22524);
   U21642 : OAI22_X1 port map( A1 => n895, A2 => n24678, B1 => n21073, B2 => 
                           n24672, ZN => n22525);
   U21643 : AOI221_X1 port map( B1 => n24690, B2 => n20071, C1 => n24684, C2 =>
                           n19521, A => n22506, ZN => n22505);
   U21644 : OAI22_X1 port map( A1 => n894, A2 => n24678, B1 => n21072, B2 => 
                           n24672, ZN => n22506);
   U21645 : AOI221_X1 port map( B1 => n24690, B2 => n20070, C1 => n24684, C2 =>
                           n19520, A => n22487, ZN => n22486);
   U21646 : OAI22_X1 port map( A1 => n893, A2 => n24678, B1 => n21071, B2 => 
                           n24672, ZN => n22487);
   U21647 : AOI221_X1 port map( B1 => n24690, B2 => n20069, C1 => n24684, C2 =>
                           n19519, A => n22468, ZN => n22467);
   U21648 : OAI22_X1 port map( A1 => n892, A2 => n24678, B1 => n21070, B2 => 
                           n24672, ZN => n22468);
   U21649 : AOI221_X1 port map( B1 => n24690, B2 => n20068, C1 => n24684, C2 =>
                           n19518, A => n22449, ZN => n22448);
   U21650 : OAI22_X1 port map( A1 => n891, A2 => n24678, B1 => n21069, B2 => 
                           n24672, ZN => n22449);
   U21651 : AOI221_X1 port map( B1 => n24690, B2 => n20067, C1 => n24684, C2 =>
                           n19517, A => n22430, ZN => n22429);
   U21652 : OAI22_X1 port map( A1 => n890, A2 => n24678, B1 => n21068, B2 => 
                           n24672, ZN => n22430);
   U21653 : AOI221_X1 port map( B1 => n24690, B2 => n20066, C1 => n24684, C2 =>
                           n19516, A => n22411, ZN => n22410);
   U21654 : OAI22_X1 port map( A1 => n889, A2 => n24678, B1 => n21067, B2 => 
                           n24672, ZN => n22411);
   U21655 : AOI221_X1 port map( B1 => n24690, B2 => n20065, C1 => n24684, C2 =>
                           n19515, A => n22392, ZN => n22391);
   U21656 : OAI22_X1 port map( A1 => n888, A2 => n24678, B1 => n21066, B2 => 
                           n24672, ZN => n22392);
   U21657 : AOI221_X1 port map( B1 => n24690, B2 => n20064, C1 => n24684, C2 =>
                           n19514, A => n22373, ZN => n22372);
   U21658 : OAI22_X1 port map( A1 => n887, A2 => n24678, B1 => n21065, B2 => 
                           n24672, ZN => n22373);
   U21659 : AOI221_X1 port map( B1 => n24690, B2 => n20063, C1 => n24684, C2 =>
                           n19513, A => n22354, ZN => n22353);
   U21660 : OAI22_X1 port map( A1 => n886, A2 => n24678, B1 => n21064, B2 => 
                           n24672, ZN => n22354);
   U21661 : AOI221_X1 port map( B1 => n24690, B2 => n20062, C1 => n24684, C2 =>
                           n19512, A => n22335, ZN => n22334);
   U21662 : OAI22_X1 port map( A1 => n885, A2 => n24678, B1 => n21063, B2 => 
                           n24672, ZN => n22335);
   U21663 : AOI221_X1 port map( B1 => n24691, B2 => n20061, C1 => n24685, C2 =>
                           n19511, A => n22316, ZN => n22315);
   U21664 : OAI22_X1 port map( A1 => n884, A2 => n24679, B1 => n21062, B2 => 
                           n24673, ZN => n22316);
   U21665 : AOI221_X1 port map( B1 => n24691, B2 => n20060, C1 => n24685, C2 =>
                           n19510, A => n22297, ZN => n22296);
   U21666 : OAI22_X1 port map( A1 => n883, A2 => n24679, B1 => n21061, B2 => 
                           n24673, ZN => n22297);
   U21667 : AOI221_X1 port map( B1 => n24691, B2 => n20059, C1 => n24685, C2 =>
                           n19509, A => n22278, ZN => n22277);
   U21668 : OAI22_X1 port map( A1 => n882, A2 => n24679, B1 => n21060, B2 => 
                           n24673, ZN => n22278);
   U21669 : AOI221_X1 port map( B1 => n24691, B2 => n20058, C1 => n24685, C2 =>
                           n19508, A => n22259, ZN => n22258);
   U21670 : OAI22_X1 port map( A1 => n881, A2 => n24679, B1 => n21059, B2 => 
                           n24673, ZN => n22259);
   U21671 : AOI221_X1 port map( B1 => n24691, B2 => n20057, C1 => n24685, C2 =>
                           n19507, A => n22240, ZN => n22239);
   U21672 : OAI22_X1 port map( A1 => n880, A2 => n24679, B1 => n21058, B2 => 
                           n24673, ZN => n22240);
   U21673 : AOI221_X1 port map( B1 => n24691, B2 => n20056, C1 => n24685, C2 =>
                           n19506, A => n22221, ZN => n22220);
   U21674 : OAI22_X1 port map( A1 => n879, A2 => n24679, B1 => n21057, B2 => 
                           n24673, ZN => n22221);
   U21675 : AOI221_X1 port map( B1 => n24691, B2 => n20055, C1 => n24685, C2 =>
                           n19505, A => n22202, ZN => n22201);
   U21676 : OAI22_X1 port map( A1 => n878, A2 => n24679, B1 => n21056, B2 => 
                           n24673, ZN => n22202);
   U21677 : AOI221_X1 port map( B1 => n24691, B2 => n20054, C1 => n24685, C2 =>
                           n19504, A => n22183, ZN => n22182);
   U21678 : OAI22_X1 port map( A1 => n877, A2 => n24679, B1 => n21055, B2 => 
                           n24673, ZN => n22183);
   U21679 : AOI221_X1 port map( B1 => n24691, B2 => n20053, C1 => n24685, C2 =>
                           n19503, A => n22164, ZN => n22163);
   U21680 : OAI22_X1 port map( A1 => n876, A2 => n24679, B1 => n21054, B2 => 
                           n24673, ZN => n22164);
   U21681 : AOI221_X1 port map( B1 => n24691, B2 => n20052, C1 => n24685, C2 =>
                           n19502, A => n22145, ZN => n22144);
   U21682 : OAI22_X1 port map( A1 => n875, A2 => n24679, B1 => n21053, B2 => 
                           n24673, ZN => n22145);
   U21683 : AOI221_X1 port map( B1 => n24691, B2 => n20051, C1 => n24685, C2 =>
                           n19501, A => n22126, ZN => n22125);
   U21684 : OAI22_X1 port map( A1 => n874, A2 => n24679, B1 => n21052, B2 => 
                           n24673, ZN => n22126);
   U21685 : AOI221_X1 port map( B1 => n24691, B2 => n20050, C1 => n24685, C2 =>
                           n19500, A => n22107, ZN => n22106);
   U21686 : OAI22_X1 port map( A1 => n873, A2 => n24679, B1 => n21051, B2 => 
                           n24673, ZN => n22107);
   U21687 : AOI221_X1 port map( B1 => n24692, B2 => n19929, C1 => n24686, C2 =>
                           n19499, A => n22088, ZN => n22087);
   U21688 : OAI22_X1 port map( A1 => n872, A2 => n24680, B1 => n20942, B2 => 
                           n24674, ZN => n22088);
   U21689 : AOI221_X1 port map( B1 => n24692, B2 => n19928, C1 => n24686, C2 =>
                           n19498, A => n22069, ZN => n22068);
   U21690 : OAI22_X1 port map( A1 => n871, A2 => n24680, B1 => n20941, B2 => 
                           n24674, ZN => n22069);
   U21691 : AOI221_X1 port map( B1 => n24692, B2 => n19927, C1 => n24686, C2 =>
                           n19497, A => n22050, ZN => n22049);
   U21692 : OAI22_X1 port map( A1 => n870, A2 => n24680, B1 => n20940, B2 => 
                           n24674, ZN => n22050);
   U21693 : AOI221_X1 port map( B1 => n24692, B2 => n19926, C1 => n24686, C2 =>
                           n19496, A => n22031, ZN => n22030);
   U21694 : OAI22_X1 port map( A1 => n869, A2 => n24680, B1 => n20939, B2 => 
                           n24674, ZN => n22031);
   U21695 : AOI221_X1 port map( B1 => n24692, B2 => n19925, C1 => n24686, C2 =>
                           n19495, A => n22012, ZN => n22011);
   U21696 : OAI22_X1 port map( A1 => n868, A2 => n24680, B1 => n20938, B2 => 
                           n24674, ZN => n22012);
   U21697 : AOI221_X1 port map( B1 => n24692, B2 => n19924, C1 => n24686, C2 =>
                           n19494, A => n21993, ZN => n21992);
   U21698 : OAI22_X1 port map( A1 => n867, A2 => n24680, B1 => n20937, B2 => 
                           n24674, ZN => n21993);
   U21699 : AOI221_X1 port map( B1 => n24692, B2 => n19923, C1 => n24686, C2 =>
                           n19493, A => n21974, ZN => n21973);
   U21700 : OAI22_X1 port map( A1 => n866, A2 => n24680, B1 => n20936, B2 => 
                           n24674, ZN => n21974);
   U21701 : AOI221_X1 port map( B1 => n24692, B2 => n19922, C1 => n24686, C2 =>
                           n19492, A => n21955, ZN => n21954);
   U21702 : OAI22_X1 port map( A1 => n865, A2 => n24680, B1 => n20935, B2 => 
                           n24674, ZN => n21955);
   U21703 : AOI221_X1 port map( B1 => n24692, B2 => n19921, C1 => n24686, C2 =>
                           n19491, A => n21936, ZN => n21935);
   U21704 : OAI22_X1 port map( A1 => n864, A2 => n24680, B1 => n20934, B2 => 
                           n24674, ZN => n21936);
   U21705 : AOI221_X1 port map( B1 => n24692, B2 => n19920, C1 => n24686, C2 =>
                           n19490, A => n21917, ZN => n21916);
   U21706 : OAI22_X1 port map( A1 => n863, A2 => n24680, B1 => n20933, B2 => 
                           n24674, ZN => n21917);
   U21707 : AOI221_X1 port map( B1 => n24692, B2 => n19919, C1 => n24686, C2 =>
                           n19489, A => n21898, ZN => n21897);
   U21708 : OAI22_X1 port map( A1 => n862, A2 => n24680, B1 => n20932, B2 => 
                           n24674, ZN => n21898);
   U21709 : AOI221_X1 port map( B1 => n24692, B2 => n19918, C1 => n24686, C2 =>
                           n19488, A => n21879, ZN => n21878);
   U21710 : OAI22_X1 port map( A1 => n861, A2 => n24680, B1 => n20931, B2 => 
                           n24674, ZN => n21879);
   U21711 : AOI221_X1 port map( B1 => n24693, B2 => n19917, C1 => n24687, C2 =>
                           n19487, A => n21860, ZN => n21859);
   U21712 : OAI22_X1 port map( A1 => n860, A2 => n24681, B1 => n20930, B2 => 
                           n24675, ZN => n21860);
   U21713 : AOI221_X1 port map( B1 => n24693, B2 => n19916, C1 => n24687, C2 =>
                           n19486, A => n21841, ZN => n21840);
   U21714 : OAI22_X1 port map( A1 => n859, A2 => n24681, B1 => n20929, B2 => 
                           n24675, ZN => n21841);
   U21715 : AOI221_X1 port map( B1 => n24693, B2 => n19915, C1 => n24687, C2 =>
                           n19485, A => n21822, ZN => n21821);
   U21716 : OAI22_X1 port map( A1 => n858, A2 => n24681, B1 => n20928, B2 => 
                           n24675, ZN => n21822);
   U21717 : AOI221_X1 port map( B1 => n24693, B2 => n19914, C1 => n24687, C2 =>
                           n19484, A => n21803, ZN => n21802);
   U21718 : OAI22_X1 port map( A1 => n857, A2 => n24681, B1 => n20927, B2 => 
                           n24675, ZN => n21803);
   U21719 : AOI221_X1 port map( B1 => n24693, B2 => n19913, C1 => n24687, C2 =>
                           n19483, A => n21784, ZN => n21783);
   U21720 : OAI22_X1 port map( A1 => n856, A2 => n24681, B1 => n20926, B2 => 
                           n24675, ZN => n21784);
   U21721 : AOI221_X1 port map( B1 => n24693, B2 => n19912, C1 => n24687, C2 =>
                           n19482, A => n21765, ZN => n21764);
   U21722 : OAI22_X1 port map( A1 => n855, A2 => n24681, B1 => n20925, B2 => 
                           n24675, ZN => n21765);
   U21723 : AOI221_X1 port map( B1 => n24693, B2 => n19911, C1 => n24687, C2 =>
                           n19481, A => n21746, ZN => n21745);
   U21724 : OAI22_X1 port map( A1 => n854, A2 => n24681, B1 => n20924, B2 => 
                           n24675, ZN => n21746);
   U21725 : AOI221_X1 port map( B1 => n24693, B2 => n19910, C1 => n24687, C2 =>
                           n19480, A => n21727, ZN => n21726);
   U21726 : OAI22_X1 port map( A1 => n853, A2 => n24681, B1 => n20923, B2 => 
                           n24675, ZN => n21727);
   U21727 : AOI221_X1 port map( B1 => n24693, B2 => n19909, C1 => n24687, C2 =>
                           n19479, A => n21708, ZN => n21707);
   U21728 : OAI22_X1 port map( A1 => n852, A2 => n24681, B1 => n20922, B2 => 
                           n24675, ZN => n21708);
   U21729 : AOI221_X1 port map( B1 => n24693, B2 => n19908, C1 => n24687, C2 =>
                           n19478, A => n21689, ZN => n21688);
   U21730 : OAI22_X1 port map( A1 => n851, A2 => n24681, B1 => n20921, B2 => 
                           n24675, ZN => n21689);
   U21731 : AOI221_X1 port map( B1 => n24693, B2 => n19907, C1 => n24687, C2 =>
                           n19477, A => n21670, ZN => n21669);
   U21732 : OAI22_X1 port map( A1 => n850, A2 => n24681, B1 => n20920, B2 => 
                           n24675, ZN => n21670);
   U21733 : AOI221_X1 port map( B1 => n24693, B2 => n19906, C1 => n24687, C2 =>
                           n19476, A => n21651, ZN => n21650);
   U21734 : OAI22_X1 port map( A1 => n849, A2 => n24681, B1 => n20919, B2 => 
                           n24675, ZN => n21651);
   U21735 : AOI221_X1 port map( B1 => n24694, B2 => n19905, C1 => n24688, C2 =>
                           n19475, A => n21632, ZN => n21631);
   U21736 : OAI22_X1 port map( A1 => n848, A2 => n24682, B1 => n20918, B2 => 
                           n24676, ZN => n21632);
   U21737 : AOI221_X1 port map( B1 => n24694, B2 => n19904, C1 => n24688, C2 =>
                           n19474, A => n21613, ZN => n21612);
   U21738 : OAI22_X1 port map( A1 => n847, A2 => n24682, B1 => n20917, B2 => 
                           n24676, ZN => n21613);
   U21739 : AOI221_X1 port map( B1 => n24694, B2 => n19903, C1 => n24688, C2 =>
                           n19473, A => n21594, ZN => n21593);
   U21740 : OAI22_X1 port map( A1 => n846, A2 => n24682, B1 => n20916, B2 => 
                           n24676, ZN => n21594);
   U21741 : AOI221_X1 port map( B1 => n24694, B2 => n19902, C1 => n24688, C2 =>
                           n19472, A => n21575, ZN => n21574);
   U21742 : OAI22_X1 port map( A1 => n845, A2 => n24682, B1 => n20915, B2 => 
                           n24676, ZN => n21575);
   U21743 : AOI221_X1 port map( B1 => n24694, B2 => n19901, C1 => n24688, C2 =>
                           n19471, A => n21556, ZN => n21555);
   U21744 : OAI22_X1 port map( A1 => n844, A2 => n24682, B1 => n20914, B2 => 
                           n24676, ZN => n21556);
   U21745 : AOI221_X1 port map( B1 => n24694, B2 => n19900, C1 => n24688, C2 =>
                           n19470, A => n21537, ZN => n21536);
   U21746 : OAI22_X1 port map( A1 => n843, A2 => n24682, B1 => n20913, B2 => 
                           n24676, ZN => n21537);
   U21747 : AOI221_X1 port map( B1 => n24694, B2 => n19899, C1 => n24688, C2 =>
                           n19469, A => n21518, ZN => n21517);
   U21748 : OAI22_X1 port map( A1 => n842, A2 => n24682, B1 => n20912, B2 => 
                           n24676, ZN => n21518);
   U21749 : AOI221_X1 port map( B1 => n24694, B2 => n19898, C1 => n24688, C2 =>
                           n19468, A => n21499, ZN => n21498);
   U21750 : OAI22_X1 port map( A1 => n841, A2 => n24682, B1 => n20911, B2 => 
                           n24676, ZN => n21499);
   U21751 : AOI221_X1 port map( B1 => n24694, B2 => n19897, C1 => n24688, C2 =>
                           n19467, A => n21480, ZN => n21479);
   U21752 : OAI22_X1 port map( A1 => n840, A2 => n24682, B1 => n20910, B2 => 
                           n24676, ZN => n21480);
   U21753 : AOI221_X1 port map( B1 => n24694, B2 => n19896, C1 => n24688, C2 =>
                           n19466, A => n21461, ZN => n21460);
   U21754 : OAI22_X1 port map( A1 => n839, A2 => n24682, B1 => n20909, B2 => 
                           n24676, ZN => n21461);
   U21755 : AOI221_X1 port map( B1 => n24694, B2 => n19895, C1 => n24688, C2 =>
                           n19465, A => n21442, ZN => n21441);
   U21756 : OAI22_X1 port map( A1 => n838, A2 => n24682, B1 => n20908, B2 => 
                           n24676, ZN => n21442);
   U21757 : AOI221_X1 port map( B1 => n24694, B2 => n19894, C1 => n24688, C2 =>
                           n19464, A => n21423, ZN => n21422);
   U21758 : OAI22_X1 port map( A1 => n837, A2 => n24682, B1 => n20907, B2 => 
                           n24676, ZN => n21423);
   U21759 : AOI221_X1 port map( B1 => n24695, B2 => n19813, C1 => n24689, C2 =>
                           n19463, A => n21404, ZN => n21403);
   U21760 : OAI22_X1 port map( A1 => n836, A2 => n24683, B1 => n20534, B2 => 
                           n24677, ZN => n21404);
   U21761 : AOI221_X1 port map( B1 => n24695, B2 => n19812, C1 => n24689, C2 =>
                           n19462, A => n21385, ZN => n21384);
   U21762 : OAI22_X1 port map( A1 => n835, A2 => n24683, B1 => n20533, B2 => 
                           n24677, ZN => n21385);
   U21763 : AOI221_X1 port map( B1 => n24695, B2 => n19811, C1 => n24689, C2 =>
                           n19461, A => n21366, ZN => n21365);
   U21764 : OAI22_X1 port map( A1 => n834, A2 => n24683, B1 => n20532, B2 => 
                           n24677, ZN => n21366);
   U21765 : AOI221_X1 port map( B1 => n24695, B2 => n19810, C1 => n24689, C2 =>
                           n19460, A => n21333, ZN => n21330);
   U21766 : OAI22_X1 port map( A1 => n833, A2 => n24683, B1 => n20531, B2 => 
                           n24677, ZN => n21333);
   U21767 : AOI221_X1 port map( B1 => n24762, B2 => n8029, C1 => n24756, C2 => 
                           n8413, A => n22541, ZN => n22534);
   U21768 : OAI22_X1 port map( A1 => n7427, A2 => n24750, B1 => n19707, B2 => 
                           n24744, ZN => n22541);
   U21769 : AOI221_X1 port map( B1 => n24762, B2 => n8028, C1 => n24756, C2 => 
                           n8412, A => n22518, ZN => n22515);
   U21770 : OAI22_X1 port map( A1 => n7425, A2 => n24750, B1 => n19706, B2 => 
                           n24744, ZN => n22518);
   U21771 : AOI221_X1 port map( B1 => n24762, B2 => n8027, C1 => n24756, C2 => 
                           n8411, A => n22499, ZN => n22496);
   U21772 : OAI22_X1 port map( A1 => n7423, A2 => n24750, B1 => n19705, B2 => 
                           n24744, ZN => n22499);
   U21773 : AOI221_X1 port map( B1 => n24762, B2 => n8026, C1 => n24756, C2 => 
                           n8410, A => n22480, ZN => n22477);
   U21774 : OAI22_X1 port map( A1 => n7421, A2 => n24750, B1 => n19704, B2 => 
                           n24744, ZN => n22480);
   U21775 : AOI221_X1 port map( B1 => n24762, B2 => n8025, C1 => n24756, C2 => 
                           n8409, A => n22461, ZN => n22458);
   U21776 : OAI22_X1 port map( A1 => n7419, A2 => n24750, B1 => n19703, B2 => 
                           n24744, ZN => n22461);
   U21777 : AOI221_X1 port map( B1 => n24762, B2 => n8024, C1 => n24756, C2 => 
                           n8408, A => n22442, ZN => n22439);
   U21778 : OAI22_X1 port map( A1 => n7417, A2 => n24750, B1 => n19702, B2 => 
                           n24744, ZN => n22442);
   U21779 : AOI221_X1 port map( B1 => n24762, B2 => n8023, C1 => n24756, C2 => 
                           n8407, A => n22423, ZN => n22420);
   U21780 : OAI22_X1 port map( A1 => n7415, A2 => n24750, B1 => n19701, B2 => 
                           n24744, ZN => n22423);
   U21781 : AOI221_X1 port map( B1 => n24762, B2 => n8022, C1 => n24756, C2 => 
                           n8406, A => n22404, ZN => n22401);
   U21782 : OAI22_X1 port map( A1 => n7413, A2 => n24750, B1 => n19700, B2 => 
                           n24744, ZN => n22404);
   U21783 : AOI221_X1 port map( B1 => n24762, B2 => n8021, C1 => n24756, C2 => 
                           n8405, A => n22385, ZN => n22382);
   U21784 : OAI22_X1 port map( A1 => n7411, A2 => n24750, B1 => n19699, B2 => 
                           n24744, ZN => n22385);
   U21785 : AOI221_X1 port map( B1 => n24762, B2 => n8020, C1 => n24756, C2 => 
                           n8404, A => n22366, ZN => n22363);
   U21786 : OAI22_X1 port map( A1 => n7409, A2 => n24750, B1 => n19698, B2 => 
                           n24744, ZN => n22366);
   U21787 : AOI221_X1 port map( B1 => n24762, B2 => n8019, C1 => n24756, C2 => 
                           n8403, A => n22347, ZN => n22344);
   U21788 : OAI22_X1 port map( A1 => n7407, A2 => n24750, B1 => n19697, B2 => 
                           n24744, ZN => n22347);
   U21789 : AOI221_X1 port map( B1 => n24762, B2 => n8018, C1 => n24756, C2 => 
                           n8402, A => n22328, ZN => n22325);
   U21790 : OAI22_X1 port map( A1 => n7405, A2 => n24750, B1 => n19696, B2 => 
                           n24744, ZN => n22328);
   U21791 : AOI221_X1 port map( B1 => n24763, B2 => n8017, C1 => n24757, C2 => 
                           n8401, A => n22309, ZN => n22306);
   U21792 : OAI22_X1 port map( A1 => n7403, A2 => n24751, B1 => n19695, B2 => 
                           n24745, ZN => n22309);
   U21793 : AOI221_X1 port map( B1 => n24763, B2 => n8016, C1 => n24757, C2 => 
                           n8400, A => n22290, ZN => n22287);
   U21794 : OAI22_X1 port map( A1 => n7401, A2 => n24751, B1 => n19694, B2 => 
                           n24745, ZN => n22290);
   U21795 : AOI221_X1 port map( B1 => n24763, B2 => n8015, C1 => n24757, C2 => 
                           n8399, A => n22271, ZN => n22268);
   U21796 : OAI22_X1 port map( A1 => n7399, A2 => n24751, B1 => n19693, B2 => 
                           n24745, ZN => n22271);
   U21797 : AOI221_X1 port map( B1 => n24763, B2 => n8014, C1 => n24757, C2 => 
                           n8398, A => n22252, ZN => n22249);
   U21798 : OAI22_X1 port map( A1 => n7397, A2 => n24751, B1 => n19692, B2 => 
                           n24745, ZN => n22252);
   U21799 : AOI221_X1 port map( B1 => n24763, B2 => n8013, C1 => n24757, C2 => 
                           n8397, A => n22233, ZN => n22230);
   U21800 : OAI22_X1 port map( A1 => n7395, A2 => n24751, B1 => n19691, B2 => 
                           n24745, ZN => n22233);
   U21801 : AOI221_X1 port map( B1 => n24763, B2 => n8012, C1 => n24757, C2 => 
                           n8396, A => n22214, ZN => n22211);
   U21802 : OAI22_X1 port map( A1 => n7393, A2 => n24751, B1 => n19690, B2 => 
                           n24745, ZN => n22214);
   U21803 : AOI221_X1 port map( B1 => n24763, B2 => n8011, C1 => n24757, C2 => 
                           n8395, A => n22195, ZN => n22192);
   U21804 : OAI22_X1 port map( A1 => n7391, A2 => n24751, B1 => n19689, B2 => 
                           n24745, ZN => n22195);
   U21805 : AOI221_X1 port map( B1 => n24763, B2 => n8010, C1 => n24757, C2 => 
                           n8394, A => n22176, ZN => n22173);
   U21806 : OAI22_X1 port map( A1 => n7389, A2 => n24751, B1 => n19688, B2 => 
                           n24745, ZN => n22176);
   U21807 : AOI221_X1 port map( B1 => n24763, B2 => n8009, C1 => n24757, C2 => 
                           n8393, A => n22157, ZN => n22154);
   U21808 : OAI22_X1 port map( A1 => n7387, A2 => n24751, B1 => n19687, B2 => 
                           n24745, ZN => n22157);
   U21809 : AOI221_X1 port map( B1 => n24763, B2 => n8008, C1 => n24757, C2 => 
                           n8392, A => n22138, ZN => n22135);
   U21810 : OAI22_X1 port map( A1 => n7385, A2 => n24751, B1 => n19686, B2 => 
                           n24745, ZN => n22138);
   U21811 : AOI221_X1 port map( B1 => n24763, B2 => n8007, C1 => n24757, C2 => 
                           n8391, A => n22119, ZN => n22116);
   U21812 : OAI22_X1 port map( A1 => n7383, A2 => n24751, B1 => n19685, B2 => 
                           n24745, ZN => n22119);
   U21813 : AOI221_X1 port map( B1 => n24763, B2 => n8006, C1 => n24757, C2 => 
                           n8390, A => n22100, ZN => n22097);
   U21814 : OAI22_X1 port map( A1 => n7381, A2 => n24751, B1 => n19684, B2 => 
                           n24745, ZN => n22100);
   U21815 : AOI221_X1 port map( B1 => n24764, B2 => n8005, C1 => n24758, C2 => 
                           n8389, A => n22081, ZN => n22078);
   U21816 : OAI22_X1 port map( A1 => n7379, A2 => n24752, B1 => n19683, B2 => 
                           n24746, ZN => n22081);
   U21817 : AOI221_X1 port map( B1 => n24764, B2 => n8004, C1 => n24758, C2 => 
                           n8388, A => n22062, ZN => n22059);
   U21818 : OAI22_X1 port map( A1 => n7377, A2 => n24752, B1 => n19682, B2 => 
                           n24746, ZN => n22062);
   U21819 : AOI221_X1 port map( B1 => n24764, B2 => n8003, C1 => n24758, C2 => 
                           n8387, A => n22043, ZN => n22040);
   U21820 : OAI22_X1 port map( A1 => n7375, A2 => n24752, B1 => n19681, B2 => 
                           n24746, ZN => n22043);
   U21821 : AOI221_X1 port map( B1 => n24764, B2 => n8002, C1 => n24758, C2 => 
                           n8386, A => n22024, ZN => n22021);
   U21822 : OAI22_X1 port map( A1 => n7373, A2 => n24752, B1 => n19680, B2 => 
                           n24746, ZN => n22024);
   U21823 : AOI221_X1 port map( B1 => n24764, B2 => n8001, C1 => n24758, C2 => 
                           n8385, A => n22005, ZN => n22002);
   U21824 : OAI22_X1 port map( A1 => n7371, A2 => n24752, B1 => n19679, B2 => 
                           n24746, ZN => n22005);
   U21825 : AOI221_X1 port map( B1 => n24764, B2 => n8000, C1 => n24758, C2 => 
                           n8384, A => n21986, ZN => n21983);
   U21826 : OAI22_X1 port map( A1 => n7369, A2 => n24752, B1 => n19678, B2 => 
                           n24746, ZN => n21986);
   U21827 : AOI221_X1 port map( B1 => n24764, B2 => n7999, C1 => n24758, C2 => 
                           n8383, A => n21967, ZN => n21964);
   U21828 : OAI22_X1 port map( A1 => n7367, A2 => n24752, B1 => n19677, B2 => 
                           n24746, ZN => n21967);
   U21829 : AOI221_X1 port map( B1 => n24764, B2 => n7998, C1 => n24758, C2 => 
                           n8382, A => n21948, ZN => n21945);
   U21830 : OAI22_X1 port map( A1 => n7365, A2 => n24752, B1 => n19676, B2 => 
                           n24746, ZN => n21948);
   U21831 : AOI221_X1 port map( B1 => n24764, B2 => n7997, C1 => n24758, C2 => 
                           n8381, A => n21929, ZN => n21926);
   U21832 : OAI22_X1 port map( A1 => n7363, A2 => n24752, B1 => n19675, B2 => 
                           n24746, ZN => n21929);
   U21833 : AOI221_X1 port map( B1 => n24764, B2 => n7996, C1 => n24758, C2 => 
                           n8380, A => n21910, ZN => n21907);
   U21834 : OAI22_X1 port map( A1 => n7361, A2 => n24752, B1 => n19674, B2 => 
                           n24746, ZN => n21910);
   U21835 : AOI221_X1 port map( B1 => n24764, B2 => n7995, C1 => n24758, C2 => 
                           n8379, A => n21891, ZN => n21888);
   U21836 : OAI22_X1 port map( A1 => n7359, A2 => n24752, B1 => n19673, B2 => 
                           n24746, ZN => n21891);
   U21837 : AOI221_X1 port map( B1 => n24764, B2 => n7994, C1 => n24758, C2 => 
                           n8378, A => n21872, ZN => n21869);
   U21838 : OAI22_X1 port map( A1 => n7357, A2 => n24752, B1 => n19672, B2 => 
                           n24746, ZN => n21872);
   U21839 : AOI221_X1 port map( B1 => n24765, B2 => n7993, C1 => n24759, C2 => 
                           n8377, A => n21853, ZN => n21850);
   U21840 : OAI22_X1 port map( A1 => n7355, A2 => n24753, B1 => n19671, B2 => 
                           n24747, ZN => n21853);
   U21841 : AOI221_X1 port map( B1 => n24765, B2 => n7992, C1 => n24759, C2 => 
                           n8376, A => n21834, ZN => n21831);
   U21842 : OAI22_X1 port map( A1 => n7353, A2 => n24753, B1 => n19670, B2 => 
                           n24747, ZN => n21834);
   U21843 : AOI221_X1 port map( B1 => n24765, B2 => n7991, C1 => n24759, C2 => 
                           n8375, A => n21815, ZN => n21812);
   U21844 : OAI22_X1 port map( A1 => n7351, A2 => n24753, B1 => n19669, B2 => 
                           n24747, ZN => n21815);
   U21845 : AOI221_X1 port map( B1 => n24765, B2 => n7990, C1 => n24759, C2 => 
                           n8374, A => n21796, ZN => n21793);
   U21846 : OAI22_X1 port map( A1 => n7349, A2 => n24753, B1 => n19668, B2 => 
                           n24747, ZN => n21796);
   U21847 : AOI221_X1 port map( B1 => n24765, B2 => n7989, C1 => n24759, C2 => 
                           n8373, A => n21777, ZN => n21774);
   U21848 : OAI22_X1 port map( A1 => n7347, A2 => n24753, B1 => n19667, B2 => 
                           n24747, ZN => n21777);
   U21849 : AOI221_X1 port map( B1 => n24765, B2 => n7988, C1 => n24759, C2 => 
                           n8372, A => n21758, ZN => n21755);
   U21850 : OAI22_X1 port map( A1 => n7345, A2 => n24753, B1 => n19666, B2 => 
                           n24747, ZN => n21758);
   U21851 : AOI221_X1 port map( B1 => n24765, B2 => n7987, C1 => n24759, C2 => 
                           n8371, A => n21739, ZN => n21736);
   U21852 : OAI22_X1 port map( A1 => n7343, A2 => n24753, B1 => n19665, B2 => 
                           n24747, ZN => n21739);
   U21853 : AOI221_X1 port map( B1 => n24765, B2 => n7986, C1 => n24759, C2 => 
                           n8370, A => n21720, ZN => n21717);
   U21854 : OAI22_X1 port map( A1 => n7341, A2 => n24753, B1 => n19664, B2 => 
                           n24747, ZN => n21720);
   U21855 : AOI221_X1 port map( B1 => n24765, B2 => n7985, C1 => n24759, C2 => 
                           n8369, A => n21701, ZN => n21698);
   U21856 : OAI22_X1 port map( A1 => n7339, A2 => n24753, B1 => n19663, B2 => 
                           n24747, ZN => n21701);
   U21857 : AOI221_X1 port map( B1 => n24765, B2 => n7984, C1 => n24759, C2 => 
                           n8368, A => n21682, ZN => n21679);
   U21858 : OAI22_X1 port map( A1 => n7337, A2 => n24753, B1 => n19662, B2 => 
                           n24747, ZN => n21682);
   U21859 : AOI221_X1 port map( B1 => n24765, B2 => n7983, C1 => n24759, C2 => 
                           n8367, A => n21663, ZN => n21660);
   U21860 : OAI22_X1 port map( A1 => n7335, A2 => n24753, B1 => n19661, B2 => 
                           n24747, ZN => n21663);
   U21861 : AOI221_X1 port map( B1 => n24765, B2 => n7982, C1 => n24759, C2 => 
                           n8366, A => n21644, ZN => n21641);
   U21862 : OAI22_X1 port map( A1 => n7333, A2 => n24753, B1 => n19660, B2 => 
                           n24747, ZN => n21644);
   U21863 : AOI221_X1 port map( B1 => n24766, B2 => n7981, C1 => n24760, C2 => 
                           n8365, A => n21625, ZN => n21622);
   U21864 : OAI22_X1 port map( A1 => n7331, A2 => n24754, B1 => n19659, B2 => 
                           n24748, ZN => n21625);
   U21865 : AOI221_X1 port map( B1 => n24766, B2 => n7980, C1 => n24760, C2 => 
                           n8364, A => n21606, ZN => n21603);
   U21866 : OAI22_X1 port map( A1 => n7329, A2 => n24754, B1 => n19658, B2 => 
                           n24748, ZN => n21606);
   U21867 : AOI221_X1 port map( B1 => n24766, B2 => n7979, C1 => n24760, C2 => 
                           n8363, A => n21587, ZN => n21584);
   U21868 : OAI22_X1 port map( A1 => n7327, A2 => n24754, B1 => n19657, B2 => 
                           n24748, ZN => n21587);
   U21869 : AOI221_X1 port map( B1 => n24766, B2 => n7978, C1 => n24760, C2 => 
                           n8362, A => n21568, ZN => n21565);
   U21870 : OAI22_X1 port map( A1 => n7325, A2 => n24754, B1 => n19656, B2 => 
                           n24748, ZN => n21568);
   U21871 : AOI221_X1 port map( B1 => n24766, B2 => n7977, C1 => n24760, C2 => 
                           n8361, A => n21549, ZN => n21546);
   U21872 : OAI22_X1 port map( A1 => n7323, A2 => n24754, B1 => n19655, B2 => 
                           n24748, ZN => n21549);
   U21873 : AOI221_X1 port map( B1 => n24766, B2 => n7976, C1 => n24760, C2 => 
                           n8360, A => n21530, ZN => n21527);
   U21874 : OAI22_X1 port map( A1 => n7321, A2 => n24754, B1 => n19654, B2 => 
                           n24748, ZN => n21530);
   U21875 : AOI221_X1 port map( B1 => n24766, B2 => n7975, C1 => n24760, C2 => 
                           n8359, A => n21511, ZN => n21508);
   U21876 : OAI22_X1 port map( A1 => n7319, A2 => n24754, B1 => n19653, B2 => 
                           n24748, ZN => n21511);
   U21877 : AOI221_X1 port map( B1 => n24766, B2 => n7974, C1 => n24760, C2 => 
                           n8358, A => n21492, ZN => n21489);
   U21878 : OAI22_X1 port map( A1 => n7317, A2 => n24754, B1 => n19652, B2 => 
                           n24748, ZN => n21492);
   U21879 : AOI221_X1 port map( B1 => n24766, B2 => n7973, C1 => n24760, C2 => 
                           n8357, A => n21473, ZN => n21470);
   U21880 : OAI22_X1 port map( A1 => n7315, A2 => n24754, B1 => n19651, B2 => 
                           n24748, ZN => n21473);
   U21881 : AOI221_X1 port map( B1 => n24766, B2 => n7972, C1 => n24760, C2 => 
                           n8356, A => n21454, ZN => n21451);
   U21882 : OAI22_X1 port map( A1 => n7313, A2 => n24754, B1 => n19650, B2 => 
                           n24748, ZN => n21454);
   U21883 : AOI221_X1 port map( B1 => n24766, B2 => n7971, C1 => n24760, C2 => 
                           n8355, A => n21435, ZN => n21432);
   U21884 : OAI22_X1 port map( A1 => n7311, A2 => n24754, B1 => n19649, B2 => 
                           n24748, ZN => n21435);
   U21885 : AOI221_X1 port map( B1 => n24766, B2 => n7970, C1 => n24760, C2 => 
                           n8354, A => n21416, ZN => n21413);
   U21886 : OAI22_X1 port map( A1 => n7309, A2 => n24754, B1 => n19648, B2 => 
                           n24748, ZN => n21416);
   U21887 : AOI221_X1 port map( B1 => n24767, B2 => n7969, C1 => n24761, C2 => 
                           n8353, A => n21397, ZN => n21394);
   U21888 : OAI22_X1 port map( A1 => n7307, A2 => n24755, B1 => n20152, B2 => 
                           n24749, ZN => n21397);
   U21889 : AOI221_X1 port map( B1 => n24767, B2 => n7968, C1 => n24761, C2 => 
                           n8352, A => n21378, ZN => n21375);
   U21890 : OAI22_X1 port map( A1 => n7305, A2 => n24755, B1 => n20151, B2 => 
                           n24749, ZN => n21378);
   U21891 : AOI221_X1 port map( B1 => n24767, B2 => n7967, C1 => n24761, C2 => 
                           n8351, A => n21359, ZN => n21356);
   U21892 : OAI22_X1 port map( A1 => n7303, A2 => n24755, B1 => n20150, B2 => 
                           n24749, ZN => n21359);
   U21893 : AOI221_X1 port map( B1 => n24767, B2 => n7966, C1 => n24761, C2 => 
                           n8350, A => n21314, ZN => n21305);
   U21894 : OAI22_X1 port map( A1 => n7301, A2 => n24755, B1 => n20149, B2 => 
                           n24749, ZN => n21314);
   U21895 : AOI221_X1 port map( B1 => n24671, B2 => n19399, C1 => n24665, C2 =>
                           n19817, A => n21405, ZN => n21402);
   U21896 : OAI22_X1 port map( A1 => n20257, A2 => n24659, B1 => n20538, B2 => 
                           n24653, ZN => n21405);
   U21897 : AOI221_X1 port map( B1 => n24671, B2 => n19398, C1 => n24665, C2 =>
                           n19816, A => n21386, ZN => n21383);
   U21898 : OAI22_X1 port map( A1 => n20256, A2 => n24659, B1 => n20537, B2 => 
                           n24653, ZN => n21386);
   U21899 : AOI221_X1 port map( B1 => n24671, B2 => n19397, C1 => n24665, C2 =>
                           n19815, A => n21367, ZN => n21364);
   U21900 : OAI22_X1 port map( A1 => n20255, A2 => n24659, B1 => n20536, B2 => 
                           n24653, ZN => n21367);
   U21901 : AOI221_X1 port map( B1 => n24671, B2 => n19396, C1 => n24665, C2 =>
                           n19814, A => n21338, ZN => n21329);
   U21902 : OAI22_X1 port map( A1 => n20254, A2 => n24659, B1 => n20535, B2 => 
                           n24653, ZN => n21338);
   U21903 : AOI221_X1 port map( B1 => n24738, B2 => n19647, C1 => n24732, C2 =>
                           n19587, A => n22544, ZN => n22533);
   U21904 : OAI22_X1 port map( A1 => n21146, A2 => n24726, B1 => n20798, B2 => 
                           n24720, ZN => n22544);
   U21905 : AOI221_X1 port map( B1 => n24738, B2 => n19646, C1 => n24732, C2 =>
                           n19586, A => n22519, ZN => n22514);
   U21906 : OAI22_X1 port map( A1 => n21145, A2 => n24726, B1 => n20797, B2 => 
                           n24720, ZN => n22519);
   U21907 : AOI221_X1 port map( B1 => n24738, B2 => n19645, C1 => n24732, C2 =>
                           n19585, A => n22500, ZN => n22495);
   U21908 : OAI22_X1 port map( A1 => n21144, A2 => n24726, B1 => n20796, B2 => 
                           n24720, ZN => n22500);
   U21909 : AOI221_X1 port map( B1 => n24738, B2 => n19644, C1 => n24732, C2 =>
                           n19584, A => n22481, ZN => n22476);
   U21910 : OAI22_X1 port map( A1 => n21143, A2 => n24726, B1 => n20795, B2 => 
                           n24720, ZN => n22481);
   U21911 : AOI221_X1 port map( B1 => n24738, B2 => n19643, C1 => n24732, C2 =>
                           n19583, A => n22462, ZN => n22457);
   U21912 : OAI22_X1 port map( A1 => n21142, A2 => n24726, B1 => n20794, B2 => 
                           n24720, ZN => n22462);
   U21913 : AOI221_X1 port map( B1 => n24738, B2 => n19642, C1 => n24732, C2 =>
                           n19582, A => n22443, ZN => n22438);
   U21914 : OAI22_X1 port map( A1 => n21141, A2 => n24726, B1 => n20793, B2 => 
                           n24720, ZN => n22443);
   U21915 : AOI221_X1 port map( B1 => n24738, B2 => n19641, C1 => n24732, C2 =>
                           n19581, A => n22424, ZN => n22419);
   U21916 : OAI22_X1 port map( A1 => n21140, A2 => n24726, B1 => n20792, B2 => 
                           n24720, ZN => n22424);
   U21917 : AOI221_X1 port map( B1 => n24738, B2 => n19640, C1 => n24732, C2 =>
                           n19580, A => n22405, ZN => n22400);
   U21918 : OAI22_X1 port map( A1 => n21139, A2 => n24726, B1 => n20791, B2 => 
                           n24720, ZN => n22405);
   U21919 : AOI221_X1 port map( B1 => n24738, B2 => n19639, C1 => n24732, C2 =>
                           n19579, A => n22386, ZN => n22381);
   U21920 : OAI22_X1 port map( A1 => n21138, A2 => n24726, B1 => n20790, B2 => 
                           n24720, ZN => n22386);
   U21921 : AOI221_X1 port map( B1 => n24738, B2 => n19638, C1 => n24732, C2 =>
                           n19578, A => n22367, ZN => n22362);
   U21922 : OAI22_X1 port map( A1 => n21137, A2 => n24726, B1 => n20789, B2 => 
                           n24720, ZN => n22367);
   U21923 : AOI221_X1 port map( B1 => n24738, B2 => n19637, C1 => n24732, C2 =>
                           n19577, A => n22348, ZN => n22343);
   U21924 : OAI22_X1 port map( A1 => n21136, A2 => n24726, B1 => n20788, B2 => 
                           n24720, ZN => n22348);
   U21925 : AOI221_X1 port map( B1 => n24738, B2 => n19636, C1 => n24732, C2 =>
                           n19576, A => n22329, ZN => n22324);
   U21926 : OAI22_X1 port map( A1 => n21135, A2 => n24726, B1 => n20787, B2 => 
                           n24720, ZN => n22329);
   U21927 : AOI221_X1 port map( B1 => n24739, B2 => n19635, C1 => n24733, C2 =>
                           n19575, A => n22310, ZN => n22305);
   U21928 : OAI22_X1 port map( A1 => n21134, A2 => n24727, B1 => n20786, B2 => 
                           n24721, ZN => n22310);
   U21929 : AOI221_X1 port map( B1 => n24739, B2 => n19634, C1 => n24733, C2 =>
                           n19574, A => n22291, ZN => n22286);
   U21930 : OAI22_X1 port map( A1 => n21133, A2 => n24727, B1 => n20785, B2 => 
                           n24721, ZN => n22291);
   U21931 : AOI221_X1 port map( B1 => n24739, B2 => n19633, C1 => n24733, C2 =>
                           n19573, A => n22272, ZN => n22267);
   U21932 : OAI22_X1 port map( A1 => n21132, A2 => n24727, B1 => n20784, B2 => 
                           n24721, ZN => n22272);
   U21933 : AOI221_X1 port map( B1 => n24739, B2 => n19632, C1 => n24733, C2 =>
                           n19572, A => n22253, ZN => n22248);
   U21934 : OAI22_X1 port map( A1 => n21131, A2 => n24727, B1 => n20783, B2 => 
                           n24721, ZN => n22253);
   U21935 : AOI221_X1 port map( B1 => n24739, B2 => n19631, C1 => n24733, C2 =>
                           n19571, A => n22234, ZN => n22229);
   U21936 : OAI22_X1 port map( A1 => n21130, A2 => n24727, B1 => n20782, B2 => 
                           n24721, ZN => n22234);
   U21937 : AOI221_X1 port map( B1 => n24739, B2 => n19630, C1 => n24733, C2 =>
                           n19570, A => n22215, ZN => n22210);
   U21938 : OAI22_X1 port map( A1 => n21129, A2 => n24727, B1 => n20781, B2 => 
                           n24721, ZN => n22215);
   U21939 : AOI221_X1 port map( B1 => n24739, B2 => n19629, C1 => n24733, C2 =>
                           n19569, A => n22196, ZN => n22191);
   U21940 : OAI22_X1 port map( A1 => n21128, A2 => n24727, B1 => n20780, B2 => 
                           n24721, ZN => n22196);
   U21941 : AOI221_X1 port map( B1 => n24739, B2 => n19628, C1 => n24733, C2 =>
                           n19568, A => n22177, ZN => n22172);
   U21942 : OAI22_X1 port map( A1 => n21127, A2 => n24727, B1 => n20779, B2 => 
                           n24721, ZN => n22177);
   U21943 : AOI221_X1 port map( B1 => n24739, B2 => n19627, C1 => n24733, C2 =>
                           n19567, A => n22158, ZN => n22153);
   U21944 : OAI22_X1 port map( A1 => n21126, A2 => n24727, B1 => n20778, B2 => 
                           n24721, ZN => n22158);
   U21945 : AOI221_X1 port map( B1 => n24739, B2 => n19626, C1 => n24733, C2 =>
                           n19566, A => n22139, ZN => n22134);
   U21946 : OAI22_X1 port map( A1 => n21125, A2 => n24727, B1 => n20777, B2 => 
                           n24721, ZN => n22139);
   U21947 : AOI221_X1 port map( B1 => n24739, B2 => n19625, C1 => n24733, C2 =>
                           n19565, A => n22120, ZN => n22115);
   U21948 : OAI22_X1 port map( A1 => n21124, A2 => n24727, B1 => n20776, B2 => 
                           n24721, ZN => n22120);
   U21949 : AOI221_X1 port map( B1 => n24739, B2 => n19624, C1 => n24733, C2 =>
                           n19564, A => n22101, ZN => n22096);
   U21950 : OAI22_X1 port map( A1 => n21123, A2 => n24727, B1 => n20775, B2 => 
                           n24721, ZN => n22101);
   U21951 : AOI221_X1 port map( B1 => n24740, B2 => n19623, C1 => n24734, C2 =>
                           n19563, A => n22082, ZN => n22077);
   U21952 : OAI22_X1 port map( A1 => n21050, A2 => n24728, B1 => n20654, B2 => 
                           n24722, ZN => n22082);
   U21953 : AOI221_X1 port map( B1 => n24740, B2 => n19622, C1 => n24734, C2 =>
                           n19562, A => n22063, ZN => n22058);
   U21954 : OAI22_X1 port map( A1 => n21049, A2 => n24728, B1 => n20653, B2 => 
                           n24722, ZN => n22063);
   U21955 : AOI221_X1 port map( B1 => n24740, B2 => n19621, C1 => n24734, C2 =>
                           n19561, A => n22044, ZN => n22039);
   U21956 : OAI22_X1 port map( A1 => n21048, A2 => n24728, B1 => n20652, B2 => 
                           n24722, ZN => n22044);
   U21957 : AOI221_X1 port map( B1 => n24740, B2 => n19620, C1 => n24734, C2 =>
                           n19560, A => n22025, ZN => n22020);
   U21958 : OAI22_X1 port map( A1 => n21047, A2 => n24728, B1 => n20651, B2 => 
                           n24722, ZN => n22025);
   U21959 : AOI221_X1 port map( B1 => n24740, B2 => n19619, C1 => n24734, C2 =>
                           n19559, A => n22006, ZN => n22001);
   U21960 : OAI22_X1 port map( A1 => n21046, A2 => n24728, B1 => n20650, B2 => 
                           n24722, ZN => n22006);
   U21961 : AOI221_X1 port map( B1 => n24740, B2 => n19618, C1 => n24734, C2 =>
                           n19558, A => n21987, ZN => n21982);
   U21962 : OAI22_X1 port map( A1 => n21045, A2 => n24728, B1 => n20649, B2 => 
                           n24722, ZN => n21987);
   U21963 : AOI221_X1 port map( B1 => n24740, B2 => n19617, C1 => n24734, C2 =>
                           n19557, A => n21968, ZN => n21963);
   U21964 : OAI22_X1 port map( A1 => n21044, A2 => n24728, B1 => n20648, B2 => 
                           n24722, ZN => n21968);
   U21965 : AOI221_X1 port map( B1 => n24740, B2 => n19616, C1 => n24734, C2 =>
                           n19556, A => n21949, ZN => n21944);
   U21966 : OAI22_X1 port map( A1 => n21043, A2 => n24728, B1 => n20647, B2 => 
                           n24722, ZN => n21949);
   U21967 : AOI221_X1 port map( B1 => n24740, B2 => n19615, C1 => n24734, C2 =>
                           n19555, A => n21930, ZN => n21925);
   U21968 : OAI22_X1 port map( A1 => n21042, A2 => n24728, B1 => n20646, B2 => 
                           n24722, ZN => n21930);
   U21969 : AOI221_X1 port map( B1 => n24740, B2 => n19614, C1 => n24734, C2 =>
                           n19554, A => n21911, ZN => n21906);
   U21970 : OAI22_X1 port map( A1 => n21041, A2 => n24728, B1 => n20645, B2 => 
                           n24722, ZN => n21911);
   U21971 : AOI221_X1 port map( B1 => n24740, B2 => n19613, C1 => n24734, C2 =>
                           n19553, A => n21892, ZN => n21887);
   U21972 : OAI22_X1 port map( A1 => n21040, A2 => n24728, B1 => n20644, B2 => 
                           n24722, ZN => n21892);
   U21973 : AOI221_X1 port map( B1 => n24740, B2 => n19612, C1 => n24734, C2 =>
                           n19552, A => n21873, ZN => n21868);
   U21974 : OAI22_X1 port map( A1 => n21039, A2 => n24728, B1 => n20643, B2 => 
                           n24722, ZN => n21873);
   U21975 : AOI221_X1 port map( B1 => n24741, B2 => n19611, C1 => n24735, C2 =>
                           n19551, A => n21854, ZN => n21849);
   U21976 : OAI22_X1 port map( A1 => n21038, A2 => n24729, B1 => n20642, B2 => 
                           n24723, ZN => n21854);
   U21977 : AOI221_X1 port map( B1 => n24741, B2 => n19610, C1 => n24735, C2 =>
                           n19550, A => n21835, ZN => n21830);
   U21978 : OAI22_X1 port map( A1 => n21037, A2 => n24729, B1 => n20641, B2 => 
                           n24723, ZN => n21835);
   U21979 : AOI221_X1 port map( B1 => n24741, B2 => n19609, C1 => n24735, C2 =>
                           n19549, A => n21816, ZN => n21811);
   U21980 : OAI22_X1 port map( A1 => n21036, A2 => n24729, B1 => n20640, B2 => 
                           n24723, ZN => n21816);
   U21981 : AOI221_X1 port map( B1 => n24741, B2 => n19608, C1 => n24735, C2 =>
                           n19548, A => n21797, ZN => n21792);
   U21982 : OAI22_X1 port map( A1 => n21035, A2 => n24729, B1 => n20639, B2 => 
                           n24723, ZN => n21797);
   U21983 : AOI221_X1 port map( B1 => n24741, B2 => n19607, C1 => n24735, C2 =>
                           n19547, A => n21778, ZN => n21773);
   U21984 : OAI22_X1 port map( A1 => n21034, A2 => n24729, B1 => n20638, B2 => 
                           n24723, ZN => n21778);
   U21985 : AOI221_X1 port map( B1 => n24741, B2 => n19606, C1 => n24735, C2 =>
                           n19546, A => n21759, ZN => n21754);
   U21986 : OAI22_X1 port map( A1 => n21033, A2 => n24729, B1 => n20637, B2 => 
                           n24723, ZN => n21759);
   U21987 : AOI221_X1 port map( B1 => n24741, B2 => n19605, C1 => n24735, C2 =>
                           n19545, A => n21740, ZN => n21735);
   U21988 : OAI22_X1 port map( A1 => n21032, A2 => n24729, B1 => n20636, B2 => 
                           n24723, ZN => n21740);
   U21989 : AOI221_X1 port map( B1 => n24741, B2 => n19604, C1 => n24735, C2 =>
                           n19544, A => n21721, ZN => n21716);
   U21990 : OAI22_X1 port map( A1 => n21031, A2 => n24729, B1 => n20635, B2 => 
                           n24723, ZN => n21721);
   U21991 : AOI221_X1 port map( B1 => n24741, B2 => n19603, C1 => n24735, C2 =>
                           n19543, A => n21702, ZN => n21697);
   U21992 : OAI22_X1 port map( A1 => n21030, A2 => n24729, B1 => n20634, B2 => 
                           n24723, ZN => n21702);
   U21993 : AOI221_X1 port map( B1 => n24741, B2 => n19602, C1 => n24735, C2 =>
                           n19542, A => n21683, ZN => n21678);
   U21994 : OAI22_X1 port map( A1 => n21029, A2 => n24729, B1 => n20633, B2 => 
                           n24723, ZN => n21683);
   U21995 : AOI221_X1 port map( B1 => n24741, B2 => n19601, C1 => n24735, C2 =>
                           n19541, A => n21664, ZN => n21659);
   U21996 : OAI22_X1 port map( A1 => n21028, A2 => n24729, B1 => n20632, B2 => 
                           n24723, ZN => n21664);
   U21997 : AOI221_X1 port map( B1 => n24741, B2 => n19600, C1 => n24735, C2 =>
                           n19540, A => n21645, ZN => n21640);
   U21998 : OAI22_X1 port map( A1 => n21027, A2 => n24729, B1 => n20631, B2 => 
                           n24723, ZN => n21645);
   U21999 : AOI221_X1 port map( B1 => n24742, B2 => n19599, C1 => n24736, C2 =>
                           n19539, A => n21626, ZN => n21621);
   U22000 : OAI22_X1 port map( A1 => n21026, A2 => n24730, B1 => n20630, B2 => 
                           n24724, ZN => n21626);
   U22001 : AOI221_X1 port map( B1 => n24742, B2 => n19598, C1 => n24736, C2 =>
                           n19538, A => n21607, ZN => n21602);
   U22002 : OAI22_X1 port map( A1 => n21025, A2 => n24730, B1 => n20629, B2 => 
                           n24724, ZN => n21607);
   U22003 : AOI221_X1 port map( B1 => n24742, B2 => n19597, C1 => n24736, C2 =>
                           n19537, A => n21588, ZN => n21583);
   U22004 : OAI22_X1 port map( A1 => n21024, A2 => n24730, B1 => n20628, B2 => 
                           n24724, ZN => n21588);
   U22005 : AOI221_X1 port map( B1 => n24742, B2 => n19596, C1 => n24736, C2 =>
                           n19536, A => n21569, ZN => n21564);
   U22006 : OAI22_X1 port map( A1 => n21023, A2 => n24730, B1 => n20627, B2 => 
                           n24724, ZN => n21569);
   U22007 : AOI221_X1 port map( B1 => n24742, B2 => n19595, C1 => n24736, C2 =>
                           n19535, A => n21550, ZN => n21545);
   U22008 : OAI22_X1 port map( A1 => n21022, A2 => n24730, B1 => n20626, B2 => 
                           n24724, ZN => n21550);
   U22009 : AOI221_X1 port map( B1 => n24742, B2 => n19594, C1 => n24736, C2 =>
                           n19534, A => n21531, ZN => n21526);
   U22010 : OAI22_X1 port map( A1 => n21021, A2 => n24730, B1 => n20625, B2 => 
                           n24724, ZN => n21531);
   U22011 : AOI221_X1 port map( B1 => n24742, B2 => n19593, C1 => n24736, C2 =>
                           n19533, A => n21512, ZN => n21507);
   U22012 : OAI22_X1 port map( A1 => n21020, A2 => n24730, B1 => n20624, B2 => 
                           n24724, ZN => n21512);
   U22013 : AOI221_X1 port map( B1 => n24742, B2 => n19592, C1 => n24736, C2 =>
                           n19532, A => n21493, ZN => n21488);
   U22014 : OAI22_X1 port map( A1 => n21019, A2 => n24730, B1 => n20623, B2 => 
                           n24724, ZN => n21493);
   U22015 : AOI221_X1 port map( B1 => n24742, B2 => n19591, C1 => n24736, C2 =>
                           n19531, A => n21474, ZN => n21469);
   U22016 : OAI22_X1 port map( A1 => n21018, A2 => n24730, B1 => n20622, B2 => 
                           n24724, ZN => n21474);
   U22017 : AOI221_X1 port map( B1 => n24742, B2 => n19590, C1 => n24736, C2 =>
                           n19530, A => n21455, ZN => n21450);
   U22018 : OAI22_X1 port map( A1 => n21017, A2 => n24730, B1 => n20621, B2 => 
                           n24724, ZN => n21455);
   U22019 : AOI221_X1 port map( B1 => n24742, B2 => n19589, C1 => n24736, C2 =>
                           n19529, A => n21436, ZN => n21431);
   U22020 : OAI22_X1 port map( A1 => n21016, A2 => n24730, B1 => n20620, B2 => 
                           n24724, ZN => n21436);
   U22021 : AOI221_X1 port map( B1 => n24742, B2 => n19588, C1 => n24736, C2 =>
                           n19528, A => n21417, ZN => n21412);
   U22022 : OAI22_X1 port map( A1 => n21015, A2 => n24730, B1 => n20619, B2 => 
                           n24724, ZN => n21417);
   U22023 : AOI221_X1 port map( B1 => n24743, B2 => n20156, C1 => n24737, C2 =>
                           n19527, A => n21398, ZN => n21393);
   U22024 : OAI22_X1 port map( A1 => n20546, A2 => n24731, B1 => n20517, B2 => 
                           n24725, ZN => n21398);
   U22025 : AOI221_X1 port map( B1 => n24647, B2 => n17652, C1 => n24641, C2 =>
                           n24208, A => n21406, ZN => n21401);
   U22026 : OAI22_X1 port map( A1 => n20525, A2 => n24635, B1 => n20542, B2 => 
                           n24629, ZN => n21406);
   U22027 : AOI221_X1 port map( B1 => n24743, B2 => n20155, C1 => n24737, C2 =>
                           n19526, A => n21379, ZN => n21374);
   U22028 : OAI22_X1 port map( A1 => n20545, A2 => n24731, B1 => n20516, B2 => 
                           n24725, ZN => n21379);
   U22029 : AOI221_X1 port map( B1 => n24647, B2 => n17655, C1 => n24641, C2 =>
                           n24209, A => n21387, ZN => n21382);
   U22030 : OAI22_X1 port map( A1 => n20524, A2 => n24635, B1 => n20541, B2 => 
                           n24629, ZN => n21387);
   U22031 : AOI221_X1 port map( B1 => n24743, B2 => n20154, C1 => n24737, C2 =>
                           n19525, A => n21360, ZN => n21355);
   U22032 : OAI22_X1 port map( A1 => n20544, A2 => n24731, B1 => n20515, B2 => 
                           n24725, ZN => n21360);
   U22033 : AOI221_X1 port map( B1 => n24647, B2 => n17658, C1 => n24641, C2 =>
                           n24210, A => n21368, ZN => n21363);
   U22034 : OAI22_X1 port map( A1 => n20523, A2 => n24635, B1 => n20540, B2 => 
                           n24629, ZN => n21368);
   U22035 : AOI221_X1 port map( B1 => n24743, B2 => n20153, C1 => n24737, C2 =>
                           n19524, A => n21319, ZN => n21304);
   U22036 : OAI22_X1 port map( A1 => n20543, A2 => n24731, B1 => n20514, B2 => 
                           n24725, ZN => n21319);
   U22037 : AOI221_X1 port map( B1 => n24647, B2 => n17661, C1 => n24641, C2 =>
                           n24211, A => n21343, ZN => n21328);
   U22038 : OAI22_X1 port map( A1 => n20522, A2 => n24635, B1 => n20539, B2 => 
                           n24629, ZN => n21343);
   U22039 : AOI221_X1 port map( B1 => n24714, B2 => n20025, C1 => n24708, C2 =>
                           n20049, A => n22547, ZN => n22532);
   U22040 : OAI22_X1 port map( A1 => n20505, A2 => n24702, B1 => n20822, B2 => 
                           n24696, ZN => n22547);
   U22041 : AOI221_X1 port map( B1 => n24618, B2 => n17540, C1 => n24612, C2 =>
                           n7709, A => n22559, ZN => n22548);
   U22042 : OAI22_X1 port map( A1 => n20445, A2 => n24606, B1 => n20397, B2 => 
                           n24600, ZN => n22559);
   U22043 : AOI221_X1 port map( B1 => n24714, B2 => n20024, C1 => n24708, C2 =>
                           n20048, A => n22520, ZN => n22513);
   U22044 : OAI22_X1 port map( A1 => n20504, A2 => n24702, B1 => n20821, B2 => 
                           n24696, ZN => n22520);
   U22045 : AOI221_X1 port map( B1 => n24618, B2 => n17543, C1 => n24612, C2 =>
                           n7708, A => n22528, ZN => n22521);
   U22046 : OAI22_X1 port map( A1 => n20444, A2 => n24606, B1 => n20396, B2 => 
                           n24600, ZN => n22528);
   U22047 : AOI221_X1 port map( B1 => n24714, B2 => n20023, C1 => n24708, C2 =>
                           n20047, A => n22501, ZN => n22494);
   U22048 : OAI22_X1 port map( A1 => n20503, A2 => n24702, B1 => n20820, B2 => 
                           n24696, ZN => n22501);
   U22049 : AOI221_X1 port map( B1 => n24618, B2 => n17546, C1 => n24612, C2 =>
                           n7707, A => n22509, ZN => n22502);
   U22050 : OAI22_X1 port map( A1 => n20443, A2 => n24606, B1 => n20395, B2 => 
                           n24600, ZN => n22509);
   U22051 : AOI221_X1 port map( B1 => n24714, B2 => n20022, C1 => n24708, C2 =>
                           n20046, A => n22482, ZN => n22475);
   U22052 : OAI22_X1 port map( A1 => n20502, A2 => n24702, B1 => n20819, B2 => 
                           n24696, ZN => n22482);
   U22053 : AOI221_X1 port map( B1 => n24618, B2 => n17549, C1 => n24612, C2 =>
                           n7706, A => n22490, ZN => n22483);
   U22054 : OAI22_X1 port map( A1 => n20442, A2 => n24606, B1 => n20394, B2 => 
                           n24600, ZN => n22490);
   U22055 : AOI221_X1 port map( B1 => n24714, B2 => n20021, C1 => n24708, C2 =>
                           n20045, A => n22463, ZN => n22456);
   U22056 : OAI22_X1 port map( A1 => n20501, A2 => n24702, B1 => n20818, B2 => 
                           n24696, ZN => n22463);
   U22057 : AOI221_X1 port map( B1 => n24618, B2 => n17552, C1 => n24612, C2 =>
                           n7705, A => n22471, ZN => n22464);
   U22058 : OAI22_X1 port map( A1 => n20441, A2 => n24606, B1 => n20393, B2 => 
                           n24600, ZN => n22471);
   U22059 : AOI221_X1 port map( B1 => n24714, B2 => n20020, C1 => n24708, C2 =>
                           n20044, A => n22444, ZN => n22437);
   U22060 : OAI22_X1 port map( A1 => n20500, A2 => n24702, B1 => n20817, B2 => 
                           n24696, ZN => n22444);
   U22061 : AOI221_X1 port map( B1 => n24618, B2 => n17555, C1 => n24612, C2 =>
                           n7704, A => n22452, ZN => n22445);
   U22062 : OAI22_X1 port map( A1 => n20440, A2 => n24606, B1 => n20392, B2 => 
                           n24600, ZN => n22452);
   U22063 : AOI221_X1 port map( B1 => n24714, B2 => n20019, C1 => n24708, C2 =>
                           n20043, A => n22425, ZN => n22418);
   U22064 : OAI22_X1 port map( A1 => n20499, A2 => n24702, B1 => n20816, B2 => 
                           n24696, ZN => n22425);
   U22065 : AOI221_X1 port map( B1 => n24618, B2 => n17558, C1 => n24612, C2 =>
                           n7703, A => n22433, ZN => n22426);
   U22066 : OAI22_X1 port map( A1 => n20439, A2 => n24606, B1 => n20391, B2 => 
                           n24600, ZN => n22433);
   U22067 : AOI221_X1 port map( B1 => n24714, B2 => n20018, C1 => n24708, C2 =>
                           n20042, A => n22406, ZN => n22399);
   U22068 : OAI22_X1 port map( A1 => n20498, A2 => n24702, B1 => n20815, B2 => 
                           n24696, ZN => n22406);
   U22069 : AOI221_X1 port map( B1 => n24618, B2 => n17561, C1 => n24612, C2 =>
                           n7702, A => n22414, ZN => n22407);
   U22070 : OAI22_X1 port map( A1 => n20438, A2 => n24606, B1 => n20390, B2 => 
                           n24600, ZN => n22414);
   U22071 : AOI221_X1 port map( B1 => n24714, B2 => n20017, C1 => n24708, C2 =>
                           n20041, A => n22387, ZN => n22380);
   U22072 : OAI22_X1 port map( A1 => n20497, A2 => n24702, B1 => n20814, B2 => 
                           n24696, ZN => n22387);
   U22073 : AOI221_X1 port map( B1 => n24618, B2 => n17564, C1 => n24612, C2 =>
                           n7701, A => n22395, ZN => n22388);
   U22074 : OAI22_X1 port map( A1 => n20437, A2 => n24606, B1 => n20389, B2 => 
                           n24600, ZN => n22395);
   U22075 : AOI221_X1 port map( B1 => n24714, B2 => n20016, C1 => n24708, C2 =>
                           n20040, A => n22368, ZN => n22361);
   U22076 : OAI22_X1 port map( A1 => n20496, A2 => n24702, B1 => n20813, B2 => 
                           n24696, ZN => n22368);
   U22077 : AOI221_X1 port map( B1 => n24618, B2 => n17567, C1 => n24612, C2 =>
                           n7700, A => n22376, ZN => n22369);
   U22078 : OAI22_X1 port map( A1 => n20436, A2 => n24606, B1 => n20388, B2 => 
                           n24600, ZN => n22376);
   U22079 : AOI221_X1 port map( B1 => n24714, B2 => n20015, C1 => n24708, C2 =>
                           n20039, A => n22349, ZN => n22342);
   U22080 : OAI22_X1 port map( A1 => n20495, A2 => n24702, B1 => n20812, B2 => 
                           n24696, ZN => n22349);
   U22081 : AOI221_X1 port map( B1 => n24618, B2 => n17570, C1 => n24612, C2 =>
                           n7699, A => n22357, ZN => n22350);
   U22082 : OAI22_X1 port map( A1 => n20435, A2 => n24606, B1 => n20387, B2 => 
                           n24600, ZN => n22357);
   U22083 : AOI221_X1 port map( B1 => n24714, B2 => n20014, C1 => n24708, C2 =>
                           n20038, A => n22330, ZN => n22323);
   U22084 : OAI22_X1 port map( A1 => n20494, A2 => n24702, B1 => n20811, B2 => 
                           n24696, ZN => n22330);
   U22085 : AOI221_X1 port map( B1 => n24618, B2 => n17573, C1 => n24612, C2 =>
                           n7698, A => n22338, ZN => n22331);
   U22086 : OAI22_X1 port map( A1 => n20434, A2 => n24606, B1 => n20386, B2 => 
                           n24600, ZN => n22338);
   U22087 : AOI221_X1 port map( B1 => n24715, B2 => n20013, C1 => n24709, C2 =>
                           n20037, A => n22311, ZN => n22304);
   U22088 : OAI22_X1 port map( A1 => n20493, A2 => n24703, B1 => n20810, B2 => 
                           n24697, ZN => n22311);
   U22089 : AOI221_X1 port map( B1 => n24619, B2 => n17576, C1 => n24613, C2 =>
                           n7697, A => n22319, ZN => n22312);
   U22090 : OAI22_X1 port map( A1 => n20433, A2 => n24607, B1 => n20385, B2 => 
                           n24601, ZN => n22319);
   U22091 : AOI221_X1 port map( B1 => n24715, B2 => n20012, C1 => n24709, C2 =>
                           n20036, A => n22292, ZN => n22285);
   U22092 : OAI22_X1 port map( A1 => n20492, A2 => n24703, B1 => n20809, B2 => 
                           n24697, ZN => n22292);
   U22093 : AOI221_X1 port map( B1 => n24619, B2 => n17579, C1 => n24613, C2 =>
                           n7696, A => n22300, ZN => n22293);
   U22094 : OAI22_X1 port map( A1 => n20432, A2 => n24607, B1 => n20384, B2 => 
                           n24601, ZN => n22300);
   U22095 : AOI221_X1 port map( B1 => n24715, B2 => n20011, C1 => n24709, C2 =>
                           n20035, A => n22273, ZN => n22266);
   U22096 : OAI22_X1 port map( A1 => n20491, A2 => n24703, B1 => n20808, B2 => 
                           n24697, ZN => n22273);
   U22097 : AOI221_X1 port map( B1 => n24619, B2 => n17582, C1 => n24613, C2 =>
                           n7695, A => n22281, ZN => n22274);
   U22098 : OAI22_X1 port map( A1 => n20431, A2 => n24607, B1 => n20383, B2 => 
                           n24601, ZN => n22281);
   U22099 : AOI221_X1 port map( B1 => n24715, B2 => n20010, C1 => n24709, C2 =>
                           n20034, A => n22254, ZN => n22247);
   U22100 : OAI22_X1 port map( A1 => n20490, A2 => n24703, B1 => n20807, B2 => 
                           n24697, ZN => n22254);
   U22101 : AOI221_X1 port map( B1 => n24619, B2 => n17585, C1 => n24613, C2 =>
                           n7694, A => n22262, ZN => n22255);
   U22102 : OAI22_X1 port map( A1 => n20430, A2 => n24607, B1 => n20382, B2 => 
                           n24601, ZN => n22262);
   U22103 : AOI221_X1 port map( B1 => n24715, B2 => n20009, C1 => n24709, C2 =>
                           n20033, A => n22235, ZN => n22228);
   U22104 : OAI22_X1 port map( A1 => n20489, A2 => n24703, B1 => n20806, B2 => 
                           n24697, ZN => n22235);
   U22105 : AOI221_X1 port map( B1 => n24619, B2 => n17588, C1 => n24613, C2 =>
                           n7693, A => n22243, ZN => n22236);
   U22106 : OAI22_X1 port map( A1 => n20429, A2 => n24607, B1 => n20381, B2 => 
                           n24601, ZN => n22243);
   U22107 : AOI221_X1 port map( B1 => n24715, B2 => n20008, C1 => n24709, C2 =>
                           n20032, A => n22216, ZN => n22209);
   U22108 : OAI22_X1 port map( A1 => n20488, A2 => n24703, B1 => n20805, B2 => 
                           n24697, ZN => n22216);
   U22109 : AOI221_X1 port map( B1 => n24619, B2 => n17591, C1 => n24613, C2 =>
                           n7692, A => n22224, ZN => n22217);
   U22110 : OAI22_X1 port map( A1 => n20428, A2 => n24607, B1 => n20380, B2 => 
                           n24601, ZN => n22224);
   U22111 : AOI221_X1 port map( B1 => n24715, B2 => n20007, C1 => n24709, C2 =>
                           n20031, A => n22197, ZN => n22190);
   U22112 : OAI22_X1 port map( A1 => n20487, A2 => n24703, B1 => n20804, B2 => 
                           n24697, ZN => n22197);
   U22113 : AOI221_X1 port map( B1 => n24619, B2 => n17594, C1 => n24613, C2 =>
                           n7691, A => n22205, ZN => n22198);
   U22114 : OAI22_X1 port map( A1 => n20427, A2 => n24607, B1 => n20379, B2 => 
                           n24601, ZN => n22205);
   U22115 : AOI221_X1 port map( B1 => n24715, B2 => n20006, C1 => n24709, C2 =>
                           n20030, A => n22178, ZN => n22171);
   U22116 : OAI22_X1 port map( A1 => n20486, A2 => n24703, B1 => n20803, B2 => 
                           n24697, ZN => n22178);
   U22117 : AOI221_X1 port map( B1 => n24619, B2 => n17597, C1 => n24613, C2 =>
                           n7690, A => n22186, ZN => n22179);
   U22118 : OAI22_X1 port map( A1 => n20426, A2 => n24607, B1 => n20378, B2 => 
                           n24601, ZN => n22186);
   U22119 : AOI221_X1 port map( B1 => n24715, B2 => n20005, C1 => n24709, C2 =>
                           n20029, A => n22159, ZN => n22152);
   U22120 : OAI22_X1 port map( A1 => n20485, A2 => n24703, B1 => n20802, B2 => 
                           n24697, ZN => n22159);
   U22121 : AOI221_X1 port map( B1 => n24619, B2 => n17600, C1 => n24613, C2 =>
                           n7689, A => n22167, ZN => n22160);
   U22122 : OAI22_X1 port map( A1 => n20425, A2 => n24607, B1 => n20377, B2 => 
                           n24601, ZN => n22167);
   U22123 : AOI221_X1 port map( B1 => n24715, B2 => n20004, C1 => n24709, C2 =>
                           n20028, A => n22140, ZN => n22133);
   U22124 : OAI22_X1 port map( A1 => n20484, A2 => n24703, B1 => n20801, B2 => 
                           n24697, ZN => n22140);
   U22125 : AOI221_X1 port map( B1 => n24619, B2 => n17603, C1 => n24613, C2 =>
                           n7688, A => n22148, ZN => n22141);
   U22126 : OAI22_X1 port map( A1 => n20424, A2 => n24607, B1 => n20376, B2 => 
                           n24601, ZN => n22148);
   U22127 : AOI221_X1 port map( B1 => n24715, B2 => n20003, C1 => n24709, C2 =>
                           n20027, A => n22121, ZN => n22114);
   U22128 : OAI22_X1 port map( A1 => n20483, A2 => n24703, B1 => n20800, B2 => 
                           n24697, ZN => n22121);
   U22129 : AOI221_X1 port map( B1 => n24619, B2 => n17606, C1 => n24613, C2 =>
                           n7687, A => n22129, ZN => n22122);
   U22130 : OAI22_X1 port map( A1 => n20423, A2 => n24607, B1 => n20375, B2 => 
                           n24601, ZN => n22129);
   U22131 : AOI221_X1 port map( B1 => n24715, B2 => n20002, C1 => n24709, C2 =>
                           n20026, A => n22102, ZN => n22095);
   U22132 : OAI22_X1 port map( A1 => n20482, A2 => n24703, B1 => n20799, B2 => 
                           n24697, ZN => n22102);
   U22133 : AOI221_X1 port map( B1 => n24619, B2 => n17609, C1 => n24613, C2 =>
                           n7686, A => n22110, ZN => n22103);
   U22134 : OAI22_X1 port map( A1 => n20422, A2 => n24607, B1 => n20374, B2 => 
                           n24601, ZN => n22110);
   U22135 : AOI221_X1 port map( B1 => n24716, B2 => n19857, C1 => n24710, C2 =>
                           n19893, A => n22083, ZN => n22076);
   U22136 : OAI22_X1 port map( A1 => n20481, A2 => n24704, B1 => n20690, B2 => 
                           n24698, ZN => n22083);
   U22137 : AOI221_X1 port map( B1 => n24620, B2 => n17612, C1 => n24614, C2 =>
                           n7685, A => n22091, ZN => n22084);
   U22138 : OAI22_X1 port map( A1 => n20373, A2 => n24608, B1 => n20301, B2 => 
                           n24602, ZN => n22091);
   U22139 : AOI221_X1 port map( B1 => n24716, B2 => n19856, C1 => n24710, C2 =>
                           n19892, A => n22064, ZN => n22057);
   U22140 : OAI22_X1 port map( A1 => n20480, A2 => n24704, B1 => n20689, B2 => 
                           n24698, ZN => n22064);
   U22141 : AOI221_X1 port map( B1 => n24620, B2 => n17615, C1 => n24614, C2 =>
                           n7684, A => n22072, ZN => n22065);
   U22142 : OAI22_X1 port map( A1 => n20372, A2 => n24608, B1 => n20300, B2 => 
                           n24602, ZN => n22072);
   U22143 : AOI221_X1 port map( B1 => n24716, B2 => n19855, C1 => n24710, C2 =>
                           n19891, A => n22045, ZN => n22038);
   U22144 : OAI22_X1 port map( A1 => n20479, A2 => n24704, B1 => n20688, B2 => 
                           n24698, ZN => n22045);
   U22145 : AOI221_X1 port map( B1 => n24620, B2 => n17618, C1 => n24614, C2 =>
                           n7683, A => n22053, ZN => n22046);
   U22146 : OAI22_X1 port map( A1 => n20371, A2 => n24608, B1 => n20299, B2 => 
                           n24602, ZN => n22053);
   U22147 : AOI221_X1 port map( B1 => n24716, B2 => n19854, C1 => n24710, C2 =>
                           n19890, A => n22026, ZN => n22019);
   U22148 : OAI22_X1 port map( A1 => n20478, A2 => n24704, B1 => n20687, B2 => 
                           n24698, ZN => n22026);
   U22149 : AOI221_X1 port map( B1 => n24620, B2 => n17621, C1 => n24614, C2 =>
                           n7682, A => n22034, ZN => n22027);
   U22150 : OAI22_X1 port map( A1 => n20370, A2 => n24608, B1 => n20298, B2 => 
                           n24602, ZN => n22034);
   U22151 : AOI221_X1 port map( B1 => n24716, B2 => n19853, C1 => n24710, C2 =>
                           n19889, A => n22007, ZN => n22000);
   U22152 : OAI22_X1 port map( A1 => n20477, A2 => n24704, B1 => n20686, B2 => 
                           n24698, ZN => n22007);
   U22153 : AOI221_X1 port map( B1 => n24620, B2 => n17624, C1 => n24614, C2 =>
                           n7681, A => n22015, ZN => n22008);
   U22154 : OAI22_X1 port map( A1 => n20369, A2 => n24608, B1 => n20297, B2 => 
                           n24602, ZN => n22015);
   U22155 : AOI221_X1 port map( B1 => n24716, B2 => n19852, C1 => n24710, C2 =>
                           n19888, A => n21988, ZN => n21981);
   U22156 : OAI22_X1 port map( A1 => n20476, A2 => n24704, B1 => n20685, B2 => 
                           n24698, ZN => n21988);
   U22157 : AOI221_X1 port map( B1 => n24620, B2 => n17471, C1 => n24614, C2 =>
                           n20144, A => n21996, ZN => n21989);
   U22158 : OAI22_X1 port map( A1 => n20368, A2 => n24608, B1 => n20296, B2 => 
                           n24602, ZN => n21996);
   U22159 : AOI221_X1 port map( B1 => n24716, B2 => n19851, C1 => n24710, C2 =>
                           n19887, A => n21969, ZN => n21962);
   U22160 : OAI22_X1 port map( A1 => n20475, A2 => n24704, B1 => n20684, B2 => 
                           n24698, ZN => n21969);
   U22161 : AOI221_X1 port map( B1 => n24620, B2 => n17474, C1 => n24614, C2 =>
                           n20143, A => n21977, ZN => n21970);
   U22162 : OAI22_X1 port map( A1 => n20367, A2 => n24608, B1 => n20295, B2 => 
                           n24602, ZN => n21977);
   U22163 : AOI221_X1 port map( B1 => n24716, B2 => n19850, C1 => n24710, C2 =>
                           n19886, A => n21950, ZN => n21943);
   U22164 : OAI22_X1 port map( A1 => n20474, A2 => n24704, B1 => n20683, B2 => 
                           n24698, ZN => n21950);
   U22165 : AOI221_X1 port map( B1 => n24620, B2 => n17477, C1 => n24614, C2 =>
                           n20142, A => n21958, ZN => n21951);
   U22166 : OAI22_X1 port map( A1 => n20366, A2 => n24608, B1 => n20294, B2 => 
                           n24602, ZN => n21958);
   U22167 : AOI221_X1 port map( B1 => n24716, B2 => n19849, C1 => n24710, C2 =>
                           n19885, A => n21931, ZN => n21924);
   U22168 : OAI22_X1 port map( A1 => n20473, A2 => n24704, B1 => n20682, B2 => 
                           n24698, ZN => n21931);
   U22169 : AOI221_X1 port map( B1 => n24620, B2 => n17480, C1 => n24614, C2 =>
                           n20141, A => n21939, ZN => n21932);
   U22170 : OAI22_X1 port map( A1 => n20365, A2 => n24608, B1 => n20293, B2 => 
                           n24602, ZN => n21939);
   U22171 : AOI221_X1 port map( B1 => n24716, B2 => n19848, C1 => n24710, C2 =>
                           n19884, A => n21912, ZN => n21905);
   U22172 : OAI22_X1 port map( A1 => n20472, A2 => n24704, B1 => n20681, B2 => 
                           n24698, ZN => n21912);
   U22173 : AOI221_X1 port map( B1 => n24620, B2 => n17483, C1 => n24614, C2 =>
                           n20140, A => n21920, ZN => n21913);
   U22174 : OAI22_X1 port map( A1 => n20364, A2 => n24608, B1 => n20292, B2 => 
                           n24602, ZN => n21920);
   U22175 : AOI221_X1 port map( B1 => n24716, B2 => n19847, C1 => n24710, C2 =>
                           n19883, A => n21893, ZN => n21886);
   U22176 : OAI22_X1 port map( A1 => n20471, A2 => n24704, B1 => n20680, B2 => 
                           n24698, ZN => n21893);
   U22177 : AOI221_X1 port map( B1 => n24620, B2 => n17486, C1 => n24614, C2 =>
                           n20139, A => n21901, ZN => n21894);
   U22178 : OAI22_X1 port map( A1 => n20363, A2 => n24608, B1 => n20291, B2 => 
                           n24602, ZN => n21901);
   U22179 : AOI221_X1 port map( B1 => n24716, B2 => n19846, C1 => n24710, C2 =>
                           n19882, A => n21874, ZN => n21867);
   U22180 : OAI22_X1 port map( A1 => n20470, A2 => n24704, B1 => n20679, B2 => 
                           n24698, ZN => n21874);
   U22181 : AOI221_X1 port map( B1 => n24620, B2 => n17489, C1 => n24614, C2 =>
                           n20133, A => n21882, ZN => n21875);
   U22182 : OAI22_X1 port map( A1 => n20362, A2 => n24608, B1 => n20290, B2 => 
                           n24602, ZN => n21882);
   U22183 : AOI221_X1 port map( B1 => n24717, B2 => n19845, C1 => n24711, C2 =>
                           n19881, A => n21855, ZN => n21848);
   U22184 : OAI22_X1 port map( A1 => n20469, A2 => n24705, B1 => n20678, B2 => 
                           n24699, ZN => n21855);
   U22185 : AOI221_X1 port map( B1 => n24621, B2 => n17492, C1 => n24615, C2 =>
                           n20138, A => n21863, ZN => n21856);
   U22186 : OAI22_X1 port map( A1 => n20361, A2 => n24609, B1 => n20289, B2 => 
                           n24603, ZN => n21863);
   U22187 : AOI221_X1 port map( B1 => n24717, B2 => n19844, C1 => n24711, C2 =>
                           n19880, A => n21836, ZN => n21829);
   U22188 : OAI22_X1 port map( A1 => n20468, A2 => n24705, B1 => n20677, B2 => 
                           n24699, ZN => n21836);
   U22189 : AOI221_X1 port map( B1 => n24621, B2 => n17495, C1 => n24615, C2 =>
                           n20137, A => n21844, ZN => n21837);
   U22190 : OAI22_X1 port map( A1 => n20360, A2 => n24609, B1 => n20288, B2 => 
                           n24603, ZN => n21844);
   U22191 : AOI221_X1 port map( B1 => n24717, B2 => n19843, C1 => n24711, C2 =>
                           n19879, A => n21817, ZN => n21810);
   U22192 : OAI22_X1 port map( A1 => n20467, A2 => n24705, B1 => n20676, B2 => 
                           n24699, ZN => n21817);
   U22193 : AOI221_X1 port map( B1 => n24621, B2 => n17498, C1 => n24615, C2 =>
                           n20136, A => n21825, ZN => n21818);
   U22194 : OAI22_X1 port map( A1 => n20359, A2 => n24609, B1 => n20287, B2 => 
                           n24603, ZN => n21825);
   U22195 : AOI221_X1 port map( B1 => n24717, B2 => n19842, C1 => n24711, C2 =>
                           n19878, A => n21798, ZN => n21791);
   U22196 : OAI22_X1 port map( A1 => n20466, A2 => n24705, B1 => n20675, B2 => 
                           n24699, ZN => n21798);
   U22197 : AOI221_X1 port map( B1 => n24621, B2 => n17501, C1 => n24615, C2 =>
                           n20132, A => n21806, ZN => n21799);
   U22198 : OAI22_X1 port map( A1 => n20358, A2 => n24609, B1 => n20286, B2 => 
                           n24603, ZN => n21806);
   U22199 : AOI221_X1 port map( B1 => n24717, B2 => n19841, C1 => n24711, C2 =>
                           n19877, A => n21779, ZN => n21772);
   U22200 : OAI22_X1 port map( A1 => n20465, A2 => n24705, B1 => n20674, B2 => 
                           n24699, ZN => n21779);
   U22201 : AOI221_X1 port map( B1 => n24621, B2 => n17504, C1 => n24615, C2 =>
                           n20135, A => n21787, ZN => n21780);
   U22202 : OAI22_X1 port map( A1 => n20357, A2 => n24609, B1 => n20285, B2 => 
                           n24603, ZN => n21787);
   U22203 : AOI221_X1 port map( B1 => n24717, B2 => n19840, C1 => n24711, C2 =>
                           n19876, A => n21760, ZN => n21753);
   U22204 : OAI22_X1 port map( A1 => n20464, A2 => n24705, B1 => n20673, B2 => 
                           n24699, ZN => n21760);
   U22205 : AOI221_X1 port map( B1 => n24621, B2 => n17507, C1 => n24615, C2 =>
                           n20131, A => n21768, ZN => n21761);
   U22206 : OAI22_X1 port map( A1 => n20356, A2 => n24609, B1 => n20284, B2 => 
                           n24603, ZN => n21768);
   U22207 : AOI221_X1 port map( B1 => n24717, B2 => n19839, C1 => n24711, C2 =>
                           n19875, A => n21741, ZN => n21734);
   U22208 : OAI22_X1 port map( A1 => n20463, A2 => n24705, B1 => n20672, B2 => 
                           n24699, ZN => n21741);
   U22209 : AOI221_X1 port map( B1 => n24621, B2 => n17510, C1 => n24615, C2 =>
                           n20134, A => n21749, ZN => n21742);
   U22210 : OAI22_X1 port map( A1 => n20355, A2 => n24609, B1 => n20283, B2 => 
                           n24603, ZN => n21749);
   U22211 : AOI221_X1 port map( B1 => n24717, B2 => n19838, C1 => n24711, C2 =>
                           n19874, A => n21722, ZN => n21715);
   U22212 : OAI22_X1 port map( A1 => n20462, A2 => n24705, B1 => n20671, B2 => 
                           n24699, ZN => n21722);
   U22213 : AOI221_X1 port map( B1 => n24621, B2 => n17513, C1 => n24615, C2 =>
                           n20130, A => n21730, ZN => n21723);
   U22214 : OAI22_X1 port map( A1 => n20354, A2 => n24609, B1 => n20282, B2 => 
                           n24603, ZN => n21730);
   U22215 : AOI221_X1 port map( B1 => n24717, B2 => n19837, C1 => n24711, C2 =>
                           n19873, A => n21703, ZN => n21696);
   U22216 : OAI22_X1 port map( A1 => n20461, A2 => n24705, B1 => n20670, B2 => 
                           n24699, ZN => n21703);
   U22217 : AOI221_X1 port map( B1 => n24621, B2 => n17516, C1 => n24615, C2 =>
                           n20129, A => n21711, ZN => n21704);
   U22218 : OAI22_X1 port map( A1 => n20353, A2 => n24609, B1 => n20281, B2 => 
                           n24603, ZN => n21711);
   U22219 : AOI221_X1 port map( B1 => n24717, B2 => n19836, C1 => n24711, C2 =>
                           n19872, A => n21684, ZN => n21677);
   U22220 : OAI22_X1 port map( A1 => n20460, A2 => n24705, B1 => n20669, B2 => 
                           n24699, ZN => n21684);
   U22221 : AOI221_X1 port map( B1 => n24621, B2 => n17519, C1 => n24615, C2 =>
                           n20128, A => n21692, ZN => n21685);
   U22222 : OAI22_X1 port map( A1 => n20352, A2 => n24609, B1 => n20280, B2 => 
                           n24603, ZN => n21692);
   U22223 : AOI221_X1 port map( B1 => n24717, B2 => n19835, C1 => n24711, C2 =>
                           n19871, A => n21665, ZN => n21658);
   U22224 : OAI22_X1 port map( A1 => n20459, A2 => n24705, B1 => n20668, B2 => 
                           n24699, ZN => n21665);
   U22225 : AOI221_X1 port map( B1 => n24621, B2 => n17522, C1 => n24615, C2 =>
                           n20127, A => n21673, ZN => n21666);
   U22226 : OAI22_X1 port map( A1 => n20351, A2 => n24609, B1 => n20279, B2 => 
                           n24603, ZN => n21673);
   U22227 : AOI221_X1 port map( B1 => n24717, B2 => n19834, C1 => n24711, C2 =>
                           n19870, A => n21646, ZN => n21639);
   U22228 : OAI22_X1 port map( A1 => n20458, A2 => n24705, B1 => n20667, B2 => 
                           n24699, ZN => n21646);
   U22229 : AOI221_X1 port map( B1 => n24621, B2 => n17525, C1 => n24615, C2 =>
                           n20126, A => n21654, ZN => n21647);
   U22230 : OAI22_X1 port map( A1 => n20350, A2 => n24609, B1 => n20278, B2 => 
                           n24603, ZN => n21654);
   U22231 : AOI221_X1 port map( B1 => n24718, B2 => n19833, C1 => n24712, C2 =>
                           n19869, A => n21627, ZN => n21620);
   U22232 : OAI22_X1 port map( A1 => n20457, A2 => n24706, B1 => n20666, B2 => 
                           n24700, ZN => n21627);
   U22233 : AOI221_X1 port map( B1 => n24622, B2 => n17528, C1 => n24616, C2 =>
                           n20125, A => n21635, ZN => n21628);
   U22234 : OAI22_X1 port map( A1 => n20349, A2 => n24610, B1 => n20277, B2 => 
                           n24604, ZN => n21635);
   U22235 : AOI221_X1 port map( B1 => n24718, B2 => n19832, C1 => n24712, C2 =>
                           n19868, A => n21608, ZN => n21601);
   U22236 : OAI22_X1 port map( A1 => n20456, A2 => n24706, B1 => n20665, B2 => 
                           n24700, ZN => n21608);
   U22237 : AOI221_X1 port map( B1 => n24622, B2 => n17531, C1 => n24616, C2 =>
                           n20124, A => n21616, ZN => n21609);
   U22238 : OAI22_X1 port map( A1 => n20348, A2 => n24610, B1 => n20276, B2 => 
                           n24604, ZN => n21616);
   U22239 : AOI221_X1 port map( B1 => n24718, B2 => n19831, C1 => n24712, C2 =>
                           n19867, A => n21589, ZN => n21582);
   U22240 : OAI22_X1 port map( A1 => n20455, A2 => n24706, B1 => n20664, B2 => 
                           n24700, ZN => n21589);
   U22241 : AOI221_X1 port map( B1 => n24622, B2 => n17534, C1 => n24616, C2 =>
                           n20123, A => n21597, ZN => n21590);
   U22242 : OAI22_X1 port map( A1 => n20347, A2 => n24610, B1 => n20275, B2 => 
                           n24604, ZN => n21597);
   U22243 : AOI221_X1 port map( B1 => n24718, B2 => n19830, C1 => n24712, C2 =>
                           n19866, A => n21570, ZN => n21563);
   U22244 : OAI22_X1 port map( A1 => n20454, A2 => n24706, B1 => n20663, B2 => 
                           n24700, ZN => n21570);
   U22245 : AOI221_X1 port map( B1 => n24622, B2 => n17537, C1 => n24616, C2 =>
                           n20122, A => n21578, ZN => n21571);
   U22246 : OAI22_X1 port map( A1 => n20346, A2 => n24610, B1 => n20274, B2 => 
                           n24604, ZN => n21578);
   U22247 : AOI221_X1 port map( B1 => n24718, B2 => n19829, C1 => n24712, C2 =>
                           n19865, A => n21551, ZN => n21544);
   U22248 : OAI22_X1 port map( A1 => n20453, A2 => n24706, B1 => n20662, B2 => 
                           n24700, ZN => n21551);
   U22249 : AOI221_X1 port map( B1 => n24622, B2 => n17627, C1 => n24616, C2 =>
                           n7657, A => n21559, ZN => n21552);
   U22250 : OAI22_X1 port map( A1 => n20345, A2 => n24610, B1 => n20273, B2 => 
                           n24604, ZN => n21559);
   U22251 : AOI221_X1 port map( B1 => n24718, B2 => n19828, C1 => n24712, C2 =>
                           n19864, A => n21532, ZN => n21525);
   U22252 : OAI22_X1 port map( A1 => n20452, A2 => n24706, B1 => n20661, B2 => 
                           n24700, ZN => n21532);
   U22253 : AOI221_X1 port map( B1 => n24622, B2 => n17630, C1 => n24616, C2 =>
                           n7656, A => n21540, ZN => n21533);
   U22254 : OAI22_X1 port map( A1 => n20344, A2 => n24610, B1 => n20272, B2 => 
                           n24604, ZN => n21540);
   U22255 : AOI221_X1 port map( B1 => n24718, B2 => n19827, C1 => n24712, C2 =>
                           n19863, A => n21513, ZN => n21506);
   U22256 : OAI22_X1 port map( A1 => n20451, A2 => n24706, B1 => n20660, B2 => 
                           n24700, ZN => n21513);
   U22257 : AOI221_X1 port map( B1 => n24622, B2 => n17633, C1 => n24616, C2 =>
                           n7655, A => n21521, ZN => n21514);
   U22258 : OAI22_X1 port map( A1 => n20343, A2 => n24610, B1 => n20271, B2 => 
                           n24604, ZN => n21521);
   U22259 : AOI221_X1 port map( B1 => n24718, B2 => n19826, C1 => n24712, C2 =>
                           n19862, A => n21494, ZN => n21487);
   U22260 : OAI22_X1 port map( A1 => n20450, A2 => n24706, B1 => n20659, B2 => 
                           n24700, ZN => n21494);
   U22261 : AOI221_X1 port map( B1 => n24622, B2 => n17636, C1 => n24616, C2 =>
                           n7654, A => n21502, ZN => n21495);
   U22262 : OAI22_X1 port map( A1 => n20342, A2 => n24610, B1 => n20270, B2 => 
                           n24604, ZN => n21502);
   U22263 : AOI221_X1 port map( B1 => n24718, B2 => n19825, C1 => n24712, C2 =>
                           n19861, A => n21475, ZN => n21468);
   U22264 : OAI22_X1 port map( A1 => n20449, A2 => n24706, B1 => n20658, B2 => 
                           n24700, ZN => n21475);
   U22265 : AOI221_X1 port map( B1 => n24622, B2 => n17639, C1 => n24616, C2 =>
                           n7653, A => n21483, ZN => n21476);
   U22266 : OAI22_X1 port map( A1 => n20341, A2 => n24610, B1 => n20269, B2 => 
                           n24604, ZN => n21483);
   U22267 : AOI221_X1 port map( B1 => n24718, B2 => n19824, C1 => n24712, C2 =>
                           n19860, A => n21456, ZN => n21449);
   U22268 : OAI22_X1 port map( A1 => n20448, A2 => n24706, B1 => n20657, B2 => 
                           n24700, ZN => n21456);
   U22269 : AOI221_X1 port map( B1 => n24622, B2 => n17642, C1 => n24616, C2 =>
                           n7652, A => n21464, ZN => n21457);
   U22270 : OAI22_X1 port map( A1 => n20340, A2 => n24610, B1 => n20268, B2 => 
                           n24604, ZN => n21464);
   U22271 : AOI221_X1 port map( B1 => n24718, B2 => n19823, C1 => n24712, C2 =>
                           n19859, A => n21437, ZN => n21430);
   U22272 : OAI22_X1 port map( A1 => n20447, A2 => n24706, B1 => n20656, B2 => 
                           n24700, ZN => n21437);
   U22273 : AOI221_X1 port map( B1 => n24622, B2 => n17645, C1 => n24616, C2 =>
                           n7651, A => n21445, ZN => n21438);
   U22274 : OAI22_X1 port map( A1 => n20339, A2 => n24610, B1 => n20267, B2 => 
                           n24604, ZN => n21445);
   U22275 : AOI221_X1 port map( B1 => n24718, B2 => n19822, C1 => n24712, C2 =>
                           n19858, A => n21418, ZN => n21411);
   U22276 : OAI22_X1 port map( A1 => n20446, A2 => n24706, B1 => n20655, B2 => 
                           n24700, ZN => n21418);
   U22277 : AOI221_X1 port map( B1 => n24622, B2 => n17648, C1 => n24616, C2 =>
                           n7650, A => n21426, ZN => n21419);
   U22278 : OAI22_X1 port map( A1 => n20338, A2 => n24610, B1 => n20266, B2 => 
                           n24604, ZN => n21426);
   U22279 : AOI221_X1 port map( B1 => n24719, B2 => n19805, C1 => n24713, C2 =>
                           n19809, A => n21399, ZN => n21392);
   U22280 : OAI22_X1 port map( A1 => n20265, A2 => n24707, B1 => n20521, B2 => 
                           n24701, ZN => n21399);
   U22281 : AOI221_X1 port map( B1 => n24623, B2 => n17651, C1 => n24617, C2 =>
                           n7649, A => n21407, ZN => n21400);
   U22282 : OAI22_X1 port map( A1 => n20261, A2 => n24611, B1 => n20253, B2 => 
                           n24605, ZN => n21407);
   U22283 : AOI221_X1 port map( B1 => n24719, B2 => n19804, C1 => n24713, C2 =>
                           n19808, A => n21380, ZN => n21373);
   U22284 : OAI22_X1 port map( A1 => n20264, A2 => n24707, B1 => n20520, B2 => 
                           n24701, ZN => n21380);
   U22285 : AOI221_X1 port map( B1 => n24623, B2 => n17654, C1 => n24617, C2 =>
                           n7648, A => n21388, ZN => n21381);
   U22286 : OAI22_X1 port map( A1 => n20260, A2 => n24611, B1 => n20252, B2 => 
                           n24605, ZN => n21388);
   U22287 : AOI221_X1 port map( B1 => n24719, B2 => n19803, C1 => n24713, C2 =>
                           n19807, A => n21361, ZN => n21354);
   U22288 : OAI22_X1 port map( A1 => n20263, A2 => n24707, B1 => n20519, B2 => 
                           n24701, ZN => n21361);
   U22289 : AOI221_X1 port map( B1 => n24623, B2 => n17657, C1 => n24617, C2 =>
                           n7647, A => n21369, ZN => n21362);
   U22290 : OAI22_X1 port map( A1 => n20259, A2 => n24611, B1 => n20251, B2 => 
                           n24605, ZN => n21369);
   U22291 : AOI221_X1 port map( B1 => n24719, B2 => n19802, C1 => n24713, C2 =>
                           n19806, A => n21324, ZN => n21303);
   U22292 : OAI22_X1 port map( A1 => n20262, A2 => n24707, B1 => n20518, B2 => 
                           n24701, ZN => n21324);
   U22293 : AOI221_X1 port map( B1 => n24623, B2 => n17660, C1 => n24617, C2 =>
                           n7646, A => n21348, ZN => n21327);
   U22294 : OAI22_X1 port map( A1 => n20258, A2 => n24611, B1 => n20250, B2 => 
                           n24605, ZN => n21348);
   U22295 : OAI221_X1 port map( B1 => n7346, B2 => n24597, C1 => n7474, C2 => 
                           n24591, A => n23016, ZN => n23015);
   U22296 : AOI22_X1 port map( A1 => n24585, A2 => n7989, B1 => n24579, B2 => 
                           n19547, ZN => n23016);
   U22297 : OAI221_X1 port map( B1 => n7344, B2 => n24597, C1 => n7472, C2 => 
                           n24591, A => n22998, ZN => n22997);
   U22298 : AOI22_X1 port map( A1 => n24585, A2 => n7988, B1 => n24579, B2 => 
                           n19546, ZN => n22998);
   U22299 : OAI221_X1 port map( B1 => n7342, B2 => n24597, C1 => n7470, C2 => 
                           n24591, A => n22980, ZN => n22979);
   U22300 : AOI22_X1 port map( A1 => n24585, A2 => n7987, B1 => n24579, B2 => 
                           n19545, ZN => n22980);
   U22301 : OAI221_X1 port map( B1 => n7340, B2 => n24597, C1 => n7468, C2 => 
                           n24591, A => n22962, ZN => n22961);
   U22302 : AOI22_X1 port map( A1 => n24585, A2 => n7986, B1 => n24579, B2 => 
                           n19544, ZN => n22962);
   U22303 : OAI221_X1 port map( B1 => n7338, B2 => n24597, C1 => n7466, C2 => 
                           n24591, A => n22944, ZN => n22943);
   U22304 : AOI22_X1 port map( A1 => n24585, A2 => n7985, B1 => n24579, B2 => 
                           n19543, ZN => n22944);
   U22305 : OAI221_X1 port map( B1 => n7336, B2 => n24597, C1 => n7464, C2 => 
                           n24591, A => n22926, ZN => n22925);
   U22306 : AOI22_X1 port map( A1 => n24585, A2 => n7984, B1 => n24579, B2 => 
                           n19542, ZN => n22926);
   U22307 : OAI221_X1 port map( B1 => n7334, B2 => n24597, C1 => n7462, C2 => 
                           n24591, A => n22908, ZN => n22907);
   U22308 : AOI22_X1 port map( A1 => n24585, A2 => n7983, B1 => n24579, B2 => 
                           n19541, ZN => n22908);
   U22309 : OAI221_X1 port map( B1 => n7332, B2 => n24597, C1 => n7460, C2 => 
                           n24591, A => n22890, ZN => n22889);
   U22310 : AOI22_X1 port map( A1 => n24585, A2 => n7982, B1 => n24579, B2 => 
                           n19540, ZN => n22890);
   U22311 : OAI221_X1 port map( B1 => n7330, B2 => n24598, C1 => n7458, C2 => 
                           n24592, A => n22872, ZN => n22871);
   U22312 : AOI22_X1 port map( A1 => n24586, A2 => n7981, B1 => n24580, B2 => 
                           n19539, ZN => n22872);
   U22313 : OAI221_X1 port map( B1 => n7328, B2 => n24598, C1 => n7456, C2 => 
                           n24592, A => n22854, ZN => n22853);
   U22314 : AOI22_X1 port map( A1 => n24586, A2 => n7980, B1 => n24580, B2 => 
                           n19538, ZN => n22854);
   U22315 : OAI221_X1 port map( B1 => n7326, B2 => n24598, C1 => n7454, C2 => 
                           n24592, A => n22836, ZN => n22835);
   U22316 : AOI22_X1 port map( A1 => n24586, A2 => n7979, B1 => n24580, B2 => 
                           n19537, ZN => n22836);
   U22317 : OAI221_X1 port map( B1 => n7324, B2 => n24598, C1 => n7452, C2 => 
                           n24592, A => n22818, ZN => n22817);
   U22318 : AOI22_X1 port map( A1 => n24586, A2 => n7978, B1 => n24580, B2 => 
                           n19536, ZN => n22818);
   U22319 : OAI221_X1 port map( B1 => n7322, B2 => n24598, C1 => n7450, C2 => 
                           n24592, A => n22800, ZN => n22799);
   U22320 : AOI22_X1 port map( A1 => n24586, A2 => n7977, B1 => n24580, B2 => 
                           n19535, ZN => n22800);
   U22321 : OAI221_X1 port map( B1 => n7320, B2 => n24598, C1 => n7448, C2 => 
                           n24592, A => n22782, ZN => n22781);
   U22322 : AOI22_X1 port map( A1 => n24586, A2 => n7976, B1 => n24580, B2 => 
                           n19534, ZN => n22782);
   U22323 : OAI221_X1 port map( B1 => n7318, B2 => n24598, C1 => n7446, C2 => 
                           n24592, A => n22764, ZN => n22763);
   U22324 : AOI22_X1 port map( A1 => n24586, A2 => n7975, B1 => n24580, B2 => 
                           n19533, ZN => n22764);
   U22325 : OAI221_X1 port map( B1 => n7316, B2 => n24598, C1 => n7444, C2 => 
                           n24592, A => n22746, ZN => n22745);
   U22326 : AOI22_X1 port map( A1 => n24586, A2 => n7974, B1 => n24580, B2 => 
                           n19532, ZN => n22746);
   U22327 : OAI221_X1 port map( B1 => n7314, B2 => n24598, C1 => n7442, C2 => 
                           n24592, A => n22728, ZN => n22727);
   U22328 : AOI22_X1 port map( A1 => n24586, A2 => n7973, B1 => n24580, B2 => 
                           n19531, ZN => n22728);
   U22329 : OAI221_X1 port map( B1 => n7312, B2 => n24598, C1 => n7440, C2 => 
                           n24592, A => n22710, ZN => n22709);
   U22330 : AOI22_X1 port map( A1 => n24586, A2 => n7972, B1 => n24580, B2 => 
                           n19530, ZN => n22710);
   U22331 : OAI221_X1 port map( B1 => n7310, B2 => n24598, C1 => n7438, C2 => 
                           n24592, A => n22692, ZN => n22691);
   U22332 : AOI22_X1 port map( A1 => n24586, A2 => n7971, B1 => n24580, B2 => 
                           n19529, ZN => n22692);
   U22333 : OAI221_X1 port map( B1 => n7308, B2 => n24598, C1 => n7436, C2 => 
                           n24592, A => n22674, ZN => n22673);
   U22334 : AOI22_X1 port map( A1 => n24586, A2 => n7970, B1 => n24580, B2 => 
                           n19528, ZN => n22674);
   U22335 : OAI221_X1 port map( B1 => n7402, B2 => n24595, C1 => n7530, C2 => 
                           n24589, A => n23520, ZN => n23519);
   U22336 : AOI22_X1 port map( A1 => n24583, A2 => n8017, B1 => n24577, B2 => 
                           n19575, ZN => n23520);
   U22337 : OAI221_X1 port map( B1 => n7400, B2 => n24595, C1 => n7528, C2 => 
                           n24589, A => n23502, ZN => n23501);
   U22338 : AOI22_X1 port map( A1 => n24583, A2 => n8016, B1 => n24577, B2 => 
                           n19574, ZN => n23502);
   U22339 : OAI221_X1 port map( B1 => n7398, B2 => n24595, C1 => n7526, C2 => 
                           n24589, A => n23484, ZN => n23483);
   U22340 : AOI22_X1 port map( A1 => n24583, A2 => n8015, B1 => n24577, B2 => 
                           n19573, ZN => n23484);
   U22341 : OAI221_X1 port map( B1 => n7396, B2 => n24595, C1 => n7524, C2 => 
                           n24589, A => n23466, ZN => n23465);
   U22342 : AOI22_X1 port map( A1 => n24583, A2 => n8014, B1 => n24577, B2 => 
                           n19572, ZN => n23466);
   U22343 : OAI221_X1 port map( B1 => n7394, B2 => n24595, C1 => n7522, C2 => 
                           n24589, A => n23448, ZN => n23447);
   U22344 : AOI22_X1 port map( A1 => n24583, A2 => n8013, B1 => n24577, B2 => 
                           n19571, ZN => n23448);
   U22345 : OAI221_X1 port map( B1 => n7392, B2 => n24595, C1 => n7520, C2 => 
                           n24589, A => n23430, ZN => n23429);
   U22346 : AOI22_X1 port map( A1 => n24583, A2 => n8012, B1 => n24577, B2 => 
                           n19570, ZN => n23430);
   U22347 : OAI221_X1 port map( B1 => n7390, B2 => n24595, C1 => n7518, C2 => 
                           n24589, A => n23412, ZN => n23411);
   U22348 : AOI22_X1 port map( A1 => n24583, A2 => n8011, B1 => n24577, B2 => 
                           n19569, ZN => n23412);
   U22349 : OAI221_X1 port map( B1 => n7388, B2 => n24595, C1 => n7516, C2 => 
                           n24589, A => n23394, ZN => n23393);
   U22350 : AOI22_X1 port map( A1 => n24583, A2 => n8010, B1 => n24577, B2 => 
                           n19568, ZN => n23394);
   U22351 : OAI221_X1 port map( B1 => n7386, B2 => n24595, C1 => n7514, C2 => 
                           n24589, A => n23376, ZN => n23375);
   U22352 : AOI22_X1 port map( A1 => n24583, A2 => n8009, B1 => n24577, B2 => 
                           n19567, ZN => n23376);
   U22353 : OAI221_X1 port map( B1 => n7384, B2 => n24595, C1 => n7512, C2 => 
                           n24589, A => n23358, ZN => n23357);
   U22354 : AOI22_X1 port map( A1 => n24583, A2 => n8008, B1 => n24577, B2 => 
                           n19566, ZN => n23358);
   U22355 : OAI221_X1 port map( B1 => n7382, B2 => n24595, C1 => n7510, C2 => 
                           n24589, A => n23340, ZN => n23339);
   U22356 : AOI22_X1 port map( A1 => n24583, A2 => n8007, B1 => n24577, B2 => 
                           n19565, ZN => n23340);
   U22357 : OAI221_X1 port map( B1 => n7380, B2 => n24595, C1 => n7508, C2 => 
                           n24589, A => n23322, ZN => n23321);
   U22358 : AOI22_X1 port map( A1 => n24583, A2 => n8006, B1 => n24577, B2 => 
                           n19564, ZN => n23322);
   U22359 : OAI221_X1 port map( B1 => n7378, B2 => n24596, C1 => n7506, C2 => 
                           n24590, A => n23304, ZN => n23303);
   U22360 : AOI22_X1 port map( A1 => n24584, A2 => n8005, B1 => n24578, B2 => 
                           n19563, ZN => n23304);
   U22361 : OAI221_X1 port map( B1 => n7376, B2 => n24596, C1 => n7504, C2 => 
                           n24590, A => n23286, ZN => n23285);
   U22362 : AOI22_X1 port map( A1 => n24584, A2 => n8004, B1 => n24578, B2 => 
                           n19562, ZN => n23286);
   U22363 : OAI221_X1 port map( B1 => n7374, B2 => n24596, C1 => n7502, C2 => 
                           n24590, A => n23268, ZN => n23267);
   U22364 : AOI22_X1 port map( A1 => n24584, A2 => n8003, B1 => n24578, B2 => 
                           n19561, ZN => n23268);
   U22365 : OAI221_X1 port map( B1 => n7372, B2 => n24596, C1 => n7500, C2 => 
                           n24590, A => n23250, ZN => n23249);
   U22366 : AOI22_X1 port map( A1 => n24584, A2 => n8002, B1 => n24578, B2 => 
                           n19560, ZN => n23250);
   U22367 : OAI221_X1 port map( B1 => n7370, B2 => n24596, C1 => n7498, C2 => 
                           n24590, A => n23232, ZN => n23231);
   U22368 : AOI22_X1 port map( A1 => n24584, A2 => n8001, B1 => n24578, B2 => 
                           n19559, ZN => n23232);
   U22369 : OAI221_X1 port map( B1 => n7368, B2 => n24596, C1 => n7496, C2 => 
                           n24590, A => n23214, ZN => n23213);
   U22370 : AOI22_X1 port map( A1 => n24584, A2 => n8000, B1 => n24578, B2 => 
                           n19558, ZN => n23214);
   U22371 : OAI221_X1 port map( B1 => n7366, B2 => n24596, C1 => n7494, C2 => 
                           n24590, A => n23196, ZN => n23195);
   U22372 : AOI22_X1 port map( A1 => n24584, A2 => n7999, B1 => n24578, B2 => 
                           n19557, ZN => n23196);
   U22373 : OAI221_X1 port map( B1 => n7364, B2 => n24596, C1 => n7492, C2 => 
                           n24590, A => n23178, ZN => n23177);
   U22374 : AOI22_X1 port map( A1 => n24584, A2 => n7998, B1 => n24578, B2 => 
                           n19556, ZN => n23178);
   U22375 : OAI221_X1 port map( B1 => n7362, B2 => n24596, C1 => n7490, C2 => 
                           n24590, A => n23160, ZN => n23159);
   U22376 : AOI22_X1 port map( A1 => n24584, A2 => n7997, B1 => n24578, B2 => 
                           n19555, ZN => n23160);
   U22377 : OAI221_X1 port map( B1 => n7360, B2 => n24596, C1 => n7488, C2 => 
                           n24590, A => n23142, ZN => n23141);
   U22378 : AOI22_X1 port map( A1 => n24584, A2 => n7996, B1 => n24578, B2 => 
                           n19554, ZN => n23142);
   U22379 : OAI221_X1 port map( B1 => n7358, B2 => n24596, C1 => n7486, C2 => 
                           n24590, A => n23124, ZN => n23123);
   U22380 : AOI22_X1 port map( A1 => n24584, A2 => n7995, B1 => n24578, B2 => 
                           n19553, ZN => n23124);
   U22381 : OAI221_X1 port map( B1 => n7356, B2 => n24596, C1 => n7484, C2 => 
                           n24590, A => n23106, ZN => n23105);
   U22382 : AOI22_X1 port map( A1 => n24584, A2 => n7994, B1 => n24578, B2 => 
                           n19552, ZN => n23106);
   U22383 : OAI221_X1 port map( B1 => n7354, B2 => n24597, C1 => n7482, C2 => 
                           n24591, A => n23088, ZN => n23087);
   U22384 : AOI22_X1 port map( A1 => n24585, A2 => n7993, B1 => n24579, B2 => 
                           n19551, ZN => n23088);
   U22385 : OAI221_X1 port map( B1 => n7352, B2 => n24597, C1 => n7480, C2 => 
                           n24591, A => n23070, ZN => n23069);
   U22386 : AOI22_X1 port map( A1 => n24585, A2 => n7992, B1 => n24579, B2 => 
                           n19550, ZN => n23070);
   U22387 : OAI221_X1 port map( B1 => n7350, B2 => n24597, C1 => n7478, C2 => 
                           n24591, A => n23052, ZN => n23051);
   U22388 : AOI22_X1 port map( A1 => n24585, A2 => n7991, B1 => n24579, B2 => 
                           n19549, ZN => n23052);
   U22389 : OAI221_X1 port map( B1 => n7348, B2 => n24597, C1 => n7476, C2 => 
                           n24591, A => n23034, ZN => n23033);
   U22390 : AOI22_X1 port map( A1 => n24585, A2 => n7990, B1 => n24579, B2 => 
                           n19548, ZN => n23034);
   U22391 : OAI221_X1 port map( B1 => n7306, B2 => n24599, C1 => n7434, C2 => 
                           n24593, A => n22656, ZN => n22655);
   U22392 : AOI22_X1 port map( A1 => n24587, A2 => n7969, B1 => n24581, B2 => 
                           n19527, ZN => n22656);
   U22393 : OAI221_X1 port map( B1 => n7304, B2 => n24599, C1 => n7432, C2 => 
                           n24593, A => n22638, ZN => n22637);
   U22394 : AOI22_X1 port map( A1 => n24587, A2 => n7968, B1 => n24581, B2 => 
                           n19526, ZN => n22638);
   U22395 : OAI221_X1 port map( B1 => n7302, B2 => n24599, C1 => n7430, C2 => 
                           n24593, A => n22620, ZN => n22619);
   U22396 : AOI22_X1 port map( A1 => n24587, A2 => n7967, B1 => n24581, B2 => 
                           n19525, ZN => n22620);
   U22397 : OAI221_X1 port map( B1 => n7300, B2 => n24599, C1 => n7428, C2 => 
                           n24593, A => n22570, ZN => n22567);
   U22398 : AOI22_X1 port map( A1 => n24587, A2 => n7966, B1 => n24581, B2 => 
                           n19524, ZN => n22570);
   U22399 : OAI221_X1 port map( B1 => n7426, B2 => n24594, C1 => n7554, C2 => 
                           n24588, A => n23736, ZN => n23735);
   U22400 : AOI22_X1 port map( A1 => n24582, A2 => n8029, B1 => n24576, B2 => 
                           n19587, ZN => n23736);
   U22401 : OAI221_X1 port map( B1 => n7424, B2 => n24594, C1 => n7552, C2 => 
                           n24588, A => n23718, ZN => n23717);
   U22402 : AOI22_X1 port map( A1 => n24582, A2 => n8028, B1 => n24576, B2 => 
                           n19586, ZN => n23718);
   U22403 : OAI221_X1 port map( B1 => n7422, B2 => n24594, C1 => n7550, C2 => 
                           n24588, A => n23700, ZN => n23699);
   U22404 : AOI22_X1 port map( A1 => n24582, A2 => n8027, B1 => n24576, B2 => 
                           n19585, ZN => n23700);
   U22405 : OAI221_X1 port map( B1 => n7420, B2 => n24594, C1 => n7548, C2 => 
                           n24588, A => n23682, ZN => n23681);
   U22406 : AOI22_X1 port map( A1 => n24582, A2 => n8026, B1 => n24576, B2 => 
                           n19584, ZN => n23682);
   U22407 : OAI221_X1 port map( B1 => n7418, B2 => n24594, C1 => n7546, C2 => 
                           n24588, A => n23664, ZN => n23663);
   U22408 : AOI22_X1 port map( A1 => n24582, A2 => n8025, B1 => n24576, B2 => 
                           n19583, ZN => n23664);
   U22409 : OAI221_X1 port map( B1 => n7416, B2 => n24594, C1 => n7544, C2 => 
                           n24588, A => n23646, ZN => n23645);
   U22410 : AOI22_X1 port map( A1 => n24582, A2 => n8024, B1 => n24576, B2 => 
                           n19582, ZN => n23646);
   U22411 : OAI221_X1 port map( B1 => n7414, B2 => n24594, C1 => n7542, C2 => 
                           n24588, A => n23628, ZN => n23627);
   U22412 : AOI22_X1 port map( A1 => n24582, A2 => n8023, B1 => n24576, B2 => 
                           n19581, ZN => n23628);
   U22413 : OAI221_X1 port map( B1 => n7412, B2 => n24594, C1 => n7540, C2 => 
                           n24588, A => n23610, ZN => n23609);
   U22414 : AOI22_X1 port map( A1 => n24582, A2 => n8022, B1 => n24576, B2 => 
                           n19580, ZN => n23610);
   U22415 : OAI221_X1 port map( B1 => n7410, B2 => n24594, C1 => n7538, C2 => 
                           n24588, A => n23592, ZN => n23591);
   U22416 : AOI22_X1 port map( A1 => n24582, A2 => n8021, B1 => n24576, B2 => 
                           n19579, ZN => n23592);
   U22417 : OAI221_X1 port map( B1 => n7408, B2 => n24594, C1 => n7536, C2 => 
                           n24588, A => n23574, ZN => n23573);
   U22418 : AOI22_X1 port map( A1 => n24582, A2 => n8020, B1 => n24576, B2 => 
                           n19578, ZN => n23574);
   U22419 : OAI221_X1 port map( B1 => n7406, B2 => n24594, C1 => n7534, C2 => 
                           n24588, A => n23556, ZN => n23555);
   U22420 : AOI22_X1 port map( A1 => n24582, A2 => n8019, B1 => n24576, B2 => 
                           n19577, ZN => n23556);
   U22421 : OAI221_X1 port map( B1 => n7404, B2 => n24594, C1 => n7532, C2 => 
                           n24588, A => n23538, ZN => n23537);
   U22422 : AOI22_X1 port map( A1 => n24582, A2 => n8018, B1 => n24576, B2 => 
                           n19576, ZN => n23538);
   U22423 : OAI22_X1 port map( A1 => n20152, A2 => n24407, B1 => n8869, B2 => 
                           n24401, ZN => n22665);
   U22424 : OAI22_X1 port map( A1 => n9124, A2 => n24431, B1 => n9125, B2 => 
                           n24425, ZN => n22664);
   U22425 : OAI22_X1 port map( A1 => n20151, A2 => n24407, B1 => n8867, B2 => 
                           n24401, ZN => n22647);
   U22426 : OAI22_X1 port map( A1 => n9122, A2 => n24431, B1 => n9123, B2 => 
                           n24425, ZN => n22646);
   U22427 : OAI22_X1 port map( A1 => n20150, A2 => n24407, B1 => n8865, B2 => 
                           n24401, ZN => n22629);
   U22428 : OAI22_X1 port map( A1 => n9120, A2 => n24431, B1 => n9121, B2 => 
                           n24425, ZN => n22628);
   U22429 : OAI22_X1 port map( A1 => n20149, A2 => n24407, B1 => n8863, B2 => 
                           n24401, ZN => n22609);
   U22430 : OAI22_X1 port map( A1 => n9118, A2 => n24431, B1 => n9119, B2 => 
                           n24425, ZN => n22604);
   U22431 : OAI22_X1 port map( A1 => n19667, A2 => n24405, B1 => n8909, B2 => 
                           n24399, ZN => n23025);
   U22432 : OAI22_X1 port map( A1 => n9164, A2 => n24429, B1 => n9165, B2 => 
                           n24423, ZN => n23024);
   U22433 : OAI22_X1 port map( A1 => n19666, A2 => n24405, B1 => n8907, B2 => 
                           n24399, ZN => n23007);
   U22434 : OAI22_X1 port map( A1 => n9162, A2 => n24429, B1 => n9163, B2 => 
                           n24423, ZN => n23006);
   U22435 : OAI22_X1 port map( A1 => n19665, A2 => n24405, B1 => n8905, B2 => 
                           n24399, ZN => n22989);
   U22436 : OAI22_X1 port map( A1 => n9160, A2 => n24429, B1 => n9161, B2 => 
                           n24423, ZN => n22988);
   U22437 : OAI22_X1 port map( A1 => n19664, A2 => n24405, B1 => n8903, B2 => 
                           n24399, ZN => n22971);
   U22438 : OAI22_X1 port map( A1 => n9158, A2 => n24429, B1 => n9159, B2 => 
                           n24423, ZN => n22970);
   U22439 : OAI22_X1 port map( A1 => n19663, A2 => n24405, B1 => n8901, B2 => 
                           n24399, ZN => n22953);
   U22440 : OAI22_X1 port map( A1 => n9156, A2 => n24429, B1 => n9157, B2 => 
                           n24423, ZN => n22952);
   U22441 : OAI22_X1 port map( A1 => n19662, A2 => n24405, B1 => n8899, B2 => 
                           n24399, ZN => n22935);
   U22442 : OAI22_X1 port map( A1 => n9154, A2 => n24429, B1 => n9155, B2 => 
                           n24423, ZN => n22934);
   U22443 : OAI22_X1 port map( A1 => n19661, A2 => n24405, B1 => n8897, B2 => 
                           n24399, ZN => n22917);
   U22444 : OAI22_X1 port map( A1 => n9152, A2 => n24429, B1 => n9153, B2 => 
                           n24423, ZN => n22916);
   U22445 : OAI22_X1 port map( A1 => n19660, A2 => n24405, B1 => n8895, B2 => 
                           n24399, ZN => n22899);
   U22446 : OAI22_X1 port map( A1 => n9150, A2 => n24429, B1 => n9151, B2 => 
                           n24423, ZN => n22898);
   U22447 : OAI22_X1 port map( A1 => n19659, A2 => n24406, B1 => n8893, B2 => 
                           n24400, ZN => n22881);
   U22448 : OAI22_X1 port map( A1 => n9148, A2 => n24430, B1 => n9149, B2 => 
                           n24424, ZN => n22880);
   U22449 : OAI22_X1 port map( A1 => n19658, A2 => n24406, B1 => n8891, B2 => 
                           n24400, ZN => n22863);
   U22450 : OAI22_X1 port map( A1 => n9146, A2 => n24430, B1 => n9147, B2 => 
                           n24424, ZN => n22862);
   U22451 : OAI22_X1 port map( A1 => n19657, A2 => n24406, B1 => n8889, B2 => 
                           n24400, ZN => n22845);
   U22452 : OAI22_X1 port map( A1 => n9144, A2 => n24430, B1 => n9145, B2 => 
                           n24424, ZN => n22844);
   U22453 : OAI22_X1 port map( A1 => n19656, A2 => n24406, B1 => n8887, B2 => 
                           n24400, ZN => n22827);
   U22454 : OAI22_X1 port map( A1 => n9142, A2 => n24430, B1 => n9143, B2 => 
                           n24424, ZN => n22826);
   U22455 : OAI22_X1 port map( A1 => n19655, A2 => n24406, B1 => n8885, B2 => 
                           n24400, ZN => n22809);
   U22456 : OAI22_X1 port map( A1 => n9140, A2 => n24430, B1 => n9141, B2 => 
                           n24424, ZN => n22808);
   U22457 : OAI22_X1 port map( A1 => n19654, A2 => n24406, B1 => n8883, B2 => 
                           n24400, ZN => n22791);
   U22458 : OAI22_X1 port map( A1 => n9138, A2 => n24430, B1 => n9139, B2 => 
                           n24424, ZN => n22790);
   U22459 : OAI22_X1 port map( A1 => n19653, A2 => n24406, B1 => n8881, B2 => 
                           n24400, ZN => n22773);
   U22460 : OAI22_X1 port map( A1 => n9136, A2 => n24430, B1 => n9137, B2 => 
                           n24424, ZN => n22772);
   U22461 : OAI22_X1 port map( A1 => n19652, A2 => n24406, B1 => n8879, B2 => 
                           n24400, ZN => n22755);
   U22462 : OAI22_X1 port map( A1 => n9134, A2 => n24430, B1 => n9135, B2 => 
                           n24424, ZN => n22754);
   U22463 : OAI22_X1 port map( A1 => n19651, A2 => n24406, B1 => n8877, B2 => 
                           n24400, ZN => n22737);
   U22464 : OAI22_X1 port map( A1 => n9132, A2 => n24430, B1 => n9133, B2 => 
                           n24424, ZN => n22736);
   U22465 : OAI22_X1 port map( A1 => n19650, A2 => n24406, B1 => n8875, B2 => 
                           n24400, ZN => n22719);
   U22466 : OAI22_X1 port map( A1 => n9130, A2 => n24430, B1 => n9131, B2 => 
                           n24424, ZN => n22718);
   U22467 : OAI22_X1 port map( A1 => n19649, A2 => n24406, B1 => n8873, B2 => 
                           n24400, ZN => n22701);
   U22468 : OAI22_X1 port map( A1 => n9128, A2 => n24430, B1 => n9129, B2 => 
                           n24424, ZN => n22700);
   U22469 : OAI22_X1 port map( A1 => n19648, A2 => n24406, B1 => n8871, B2 => 
                           n24400, ZN => n22683);
   U22470 : OAI22_X1 port map( A1 => n9126, A2 => n24430, B1 => n9127, B2 => 
                           n24424, ZN => n22682);
   U22471 : OAI22_X1 port map( A1 => n19707, A2 => n24402, B1 => n8989, B2 => 
                           n24396, ZN => n23763);
   U22472 : OAI22_X1 port map( A1 => n9244, A2 => n24426, B1 => n9245, B2 => 
                           n24420, ZN => n23762);
   U22473 : OAI22_X1 port map( A1 => n19706, A2 => n24402, B1 => n8987, B2 => 
                           n24396, ZN => n23727);
   U22474 : OAI22_X1 port map( A1 => n9242, A2 => n24426, B1 => n9243, B2 => 
                           n24420, ZN => n23726);
   U22475 : OAI22_X1 port map( A1 => n19705, A2 => n24402, B1 => n8985, B2 => 
                           n24396, ZN => n23709);
   U22476 : OAI22_X1 port map( A1 => n9240, A2 => n24426, B1 => n9241, B2 => 
                           n24420, ZN => n23708);
   U22477 : OAI22_X1 port map( A1 => n19704, A2 => n24402, B1 => n8983, B2 => 
                           n24396, ZN => n23691);
   U22478 : OAI22_X1 port map( A1 => n9238, A2 => n24426, B1 => n9239, B2 => 
                           n24420, ZN => n23690);
   U22479 : OAI22_X1 port map( A1 => n19703, A2 => n24402, B1 => n8981, B2 => 
                           n24396, ZN => n23673);
   U22480 : OAI22_X1 port map( A1 => n9236, A2 => n24426, B1 => n9237, B2 => 
                           n24420, ZN => n23672);
   U22481 : OAI22_X1 port map( A1 => n19702, A2 => n24402, B1 => n8979, B2 => 
                           n24396, ZN => n23655);
   U22482 : OAI22_X1 port map( A1 => n9234, A2 => n24426, B1 => n9235, B2 => 
                           n24420, ZN => n23654);
   U22483 : OAI22_X1 port map( A1 => n19701, A2 => n24402, B1 => n8977, B2 => 
                           n24396, ZN => n23637);
   U22484 : OAI22_X1 port map( A1 => n9232, A2 => n24426, B1 => n9233, B2 => 
                           n24420, ZN => n23636);
   U22485 : OAI22_X1 port map( A1 => n19700, A2 => n24402, B1 => n8975, B2 => 
                           n24396, ZN => n23619);
   U22486 : OAI22_X1 port map( A1 => n9230, A2 => n24426, B1 => n9231, B2 => 
                           n24420, ZN => n23618);
   U22487 : OAI22_X1 port map( A1 => n19699, A2 => n24402, B1 => n8973, B2 => 
                           n24396, ZN => n23601);
   U22488 : OAI22_X1 port map( A1 => n9228, A2 => n24426, B1 => n9229, B2 => 
                           n24420, ZN => n23600);
   U22489 : OAI22_X1 port map( A1 => n19698, A2 => n24402, B1 => n8971, B2 => 
                           n24396, ZN => n23583);
   U22490 : OAI22_X1 port map( A1 => n9226, A2 => n24426, B1 => n9227, B2 => 
                           n24420, ZN => n23582);
   U22491 : OAI22_X1 port map( A1 => n19697, A2 => n24402, B1 => n8969, B2 => 
                           n24396, ZN => n23565);
   U22492 : OAI22_X1 port map( A1 => n9224, A2 => n24426, B1 => n9225, B2 => 
                           n24420, ZN => n23564);
   U22493 : OAI22_X1 port map( A1 => n19696, A2 => n24402, B1 => n8967, B2 => 
                           n24396, ZN => n23547);
   U22494 : OAI22_X1 port map( A1 => n9222, A2 => n24426, B1 => n9223, B2 => 
                           n24420, ZN => n23546);
   U22495 : OAI22_X1 port map( A1 => n19695, A2 => n24403, B1 => n8965, B2 => 
                           n24397, ZN => n23529);
   U22496 : OAI22_X1 port map( A1 => n9220, A2 => n24427, B1 => n9221, B2 => 
                           n24421, ZN => n23528);
   U22497 : OAI22_X1 port map( A1 => n19694, A2 => n24403, B1 => n8963, B2 => 
                           n24397, ZN => n23511);
   U22498 : OAI22_X1 port map( A1 => n9218, A2 => n24427, B1 => n9219, B2 => 
                           n24421, ZN => n23510);
   U22499 : OAI22_X1 port map( A1 => n19693, A2 => n24403, B1 => n8961, B2 => 
                           n24397, ZN => n23493);
   U22500 : OAI22_X1 port map( A1 => n9216, A2 => n24427, B1 => n9217, B2 => 
                           n24421, ZN => n23492);
   U22501 : OAI22_X1 port map( A1 => n19692, A2 => n24403, B1 => n8959, B2 => 
                           n24397, ZN => n23475);
   U22502 : OAI22_X1 port map( A1 => n9214, A2 => n24427, B1 => n9215, B2 => 
                           n24421, ZN => n23474);
   U22503 : OAI22_X1 port map( A1 => n19691, A2 => n24403, B1 => n8957, B2 => 
                           n24397, ZN => n23457);
   U22504 : OAI22_X1 port map( A1 => n9212, A2 => n24427, B1 => n9213, B2 => 
                           n24421, ZN => n23456);
   U22505 : OAI22_X1 port map( A1 => n19690, A2 => n24403, B1 => n8955, B2 => 
                           n24397, ZN => n23439);
   U22506 : OAI22_X1 port map( A1 => n9210, A2 => n24427, B1 => n9211, B2 => 
                           n24421, ZN => n23438);
   U22507 : OAI22_X1 port map( A1 => n19689, A2 => n24403, B1 => n8953, B2 => 
                           n24397, ZN => n23421);
   U22508 : OAI22_X1 port map( A1 => n9208, A2 => n24427, B1 => n9209, B2 => 
                           n24421, ZN => n23420);
   U22509 : OAI22_X1 port map( A1 => n19688, A2 => n24403, B1 => n8951, B2 => 
                           n24397, ZN => n23403);
   U22510 : OAI22_X1 port map( A1 => n9206, A2 => n24427, B1 => n9207, B2 => 
                           n24421, ZN => n23402);
   U22511 : OAI22_X1 port map( A1 => n19687, A2 => n24403, B1 => n8949, B2 => 
                           n24397, ZN => n23385);
   U22512 : OAI22_X1 port map( A1 => n9204, A2 => n24427, B1 => n9205, B2 => 
                           n24421, ZN => n23384);
   U22513 : OAI22_X1 port map( A1 => n19686, A2 => n24403, B1 => n8947, B2 => 
                           n24397, ZN => n23367);
   U22514 : OAI22_X1 port map( A1 => n9202, A2 => n24427, B1 => n9203, B2 => 
                           n24421, ZN => n23366);
   U22515 : OAI22_X1 port map( A1 => n19685, A2 => n24403, B1 => n8945, B2 => 
                           n24397, ZN => n23349);
   U22516 : OAI22_X1 port map( A1 => n9200, A2 => n24427, B1 => n9201, B2 => 
                           n24421, ZN => n23348);
   U22517 : OAI22_X1 port map( A1 => n19684, A2 => n24403, B1 => n8943, B2 => 
                           n24397, ZN => n23331);
   U22518 : OAI22_X1 port map( A1 => n9198, A2 => n24427, B1 => n9199, B2 => 
                           n24421, ZN => n23330);
   U22519 : OAI22_X1 port map( A1 => n19683, A2 => n24404, B1 => n8941, B2 => 
                           n24398, ZN => n23313);
   U22520 : OAI22_X1 port map( A1 => n9196, A2 => n24428, B1 => n9197, B2 => 
                           n24422, ZN => n23312);
   U22521 : OAI22_X1 port map( A1 => n19682, A2 => n24404, B1 => n8939, B2 => 
                           n24398, ZN => n23295);
   U22522 : OAI22_X1 port map( A1 => n9194, A2 => n24428, B1 => n9195, B2 => 
                           n24422, ZN => n23294);
   U22523 : OAI22_X1 port map( A1 => n19681, A2 => n24404, B1 => n8937, B2 => 
                           n24398, ZN => n23277);
   U22524 : OAI22_X1 port map( A1 => n9192, A2 => n24428, B1 => n9193, B2 => 
                           n24422, ZN => n23276);
   U22525 : OAI22_X1 port map( A1 => n19680, A2 => n24404, B1 => n8935, B2 => 
                           n24398, ZN => n23259);
   U22526 : OAI22_X1 port map( A1 => n9190, A2 => n24428, B1 => n9191, B2 => 
                           n24422, ZN => n23258);
   U22527 : OAI22_X1 port map( A1 => n19679, A2 => n24404, B1 => n8933, B2 => 
                           n24398, ZN => n23241);
   U22528 : OAI22_X1 port map( A1 => n9188, A2 => n24428, B1 => n9189, B2 => 
                           n24422, ZN => n23240);
   U22529 : OAI22_X1 port map( A1 => n19678, A2 => n24404, B1 => n8931, B2 => 
                           n24398, ZN => n23223);
   U22530 : OAI22_X1 port map( A1 => n9186, A2 => n24428, B1 => n9187, B2 => 
                           n24422, ZN => n23222);
   U22531 : OAI22_X1 port map( A1 => n19677, A2 => n24404, B1 => n8929, B2 => 
                           n24398, ZN => n23205);
   U22532 : OAI22_X1 port map( A1 => n9184, A2 => n24428, B1 => n9185, B2 => 
                           n24422, ZN => n23204);
   U22533 : OAI22_X1 port map( A1 => n19676, A2 => n24404, B1 => n8927, B2 => 
                           n24398, ZN => n23187);
   U22534 : OAI22_X1 port map( A1 => n9182, A2 => n24428, B1 => n9183, B2 => 
                           n24422, ZN => n23186);
   U22535 : OAI22_X1 port map( A1 => n19675, A2 => n24404, B1 => n8925, B2 => 
                           n24398, ZN => n23169);
   U22536 : OAI22_X1 port map( A1 => n9180, A2 => n24428, B1 => n9181, B2 => 
                           n24422, ZN => n23168);
   U22537 : OAI22_X1 port map( A1 => n19674, A2 => n24404, B1 => n8923, B2 => 
                           n24398, ZN => n23151);
   U22538 : OAI22_X1 port map( A1 => n9178, A2 => n24428, B1 => n9179, B2 => 
                           n24422, ZN => n23150);
   U22539 : OAI22_X1 port map( A1 => n19673, A2 => n24404, B1 => n8921, B2 => 
                           n24398, ZN => n23133);
   U22540 : OAI22_X1 port map( A1 => n9176, A2 => n24428, B1 => n9177, B2 => 
                           n24422, ZN => n23132);
   U22541 : OAI22_X1 port map( A1 => n19672, A2 => n24404, B1 => n8919, B2 => 
                           n24398, ZN => n23115);
   U22542 : OAI22_X1 port map( A1 => n9174, A2 => n24428, B1 => n9175, B2 => 
                           n24422, ZN => n23114);
   U22543 : OAI22_X1 port map( A1 => n19671, A2 => n24405, B1 => n8917, B2 => 
                           n24399, ZN => n23097);
   U22544 : OAI22_X1 port map( A1 => n9172, A2 => n24429, B1 => n9173, B2 => 
                           n24423, ZN => n23096);
   U22545 : OAI22_X1 port map( A1 => n19670, A2 => n24405, B1 => n8915, B2 => 
                           n24399, ZN => n23079);
   U22546 : OAI22_X1 port map( A1 => n9170, A2 => n24429, B1 => n9171, B2 => 
                           n24423, ZN => n23078);
   U22547 : OAI22_X1 port map( A1 => n19669, A2 => n24405, B1 => n8913, B2 => 
                           n24399, ZN => n23061);
   U22548 : OAI22_X1 port map( A1 => n9168, A2 => n24429, B1 => n9169, B2 => 
                           n24423, ZN => n23060);
   U22549 : OAI22_X1 port map( A1 => n19668, A2 => n24405, B1 => n8911, B2 => 
                           n24399, ZN => n23043);
   U22550 : OAI22_X1 port map( A1 => n9166, A2 => n24429, B1 => n9167, B2 => 
                           n24423, ZN => n23042);
   U22551 : OAI22_X1 port map( A1 => n88, A2 => n24495, B1 => n20710, B2 => 
                           n24489, ZN => n23023);
   U22552 : OAI22_X1 port map( A1 => n87, A2 => n24495, B1 => n20709, B2 => 
                           n24489, ZN => n23005);
   U22553 : OAI22_X1 port map( A1 => n86, A2 => n24495, B1 => n20708, B2 => 
                           n24489, ZN => n22987);
   U22554 : OAI22_X1 port map( A1 => n85, A2 => n24495, B1 => n20707, B2 => 
                           n24489, ZN => n22969);
   U22555 : OAI22_X1 port map( A1 => n84, A2 => n24495, B1 => n20706, B2 => 
                           n24489, ZN => n22951);
   U22556 : OAI22_X1 port map( A1 => n83, A2 => n24495, B1 => n20705, B2 => 
                           n24489, ZN => n22933);
   U22557 : OAI22_X1 port map( A1 => n82, A2 => n24495, B1 => n20704, B2 => 
                           n24489, ZN => n22915);
   U22558 : OAI22_X1 port map( A1 => n81, A2 => n24495, B1 => n20703, B2 => 
                           n24489, ZN => n22897);
   U22559 : OAI22_X1 port map( A1 => n80, A2 => n24496, B1 => n20702, B2 => 
                           n24490, ZN => n22879);
   U22560 : OAI22_X1 port map( A1 => n79, A2 => n24496, B1 => n20701, B2 => 
                           n24490, ZN => n22861);
   U22561 : OAI22_X1 port map( A1 => n78, A2 => n24496, B1 => n20700, B2 => 
                           n24490, ZN => n22843);
   U22562 : OAI22_X1 port map( A1 => n77, A2 => n24496, B1 => n20699, B2 => 
                           n24490, ZN => n22825);
   U22563 : OAI22_X1 port map( A1 => n99, A2 => n24494, B1 => n20721, B2 => 
                           n24488, ZN => n23221);
   U22564 : OAI22_X1 port map( A1 => n98, A2 => n24494, B1 => n20720, B2 => 
                           n24488, ZN => n23203);
   U22565 : OAI22_X1 port map( A1 => n97, A2 => n24494, B1 => n20719, B2 => 
                           n24488, ZN => n23185);
   U22566 : OAI22_X1 port map( A1 => n96, A2 => n24494, B1 => n20718, B2 => 
                           n24488, ZN => n23167);
   U22567 : OAI22_X1 port map( A1 => n95, A2 => n24494, B1 => n20717, B2 => 
                           n24488, ZN => n23149);
   U22568 : OAI22_X1 port map( A1 => n94, A2 => n24494, B1 => n20716, B2 => 
                           n24488, ZN => n23131);
   U22569 : OAI22_X1 port map( A1 => n93, A2 => n24494, B1 => n20715, B2 => 
                           n24488, ZN => n23113);
   U22570 : OAI22_X1 port map( A1 => n92, A2 => n24495, B1 => n20714, B2 => 
                           n24489, ZN => n23095);
   U22571 : OAI22_X1 port map( A1 => n91, A2 => n24495, B1 => n20713, B2 => 
                           n24489, ZN => n23077);
   U22572 : OAI22_X1 port map( A1 => n90, A2 => n24495, B1 => n20712, B2 => 
                           n24489, ZN => n23059);
   U22573 : OAI22_X1 port map( A1 => n89, A2 => n24495, B1 => n20711, B2 => 
                           n24489, ZN => n23041);
   U22574 : AOI221_X1 port map( B1 => n24666, B2 => n24272, C1 => n24660, C2 =>
                           n24148, A => n22555, ZN => n22550);
   U22575 : OAI22_X1 port map( A1 => n20421, A2 => n24654, B1 => n21098, B2 => 
                           n24648, ZN => n22555);
   U22576 : AOI221_X1 port map( B1 => n24642, B2 => n17541, C1 => n24636, C2 =>
                           n24212, A => n22556, ZN => n22549);
   U22577 : OAI22_X1 port map( A1 => n20846, A2 => n24630, B1 => n21122, B2 => 
                           n24624, ZN => n22556);
   U22578 : AOI221_X1 port map( B1 => n24666, B2 => n24273, C1 => n24660, C2 =>
                           n24149, A => n22526, ZN => n22523);
   U22579 : OAI22_X1 port map( A1 => n20420, A2 => n24654, B1 => n21097, B2 => 
                           n24648, ZN => n22526);
   U22580 : AOI221_X1 port map( B1 => n24642, B2 => n17544, C1 => n24636, C2 =>
                           n24213, A => n22527, ZN => n22522);
   U22581 : OAI22_X1 port map( A1 => n20845, A2 => n24630, B1 => n21121, B2 => 
                           n24624, ZN => n22527);
   U22582 : AOI221_X1 port map( B1 => n24666, B2 => n24274, C1 => n24660, C2 =>
                           n24150, A => n22507, ZN => n22504);
   U22583 : OAI22_X1 port map( A1 => n20419, A2 => n24654, B1 => n21096, B2 => 
                           n24648, ZN => n22507);
   U22584 : AOI221_X1 port map( B1 => n24642, B2 => n17547, C1 => n24636, C2 =>
                           n24214, A => n22508, ZN => n22503);
   U22585 : OAI22_X1 port map( A1 => n20844, A2 => n24630, B1 => n21120, B2 => 
                           n24624, ZN => n22508);
   U22586 : AOI221_X1 port map( B1 => n24666, B2 => n24275, C1 => n24660, C2 =>
                           n24151, A => n22488, ZN => n22485);
   U22587 : OAI22_X1 port map( A1 => n20418, A2 => n24654, B1 => n21095, B2 => 
                           n24648, ZN => n22488);
   U22588 : AOI221_X1 port map( B1 => n24642, B2 => n17550, C1 => n24636, C2 =>
                           n24215, A => n22489, ZN => n22484);
   U22589 : OAI22_X1 port map( A1 => n20843, A2 => n24630, B1 => n21119, B2 => 
                           n24624, ZN => n22489);
   U22590 : AOI221_X1 port map( B1 => n24666, B2 => n24276, C1 => n24660, C2 =>
                           n24152, A => n22469, ZN => n22466);
   U22591 : OAI22_X1 port map( A1 => n20417, A2 => n24654, B1 => n21094, B2 => 
                           n24648, ZN => n22469);
   U22592 : AOI221_X1 port map( B1 => n24642, B2 => n17553, C1 => n24636, C2 =>
                           n24216, A => n22470, ZN => n22465);
   U22593 : OAI22_X1 port map( A1 => n20842, A2 => n24630, B1 => n21118, B2 => 
                           n24624, ZN => n22470);
   U22594 : AOI221_X1 port map( B1 => n24666, B2 => n24277, C1 => n24660, C2 =>
                           n24153, A => n22450, ZN => n22447);
   U22595 : OAI22_X1 port map( A1 => n20416, A2 => n24654, B1 => n21093, B2 => 
                           n24648, ZN => n22450);
   U22596 : AOI221_X1 port map( B1 => n24642, B2 => n17556, C1 => n24636, C2 =>
                           n24217, A => n22451, ZN => n22446);
   U22597 : OAI22_X1 port map( A1 => n20841, A2 => n24630, B1 => n21117, B2 => 
                           n24624, ZN => n22451);
   U22598 : AOI221_X1 port map( B1 => n24666, B2 => n24278, C1 => n24660, C2 =>
                           n24154, A => n22431, ZN => n22428);
   U22599 : OAI22_X1 port map( A1 => n20415, A2 => n24654, B1 => n21092, B2 => 
                           n24648, ZN => n22431);
   U22600 : AOI221_X1 port map( B1 => n24642, B2 => n17559, C1 => n24636, C2 =>
                           n24218, A => n22432, ZN => n22427);
   U22601 : OAI22_X1 port map( A1 => n20840, A2 => n24630, B1 => n21116, B2 => 
                           n24624, ZN => n22432);
   U22602 : AOI221_X1 port map( B1 => n24666, B2 => n24279, C1 => n24660, C2 =>
                           n24155, A => n22412, ZN => n22409);
   U22603 : OAI22_X1 port map( A1 => n20414, A2 => n24654, B1 => n21091, B2 => 
                           n24648, ZN => n22412);
   U22604 : AOI221_X1 port map( B1 => n24642, B2 => n17562, C1 => n24636, C2 =>
                           n24219, A => n22413, ZN => n22408);
   U22605 : OAI22_X1 port map( A1 => n20839, A2 => n24630, B1 => n21115, B2 => 
                           n24624, ZN => n22413);
   U22606 : AOI221_X1 port map( B1 => n24666, B2 => n24280, C1 => n24660, C2 =>
                           n24156, A => n22393, ZN => n22390);
   U22607 : OAI22_X1 port map( A1 => n20413, A2 => n24654, B1 => n21090, B2 => 
                           n24648, ZN => n22393);
   U22608 : AOI221_X1 port map( B1 => n24642, B2 => n17565, C1 => n24636, C2 =>
                           n24220, A => n22394, ZN => n22389);
   U22609 : OAI22_X1 port map( A1 => n20838, A2 => n24630, B1 => n21114, B2 => 
                           n24624, ZN => n22394);
   U22610 : AOI221_X1 port map( B1 => n24666, B2 => n24281, C1 => n24660, C2 =>
                           n24157, A => n22374, ZN => n22371);
   U22611 : OAI22_X1 port map( A1 => n20412, A2 => n24654, B1 => n21089, B2 => 
                           n24648, ZN => n22374);
   U22612 : AOI221_X1 port map( B1 => n24642, B2 => n17568, C1 => n24636, C2 =>
                           n24221, A => n22375, ZN => n22370);
   U22613 : OAI22_X1 port map( A1 => n20837, A2 => n24630, B1 => n21113, B2 => 
                           n24624, ZN => n22375);
   U22614 : AOI221_X1 port map( B1 => n24666, B2 => n24282, C1 => n24660, C2 =>
                           n24158, A => n22355, ZN => n22352);
   U22615 : OAI22_X1 port map( A1 => n20411, A2 => n24654, B1 => n21088, B2 => 
                           n24648, ZN => n22355);
   U22616 : AOI221_X1 port map( B1 => n24642, B2 => n17571, C1 => n24636, C2 =>
                           n24222, A => n22356, ZN => n22351);
   U22617 : OAI22_X1 port map( A1 => n20836, A2 => n24630, B1 => n21112, B2 => 
                           n24624, ZN => n22356);
   U22618 : AOI221_X1 port map( B1 => n24666, B2 => n24283, C1 => n24660, C2 =>
                           n24159, A => n22336, ZN => n22333);
   U22619 : OAI22_X1 port map( A1 => n20410, A2 => n24654, B1 => n21087, B2 => 
                           n24648, ZN => n22336);
   U22620 : AOI221_X1 port map( B1 => n24642, B2 => n17574, C1 => n24636, C2 =>
                           n24223, A => n22337, ZN => n22332);
   U22621 : OAI22_X1 port map( A1 => n20835, A2 => n24630, B1 => n21111, B2 => 
                           n24624, ZN => n22337);
   U22622 : AOI221_X1 port map( B1 => n24667, B2 => n24284, C1 => n24661, C2 =>
                           n24160, A => n22317, ZN => n22314);
   U22623 : OAI22_X1 port map( A1 => n20409, A2 => n24655, B1 => n21086, B2 => 
                           n24649, ZN => n22317);
   U22624 : AOI221_X1 port map( B1 => n24643, B2 => n17577, C1 => n24637, C2 =>
                           n24224, A => n22318, ZN => n22313);
   U22625 : OAI22_X1 port map( A1 => n20834, A2 => n24631, B1 => n21110, B2 => 
                           n24625, ZN => n22318);
   U22626 : AOI221_X1 port map( B1 => n24667, B2 => n24285, C1 => n24661, C2 =>
                           n24161, A => n22298, ZN => n22295);
   U22627 : OAI22_X1 port map( A1 => n20408, A2 => n24655, B1 => n21085, B2 => 
                           n24649, ZN => n22298);
   U22628 : AOI221_X1 port map( B1 => n24643, B2 => n17580, C1 => n24637, C2 =>
                           n24225, A => n22299, ZN => n22294);
   U22629 : OAI22_X1 port map( A1 => n20833, A2 => n24631, B1 => n21109, B2 => 
                           n24625, ZN => n22299);
   U22630 : AOI221_X1 port map( B1 => n24667, B2 => n24286, C1 => n24661, C2 =>
                           n24162, A => n22279, ZN => n22276);
   U22631 : OAI22_X1 port map( A1 => n20407, A2 => n24655, B1 => n21084, B2 => 
                           n24649, ZN => n22279);
   U22632 : AOI221_X1 port map( B1 => n24643, B2 => n17583, C1 => n24637, C2 =>
                           n24226, A => n22280, ZN => n22275);
   U22633 : OAI22_X1 port map( A1 => n20832, A2 => n24631, B1 => n21108, B2 => 
                           n24625, ZN => n22280);
   U22634 : AOI221_X1 port map( B1 => n24667, B2 => n24287, C1 => n24661, C2 =>
                           n24163, A => n22260, ZN => n22257);
   U22635 : OAI22_X1 port map( A1 => n20406, A2 => n24655, B1 => n21083, B2 => 
                           n24649, ZN => n22260);
   U22636 : AOI221_X1 port map( B1 => n24643, B2 => n17586, C1 => n24637, C2 =>
                           n24227, A => n22261, ZN => n22256);
   U22637 : OAI22_X1 port map( A1 => n20831, A2 => n24631, B1 => n21107, B2 => 
                           n24625, ZN => n22261);
   U22638 : AOI221_X1 port map( B1 => n24667, B2 => n24288, C1 => n24661, C2 =>
                           n24164, A => n22241, ZN => n22238);
   U22639 : OAI22_X1 port map( A1 => n20405, A2 => n24655, B1 => n21082, B2 => 
                           n24649, ZN => n22241);
   U22640 : AOI221_X1 port map( B1 => n24643, B2 => n17589, C1 => n24637, C2 =>
                           n24228, A => n22242, ZN => n22237);
   U22641 : OAI22_X1 port map( A1 => n20830, A2 => n24631, B1 => n21106, B2 => 
                           n24625, ZN => n22242);
   U22642 : AOI221_X1 port map( B1 => n24667, B2 => n24289, C1 => n24661, C2 =>
                           n24165, A => n22222, ZN => n22219);
   U22643 : OAI22_X1 port map( A1 => n20404, A2 => n24655, B1 => n21081, B2 => 
                           n24649, ZN => n22222);
   U22644 : AOI221_X1 port map( B1 => n24643, B2 => n17592, C1 => n24637, C2 =>
                           n24229, A => n22223, ZN => n22218);
   U22645 : OAI22_X1 port map( A1 => n20829, A2 => n24631, B1 => n21105, B2 => 
                           n24625, ZN => n22223);
   U22646 : AOI221_X1 port map( B1 => n24667, B2 => n24290, C1 => n24661, C2 =>
                           n24166, A => n22203, ZN => n22200);
   U22647 : OAI22_X1 port map( A1 => n20403, A2 => n24655, B1 => n21080, B2 => 
                           n24649, ZN => n22203);
   U22648 : AOI221_X1 port map( B1 => n24643, B2 => n17595, C1 => n24637, C2 =>
                           n24230, A => n22204, ZN => n22199);
   U22649 : OAI22_X1 port map( A1 => n20828, A2 => n24631, B1 => n21104, B2 => 
                           n24625, ZN => n22204);
   U22650 : AOI221_X1 port map( B1 => n24667, B2 => n24291, C1 => n24661, C2 =>
                           n24167, A => n22184, ZN => n22181);
   U22651 : OAI22_X1 port map( A1 => n20402, A2 => n24655, B1 => n21079, B2 => 
                           n24649, ZN => n22184);
   U22652 : AOI221_X1 port map( B1 => n24643, B2 => n17598, C1 => n24637, C2 =>
                           n24231, A => n22185, ZN => n22180);
   U22653 : OAI22_X1 port map( A1 => n20827, A2 => n24631, B1 => n21103, B2 => 
                           n24625, ZN => n22185);
   U22654 : AOI221_X1 port map( B1 => n24667, B2 => n24292, C1 => n24661, C2 =>
                           n24168, A => n22165, ZN => n22162);
   U22655 : OAI22_X1 port map( A1 => n20401, A2 => n24655, B1 => n21078, B2 => 
                           n24649, ZN => n22165);
   U22656 : AOI221_X1 port map( B1 => n24643, B2 => n17601, C1 => n24637, C2 =>
                           n24232, A => n22166, ZN => n22161);
   U22657 : OAI22_X1 port map( A1 => n20826, A2 => n24631, B1 => n21102, B2 => 
                           n24625, ZN => n22166);
   U22658 : AOI221_X1 port map( B1 => n24667, B2 => n24293, C1 => n24661, C2 =>
                           n24169, A => n22146, ZN => n22143);
   U22659 : OAI22_X1 port map( A1 => n20400, A2 => n24655, B1 => n21077, B2 => 
                           n24649, ZN => n22146);
   U22660 : AOI221_X1 port map( B1 => n24643, B2 => n17604, C1 => n24637, C2 =>
                           n24233, A => n22147, ZN => n22142);
   U22661 : OAI22_X1 port map( A1 => n20825, A2 => n24631, B1 => n21101, B2 => 
                           n24625, ZN => n22147);
   U22662 : AOI221_X1 port map( B1 => n24667, B2 => n24294, C1 => n24661, C2 =>
                           n24170, A => n22127, ZN => n22124);
   U22663 : OAI22_X1 port map( A1 => n20399, A2 => n24655, B1 => n21076, B2 => 
                           n24649, ZN => n22127);
   U22664 : AOI221_X1 port map( B1 => n24643, B2 => n17607, C1 => n24637, C2 =>
                           n24234, A => n22128, ZN => n22123);
   U22665 : OAI22_X1 port map( A1 => n20824, A2 => n24631, B1 => n21100, B2 => 
                           n24625, ZN => n22128);
   U22666 : AOI221_X1 port map( B1 => n24667, B2 => n24295, C1 => n24661, C2 =>
                           n24171, A => n22108, ZN => n22105);
   U22667 : OAI22_X1 port map( A1 => n20398, A2 => n24655, B1 => n21075, B2 => 
                           n24649, ZN => n22108);
   U22668 : AOI221_X1 port map( B1 => n24643, B2 => n17610, C1 => n24637, C2 =>
                           n24235, A => n22109, ZN => n22104);
   U22669 : OAI22_X1 port map( A1 => n20823, A2 => n24631, B1 => n21099, B2 => 
                           n24625, ZN => n22109);
   U22670 : AOI221_X1 port map( B1 => n24668, B2 => n24296, C1 => n24662, C2 =>
                           n24172, A => n22089, ZN => n22086);
   U22671 : OAI22_X1 port map( A1 => n20337, A2 => n24656, B1 => n20978, B2 => 
                           n24650, ZN => n22089);
   U22672 : AOI221_X1 port map( B1 => n24644, B2 => n17613, C1 => n24638, C2 =>
                           n24236, A => n22090, ZN => n22085);
   U22673 : OAI22_X1 port map( A1 => n20726, A2 => n24632, B1 => n21014, B2 => 
                           n24626, ZN => n22090);
   U22674 : AOI221_X1 port map( B1 => n24668, B2 => n24297, C1 => n24662, C2 =>
                           n24173, A => n22070, ZN => n22067);
   U22675 : OAI22_X1 port map( A1 => n20336, A2 => n24656, B1 => n20977, B2 => 
                           n24650, ZN => n22070);
   U22676 : AOI221_X1 port map( B1 => n24644, B2 => n17616, C1 => n24638, C2 =>
                           n24237, A => n22071, ZN => n22066);
   U22677 : OAI22_X1 port map( A1 => n20725, A2 => n24632, B1 => n21013, B2 => 
                           n24626, ZN => n22071);
   U22678 : AOI221_X1 port map( B1 => n24668, B2 => n24298, C1 => n24662, C2 =>
                           n24174, A => n22051, ZN => n22048);
   U22679 : OAI22_X1 port map( A1 => n20335, A2 => n24656, B1 => n20976, B2 => 
                           n24650, ZN => n22051);
   U22680 : AOI221_X1 port map( B1 => n24644, B2 => n17619, C1 => n24638, C2 =>
                           n24238, A => n22052, ZN => n22047);
   U22681 : OAI22_X1 port map( A1 => n20724, A2 => n24632, B1 => n21012, B2 => 
                           n24626, ZN => n22052);
   U22682 : AOI221_X1 port map( B1 => n24668, B2 => n24299, C1 => n24662, C2 =>
                           n24175, A => n22032, ZN => n22029);
   U22683 : OAI22_X1 port map( A1 => n20334, A2 => n24656, B1 => n20975, B2 => 
                           n24650, ZN => n22032);
   U22684 : AOI221_X1 port map( B1 => n24644, B2 => n17622, C1 => n24638, C2 =>
                           n24239, A => n22033, ZN => n22028);
   U22685 : OAI22_X1 port map( A1 => n20723, A2 => n24632, B1 => n21011, B2 => 
                           n24626, ZN => n22033);
   U22686 : AOI221_X1 port map( B1 => n24668, B2 => n24300, C1 => n24662, C2 =>
                           n24176, A => n22013, ZN => n22010);
   U22687 : OAI22_X1 port map( A1 => n20333, A2 => n24656, B1 => n20974, B2 => 
                           n24650, ZN => n22013);
   U22688 : AOI221_X1 port map( B1 => n24644, B2 => n17625, C1 => n24638, C2 =>
                           n24240, A => n22014, ZN => n22009);
   U22689 : OAI22_X1 port map( A1 => n20722, A2 => n24632, B1 => n21010, B2 => 
                           n24626, ZN => n22014);
   U22690 : AOI221_X1 port map( B1 => n24668, B2 => n24301, C1 => n24662, C2 =>
                           n24177, A => n21994, ZN => n21991);
   U22691 : OAI22_X1 port map( A1 => n20332, A2 => n24656, B1 => n20973, B2 => 
                           n24650, ZN => n21994);
   U22692 : AOI221_X1 port map( B1 => n24644, B2 => n17472, C1 => n24638, C2 =>
                           n24241, A => n21995, ZN => n21990);
   U22693 : OAI22_X1 port map( A1 => n20721, A2 => n24632, B1 => n21009, B2 => 
                           n24626, ZN => n21995);
   U22694 : AOI221_X1 port map( B1 => n24668, B2 => n24302, C1 => n24662, C2 =>
                           n24178, A => n21975, ZN => n21972);
   U22695 : OAI22_X1 port map( A1 => n20331, A2 => n24656, B1 => n20972, B2 => 
                           n24650, ZN => n21975);
   U22696 : AOI221_X1 port map( B1 => n24644, B2 => n17475, C1 => n24638, C2 =>
                           n24242, A => n21976, ZN => n21971);
   U22697 : OAI22_X1 port map( A1 => n20720, A2 => n24632, B1 => n21008, B2 => 
                           n24626, ZN => n21976);
   U22698 : AOI221_X1 port map( B1 => n24668, B2 => n24303, C1 => n24662, C2 =>
                           n24179, A => n21956, ZN => n21953);
   U22699 : OAI22_X1 port map( A1 => n20330, A2 => n24656, B1 => n20971, B2 => 
                           n24650, ZN => n21956);
   U22700 : AOI221_X1 port map( B1 => n24644, B2 => n17478, C1 => n24638, C2 =>
                           n24243, A => n21957, ZN => n21952);
   U22701 : OAI22_X1 port map( A1 => n20719, A2 => n24632, B1 => n21007, B2 => 
                           n24626, ZN => n21957);
   U22702 : AOI221_X1 port map( B1 => n24668, B2 => n24304, C1 => n24662, C2 =>
                           n24180, A => n21937, ZN => n21934);
   U22703 : OAI22_X1 port map( A1 => n20329, A2 => n24656, B1 => n20970, B2 => 
                           n24650, ZN => n21937);
   U22704 : AOI221_X1 port map( B1 => n24644, B2 => n17481, C1 => n24638, C2 =>
                           n24244, A => n21938, ZN => n21933);
   U22705 : OAI22_X1 port map( A1 => n20718, A2 => n24632, B1 => n21006, B2 => 
                           n24626, ZN => n21938);
   U22706 : AOI221_X1 port map( B1 => n24668, B2 => n24305, C1 => n24662, C2 =>
                           n24181, A => n21918, ZN => n21915);
   U22707 : OAI22_X1 port map( A1 => n20328, A2 => n24656, B1 => n20969, B2 => 
                           n24650, ZN => n21918);
   U22708 : AOI221_X1 port map( B1 => n24644, B2 => n17484, C1 => n24638, C2 =>
                           n24245, A => n21919, ZN => n21914);
   U22709 : OAI22_X1 port map( A1 => n20717, A2 => n24632, B1 => n21005, B2 => 
                           n24626, ZN => n21919);
   U22710 : AOI221_X1 port map( B1 => n24668, B2 => n24306, C1 => n24662, C2 =>
                           n24182, A => n21899, ZN => n21896);
   U22711 : OAI22_X1 port map( A1 => n20327, A2 => n24656, B1 => n20968, B2 => 
                           n24650, ZN => n21899);
   U22712 : AOI221_X1 port map( B1 => n24644, B2 => n17487, C1 => n24638, C2 =>
                           n24246, A => n21900, ZN => n21895);
   U22713 : OAI22_X1 port map( A1 => n20716, A2 => n24632, B1 => n21004, B2 => 
                           n24626, ZN => n21900);
   U22714 : AOI221_X1 port map( B1 => n24668, B2 => n24307, C1 => n24662, C2 =>
                           n24183, A => n21880, ZN => n21877);
   U22715 : OAI22_X1 port map( A1 => n20326, A2 => n24656, B1 => n20967, B2 => 
                           n24650, ZN => n21880);
   U22716 : AOI221_X1 port map( B1 => n24644, B2 => n17490, C1 => n24638, C2 =>
                           n24247, A => n21881, ZN => n21876);
   U22717 : OAI22_X1 port map( A1 => n20715, A2 => n24632, B1 => n21003, B2 => 
                           n24626, ZN => n21881);
   U22718 : AOI221_X1 port map( B1 => n24669, B2 => n24308, C1 => n24663, C2 =>
                           n24184, A => n21861, ZN => n21858);
   U22719 : OAI22_X1 port map( A1 => n20325, A2 => n24657, B1 => n20966, B2 => 
                           n24651, ZN => n21861);
   U22720 : AOI221_X1 port map( B1 => n24645, B2 => n17493, C1 => n24639, C2 =>
                           n24248, A => n21862, ZN => n21857);
   U22721 : OAI22_X1 port map( A1 => n20714, A2 => n24633, B1 => n21002, B2 => 
                           n24627, ZN => n21862);
   U22722 : AOI221_X1 port map( B1 => n24669, B2 => n24309, C1 => n24663, C2 =>
                           n24185, A => n21842, ZN => n21839);
   U22723 : OAI22_X1 port map( A1 => n20324, A2 => n24657, B1 => n20965, B2 => 
                           n24651, ZN => n21842);
   U22724 : AOI221_X1 port map( B1 => n24645, B2 => n17496, C1 => n24639, C2 =>
                           n24249, A => n21843, ZN => n21838);
   U22725 : OAI22_X1 port map( A1 => n20713, A2 => n24633, B1 => n21001, B2 => 
                           n24627, ZN => n21843);
   U22726 : AOI221_X1 port map( B1 => n24669, B2 => n24310, C1 => n24663, C2 =>
                           n24186, A => n21823, ZN => n21820);
   U22727 : OAI22_X1 port map( A1 => n20323, A2 => n24657, B1 => n20964, B2 => 
                           n24651, ZN => n21823);
   U22728 : AOI221_X1 port map( B1 => n24645, B2 => n17499, C1 => n24639, C2 =>
                           n24250, A => n21824, ZN => n21819);
   U22729 : OAI22_X1 port map( A1 => n20712, A2 => n24633, B1 => n21000, B2 => 
                           n24627, ZN => n21824);
   U22730 : AOI221_X1 port map( B1 => n24669, B2 => n24311, C1 => n24663, C2 =>
                           n24187, A => n21804, ZN => n21801);
   U22731 : OAI22_X1 port map( A1 => n20322, A2 => n24657, B1 => n20963, B2 => 
                           n24651, ZN => n21804);
   U22732 : AOI221_X1 port map( B1 => n24645, B2 => n17502, C1 => n24639, C2 =>
                           n24251, A => n21805, ZN => n21800);
   U22733 : OAI22_X1 port map( A1 => n20711, A2 => n24633, B1 => n20999, B2 => 
                           n24627, ZN => n21805);
   U22734 : AOI221_X1 port map( B1 => n24669, B2 => n24312, C1 => n24663, C2 =>
                           n24188, A => n21785, ZN => n21782);
   U22735 : OAI22_X1 port map( A1 => n20321, A2 => n24657, B1 => n20962, B2 => 
                           n24651, ZN => n21785);
   U22736 : AOI221_X1 port map( B1 => n24645, B2 => n17505, C1 => n24639, C2 =>
                           n24252, A => n21786, ZN => n21781);
   U22737 : OAI22_X1 port map( A1 => n20710, A2 => n24633, B1 => n20998, B2 => 
                           n24627, ZN => n21786);
   U22738 : AOI221_X1 port map( B1 => n24669, B2 => n24313, C1 => n24663, C2 =>
                           n24189, A => n21766, ZN => n21763);
   U22739 : OAI22_X1 port map( A1 => n20320, A2 => n24657, B1 => n20961, B2 => 
                           n24651, ZN => n21766);
   U22740 : AOI221_X1 port map( B1 => n24645, B2 => n17508, C1 => n24639, C2 =>
                           n24253, A => n21767, ZN => n21762);
   U22741 : OAI22_X1 port map( A1 => n20709, A2 => n24633, B1 => n20997, B2 => 
                           n24627, ZN => n21767);
   U22742 : AOI221_X1 port map( B1 => n24669, B2 => n24314, C1 => n24663, C2 =>
                           n24190, A => n21747, ZN => n21744);
   U22743 : OAI22_X1 port map( A1 => n20319, A2 => n24657, B1 => n20960, B2 => 
                           n24651, ZN => n21747);
   U22744 : AOI221_X1 port map( B1 => n24645, B2 => n17511, C1 => n24639, C2 =>
                           n24254, A => n21748, ZN => n21743);
   U22745 : OAI22_X1 port map( A1 => n20708, A2 => n24633, B1 => n20996, B2 => 
                           n24627, ZN => n21748);
   U22746 : AOI221_X1 port map( B1 => n24669, B2 => n24315, C1 => n24663, C2 =>
                           n24191, A => n21728, ZN => n21725);
   U22747 : OAI22_X1 port map( A1 => n20318, A2 => n24657, B1 => n20959, B2 => 
                           n24651, ZN => n21728);
   U22748 : AOI221_X1 port map( B1 => n24645, B2 => n17514, C1 => n24639, C2 =>
                           n24255, A => n21729, ZN => n21724);
   U22749 : OAI22_X1 port map( A1 => n20707, A2 => n24633, B1 => n20995, B2 => 
                           n24627, ZN => n21729);
   U22750 : AOI221_X1 port map( B1 => n24669, B2 => n24316, C1 => n24663, C2 =>
                           n24192, A => n21709, ZN => n21706);
   U22751 : OAI22_X1 port map( A1 => n20317, A2 => n24657, B1 => n20958, B2 => 
                           n24651, ZN => n21709);
   U22752 : AOI221_X1 port map( B1 => n24645, B2 => n17517, C1 => n24639, C2 =>
                           n24256, A => n21710, ZN => n21705);
   U22753 : OAI22_X1 port map( A1 => n20706, A2 => n24633, B1 => n20994, B2 => 
                           n24627, ZN => n21710);
   U22754 : AOI221_X1 port map( B1 => n24669, B2 => n24317, C1 => n24663, C2 =>
                           n24193, A => n21690, ZN => n21687);
   U22755 : OAI22_X1 port map( A1 => n20316, A2 => n24657, B1 => n20957, B2 => 
                           n24651, ZN => n21690);
   U22756 : AOI221_X1 port map( B1 => n24645, B2 => n17520, C1 => n24639, C2 =>
                           n24257, A => n21691, ZN => n21686);
   U22757 : OAI22_X1 port map( A1 => n20705, A2 => n24633, B1 => n20993, B2 => 
                           n24627, ZN => n21691);
   U22758 : AOI221_X1 port map( B1 => n24669, B2 => n24318, C1 => n24663, C2 =>
                           n24194, A => n21671, ZN => n21668);
   U22759 : OAI22_X1 port map( A1 => n20315, A2 => n24657, B1 => n20956, B2 => 
                           n24651, ZN => n21671);
   U22760 : AOI221_X1 port map( B1 => n24645, B2 => n17523, C1 => n24639, C2 =>
                           n24258, A => n21672, ZN => n21667);
   U22761 : OAI22_X1 port map( A1 => n20704, A2 => n24633, B1 => n20992, B2 => 
                           n24627, ZN => n21672);
   U22762 : AOI221_X1 port map( B1 => n24669, B2 => n24319, C1 => n24663, C2 =>
                           n24195, A => n21652, ZN => n21649);
   U22763 : OAI22_X1 port map( A1 => n20314, A2 => n24657, B1 => n20955, B2 => 
                           n24651, ZN => n21652);
   U22764 : AOI221_X1 port map( B1 => n24645, B2 => n17526, C1 => n24639, C2 =>
                           n24259, A => n21653, ZN => n21648);
   U22765 : OAI22_X1 port map( A1 => n20703, A2 => n24633, B1 => n20991, B2 => 
                           n24627, ZN => n21653);
   U22766 : AOI221_X1 port map( B1 => n24670, B2 => n24320, C1 => n24664, C2 =>
                           n24196, A => n21633, ZN => n21630);
   U22767 : OAI22_X1 port map( A1 => n20313, A2 => n24658, B1 => n20954, B2 => 
                           n24652, ZN => n21633);
   U22768 : AOI221_X1 port map( B1 => n24646, B2 => n17529, C1 => n24640, C2 =>
                           n24260, A => n21634, ZN => n21629);
   U22769 : OAI22_X1 port map( A1 => n20702, A2 => n24634, B1 => n20990, B2 => 
                           n24628, ZN => n21634);
   U22770 : AOI221_X1 port map( B1 => n24670, B2 => n24321, C1 => n24664, C2 =>
                           n24197, A => n21614, ZN => n21611);
   U22771 : OAI22_X1 port map( A1 => n20312, A2 => n24658, B1 => n20953, B2 => 
                           n24652, ZN => n21614);
   U22772 : AOI221_X1 port map( B1 => n24646, B2 => n17532, C1 => n24640, C2 =>
                           n24261, A => n21615, ZN => n21610);
   U22773 : OAI22_X1 port map( A1 => n20701, A2 => n24634, B1 => n20989, B2 => 
                           n24628, ZN => n21615);
   U22774 : AOI221_X1 port map( B1 => n24670, B2 => n24322, C1 => n24664, C2 =>
                           n24198, A => n21595, ZN => n21592);
   U22775 : OAI22_X1 port map( A1 => n20311, A2 => n24658, B1 => n20952, B2 => 
                           n24652, ZN => n21595);
   U22776 : AOI221_X1 port map( B1 => n24646, B2 => n17535, C1 => n24640, C2 =>
                           n24262, A => n21596, ZN => n21591);
   U22777 : OAI22_X1 port map( A1 => n20700, A2 => n24634, B1 => n20988, B2 => 
                           n24628, ZN => n21596);
   U22778 : AOI221_X1 port map( B1 => n24670, B2 => n24323, C1 => n24664, C2 =>
                           n24199, A => n21576, ZN => n21573);
   U22779 : OAI22_X1 port map( A1 => n20310, A2 => n24658, B1 => n20951, B2 => 
                           n24652, ZN => n21576);
   U22780 : AOI221_X1 port map( B1 => n24646, B2 => n17538, C1 => n24640, C2 =>
                           n24263, A => n21577, ZN => n21572);
   U22781 : OAI22_X1 port map( A1 => n20699, A2 => n24634, B1 => n20987, B2 => 
                           n24628, ZN => n21577);
   U22782 : AOI221_X1 port map( B1 => n24670, B2 => n24324, C1 => n24664, C2 =>
                           n24200, A => n21557, ZN => n21554);
   U22783 : OAI22_X1 port map( A1 => n20309, A2 => n24658, B1 => n20950, B2 => 
                           n24652, ZN => n21557);
   U22784 : AOI221_X1 port map( B1 => n24646, B2 => n17628, C1 => n24640, C2 =>
                           n24264, A => n21558, ZN => n21553);
   U22785 : OAI22_X1 port map( A1 => n20698, A2 => n24634, B1 => n20986, B2 => 
                           n24628, ZN => n21558);
   U22786 : AOI221_X1 port map( B1 => n24670, B2 => n24325, C1 => n24664, C2 =>
                           n24201, A => n21538, ZN => n21535);
   U22787 : OAI22_X1 port map( A1 => n20308, A2 => n24658, B1 => n20949, B2 => 
                           n24652, ZN => n21538);
   U22788 : AOI221_X1 port map( B1 => n24646, B2 => n17631, C1 => n24640, C2 =>
                           n24265, A => n21539, ZN => n21534);
   U22789 : OAI22_X1 port map( A1 => n20697, A2 => n24634, B1 => n20985, B2 => 
                           n24628, ZN => n21539);
   U22790 : AOI221_X1 port map( B1 => n24670, B2 => n24326, C1 => n24664, C2 =>
                           n24202, A => n21519, ZN => n21516);
   U22791 : OAI22_X1 port map( A1 => n20307, A2 => n24658, B1 => n20948, B2 => 
                           n24652, ZN => n21519);
   U22792 : AOI221_X1 port map( B1 => n24646, B2 => n17634, C1 => n24640, C2 =>
                           n24266, A => n21520, ZN => n21515);
   U22793 : OAI22_X1 port map( A1 => n20696, A2 => n24634, B1 => n20984, B2 => 
                           n24628, ZN => n21520);
   U22794 : AOI221_X1 port map( B1 => n24670, B2 => n24327, C1 => n24664, C2 =>
                           n24203, A => n21500, ZN => n21497);
   U22795 : OAI22_X1 port map( A1 => n20306, A2 => n24658, B1 => n20947, B2 => 
                           n24652, ZN => n21500);
   U22796 : AOI221_X1 port map( B1 => n24646, B2 => n17637, C1 => n24640, C2 =>
                           n24267, A => n21501, ZN => n21496);
   U22797 : OAI22_X1 port map( A1 => n20695, A2 => n24634, B1 => n20983, B2 => 
                           n24628, ZN => n21501);
   U22798 : AOI221_X1 port map( B1 => n24670, B2 => n24328, C1 => n24664, C2 =>
                           n24204, A => n21481, ZN => n21478);
   U22799 : OAI22_X1 port map( A1 => n20305, A2 => n24658, B1 => n20946, B2 => 
                           n24652, ZN => n21481);
   U22800 : AOI221_X1 port map( B1 => n24646, B2 => n17640, C1 => n24640, C2 =>
                           n24268, A => n21482, ZN => n21477);
   U22801 : OAI22_X1 port map( A1 => n20694, A2 => n24634, B1 => n20982, B2 => 
                           n24628, ZN => n21482);
   U22802 : AOI221_X1 port map( B1 => n24670, B2 => n24329, C1 => n24664, C2 =>
                           n24205, A => n21462, ZN => n21459);
   U22803 : OAI22_X1 port map( A1 => n20304, A2 => n24658, B1 => n20945, B2 => 
                           n24652, ZN => n21462);
   U22804 : AOI221_X1 port map( B1 => n24646, B2 => n17643, C1 => n24640, C2 =>
                           n24269, A => n21463, ZN => n21458);
   U22805 : OAI22_X1 port map( A1 => n20693, A2 => n24634, B1 => n20981, B2 => 
                           n24628, ZN => n21463);
   U22806 : AOI221_X1 port map( B1 => n24670, B2 => n24330, C1 => n24664, C2 =>
                           n24206, A => n21443, ZN => n21440);
   U22807 : OAI22_X1 port map( A1 => n20303, A2 => n24658, B1 => n20944, B2 => 
                           n24652, ZN => n21443);
   U22808 : AOI221_X1 port map( B1 => n24646, B2 => n17646, C1 => n24640, C2 =>
                           n24270, A => n21444, ZN => n21439);
   U22809 : OAI22_X1 port map( A1 => n20692, A2 => n24634, B1 => n20980, B2 => 
                           n24628, ZN => n21444);
   U22810 : AOI221_X1 port map( B1 => n24670, B2 => n24331, C1 => n24664, C2 =>
                           n24207, A => n21424, ZN => n21421);
   U22811 : OAI22_X1 port map( A1 => n20302, A2 => n24658, B1 => n20943, B2 => 
                           n24652, ZN => n21424);
   U22812 : AOI221_X1 port map( B1 => n24646, B2 => n17649, C1 => n24640, C2 =>
                           n24271, A => n21425, ZN => n21420);
   U22813 : OAI22_X1 port map( A1 => n20691, A2 => n24634, B1 => n20979, B2 => 
                           n24628, ZN => n21425);
   U22814 : OAI22_X1 port map( A1 => n24824, A2 => n20213, B1 => n24818, B2 => 
                           n25467, ZN => n5100);
   U22815 : OAI22_X1 port map( A1 => n24824, A2 => n20212, B1 => n24818, B2 => 
                           n25470, ZN => n5101);
   U22816 : OAI22_X1 port map( A1 => n24824, A2 => n20211, B1 => n24818, B2 => 
                           n25473, ZN => n5102);
   U22817 : OAI22_X1 port map( A1 => n24824, A2 => n20210, B1 => n24818, B2 => 
                           n25476, ZN => n5103);
   U22818 : OAI22_X1 port map( A1 => n24823, A2 => n20209, B1 => n24818, B2 => 
                           n25479, ZN => n5104);
   U22819 : OAI22_X1 port map( A1 => n24823, A2 => n20208, B1 => n24818, B2 => 
                           n25482, ZN => n5105);
   U22820 : OAI22_X1 port map( A1 => n24823, A2 => n20207, B1 => n24818, B2 => 
                           n25485, ZN => n5106);
   U22821 : OAI22_X1 port map( A1 => n24823, A2 => n20206, B1 => n24818, B2 => 
                           n25488, ZN => n5107);
   U22822 : OAI22_X1 port map( A1 => n24823, A2 => n20205, B1 => n24818, B2 => 
                           n25491, ZN => n5108);
   U22823 : OAI22_X1 port map( A1 => n24822, A2 => n20204, B1 => n24818, B2 => 
                           n25494, ZN => n5109);
   U22824 : OAI22_X1 port map( A1 => n24822, A2 => n20203, B1 => n24818, B2 => 
                           n25497, ZN => n5110);
   U22825 : OAI22_X1 port map( A1 => n24822, A2 => n20202, B1 => n24818, B2 => 
                           n25500, ZN => n5111);
   U22826 : OAI22_X1 port map( A1 => n24822, A2 => n20201, B1 => n24817, B2 => 
                           n25503, ZN => n5112);
   U22827 : OAI22_X1 port map( A1 => n24822, A2 => n20200, B1 => n24817, B2 => 
                           n25506, ZN => n5113);
   U22828 : OAI22_X1 port map( A1 => n24821, A2 => n20199, B1 => n24817, B2 => 
                           n25509, ZN => n5114);
   U22829 : OAI22_X1 port map( A1 => n24821, A2 => n20198, B1 => n24817, B2 => 
                           n25512, ZN => n5115);
   U22830 : OAI22_X1 port map( A1 => n24821, A2 => n20197, B1 => n24817, B2 => 
                           n25515, ZN => n5116);
   U22831 : OAI22_X1 port map( A1 => n24821, A2 => n20196, B1 => n24817, B2 => 
                           n25518, ZN => n5117);
   U22832 : OAI22_X1 port map( A1 => n24821, A2 => n20195, B1 => n24817, B2 => 
                           n25521, ZN => n5118);
   U22833 : OAI22_X1 port map( A1 => n24820, A2 => n20194, B1 => n24817, B2 => 
                           n25524, ZN => n5119);
   U22834 : OAI22_X1 port map( A1 => n24820, A2 => n20193, B1 => n24817, B2 => 
                           n25527, ZN => n5120);
   U22835 : OAI22_X1 port map( A1 => n24820, A2 => n20192, B1 => n24817, B2 => 
                           n25530, ZN => n5121);
   U22836 : OAI22_X1 port map( A1 => n24820, A2 => n20191, B1 => n24817, B2 => 
                           n25533, ZN => n5122);
   U22837 : OAI22_X1 port map( A1 => n24820, A2 => n20190, B1 => n24817, B2 => 
                           n25553, ZN => n5123);
   U22838 : AOI22_X1 port map( A1 => n24561, A2 => n8053, B1 => n24555, B2 => 
                           n8245, ZN => n23017);
   U22839 : AOI22_X1 port map( A1 => n24537, A2 => n8309, B1 => n24531, B2 => 
                           n23936, ZN => n23018);
   U22840 : AOI22_X1 port map( A1 => n24561, A2 => n8052, B1 => n24555, B2 => 
                           n8244, ZN => n22999);
   U22841 : AOI22_X1 port map( A1 => n24537, A2 => n8308, B1 => n24531, B2 => 
                           n23938, ZN => n23000);
   U22842 : AOI22_X1 port map( A1 => n24561, A2 => n8051, B1 => n24555, B2 => 
                           n8243, ZN => n22981);
   U22843 : AOI22_X1 port map( A1 => n24537, A2 => n8307, B1 => n24531, B2 => 
                           n23940, ZN => n22982);
   U22844 : AOI22_X1 port map( A1 => n24561, A2 => n8050, B1 => n24555, B2 => 
                           n8242, ZN => n22963);
   U22845 : AOI22_X1 port map( A1 => n24537, A2 => n8306, B1 => n24531, B2 => 
                           n23942, ZN => n22964);
   U22846 : AOI22_X1 port map( A1 => n24561, A2 => n8049, B1 => n24555, B2 => 
                           n8241, ZN => n22945);
   U22847 : AOI22_X1 port map( A1 => n24537, A2 => n8305, B1 => n24531, B2 => 
                           n23944, ZN => n22946);
   U22848 : AOI22_X1 port map( A1 => n24561, A2 => n8048, B1 => n24555, B2 => 
                           n8240, ZN => n22927);
   U22849 : AOI22_X1 port map( A1 => n24537, A2 => n8304, B1 => n24531, B2 => 
                           n23946, ZN => n22928);
   U22850 : AOI22_X1 port map( A1 => n24561, A2 => n8047, B1 => n24555, B2 => 
                           n8239, ZN => n22909);
   U22851 : AOI22_X1 port map( A1 => n24537, A2 => n8303, B1 => n24531, B2 => 
                           n23948, ZN => n22910);
   U22852 : AOI22_X1 port map( A1 => n24561, A2 => n8046, B1 => n24555, B2 => 
                           n8238, ZN => n22891);
   U22853 : AOI22_X1 port map( A1 => n24537, A2 => n8302, B1 => n24531, B2 => 
                           n23950, ZN => n22892);
   U22854 : AOI22_X1 port map( A1 => n24562, A2 => n8045, B1 => n24556, B2 => 
                           n8237, ZN => n22873);
   U22855 : AOI22_X1 port map( A1 => n24538, A2 => n8301, B1 => n24532, B2 => 
                           n23952, ZN => n22874);
   U22856 : AOI22_X1 port map( A1 => n24562, A2 => n8044, B1 => n24556, B2 => 
                           n8236, ZN => n22855);
   U22857 : AOI22_X1 port map( A1 => n24538, A2 => n8300, B1 => n24532, B2 => 
                           n23953, ZN => n22856);
   U22858 : AOI22_X1 port map( A1 => n24562, A2 => n8043, B1 => n24556, B2 => 
                           n8235, ZN => n22837);
   U22859 : AOI22_X1 port map( A1 => n24538, A2 => n8299, B1 => n24532, B2 => 
                           n23954, ZN => n22838);
   U22860 : AOI22_X1 port map( A1 => n24562, A2 => n8042, B1 => n24556, B2 => 
                           n8234, ZN => n22819);
   U22861 : AOI22_X1 port map( A1 => n24538, A2 => n8298, B1 => n24532, B2 => 
                           n23955, ZN => n22820);
   U22862 : AOI22_X1 port map( A1 => n24562, A2 => n8041, B1 => n24556, B2 => 
                           n8233, ZN => n22801);
   U22863 : AOI22_X1 port map( A1 => n24538, A2 => n8297, B1 => n24532, B2 => 
                           n23956, ZN => n22802);
   U22864 : AOI22_X1 port map( A1 => n24562, A2 => n8040, B1 => n24556, B2 => 
                           n8232, ZN => n22783);
   U22865 : AOI22_X1 port map( A1 => n24538, A2 => n8296, B1 => n24532, B2 => 
                           n23957, ZN => n22784);
   U22866 : AOI22_X1 port map( A1 => n24562, A2 => n8039, B1 => n24556, B2 => 
                           n8231, ZN => n22765);
   U22867 : AOI22_X1 port map( A1 => n24538, A2 => n8295, B1 => n24532, B2 => 
                           n23958, ZN => n22766);
   U22868 : AOI22_X1 port map( A1 => n24562, A2 => n8038, B1 => n24556, B2 => 
                           n8230, ZN => n22747);
   U22869 : AOI22_X1 port map( A1 => n24538, A2 => n8294, B1 => n24532, B2 => 
                           n23959, ZN => n22748);
   U22870 : AOI22_X1 port map( A1 => n24562, A2 => n8037, B1 => n24556, B2 => 
                           n8229, ZN => n22729);
   U22871 : AOI22_X1 port map( A1 => n24538, A2 => n8293, B1 => n24532, B2 => 
                           n23960, ZN => n22730);
   U22872 : AOI22_X1 port map( A1 => n24562, A2 => n8036, B1 => n24556, B2 => 
                           n8228, ZN => n22711);
   U22873 : AOI22_X1 port map( A1 => n24538, A2 => n8292, B1 => n24532, B2 => 
                           n23961, ZN => n22712);
   U22874 : AOI22_X1 port map( A1 => n24562, A2 => n8035, B1 => n24556, B2 => 
                           n8227, ZN => n22693);
   U22875 : AOI22_X1 port map( A1 => n24538, A2 => n8291, B1 => n24532, B2 => 
                           n23962, ZN => n22694);
   U22876 : AOI22_X1 port map( A1 => n24562, A2 => n8034, B1 => n24556, B2 => 
                           n8226, ZN => n22675);
   U22877 : AOI22_X1 port map( A1 => n24538, A2 => n8290, B1 => n24532, B2 => 
                           n23963, ZN => n22676);
   U22878 : AOI22_X1 port map( A1 => n24563, A2 => n8033, B1 => n24557, B2 => 
                           n8225, ZN => n22657);
   U22879 : AOI22_X1 port map( A1 => n24539, A2 => n8289, B1 => n24533, B2 => 
                           n23964, ZN => n22658);
   U22880 : AOI22_X1 port map( A1 => n24563, A2 => n8032, B1 => n24557, B2 => 
                           n8224, ZN => n22639);
   U22881 : AOI22_X1 port map( A1 => n24539, A2 => n8288, B1 => n24533, B2 => 
                           n23965, ZN => n22640);
   U22882 : AOI22_X1 port map( A1 => n24563, A2 => n8031, B1 => n24557, B2 => 
                           n8223, ZN => n22621);
   U22883 : AOI22_X1 port map( A1 => n24539, A2 => n8287, B1 => n24533, B2 => 
                           n23966, ZN => n22622);
   U22884 : AOI22_X1 port map( A1 => n24563, A2 => n8030, B1 => n24557, B2 => 
                           n8222, ZN => n22575);
   U22885 : AOI22_X1 port map( A1 => n24539, A2 => n8286, B1 => n24533, B2 => 
                           n23967, ZN => n22580);
   U22886 : AOI22_X1 port map( A1 => n24558, A2 => n8093, B1 => n24552, B2 => 
                           n8285, ZN => n23743);
   U22887 : AOI22_X1 port map( A1 => n24534, A2 => n8349, B1 => n24528, B2 => 
                           n23856, ZN => n23746);
   U22888 : AOI22_X1 port map( A1 => n24558, A2 => n8092, B1 => n24552, B2 => 
                           n8284, ZN => n23719);
   U22889 : AOI22_X1 port map( A1 => n24534, A2 => n8348, B1 => n24528, B2 => 
                           n23858, ZN => n23720);
   U22890 : AOI22_X1 port map( A1 => n24558, A2 => n8091, B1 => n24552, B2 => 
                           n8283, ZN => n23701);
   U22891 : AOI22_X1 port map( A1 => n24534, A2 => n8347, B1 => n24528, B2 => 
                           n23860, ZN => n23702);
   U22892 : AOI22_X1 port map( A1 => n24558, A2 => n8090, B1 => n24552, B2 => 
                           n8282, ZN => n23683);
   U22893 : AOI22_X1 port map( A1 => n24534, A2 => n8346, B1 => n24528, B2 => 
                           n23862, ZN => n23684);
   U22894 : AOI22_X1 port map( A1 => n24558, A2 => n8089, B1 => n24552, B2 => 
                           n8281, ZN => n23665);
   U22895 : AOI22_X1 port map( A1 => n24534, A2 => n8345, B1 => n24528, B2 => 
                           n23864, ZN => n23666);
   U22896 : AOI22_X1 port map( A1 => n24558, A2 => n8088, B1 => n24552, B2 => 
                           n8280, ZN => n23647);
   U22897 : AOI22_X1 port map( A1 => n24534, A2 => n8344, B1 => n24528, B2 => 
                           n23866, ZN => n23648);
   U22898 : AOI22_X1 port map( A1 => n24558, A2 => n8087, B1 => n24552, B2 => 
                           n8279, ZN => n23629);
   U22899 : AOI22_X1 port map( A1 => n24534, A2 => n8343, B1 => n24528, B2 => 
                           n23868, ZN => n23630);
   U22900 : AOI22_X1 port map( A1 => n24558, A2 => n8086, B1 => n24552, B2 => 
                           n8278, ZN => n23611);
   U22901 : AOI22_X1 port map( A1 => n24534, A2 => n8342, B1 => n24528, B2 => 
                           n23870, ZN => n23612);
   U22902 : AOI22_X1 port map( A1 => n24558, A2 => n8085, B1 => n24552, B2 => 
                           n8277, ZN => n23593);
   U22903 : AOI22_X1 port map( A1 => n24534, A2 => n8341, B1 => n24528, B2 => 
                           n23872, ZN => n23594);
   U22904 : AOI22_X1 port map( A1 => n24558, A2 => n8084, B1 => n24552, B2 => 
                           n8276, ZN => n23575);
   U22905 : AOI22_X1 port map( A1 => n24534, A2 => n8340, B1 => n24528, B2 => 
                           n23874, ZN => n23576);
   U22906 : AOI22_X1 port map( A1 => n24558, A2 => n8083, B1 => n24552, B2 => 
                           n8275, ZN => n23557);
   U22907 : AOI22_X1 port map( A1 => n24534, A2 => n8339, B1 => n24528, B2 => 
                           n23876, ZN => n23558);
   U22908 : AOI22_X1 port map( A1 => n24558, A2 => n8082, B1 => n24552, B2 => 
                           n8274, ZN => n23539);
   U22909 : AOI22_X1 port map( A1 => n24534, A2 => n8338, B1 => n24528, B2 => 
                           n23878, ZN => n23540);
   U22910 : AOI22_X1 port map( A1 => n24559, A2 => n8081, B1 => n24553, B2 => 
                           n8273, ZN => n23521);
   U22911 : AOI22_X1 port map( A1 => n24535, A2 => n8337, B1 => n24529, B2 => 
                           n23880, ZN => n23522);
   U22912 : AOI22_X1 port map( A1 => n24559, A2 => n8080, B1 => n24553, B2 => 
                           n8272, ZN => n23503);
   U22913 : AOI22_X1 port map( A1 => n24535, A2 => n8336, B1 => n24529, B2 => 
                           n23882, ZN => n23504);
   U22914 : AOI22_X1 port map( A1 => n24559, A2 => n8079, B1 => n24553, B2 => 
                           n8271, ZN => n23485);
   U22915 : AOI22_X1 port map( A1 => n24535, A2 => n8335, B1 => n24529, B2 => 
                           n23884, ZN => n23486);
   U22916 : AOI22_X1 port map( A1 => n24559, A2 => n8078, B1 => n24553, B2 => 
                           n8270, ZN => n23467);
   U22917 : AOI22_X1 port map( A1 => n24535, A2 => n8334, B1 => n24529, B2 => 
                           n23886, ZN => n23468);
   U22918 : AOI22_X1 port map( A1 => n24559, A2 => n8077, B1 => n24553, B2 => 
                           n8269, ZN => n23449);
   U22919 : AOI22_X1 port map( A1 => n24535, A2 => n8333, B1 => n24529, B2 => 
                           n23888, ZN => n23450);
   U22920 : AOI22_X1 port map( A1 => n24559, A2 => n8076, B1 => n24553, B2 => 
                           n8268, ZN => n23431);
   U22921 : AOI22_X1 port map( A1 => n24535, A2 => n8332, B1 => n24529, B2 => 
                           n23890, ZN => n23432);
   U22922 : AOI22_X1 port map( A1 => n24559, A2 => n8075, B1 => n24553, B2 => 
                           n8267, ZN => n23413);
   U22923 : AOI22_X1 port map( A1 => n24535, A2 => n8331, B1 => n24529, B2 => 
                           n23892, ZN => n23414);
   U22924 : AOI22_X1 port map( A1 => n24559, A2 => n8074, B1 => n24553, B2 => 
                           n8266, ZN => n23395);
   U22925 : AOI22_X1 port map( A1 => n24535, A2 => n8330, B1 => n24529, B2 => 
                           n23894, ZN => n23396);
   U22926 : AOI22_X1 port map( A1 => n24559, A2 => n8073, B1 => n24553, B2 => 
                           n8265, ZN => n23377);
   U22927 : AOI22_X1 port map( A1 => n24535, A2 => n8329, B1 => n24529, B2 => 
                           n23896, ZN => n23378);
   U22928 : AOI22_X1 port map( A1 => n24559, A2 => n8072, B1 => n24553, B2 => 
                           n8264, ZN => n23359);
   U22929 : AOI22_X1 port map( A1 => n24535, A2 => n8328, B1 => n24529, B2 => 
                           n23898, ZN => n23360);
   U22930 : AOI22_X1 port map( A1 => n24559, A2 => n8071, B1 => n24553, B2 => 
                           n8263, ZN => n23341);
   U22931 : AOI22_X1 port map( A1 => n24535, A2 => n8327, B1 => n24529, B2 => 
                           n23900, ZN => n23342);
   U22932 : AOI22_X1 port map( A1 => n24559, A2 => n8070, B1 => n24553, B2 => 
                           n8262, ZN => n23323);
   U22933 : AOI22_X1 port map( A1 => n24535, A2 => n8326, B1 => n24529, B2 => 
                           n23902, ZN => n23324);
   U22934 : AOI22_X1 port map( A1 => n24560, A2 => n8069, B1 => n24554, B2 => 
                           n8261, ZN => n23305);
   U22935 : AOI22_X1 port map( A1 => n24536, A2 => n8325, B1 => n24530, B2 => 
                           n23904, ZN => n23306);
   U22936 : AOI22_X1 port map( A1 => n24560, A2 => n8068, B1 => n24554, B2 => 
                           n8260, ZN => n23287);
   U22937 : AOI22_X1 port map( A1 => n24536, A2 => n8324, B1 => n24530, B2 => 
                           n23906, ZN => n23288);
   U22938 : AOI22_X1 port map( A1 => n24560, A2 => n8067, B1 => n24554, B2 => 
                           n8259, ZN => n23269);
   U22939 : AOI22_X1 port map( A1 => n24536, A2 => n8323, B1 => n24530, B2 => 
                           n23908, ZN => n23270);
   U22940 : AOI22_X1 port map( A1 => n24560, A2 => n8066, B1 => n24554, B2 => 
                           n8258, ZN => n23251);
   U22941 : AOI22_X1 port map( A1 => n24536, A2 => n8322, B1 => n24530, B2 => 
                           n23910, ZN => n23252);
   U22942 : AOI22_X1 port map( A1 => n24560, A2 => n8065, B1 => n24554, B2 => 
                           n8257, ZN => n23233);
   U22943 : AOI22_X1 port map( A1 => n24536, A2 => n8321, B1 => n24530, B2 => 
                           n23912, ZN => n23234);
   U22944 : AOI22_X1 port map( A1 => n24560, A2 => n8064, B1 => n24554, B2 => 
                           n8256, ZN => n23215);
   U22945 : AOI22_X1 port map( A1 => n24536, A2 => n8320, B1 => n24530, B2 => 
                           n23914, ZN => n23216);
   U22946 : AOI22_X1 port map( A1 => n24560, A2 => n8063, B1 => n24554, B2 => 
                           n8255, ZN => n23197);
   U22947 : AOI22_X1 port map( A1 => n24536, A2 => n8319, B1 => n24530, B2 => 
                           n23916, ZN => n23198);
   U22948 : AOI22_X1 port map( A1 => n24560, A2 => n8062, B1 => n24554, B2 => 
                           n8254, ZN => n23179);
   U22949 : AOI22_X1 port map( A1 => n24536, A2 => n8318, B1 => n24530, B2 => 
                           n23918, ZN => n23180);
   U22950 : AOI22_X1 port map( A1 => n24560, A2 => n8061, B1 => n24554, B2 => 
                           n8253, ZN => n23161);
   U22951 : AOI22_X1 port map( A1 => n24536, A2 => n8317, B1 => n24530, B2 => 
                           n23920, ZN => n23162);
   U22952 : AOI22_X1 port map( A1 => n24560, A2 => n8060, B1 => n24554, B2 => 
                           n8252, ZN => n23143);
   U22953 : AOI22_X1 port map( A1 => n24536, A2 => n8316, B1 => n24530, B2 => 
                           n23922, ZN => n23144);
   U22954 : AOI22_X1 port map( A1 => n24560, A2 => n8059, B1 => n24554, B2 => 
                           n8251, ZN => n23125);
   U22955 : AOI22_X1 port map( A1 => n24536, A2 => n8315, B1 => n24530, B2 => 
                           n23924, ZN => n23126);
   U22956 : AOI22_X1 port map( A1 => n24560, A2 => n8058, B1 => n24554, B2 => 
                           n8250, ZN => n23107);
   U22957 : AOI22_X1 port map( A1 => n24536, A2 => n8314, B1 => n24530, B2 => 
                           n23926, ZN => n23108);
   U22958 : AOI22_X1 port map( A1 => n24561, A2 => n8057, B1 => n24555, B2 => 
                           n8249, ZN => n23089);
   U22959 : AOI22_X1 port map( A1 => n24537, A2 => n8313, B1 => n24531, B2 => 
                           n23928, ZN => n23090);
   U22960 : AOI22_X1 port map( A1 => n24561, A2 => n8056, B1 => n24555, B2 => 
                           n8248, ZN => n23071);
   U22961 : AOI22_X1 port map( A1 => n24537, A2 => n8312, B1 => n24531, B2 => 
                           n23930, ZN => n23072);
   U22962 : AOI22_X1 port map( A1 => n24561, A2 => n8055, B1 => n24555, B2 => 
                           n8247, ZN => n23053);
   U22963 : AOI22_X1 port map( A1 => n24537, A2 => n8311, B1 => n24531, B2 => 
                           n23932, ZN => n23054);
   U22964 : AOI22_X1 port map( A1 => n24561, A2 => n8054, B1 => n24555, B2 => 
                           n8246, ZN => n23035);
   U22965 : AOI22_X1 port map( A1 => n24537, A2 => n8310, B1 => n24531, B2 => 
                           n23934, ZN => n23036);
   U22966 : OAI22_X1 port map( A1 => n24831, A2 => n20249, B1 => n24819, B2 => 
                           n25359, ZN => n5064);
   U22967 : OAI22_X1 port map( A1 => n24831, A2 => n20248, B1 => n24819, B2 => 
                           n25362, ZN => n5065);
   U22968 : OAI22_X1 port map( A1 => n24831, A2 => n20247, B1 => n24819, B2 => 
                           n25365, ZN => n5066);
   U22969 : OAI22_X1 port map( A1 => n24831, A2 => n20246, B1 => n24819, B2 => 
                           n25368, ZN => n5067);
   U22970 : OAI22_X1 port map( A1 => n24831, A2 => n20245, B1 => n24819, B2 => 
                           n25371, ZN => n5068);
   U22971 : OAI22_X1 port map( A1 => n24830, A2 => n20244, B1 => n24819, B2 => 
                           n25374, ZN => n5069);
   U22972 : OAI22_X1 port map( A1 => n24830, A2 => n20243, B1 => n24819, B2 => 
                           n25377, ZN => n5070);
   U22973 : OAI22_X1 port map( A1 => n24830, A2 => n20242, B1 => n24819, B2 => 
                           n25380, ZN => n5071);
   U22974 : OAI22_X1 port map( A1 => n24830, A2 => n20241, B1 => n24819, B2 => 
                           n25383, ZN => n5072);
   U22975 : OAI22_X1 port map( A1 => n24830, A2 => n20240, B1 => n24819, B2 => 
                           n25386, ZN => n5073);
   U22976 : OAI22_X1 port map( A1 => n24829, A2 => n20239, B1 => n24819, B2 => 
                           n25389, ZN => n5074);
   U22977 : OAI22_X1 port map( A1 => n24829, A2 => n20238, B1 => n24819, B2 => 
                           n25392, ZN => n5075);
   U22978 : OAI22_X1 port map( A1 => n24829, A2 => n20237, B1 => n24817, B2 => 
                           n25395, ZN => n5076);
   U22979 : OAI22_X1 port map( A1 => n24829, A2 => n20236, B1 => n24819, B2 => 
                           n25398, ZN => n5077);
   U22980 : OAI22_X1 port map( A1 => n24829, A2 => n20235, B1 => n24818, B2 => 
                           n25401, ZN => n5078);
   U22981 : OAI22_X1 port map( A1 => n24828, A2 => n20234, B1 => n24817, B2 => 
                           n25404, ZN => n5079);
   U22982 : OAI22_X1 port map( A1 => n24828, A2 => n20233, B1 => n24819, B2 => 
                           n25407, ZN => n5080);
   U22983 : OAI22_X1 port map( A1 => n24828, A2 => n20232, B1 => n24818, B2 => 
                           n25410, ZN => n5081);
   U22984 : OAI22_X1 port map( A1 => n24828, A2 => n20231, B1 => n24817, B2 => 
                           n25413, ZN => n5082);
   U22985 : OAI22_X1 port map( A1 => n24828, A2 => n20230, B1 => n24819, B2 => 
                           n25416, ZN => n5083);
   U22986 : OAI22_X1 port map( A1 => n24827, A2 => n20229, B1 => n24818, B2 => 
                           n25419, ZN => n5084);
   U22987 : OAI22_X1 port map( A1 => n24827, A2 => n20228, B1 => n24817, B2 => 
                           n25422, ZN => n5085);
   U22988 : OAI22_X1 port map( A1 => n24827, A2 => n20227, B1 => n24819, B2 => 
                           n25425, ZN => n5086);
   U22989 : OAI22_X1 port map( A1 => n24827, A2 => n20226, B1 => n24818, B2 => 
                           n25428, ZN => n5087);
   U22990 : OAI22_X1 port map( A1 => n24827, A2 => n20225, B1 => n24818, B2 => 
                           n25431, ZN => n5088);
   U22991 : OAI22_X1 port map( A1 => n24826, A2 => n20224, B1 => n24817, B2 => 
                           n25434, ZN => n5089);
   U22992 : OAI22_X1 port map( A1 => n24826, A2 => n20223, B1 => n24819, B2 => 
                           n25437, ZN => n5090);
   U22993 : OAI22_X1 port map( A1 => n24826, A2 => n20222, B1 => n24818, B2 => 
                           n25440, ZN => n5091);
   U22994 : OAI22_X1 port map( A1 => n24826, A2 => n20221, B1 => n24818, B2 => 
                           n25443, ZN => n5092);
   U22995 : OAI22_X1 port map( A1 => n24826, A2 => n20220, B1 => n24817, B2 => 
                           n25446, ZN => n5093);
   U22996 : OAI22_X1 port map( A1 => n24825, A2 => n20219, B1 => n24819, B2 => 
                           n25449, ZN => n5094);
   U22997 : OAI22_X1 port map( A1 => n24825, A2 => n20218, B1 => n24817, B2 => 
                           n25452, ZN => n5095);
   U22998 : OAI22_X1 port map( A1 => n24825, A2 => n20217, B1 => n24818, B2 => 
                           n25455, ZN => n5096);
   U22999 : OAI22_X1 port map( A1 => n24825, A2 => n20216, B1 => n24817, B2 => 
                           n25458, ZN => n5097);
   U23000 : OAI22_X1 port map( A1 => n24825, A2 => n20215, B1 => n24819, B2 => 
                           n25461, ZN => n5098);
   U23001 : OAI22_X1 port map( A1 => n24824, A2 => n20214, B1 => n24819, B2 => 
                           n25464, ZN => n5099);
   U23002 : OAI22_X1 port map( A1 => n24832, A2 => n20526, B1 => n24818, B2 => 
                           n25347, ZN => n5060);
   U23003 : OAI22_X1 port map( A1 => n24832, A2 => n20189, B1 => n24817, B2 => 
                           n25350, ZN => n5061);
   U23004 : OAI22_X1 port map( A1 => n24832, A2 => n20188, B1 => n24819, B2 => 
                           n25353, ZN => n5062);
   U23005 : OAI22_X1 port map( A1 => n24832, A2 => n20187, B1 => n24818, B2 => 
                           n25356, ZN => n5063);
   U23006 : OAI22_X1 port map( A1 => n25337, A2 => n25450, B1 => n93, B2 => 
                           n25327, ZN => n7015);
   U23007 : OAI22_X1 port map( A1 => n25337, A2 => n25462, B1 => n89, B2 => 
                           n21255, ZN => n7019);
   U23008 : OAI22_X1 port map( A1 => n25338, A2 => n25468, B1 => n87, B2 => 
                           n25327, ZN => n7021);
   U23009 : OAI22_X1 port map( A1 => n25338, A2 => n25474, B1 => n85, B2 => 
                           n21255, ZN => n7023);
   U23010 : OAI22_X1 port map( A1 => n25338, A2 => n25477, B1 => n84, B2 => 
                           n25327, ZN => n7024);
   U23011 : OAI22_X1 port map( A1 => n25339, A2 => n25480, B1 => n83, B2 => 
                           n21255, ZN => n7025);
   U23012 : OAI22_X1 port map( A1 => n25339, A2 => n25483, B1 => n82, B2 => 
                           n25327, ZN => n7026);
   U23013 : OAI22_X1 port map( A1 => n25339, A2 => n25486, B1 => n81, B2 => 
                           n21255, ZN => n7027);
   U23014 : OAI22_X1 port map( A1 => n25339, A2 => n25489, B1 => n80, B2 => 
                           n25327, ZN => n7028);
   U23015 : OAI22_X1 port map( A1 => n25339, A2 => n25492, B1 => n79, B2 => 
                           n21255, ZN => n7029);
   U23016 : OAI22_X1 port map( A1 => n25340, A2 => n25495, B1 => n78, B2 => 
                           n25327, ZN => n7030);
   U23017 : OAI22_X1 port map( A1 => n25340, A2 => n25498, B1 => n77, B2 => 
                           n21255, ZN => n7031);
   U23018 : OAI22_X1 port map( A1 => n25262, A2 => n25345, B1 => n17410, B2 => 
                           n25260, ZN => n6724);
   U23019 : OAI22_X1 port map( A1 => n25262, A2 => n25348, B1 => n17407, B2 => 
                           n25260, ZN => n6725);
   U23020 : OAI22_X1 port map( A1 => n25262, A2 => n25351, B1 => n17404, B2 => 
                           n25260, ZN => n6726);
   U23021 : OAI22_X1 port map( A1 => n25262, A2 => n25354, B1 => n17401, B2 => 
                           n25260, ZN => n6727);
   U23022 : OAI22_X1 port map( A1 => n25262, A2 => n25357, B1 => n17398, B2 => 
                           n25260, ZN => n6728);
   U23023 : OAI22_X1 port map( A1 => n25263, A2 => n25360, B1 => n17395, B2 => 
                           n25260, ZN => n6729);
   U23024 : OAI22_X1 port map( A1 => n25263, A2 => n25363, B1 => n17392, B2 => 
                           n25260, ZN => n6730);
   U23025 : OAI22_X1 port map( A1 => n25263, A2 => n25366, B1 => n17389, B2 => 
                           n25260, ZN => n6731);
   U23026 : OAI22_X1 port map( A1 => n25263, A2 => n25369, B1 => n17386, B2 => 
                           n25260, ZN => n6732);
   U23027 : OAI22_X1 port map( A1 => n25263, A2 => n25372, B1 => n17383, B2 => 
                           n25260, ZN => n6733);
   U23028 : OAI22_X1 port map( A1 => n25264, A2 => n25375, B1 => n17380, B2 => 
                           n25260, ZN => n6734);
   U23029 : OAI22_X1 port map( A1 => n25264, A2 => n25378, B1 => n17377, B2 => 
                           n25260, ZN => n6735);
   U23030 : OAI22_X1 port map( A1 => n25264, A2 => n25381, B1 => n17374, B2 => 
                           n25261, ZN => n6736);
   U23031 : OAI22_X1 port map( A1 => n25264, A2 => n25384, B1 => n17371, B2 => 
                           n25261, ZN => n6737);
   U23032 : OAI22_X1 port map( A1 => n25264, A2 => n25387, B1 => n17368, B2 => 
                           n25261, ZN => n6738);
   U23033 : OAI22_X1 port map( A1 => n25265, A2 => n25390, B1 => n17365, B2 => 
                           n25261, ZN => n6739);
   U23034 : OAI22_X1 port map( A1 => n25265, A2 => n25393, B1 => n17362, B2 => 
                           n25261, ZN => n6740);
   U23035 : OAI22_X1 port map( A1 => n25265, A2 => n25396, B1 => n17359, B2 => 
                           n25261, ZN => n6741);
   U23036 : OAI22_X1 port map( A1 => n25265, A2 => n25399, B1 => n17356, B2 => 
                           n25261, ZN => n6742);
   U23037 : OAI22_X1 port map( A1 => n25265, A2 => n25402, B1 => n17353, B2 => 
                           n25261, ZN => n6743);
   U23038 : OAI22_X1 port map( A1 => n25266, A2 => n25405, B1 => n17350, B2 => 
                           n25261, ZN => n6744);
   U23039 : OAI22_X1 port map( A1 => n25266, A2 => n25408, B1 => n17347, B2 => 
                           n25261, ZN => n6745);
   U23040 : OAI22_X1 port map( A1 => n25266, A2 => n25411, B1 => n17344, B2 => 
                           n25261, ZN => n6746);
   U23041 : OAI22_X1 port map( A1 => n25266, A2 => n25414, B1 => n17341, B2 => 
                           n25261, ZN => n6747);
   U23042 : OAI22_X1 port map( A1 => n25177, A2 => n25345, B1 => n7554, B2 => 
                           n25175, ZN => n6404);
   U23043 : OAI22_X1 port map( A1 => n25177, A2 => n25348, B1 => n7552, B2 => 
                           n25175, ZN => n6405);
   U23044 : OAI22_X1 port map( A1 => n25177, A2 => n25351, B1 => n7550, B2 => 
                           n25175, ZN => n6406);
   U23045 : OAI22_X1 port map( A1 => n25177, A2 => n25354, B1 => n7548, B2 => 
                           n25175, ZN => n6407);
   U23046 : OAI22_X1 port map( A1 => n25177, A2 => n25357, B1 => n7546, B2 => 
                           n25175, ZN => n6408);
   U23047 : OAI22_X1 port map( A1 => n25178, A2 => n25360, B1 => n7544, B2 => 
                           n25175, ZN => n6409);
   U23048 : OAI22_X1 port map( A1 => n25178, A2 => n25363, B1 => n7542, B2 => 
                           n25175, ZN => n6410);
   U23049 : OAI22_X1 port map( A1 => n25178, A2 => n25366, B1 => n7540, B2 => 
                           n25175, ZN => n6411);
   U23050 : OAI22_X1 port map( A1 => n25178, A2 => n25369, B1 => n7538, B2 => 
                           n25175, ZN => n6412);
   U23051 : OAI22_X1 port map( A1 => n25178, A2 => n25372, B1 => n7536, B2 => 
                           n25175, ZN => n6413);
   U23052 : OAI22_X1 port map( A1 => n25179, A2 => n25375, B1 => n7534, B2 => 
                           n25175, ZN => n6414);
   U23053 : OAI22_X1 port map( A1 => n25179, A2 => n25378, B1 => n7532, B2 => 
                           n25175, ZN => n6415);
   U23054 : OAI22_X1 port map( A1 => n25179, A2 => n25381, B1 => n7530, B2 => 
                           n25176, ZN => n6416);
   U23055 : OAI22_X1 port map( A1 => n25179, A2 => n25384, B1 => n7528, B2 => 
                           n25176, ZN => n6417);
   U23056 : OAI22_X1 port map( A1 => n25179, A2 => n25387, B1 => n7526, B2 => 
                           n25176, ZN => n6418);
   U23057 : OAI22_X1 port map( A1 => n25180, A2 => n25390, B1 => n7524, B2 => 
                           n25176, ZN => n6419);
   U23058 : OAI22_X1 port map( A1 => n25180, A2 => n25393, B1 => n7522, B2 => 
                           n25176, ZN => n6420);
   U23059 : OAI22_X1 port map( A1 => n25180, A2 => n25396, B1 => n7520, B2 => 
                           n25176, ZN => n6421);
   U23060 : OAI22_X1 port map( A1 => n25180, A2 => n25399, B1 => n7518, B2 => 
                           n25176, ZN => n6422);
   U23061 : OAI22_X1 port map( A1 => n25180, A2 => n25402, B1 => n7516, B2 => 
                           n25176, ZN => n6423);
   U23062 : OAI22_X1 port map( A1 => n25181, A2 => n25405, B1 => n7514, B2 => 
                           n25176, ZN => n6424);
   U23063 : OAI22_X1 port map( A1 => n25181, A2 => n25408, B1 => n7512, B2 => 
                           n25176, ZN => n6425);
   U23064 : OAI22_X1 port map( A1 => n25181, A2 => n25411, B1 => n7510, B2 => 
                           n25176, ZN => n6426);
   U23065 : OAI22_X1 port map( A1 => n25181, A2 => n25414, B1 => n7508, B2 => 
                           n25176, ZN => n6427);
   U23066 : OAI22_X1 port map( A1 => n25092, A2 => n25346, B1 => n7426, B2 => 
                           n25090, ZN => n6084);
   U23067 : OAI22_X1 port map( A1 => n25092, A2 => n25349, B1 => n7424, B2 => 
                           n25090, ZN => n6085);
   U23068 : OAI22_X1 port map( A1 => n25092, A2 => n25352, B1 => n7422, B2 => 
                           n25090, ZN => n6086);
   U23069 : OAI22_X1 port map( A1 => n25092, A2 => n25355, B1 => n7420, B2 => 
                           n25090, ZN => n6087);
   U23070 : OAI22_X1 port map( A1 => n25092, A2 => n25358, B1 => n7418, B2 => 
                           n25090, ZN => n6088);
   U23071 : OAI22_X1 port map( A1 => n25093, A2 => n25361, B1 => n7416, B2 => 
                           n25090, ZN => n6089);
   U23072 : OAI22_X1 port map( A1 => n25093, A2 => n25364, B1 => n7414, B2 => 
                           n25090, ZN => n6090);
   U23073 : OAI22_X1 port map( A1 => n25093, A2 => n25367, B1 => n7412, B2 => 
                           n25090, ZN => n6091);
   U23074 : OAI22_X1 port map( A1 => n25093, A2 => n25370, B1 => n7410, B2 => 
                           n25090, ZN => n6092);
   U23075 : OAI22_X1 port map( A1 => n25093, A2 => n25373, B1 => n7408, B2 => 
                           n25090, ZN => n6093);
   U23076 : OAI22_X1 port map( A1 => n25094, A2 => n25376, B1 => n7406, B2 => 
                           n25090, ZN => n6094);
   U23077 : OAI22_X1 port map( A1 => n25094, A2 => n25379, B1 => n7404, B2 => 
                           n25090, ZN => n6095);
   U23078 : OAI22_X1 port map( A1 => n25094, A2 => n25382, B1 => n7402, B2 => 
                           n25091, ZN => n6096);
   U23079 : OAI22_X1 port map( A1 => n25094, A2 => n25385, B1 => n7400, B2 => 
                           n25091, ZN => n6097);
   U23080 : OAI22_X1 port map( A1 => n25094, A2 => n25388, B1 => n7398, B2 => 
                           n25091, ZN => n6098);
   U23081 : OAI22_X1 port map( A1 => n25095, A2 => n25391, B1 => n7396, B2 => 
                           n25091, ZN => n6099);
   U23082 : OAI22_X1 port map( A1 => n25095, A2 => n25394, B1 => n7394, B2 => 
                           n25091, ZN => n6100);
   U23083 : OAI22_X1 port map( A1 => n25095, A2 => n25397, B1 => n7392, B2 => 
                           n25091, ZN => n6101);
   U23084 : OAI22_X1 port map( A1 => n25095, A2 => n25400, B1 => n7390, B2 => 
                           n25091, ZN => n6102);
   U23085 : OAI22_X1 port map( A1 => n25095, A2 => n25403, B1 => n7388, B2 => 
                           n25091, ZN => n6103);
   U23086 : OAI22_X1 port map( A1 => n25096, A2 => n25406, B1 => n7386, B2 => 
                           n25091, ZN => n6104);
   U23087 : OAI22_X1 port map( A1 => n25096, A2 => n25409, B1 => n7384, B2 => 
                           n25091, ZN => n6105);
   U23088 : OAI22_X1 port map( A1 => n25096, A2 => n25412, B1 => n7382, B2 => 
                           n25091, ZN => n6106);
   U23089 : OAI22_X1 port map( A1 => n25096, A2 => n25415, B1 => n7380, B2 => 
                           n25091, ZN => n6107);
   U23090 : OAI22_X1 port map( A1 => n25041, A2 => n25346, B1 => n8861, B2 => 
                           n25039, ZN => n5892);
   U23091 : OAI22_X1 port map( A1 => n25041, A2 => n25349, B1 => n8859, B2 => 
                           n25039, ZN => n5893);
   U23092 : OAI22_X1 port map( A1 => n25041, A2 => n25352, B1 => n8857, B2 => 
                           n25039, ZN => n5894);
   U23093 : OAI22_X1 port map( A1 => n25041, A2 => n25355, B1 => n8855, B2 => 
                           n25039, ZN => n5895);
   U23094 : OAI22_X1 port map( A1 => n25041, A2 => n25358, B1 => n8853, B2 => 
                           n25039, ZN => n5896);
   U23095 : OAI22_X1 port map( A1 => n25042, A2 => n25361, B1 => n8851, B2 => 
                           n25039, ZN => n5897);
   U23096 : OAI22_X1 port map( A1 => n25042, A2 => n25364, B1 => n8849, B2 => 
                           n25039, ZN => n5898);
   U23097 : OAI22_X1 port map( A1 => n25042, A2 => n25367, B1 => n8847, B2 => 
                           n25039, ZN => n5899);
   U23098 : OAI22_X1 port map( A1 => n25042, A2 => n25370, B1 => n8845, B2 => 
                           n25039, ZN => n5900);
   U23099 : OAI22_X1 port map( A1 => n25042, A2 => n25373, B1 => n8843, B2 => 
                           n25039, ZN => n5901);
   U23100 : OAI22_X1 port map( A1 => n25043, A2 => n25376, B1 => n8841, B2 => 
                           n25039, ZN => n5902);
   U23101 : OAI22_X1 port map( A1 => n25043, A2 => n25379, B1 => n8839, B2 => 
                           n25039, ZN => n5903);
   U23102 : OAI22_X1 port map( A1 => n25043, A2 => n25382, B1 => n8837, B2 => 
                           n25040, ZN => n5904);
   U23103 : OAI22_X1 port map( A1 => n25043, A2 => n25385, B1 => n8835, B2 => 
                           n25040, ZN => n5905);
   U23104 : OAI22_X1 port map( A1 => n25043, A2 => n25388, B1 => n8833, B2 => 
                           n25040, ZN => n5906);
   U23105 : OAI22_X1 port map( A1 => n25044, A2 => n25391, B1 => n8831, B2 => 
                           n25040, ZN => n5907);
   U23106 : OAI22_X1 port map( A1 => n25044, A2 => n25394, B1 => n8829, B2 => 
                           n25040, ZN => n5908);
   U23107 : OAI22_X1 port map( A1 => n25044, A2 => n25397, B1 => n8827, B2 => 
                           n25040, ZN => n5909);
   U23108 : OAI22_X1 port map( A1 => n25044, A2 => n25400, B1 => n8825, B2 => 
                           n25040, ZN => n5910);
   U23109 : OAI22_X1 port map( A1 => n25044, A2 => n25403, B1 => n8823, B2 => 
                           n25040, ZN => n5911);
   U23110 : OAI22_X1 port map( A1 => n25045, A2 => n25406, B1 => n8821, B2 => 
                           n25040, ZN => n5912);
   U23111 : OAI22_X1 port map( A1 => n25045, A2 => n25409, B1 => n8819, B2 => 
                           n25040, ZN => n5913);
   U23112 : OAI22_X1 port map( A1 => n25045, A2 => n25412, B1 => n8817, B2 => 
                           n25040, ZN => n5914);
   U23113 : OAI22_X1 port map( A1 => n25045, A2 => n25415, B1 => n8815, B2 => 
                           n25040, ZN => n5915);
   U23114 : OAI22_X1 port map( A1 => n25024, A2 => n25346, B1 => n8989, B2 => 
                           n25022, ZN => n5828);
   U23115 : OAI22_X1 port map( A1 => n25024, A2 => n25349, B1 => n8987, B2 => 
                           n25022, ZN => n5829);
   U23116 : OAI22_X1 port map( A1 => n25024, A2 => n25352, B1 => n8985, B2 => 
                           n25022, ZN => n5830);
   U23117 : OAI22_X1 port map( A1 => n25024, A2 => n25355, B1 => n8983, B2 => 
                           n25022, ZN => n5831);
   U23118 : OAI22_X1 port map( A1 => n25024, A2 => n25358, B1 => n8981, B2 => 
                           n25022, ZN => n5832);
   U23119 : OAI22_X1 port map( A1 => n25025, A2 => n25361, B1 => n8979, B2 => 
                           n25022, ZN => n5833);
   U23120 : OAI22_X1 port map( A1 => n25025, A2 => n25364, B1 => n8977, B2 => 
                           n25022, ZN => n5834);
   U23121 : OAI22_X1 port map( A1 => n25025, A2 => n25367, B1 => n8975, B2 => 
                           n25022, ZN => n5835);
   U23122 : OAI22_X1 port map( A1 => n25025, A2 => n25370, B1 => n8973, B2 => 
                           n25022, ZN => n5836);
   U23123 : OAI22_X1 port map( A1 => n25025, A2 => n25373, B1 => n8971, B2 => 
                           n25022, ZN => n5837);
   U23124 : OAI22_X1 port map( A1 => n25026, A2 => n25376, B1 => n8969, B2 => 
                           n25022, ZN => n5838);
   U23125 : OAI22_X1 port map( A1 => n25026, A2 => n25379, B1 => n8967, B2 => 
                           n25022, ZN => n5839);
   U23126 : OAI22_X1 port map( A1 => n25026, A2 => n25382, B1 => n8965, B2 => 
                           n25023, ZN => n5840);
   U23127 : OAI22_X1 port map( A1 => n25026, A2 => n25385, B1 => n8963, B2 => 
                           n25023, ZN => n5841);
   U23128 : OAI22_X1 port map( A1 => n25026, A2 => n25388, B1 => n8961, B2 => 
                           n25023, ZN => n5842);
   U23129 : OAI22_X1 port map( A1 => n25027, A2 => n25391, B1 => n8959, B2 => 
                           n25023, ZN => n5843);
   U23130 : OAI22_X1 port map( A1 => n25027, A2 => n25394, B1 => n8957, B2 => 
                           n25023, ZN => n5844);
   U23131 : OAI22_X1 port map( A1 => n25027, A2 => n25397, B1 => n8955, B2 => 
                           n25023, ZN => n5845);
   U23132 : OAI22_X1 port map( A1 => n25027, A2 => n25400, B1 => n8953, B2 => 
                           n25023, ZN => n5846);
   U23133 : OAI22_X1 port map( A1 => n25027, A2 => n25403, B1 => n8951, B2 => 
                           n25023, ZN => n5847);
   U23134 : OAI22_X1 port map( A1 => n25028, A2 => n25406, B1 => n8949, B2 => 
                           n25023, ZN => n5848);
   U23135 : OAI22_X1 port map( A1 => n25028, A2 => n25409, B1 => n8947, B2 => 
                           n25023, ZN => n5849);
   U23136 : OAI22_X1 port map( A1 => n25028, A2 => n25412, B1 => n8945, B2 => 
                           n25023, ZN => n5850);
   U23137 : OAI22_X1 port map( A1 => n25028, A2 => n25415, B1 => n8943, B2 => 
                           n25023, ZN => n5851);
   U23138 : OAI22_X1 port map( A1 => n24854, A2 => n25347, B1 => n8988, B2 => 
                           n24852, ZN => n5188);
   U23139 : OAI22_X1 port map( A1 => n24854, A2 => n25350, B1 => n8986, B2 => 
                           n24852, ZN => n5189);
   U23140 : OAI22_X1 port map( A1 => n24854, A2 => n25353, B1 => n8984, B2 => 
                           n24852, ZN => n5190);
   U23141 : OAI22_X1 port map( A1 => n24854, A2 => n25356, B1 => n8982, B2 => 
                           n24852, ZN => n5191);
   U23142 : OAI22_X1 port map( A1 => n24854, A2 => n25359, B1 => n8980, B2 => 
                           n24852, ZN => n5192);
   U23143 : OAI22_X1 port map( A1 => n24855, A2 => n25362, B1 => n8978, B2 => 
                           n24852, ZN => n5193);
   U23144 : OAI22_X1 port map( A1 => n24855, A2 => n25365, B1 => n8976, B2 => 
                           n24852, ZN => n5194);
   U23145 : OAI22_X1 port map( A1 => n24855, A2 => n25368, B1 => n8974, B2 => 
                           n24852, ZN => n5195);
   U23146 : OAI22_X1 port map( A1 => n24855, A2 => n25371, B1 => n8972, B2 => 
                           n24852, ZN => n5196);
   U23147 : OAI22_X1 port map( A1 => n24855, A2 => n25374, B1 => n8970, B2 => 
                           n24852, ZN => n5197);
   U23148 : OAI22_X1 port map( A1 => n24856, A2 => n25377, B1 => n8968, B2 => 
                           n24852, ZN => n5198);
   U23149 : OAI22_X1 port map( A1 => n24856, A2 => n25380, B1 => n8966, B2 => 
                           n24852, ZN => n5199);
   U23150 : OAI22_X1 port map( A1 => n24856, A2 => n25383, B1 => n8964, B2 => 
                           n24853, ZN => n5200);
   U23151 : OAI22_X1 port map( A1 => n24856, A2 => n25386, B1 => n8962, B2 => 
                           n24853, ZN => n5201);
   U23152 : OAI22_X1 port map( A1 => n24856, A2 => n25389, B1 => n8960, B2 => 
                           n24853, ZN => n5202);
   U23153 : OAI22_X1 port map( A1 => n24857, A2 => n25392, B1 => n8958, B2 => 
                           n24853, ZN => n5203);
   U23154 : OAI22_X1 port map( A1 => n24857, A2 => n25395, B1 => n8956, B2 => 
                           n24853, ZN => n5204);
   U23155 : OAI22_X1 port map( A1 => n24857, A2 => n25398, B1 => n8954, B2 => 
                           n24853, ZN => n5205);
   U23156 : OAI22_X1 port map( A1 => n24857, A2 => n25401, B1 => n8952, B2 => 
                           n24853, ZN => n5206);
   U23157 : OAI22_X1 port map( A1 => n24857, A2 => n25404, B1 => n8950, B2 => 
                           n24853, ZN => n5207);
   U23158 : OAI22_X1 port map( A1 => n24858, A2 => n25407, B1 => n8948, B2 => 
                           n24853, ZN => n5208);
   U23159 : OAI22_X1 port map( A1 => n24858, A2 => n25410, B1 => n8946, B2 => 
                           n24853, ZN => n5209);
   U23160 : OAI22_X1 port map( A1 => n24858, A2 => n25413, B1 => n8944, B2 => 
                           n24853, ZN => n5210);
   U23161 : OAI22_X1 port map( A1 => n24858, A2 => n25416, B1 => n8942, B2 => 
                           n24853, ZN => n5211);
   U23162 : OAI22_X1 port map( A1 => n24922, A2 => n25347, B1 => n7427, B2 => 
                           n24920, ZN => n5444);
   U23163 : OAI22_X1 port map( A1 => n24922, A2 => n25350, B1 => n7425, B2 => 
                           n24920, ZN => n5445);
   U23164 : OAI22_X1 port map( A1 => n24922, A2 => n25353, B1 => n7423, B2 => 
                           n24920, ZN => n5446);
   U23165 : OAI22_X1 port map( A1 => n24922, A2 => n25356, B1 => n7421, B2 => 
                           n24920, ZN => n5447);
   U23166 : OAI22_X1 port map( A1 => n24922, A2 => n25359, B1 => n7419, B2 => 
                           n24920, ZN => n5448);
   U23167 : OAI22_X1 port map( A1 => n24923, A2 => n25362, B1 => n7417, B2 => 
                           n24920, ZN => n5449);
   U23168 : OAI22_X1 port map( A1 => n24923, A2 => n25365, B1 => n7415, B2 => 
                           n24920, ZN => n5450);
   U23169 : OAI22_X1 port map( A1 => n24923, A2 => n25368, B1 => n7413, B2 => 
                           n24920, ZN => n5451);
   U23170 : OAI22_X1 port map( A1 => n24923, A2 => n25371, B1 => n7411, B2 => 
                           n24920, ZN => n5452);
   U23171 : OAI22_X1 port map( A1 => n24923, A2 => n25374, B1 => n7409, B2 => 
                           n24920, ZN => n5453);
   U23172 : OAI22_X1 port map( A1 => n24924, A2 => n25377, B1 => n7407, B2 => 
                           n24920, ZN => n5454);
   U23173 : OAI22_X1 port map( A1 => n24924, A2 => n25380, B1 => n7405, B2 => 
                           n24920, ZN => n5455);
   U23174 : OAI22_X1 port map( A1 => n24924, A2 => n25383, B1 => n7403, B2 => 
                           n24921, ZN => n5456);
   U23175 : OAI22_X1 port map( A1 => n24924, A2 => n25386, B1 => n7401, B2 => 
                           n24921, ZN => n5457);
   U23176 : OAI22_X1 port map( A1 => n24924, A2 => n25389, B1 => n7399, B2 => 
                           n24921, ZN => n5458);
   U23177 : OAI22_X1 port map( A1 => n24925, A2 => n25392, B1 => n7397, B2 => 
                           n24921, ZN => n5459);
   U23178 : OAI22_X1 port map( A1 => n24925, A2 => n25395, B1 => n7395, B2 => 
                           n24921, ZN => n5460);
   U23179 : OAI22_X1 port map( A1 => n24925, A2 => n25398, B1 => n7393, B2 => 
                           n24921, ZN => n5461);
   U23180 : OAI22_X1 port map( A1 => n24925, A2 => n25401, B1 => n7391, B2 => 
                           n24921, ZN => n5462);
   U23181 : OAI22_X1 port map( A1 => n24925, A2 => n25404, B1 => n7389, B2 => 
                           n24921, ZN => n5463);
   U23182 : OAI22_X1 port map( A1 => n24926, A2 => n25407, B1 => n7387, B2 => 
                           n24921, ZN => n5464);
   U23183 : OAI22_X1 port map( A1 => n24926, A2 => n25410, B1 => n7385, B2 => 
                           n24921, ZN => n5465);
   U23184 : OAI22_X1 port map( A1 => n24926, A2 => n25413, B1 => n7383, B2 => 
                           n24921, ZN => n5466);
   U23185 : OAI22_X1 port map( A1 => n24926, A2 => n25416, B1 => n7381, B2 => 
                           n24921, ZN => n5467);
   U23186 : OAI22_X1 port map( A1 => n24956, A2 => n25346, B1 => n9245, B2 => 
                           n24954, ZN => n5572);
   U23187 : OAI22_X1 port map( A1 => n24956, A2 => n25349, B1 => n9243, B2 => 
                           n24954, ZN => n5573);
   U23188 : OAI22_X1 port map( A1 => n24956, A2 => n25352, B1 => n9241, B2 => 
                           n24954, ZN => n5574);
   U23189 : OAI22_X1 port map( A1 => n24956, A2 => n25355, B1 => n9239, B2 => 
                           n24954, ZN => n5575);
   U23190 : OAI22_X1 port map( A1 => n24956, A2 => n25358, B1 => n9237, B2 => 
                           n24954, ZN => n5576);
   U23191 : OAI22_X1 port map( A1 => n24957, A2 => n25361, B1 => n9235, B2 => 
                           n24954, ZN => n5577);
   U23192 : OAI22_X1 port map( A1 => n24957, A2 => n25364, B1 => n9233, B2 => 
                           n24954, ZN => n5578);
   U23193 : OAI22_X1 port map( A1 => n24957, A2 => n25367, B1 => n9231, B2 => 
                           n24954, ZN => n5579);
   U23194 : OAI22_X1 port map( A1 => n24957, A2 => n25370, B1 => n9229, B2 => 
                           n24954, ZN => n5580);
   U23195 : OAI22_X1 port map( A1 => n24957, A2 => n25373, B1 => n9227, B2 => 
                           n24954, ZN => n5581);
   U23196 : OAI22_X1 port map( A1 => n24958, A2 => n25376, B1 => n9225, B2 => 
                           n24954, ZN => n5582);
   U23197 : OAI22_X1 port map( A1 => n24958, A2 => n25379, B1 => n9223, B2 => 
                           n24954, ZN => n5583);
   U23198 : OAI22_X1 port map( A1 => n24958, A2 => n25382, B1 => n9221, B2 => 
                           n24955, ZN => n5584);
   U23199 : OAI22_X1 port map( A1 => n24958, A2 => n25385, B1 => n9219, B2 => 
                           n24955, ZN => n5585);
   U23200 : OAI22_X1 port map( A1 => n24958, A2 => n25388, B1 => n9217, B2 => 
                           n24955, ZN => n5586);
   U23201 : OAI22_X1 port map( A1 => n24959, A2 => n25391, B1 => n9215, B2 => 
                           n24955, ZN => n5587);
   U23202 : OAI22_X1 port map( A1 => n24959, A2 => n25394, B1 => n9213, B2 => 
                           n24955, ZN => n5588);
   U23203 : OAI22_X1 port map( A1 => n24959, A2 => n25397, B1 => n9211, B2 => 
                           n24955, ZN => n5589);
   U23204 : OAI22_X1 port map( A1 => n24959, A2 => n25400, B1 => n9209, B2 => 
                           n24955, ZN => n5590);
   U23205 : OAI22_X1 port map( A1 => n24959, A2 => n25403, B1 => n9207, B2 => 
                           n24955, ZN => n5591);
   U23206 : OAI22_X1 port map( A1 => n24960, A2 => n25406, B1 => n9205, B2 => 
                           n24955, ZN => n5592);
   U23207 : OAI22_X1 port map( A1 => n24960, A2 => n25409, B1 => n9203, B2 => 
                           n24955, ZN => n5593);
   U23208 : OAI22_X1 port map( A1 => n24960, A2 => n25412, B1 => n9201, B2 => 
                           n24955, ZN => n5594);
   U23209 : OAI22_X1 port map( A1 => n24960, A2 => n25415, B1 => n9199, B2 => 
                           n24955, ZN => n5595);
   U23210 : OAI22_X1 port map( A1 => n24973, A2 => n25346, B1 => n7555, B2 => 
                           n24971, ZN => n5636);
   U23211 : OAI22_X1 port map( A1 => n24973, A2 => n25349, B1 => n7553, B2 => 
                           n24971, ZN => n5637);
   U23212 : OAI22_X1 port map( A1 => n24973, A2 => n25352, B1 => n7551, B2 => 
                           n24971, ZN => n5638);
   U23213 : OAI22_X1 port map( A1 => n24973, A2 => n25355, B1 => n7549, B2 => 
                           n24971, ZN => n5639);
   U23214 : OAI22_X1 port map( A1 => n24973, A2 => n25358, B1 => n7547, B2 => 
                           n24971, ZN => n5640);
   U23215 : OAI22_X1 port map( A1 => n24974, A2 => n25361, B1 => n7545, B2 => 
                           n24971, ZN => n5641);
   U23216 : OAI22_X1 port map( A1 => n24974, A2 => n25364, B1 => n7543, B2 => 
                           n24971, ZN => n5642);
   U23217 : OAI22_X1 port map( A1 => n24974, A2 => n25367, B1 => n7541, B2 => 
                           n24971, ZN => n5643);
   U23218 : OAI22_X1 port map( A1 => n24974, A2 => n25370, B1 => n7539, B2 => 
                           n24971, ZN => n5644);
   U23219 : OAI22_X1 port map( A1 => n24974, A2 => n25373, B1 => n7537, B2 => 
                           n24971, ZN => n5645);
   U23220 : OAI22_X1 port map( A1 => n24975, A2 => n25376, B1 => n7535, B2 => 
                           n24971, ZN => n5646);
   U23221 : OAI22_X1 port map( A1 => n24975, A2 => n25379, B1 => n7533, B2 => 
                           n24971, ZN => n5647);
   U23222 : OAI22_X1 port map( A1 => n24975, A2 => n25382, B1 => n7531, B2 => 
                           n24972, ZN => n5648);
   U23223 : OAI22_X1 port map( A1 => n24975, A2 => n25385, B1 => n7529, B2 => 
                           n24972, ZN => n5649);
   U23224 : OAI22_X1 port map( A1 => n24975, A2 => n25388, B1 => n7527, B2 => 
                           n24972, ZN => n5650);
   U23225 : OAI22_X1 port map( A1 => n24976, A2 => n25391, B1 => n7525, B2 => 
                           n24972, ZN => n5651);
   U23226 : OAI22_X1 port map( A1 => n24976, A2 => n25394, B1 => n7523, B2 => 
                           n24972, ZN => n5652);
   U23227 : OAI22_X1 port map( A1 => n24976, A2 => n25397, B1 => n7521, B2 => 
                           n24972, ZN => n5653);
   U23228 : OAI22_X1 port map( A1 => n24976, A2 => n25400, B1 => n7519, B2 => 
                           n24972, ZN => n5654);
   U23229 : OAI22_X1 port map( A1 => n24976, A2 => n25403, B1 => n7517, B2 => 
                           n24972, ZN => n5655);
   U23230 : OAI22_X1 port map( A1 => n24977, A2 => n25406, B1 => n7515, B2 => 
                           n24972, ZN => n5656);
   U23231 : OAI22_X1 port map( A1 => n24977, A2 => n25409, B1 => n7513, B2 => 
                           n24972, ZN => n5657);
   U23232 : OAI22_X1 port map( A1 => n24977, A2 => n25412, B1 => n7511, B2 => 
                           n24972, ZN => n5658);
   U23233 : OAI22_X1 port map( A1 => n24977, A2 => n25415, B1 => n7509, B2 => 
                           n24972, ZN => n5659);
   U23234 : OAI22_X1 port map( A1 => n25109, A2 => n25346, B1 => n9116, B2 => 
                           n25107, ZN => n6148);
   U23235 : OAI22_X1 port map( A1 => n25109, A2 => n25349, B1 => n9114, B2 => 
                           n25107, ZN => n6149);
   U23236 : OAI22_X1 port map( A1 => n25109, A2 => n25352, B1 => n9112, B2 => 
                           n25107, ZN => n6150);
   U23237 : OAI22_X1 port map( A1 => n25109, A2 => n25355, B1 => n9110, B2 => 
                           n25107, ZN => n6151);
   U23238 : OAI22_X1 port map( A1 => n25109, A2 => n25358, B1 => n9108, B2 => 
                           n25107, ZN => n6152);
   U23239 : OAI22_X1 port map( A1 => n25110, A2 => n25361, B1 => n9106, B2 => 
                           n25107, ZN => n6153);
   U23240 : OAI22_X1 port map( A1 => n25110, A2 => n25364, B1 => n9104, B2 => 
                           n25107, ZN => n6154);
   U23241 : OAI22_X1 port map( A1 => n25110, A2 => n25367, B1 => n9102, B2 => 
                           n25107, ZN => n6155);
   U23242 : OAI22_X1 port map( A1 => n25110, A2 => n25370, B1 => n9100, B2 => 
                           n25107, ZN => n6156);
   U23243 : OAI22_X1 port map( A1 => n25110, A2 => n25373, B1 => n9098, B2 => 
                           n25107, ZN => n6157);
   U23244 : OAI22_X1 port map( A1 => n25111, A2 => n25376, B1 => n9096, B2 => 
                           n25107, ZN => n6158);
   U23245 : OAI22_X1 port map( A1 => n25111, A2 => n25379, B1 => n9094, B2 => 
                           n25107, ZN => n6159);
   U23246 : OAI22_X1 port map( A1 => n25111, A2 => n25382, B1 => n9092, B2 => 
                           n25108, ZN => n6160);
   U23247 : OAI22_X1 port map( A1 => n25111, A2 => n25385, B1 => n9090, B2 => 
                           n25108, ZN => n6161);
   U23248 : OAI22_X1 port map( A1 => n25111, A2 => n25388, B1 => n9088, B2 => 
                           n25108, ZN => n6162);
   U23249 : OAI22_X1 port map( A1 => n25112, A2 => n25391, B1 => n9086, B2 => 
                           n25108, ZN => n6163);
   U23250 : OAI22_X1 port map( A1 => n25112, A2 => n25394, B1 => n9084, B2 => 
                           n25108, ZN => n6164);
   U23251 : OAI22_X1 port map( A1 => n25112, A2 => n25397, B1 => n9082, B2 => 
                           n25108, ZN => n6165);
   U23252 : OAI22_X1 port map( A1 => n25112, A2 => n25400, B1 => n9080, B2 => 
                           n25108, ZN => n6166);
   U23253 : OAI22_X1 port map( A1 => n25112, A2 => n25403, B1 => n9078, B2 => 
                           n25108, ZN => n6167);
   U23254 : OAI22_X1 port map( A1 => n25113, A2 => n25406, B1 => n9076, B2 => 
                           n25108, ZN => n6168);
   U23255 : OAI22_X1 port map( A1 => n25113, A2 => n25409, B1 => n9074, B2 => 
                           n25108, ZN => n6169);
   U23256 : OAI22_X1 port map( A1 => n25113, A2 => n25412, B1 => n9072, B2 => 
                           n25108, ZN => n6170);
   U23257 : OAI22_X1 port map( A1 => n25113, A2 => n25415, B1 => n9070, B2 => 
                           n25108, ZN => n6171);
   U23258 : OAI22_X1 port map( A1 => n25126, A2 => n25346, B1 => n896, B2 => 
                           n25124, ZN => n6212);
   U23259 : OAI22_X1 port map( A1 => n25126, A2 => n25349, B1 => n895, B2 => 
                           n25124, ZN => n6213);
   U23260 : OAI22_X1 port map( A1 => n25126, A2 => n25352, B1 => n894, B2 => 
                           n25124, ZN => n6214);
   U23261 : OAI22_X1 port map( A1 => n25126, A2 => n25355, B1 => n893, B2 => 
                           n25124, ZN => n6215);
   U23262 : OAI22_X1 port map( A1 => n25126, A2 => n25358, B1 => n892, B2 => 
                           n25124, ZN => n6216);
   U23263 : OAI22_X1 port map( A1 => n25127, A2 => n25361, B1 => n891, B2 => 
                           n25124, ZN => n6217);
   U23264 : OAI22_X1 port map( A1 => n25127, A2 => n25364, B1 => n890, B2 => 
                           n25124, ZN => n6218);
   U23265 : OAI22_X1 port map( A1 => n25127, A2 => n25367, B1 => n889, B2 => 
                           n25124, ZN => n6219);
   U23266 : OAI22_X1 port map( A1 => n25127, A2 => n25370, B1 => n888, B2 => 
                           n25124, ZN => n6220);
   U23267 : OAI22_X1 port map( A1 => n25127, A2 => n25373, B1 => n887, B2 => 
                           n25124, ZN => n6221);
   U23268 : OAI22_X1 port map( A1 => n25128, A2 => n25376, B1 => n886, B2 => 
                           n25124, ZN => n6222);
   U23269 : OAI22_X1 port map( A1 => n25128, A2 => n25379, B1 => n885, B2 => 
                           n25124, ZN => n6223);
   U23270 : OAI22_X1 port map( A1 => n25128, A2 => n25382, B1 => n884, B2 => 
                           n25125, ZN => n6224);
   U23271 : OAI22_X1 port map( A1 => n25128, A2 => n25385, B1 => n883, B2 => 
                           n25125, ZN => n6225);
   U23272 : OAI22_X1 port map( A1 => n25128, A2 => n25388, B1 => n882, B2 => 
                           n25125, ZN => n6226);
   U23273 : OAI22_X1 port map( A1 => n25129, A2 => n25391, B1 => n881, B2 => 
                           n25125, ZN => n6227);
   U23274 : OAI22_X1 port map( A1 => n25129, A2 => n25394, B1 => n880, B2 => 
                           n25125, ZN => n6228);
   U23275 : OAI22_X1 port map( A1 => n25129, A2 => n25397, B1 => n879, B2 => 
                           n25125, ZN => n6229);
   U23276 : OAI22_X1 port map( A1 => n25129, A2 => n25400, B1 => n878, B2 => 
                           n25125, ZN => n6230);
   U23277 : OAI22_X1 port map( A1 => n25129, A2 => n25403, B1 => n877, B2 => 
                           n25125, ZN => n6231);
   U23278 : OAI22_X1 port map( A1 => n25130, A2 => n25406, B1 => n876, B2 => 
                           n25125, ZN => n6232);
   U23279 : OAI22_X1 port map( A1 => n25130, A2 => n25409, B1 => n875, B2 => 
                           n25125, ZN => n6233);
   U23280 : OAI22_X1 port map( A1 => n25130, A2 => n25412, B1 => n874, B2 => 
                           n25125, ZN => n6234);
   U23281 : OAI22_X1 port map( A1 => n25130, A2 => n25415, B1 => n873, B2 => 
                           n25125, ZN => n6235);
   U23282 : OAI22_X1 port map( A1 => n25160, A2 => n25345, B1 => n9244, B2 => 
                           n25158, ZN => n6340);
   U23283 : OAI22_X1 port map( A1 => n25160, A2 => n25348, B1 => n9242, B2 => 
                           n25158, ZN => n6341);
   U23284 : OAI22_X1 port map( A1 => n25160, A2 => n25351, B1 => n9240, B2 => 
                           n25158, ZN => n6342);
   U23285 : OAI22_X1 port map( A1 => n25160, A2 => n25354, B1 => n9238, B2 => 
                           n25158, ZN => n6343);
   U23286 : OAI22_X1 port map( A1 => n25160, A2 => n25357, B1 => n9236, B2 => 
                           n25158, ZN => n6344);
   U23287 : OAI22_X1 port map( A1 => n25161, A2 => n25360, B1 => n9234, B2 => 
                           n25158, ZN => n6345);
   U23288 : OAI22_X1 port map( A1 => n25161, A2 => n25363, B1 => n9232, B2 => 
                           n25158, ZN => n6346);
   U23289 : OAI22_X1 port map( A1 => n25161, A2 => n25366, B1 => n9230, B2 => 
                           n25158, ZN => n6347);
   U23290 : OAI22_X1 port map( A1 => n25161, A2 => n25369, B1 => n9228, B2 => 
                           n25158, ZN => n6348);
   U23291 : OAI22_X1 port map( A1 => n25161, A2 => n25372, B1 => n9226, B2 => 
                           n25158, ZN => n6349);
   U23292 : OAI22_X1 port map( A1 => n25162, A2 => n25375, B1 => n9224, B2 => 
                           n25158, ZN => n6350);
   U23293 : OAI22_X1 port map( A1 => n25162, A2 => n25378, B1 => n9222, B2 => 
                           n25158, ZN => n6351);
   U23294 : OAI22_X1 port map( A1 => n25162, A2 => n25381, B1 => n9220, B2 => 
                           n25159, ZN => n6352);
   U23295 : OAI22_X1 port map( A1 => n25162, A2 => n25384, B1 => n9218, B2 => 
                           n25159, ZN => n6353);
   U23296 : OAI22_X1 port map( A1 => n25162, A2 => n25387, B1 => n9216, B2 => 
                           n25159, ZN => n6354);
   U23297 : OAI22_X1 port map( A1 => n25163, A2 => n25390, B1 => n9214, B2 => 
                           n25159, ZN => n6355);
   U23298 : OAI22_X1 port map( A1 => n25163, A2 => n25393, B1 => n9212, B2 => 
                           n25159, ZN => n6356);
   U23299 : OAI22_X1 port map( A1 => n25163, A2 => n25396, B1 => n9210, B2 => 
                           n25159, ZN => n6357);
   U23300 : OAI22_X1 port map( A1 => n25163, A2 => n25399, B1 => n9208, B2 => 
                           n25159, ZN => n6358);
   U23301 : OAI22_X1 port map( A1 => n25163, A2 => n25402, B1 => n9206, B2 => 
                           n25159, ZN => n6359);
   U23302 : OAI22_X1 port map( A1 => n25164, A2 => n25405, B1 => n9204, B2 => 
                           n25159, ZN => n6360);
   U23303 : OAI22_X1 port map( A1 => n25164, A2 => n25408, B1 => n9202, B2 => 
                           n25159, ZN => n6361);
   U23304 : OAI22_X1 port map( A1 => n25164, A2 => n25411, B1 => n9200, B2 => 
                           n25159, ZN => n6362);
   U23305 : OAI22_X1 port map( A1 => n25164, A2 => n25414, B1 => n9198, B2 => 
                           n25159, ZN => n6363);
   U23306 : OAI22_X1 port map( A1 => n25335, A2 => n25432, B1 => n99, B2 => 
                           n21255, ZN => n7009);
   U23307 : OAI22_X1 port map( A1 => n25336, A2 => n25435, B1 => n98, B2 => 
                           n25327, ZN => n7010);
   U23308 : OAI22_X1 port map( A1 => n25336, A2 => n25438, B1 => n97, B2 => 
                           n21255, ZN => n7011);
   U23309 : OAI22_X1 port map( A1 => n25336, A2 => n25441, B1 => n96, B2 => 
                           n25327, ZN => n7012);
   U23310 : OAI22_X1 port map( A1 => n25336, A2 => n25444, B1 => n95, B2 => 
                           n21255, ZN => n7013);
   U23311 : OAI22_X1 port map( A1 => n25336, A2 => n25447, B1 => n94, B2 => 
                           n25327, ZN => n7014);
   U23312 : OAI22_X1 port map( A1 => n25337, A2 => n25453, B1 => n92, B2 => 
                           n21255, ZN => n7016);
   U23313 : OAI22_X1 port map( A1 => n25337, A2 => n25456, B1 => n91, B2 => 
                           n25327, ZN => n7017);
   U23314 : OAI22_X1 port map( A1 => n25337, A2 => n25459, B1 => n90, B2 => 
                           n25327, ZN => n7018);
   U23315 : OAI22_X1 port map( A1 => n25338, A2 => n25465, B1 => n88, B2 => 
                           n25327, ZN => n7020);
   U23316 : OAI22_X1 port map( A1 => n25338, A2 => n25471, B1 => n86, B2 => 
                           n25329, ZN => n7022);
   U23317 : OAI22_X1 port map( A1 => n25096, A2 => n25418, B1 => n7378, B2 => 
                           n25090, ZN => n6108);
   U23318 : OAI22_X1 port map( A1 => n25097, A2 => n25421, B1 => n7376, B2 => 
                           n25091, ZN => n6109);
   U23319 : OAI22_X1 port map( A1 => n25097, A2 => n25424, B1 => n7374, B2 => 
                           n25089, ZN => n6110);
   U23320 : OAI22_X1 port map( A1 => n25097, A2 => n25427, B1 => n7372, B2 => 
                           n25090, ZN => n6111);
   U23321 : OAI22_X1 port map( A1 => n25097, A2 => n25430, B1 => n7370, B2 => 
                           n25091, ZN => n6112);
   U23322 : OAI22_X1 port map( A1 => n25097, A2 => n25433, B1 => n7368, B2 => 
                           n25089, ZN => n6113);
   U23323 : OAI22_X1 port map( A1 => n25098, A2 => n25436, B1 => n7366, B2 => 
                           n25090, ZN => n6114);
   U23324 : OAI22_X1 port map( A1 => n25098, A2 => n25439, B1 => n7364, B2 => 
                           n25091, ZN => n6115);
   U23325 : OAI22_X1 port map( A1 => n25098, A2 => n25442, B1 => n7362, B2 => 
                           n25089, ZN => n6116);
   U23326 : OAI22_X1 port map( A1 => n25098, A2 => n25445, B1 => n7360, B2 => 
                           n25090, ZN => n6117);
   U23327 : OAI22_X1 port map( A1 => n25098, A2 => n25448, B1 => n7358, B2 => 
                           n25091, ZN => n6118);
   U23328 : OAI22_X1 port map( A1 => n25099, A2 => n25451, B1 => n7356, B2 => 
                           n25089, ZN => n6119);
   U23329 : OAI22_X1 port map( A1 => n25099, A2 => n25454, B1 => n7354, B2 => 
                           n21278, ZN => n6120);
   U23330 : OAI22_X1 port map( A1 => n25099, A2 => n25457, B1 => n7352, B2 => 
                           n25089, ZN => n6121);
   U23331 : OAI22_X1 port map( A1 => n25099, A2 => n25460, B1 => n7350, B2 => 
                           n21278, ZN => n6122);
   U23332 : OAI22_X1 port map( A1 => n25099, A2 => n25463, B1 => n7348, B2 => 
                           n25089, ZN => n6123);
   U23333 : OAI22_X1 port map( A1 => n25100, A2 => n25466, B1 => n7346, B2 => 
                           n21278, ZN => n6124);
   U23334 : OAI22_X1 port map( A1 => n25100, A2 => n25469, B1 => n7344, B2 => 
                           n25089, ZN => n6125);
   U23335 : OAI22_X1 port map( A1 => n25100, A2 => n25472, B1 => n7342, B2 => 
                           n25090, ZN => n6126);
   U23336 : OAI22_X1 port map( A1 => n25100, A2 => n25475, B1 => n7340, B2 => 
                           n25091, ZN => n6127);
   U23337 : OAI22_X1 port map( A1 => n25100, A2 => n25478, B1 => n7338, B2 => 
                           n25089, ZN => n6128);
   U23338 : OAI22_X1 port map( A1 => n25101, A2 => n25481, B1 => n7336, B2 => 
                           n25089, ZN => n6129);
   U23339 : OAI22_X1 port map( A1 => n25101, A2 => n25484, B1 => n7334, B2 => 
                           n25090, ZN => n6130);
   U23340 : OAI22_X1 port map( A1 => n25101, A2 => n25487, B1 => n7332, B2 => 
                           n25091, ZN => n6131);
   U23341 : OAI22_X1 port map( A1 => n25101, A2 => n25490, B1 => n7330, B2 => 
                           n25089, ZN => n6132);
   U23342 : OAI22_X1 port map( A1 => n25101, A2 => n25493, B1 => n7328, B2 => 
                           n25089, ZN => n6133);
   U23343 : OAI22_X1 port map( A1 => n25102, A2 => n25496, B1 => n7326, B2 => 
                           n21278, ZN => n6134);
   U23344 : OAI22_X1 port map( A1 => n25102, A2 => n25499, B1 => n7324, B2 => 
                           n25089, ZN => n6135);
   U23345 : OAI22_X1 port map( A1 => n25102, A2 => n25502, B1 => n7322, B2 => 
                           n21278, ZN => n6136);
   U23346 : OAI22_X1 port map( A1 => n25102, A2 => n25505, B1 => n7320, B2 => 
                           n25089, ZN => n6137);
   U23347 : OAI22_X1 port map( A1 => n25102, A2 => n25508, B1 => n7318, B2 => 
                           n21278, ZN => n6138);
   U23348 : OAI22_X1 port map( A1 => n25103, A2 => n25511, B1 => n7316, B2 => 
                           n25089, ZN => n6139);
   U23349 : OAI22_X1 port map( A1 => n25103, A2 => n25514, B1 => n7314, B2 => 
                           n21278, ZN => n6140);
   U23350 : OAI22_X1 port map( A1 => n25103, A2 => n25517, B1 => n7312, B2 => 
                           n25089, ZN => n6141);
   U23351 : OAI22_X1 port map( A1 => n25103, A2 => n25520, B1 => n7310, B2 => 
                           n21278, ZN => n6142);
   U23352 : OAI22_X1 port map( A1 => n25103, A2 => n25523, B1 => n7308, B2 => 
                           n25089, ZN => n6143);
   U23353 : OAI22_X1 port map( A1 => n25104, A2 => n25526, B1 => n7306, B2 => 
                           n21278, ZN => n6144);
   U23354 : OAI22_X1 port map( A1 => n25104, A2 => n25529, B1 => n7304, B2 => 
                           n21278, ZN => n6145);
   U23355 : OAI22_X1 port map( A1 => n25104, A2 => n25532, B1 => n7302, B2 => 
                           n25089, ZN => n6146);
   U23356 : OAI22_X1 port map( A1 => n25104, A2 => n25552, B1 => n7300, B2 => 
                           n21278, ZN => n6147);
   U23357 : OAI22_X1 port map( A1 => n25266, A2 => n25417, B1 => n17338, B2 => 
                           n25260, ZN => n6748);
   U23358 : OAI22_X1 port map( A1 => n25267, A2 => n25420, B1 => n17335, B2 => 
                           n25261, ZN => n6749);
   U23359 : OAI22_X1 port map( A1 => n25267, A2 => n25423, B1 => n17332, B2 => 
                           n25259, ZN => n6750);
   U23360 : OAI22_X1 port map( A1 => n25267, A2 => n25426, B1 => n17329, B2 => 
                           n25260, ZN => n6751);
   U23361 : OAI22_X1 port map( A1 => n25267, A2 => n25429, B1 => n17326, B2 => 
                           n25261, ZN => n6752);
   U23362 : OAI22_X1 port map( A1 => n25267, A2 => n25432, B1 => n17323, B2 => 
                           n25259, ZN => n6753);
   U23363 : OAI22_X1 port map( A1 => n25268, A2 => n25435, B1 => n17320, B2 => 
                           n25260, ZN => n6754);
   U23364 : OAI22_X1 port map( A1 => n25268, A2 => n25438, B1 => n17317, B2 => 
                           n25261, ZN => n6755);
   U23365 : OAI22_X1 port map( A1 => n25268, A2 => n25441, B1 => n17314, B2 => 
                           n25259, ZN => n6756);
   U23366 : OAI22_X1 port map( A1 => n25268, A2 => n25444, B1 => n17311, B2 => 
                           n25260, ZN => n6757);
   U23367 : OAI22_X1 port map( A1 => n25268, A2 => n25447, B1 => n17308, B2 => 
                           n25261, ZN => n6758);
   U23368 : OAI22_X1 port map( A1 => n25269, A2 => n25450, B1 => n17305, B2 => 
                           n25259, ZN => n6759);
   U23369 : OAI22_X1 port map( A1 => n25269, A2 => n25453, B1 => n17302, B2 => 
                           n21263, ZN => n6760);
   U23370 : OAI22_X1 port map( A1 => n25269, A2 => n25456, B1 => n17299, B2 => 
                           n25259, ZN => n6761);
   U23371 : OAI22_X1 port map( A1 => n25269, A2 => n25459, B1 => n17296, B2 => 
                           n21263, ZN => n6762);
   U23372 : OAI22_X1 port map( A1 => n25269, A2 => n25462, B1 => n17293, B2 => 
                           n25259, ZN => n6763);
   U23373 : OAI22_X1 port map( A1 => n25270, A2 => n25465, B1 => n17290, B2 => 
                           n21263, ZN => n6764);
   U23374 : OAI22_X1 port map( A1 => n25270, A2 => n25468, B1 => n17287, B2 => 
                           n25259, ZN => n6765);
   U23375 : OAI22_X1 port map( A1 => n25270, A2 => n25471, B1 => n17284, B2 => 
                           n25260, ZN => n6766);
   U23376 : OAI22_X1 port map( A1 => n25270, A2 => n25474, B1 => n17281, B2 => 
                           n25261, ZN => n6767);
   U23377 : OAI22_X1 port map( A1 => n25270, A2 => n25477, B1 => n17278, B2 => 
                           n25259, ZN => n6768);
   U23378 : OAI22_X1 port map( A1 => n25271, A2 => n25480, B1 => n17275, B2 => 
                           n25259, ZN => n6769);
   U23379 : OAI22_X1 port map( A1 => n25271, A2 => n25483, B1 => n17272, B2 => 
                           n25260, ZN => n6770);
   U23380 : OAI22_X1 port map( A1 => n25271, A2 => n25486, B1 => n17269, B2 => 
                           n25261, ZN => n6771);
   U23381 : OAI22_X1 port map( A1 => n25271, A2 => n25489, B1 => n17266, B2 => 
                           n25259, ZN => n6772);
   U23382 : OAI22_X1 port map( A1 => n25271, A2 => n25492, B1 => n17263, B2 => 
                           n25259, ZN => n6773);
   U23383 : OAI22_X1 port map( A1 => n25272, A2 => n25495, B1 => n17260, B2 => 
                           n21263, ZN => n6774);
   U23384 : OAI22_X1 port map( A1 => n25272, A2 => n25498, B1 => n17257, B2 => 
                           n25259, ZN => n6775);
   U23385 : OAI22_X1 port map( A1 => n25272, A2 => n25501, B1 => n17254, B2 => 
                           n21263, ZN => n6776);
   U23386 : OAI22_X1 port map( A1 => n25272, A2 => n25504, B1 => n17251, B2 => 
                           n25259, ZN => n6777);
   U23387 : OAI22_X1 port map( A1 => n25272, A2 => n25507, B1 => n17248, B2 => 
                           n21263, ZN => n6778);
   U23388 : OAI22_X1 port map( A1 => n25273, A2 => n25510, B1 => n17245, B2 => 
                           n25259, ZN => n6779);
   U23389 : OAI22_X1 port map( A1 => n25273, A2 => n25513, B1 => n17242, B2 => 
                           n21263, ZN => n6780);
   U23390 : OAI22_X1 port map( A1 => n25273, A2 => n25516, B1 => n17239, B2 => 
                           n25259, ZN => n6781);
   U23391 : OAI22_X1 port map( A1 => n25273, A2 => n25519, B1 => n17236, B2 => 
                           n21263, ZN => n6782);
   U23392 : OAI22_X1 port map( A1 => n25273, A2 => n25522, B1 => n17233, B2 => 
                           n25259, ZN => n6783);
   U23393 : OAI22_X1 port map( A1 => n25181, A2 => n25417, B1 => n7506, B2 => 
                           n25175, ZN => n6428);
   U23394 : OAI22_X1 port map( A1 => n25182, A2 => n25420, B1 => n7504, B2 => 
                           n25176, ZN => n6429);
   U23395 : OAI22_X1 port map( A1 => n25182, A2 => n25423, B1 => n7502, B2 => 
                           n25174, ZN => n6430);
   U23396 : OAI22_X1 port map( A1 => n25182, A2 => n25426, B1 => n7500, B2 => 
                           n25175, ZN => n6431);
   U23397 : OAI22_X1 port map( A1 => n25182, A2 => n25429, B1 => n7498, B2 => 
                           n25176, ZN => n6432);
   U23398 : OAI22_X1 port map( A1 => n25182, A2 => n25432, B1 => n7496, B2 => 
                           n25174, ZN => n6433);
   U23399 : OAI22_X1 port map( A1 => n25183, A2 => n25435, B1 => n7494, B2 => 
                           n25175, ZN => n6434);
   U23400 : OAI22_X1 port map( A1 => n25183, A2 => n25438, B1 => n7492, B2 => 
                           n25176, ZN => n6435);
   U23401 : OAI22_X1 port map( A1 => n25183, A2 => n25441, B1 => n7490, B2 => 
                           n25174, ZN => n6436);
   U23402 : OAI22_X1 port map( A1 => n25183, A2 => n25444, B1 => n7488, B2 => 
                           n25175, ZN => n6437);
   U23403 : OAI22_X1 port map( A1 => n25183, A2 => n25447, B1 => n7486, B2 => 
                           n25176, ZN => n6438);
   U23404 : OAI22_X1 port map( A1 => n25184, A2 => n25450, B1 => n7484, B2 => 
                           n25174, ZN => n6439);
   U23405 : OAI22_X1 port map( A1 => n25184, A2 => n25453, B1 => n7482, B2 => 
                           n21273, ZN => n6440);
   U23406 : OAI22_X1 port map( A1 => n25184, A2 => n25456, B1 => n7480, B2 => 
                           n25174, ZN => n6441);
   U23407 : OAI22_X1 port map( A1 => n25184, A2 => n25459, B1 => n7478, B2 => 
                           n21273, ZN => n6442);
   U23408 : OAI22_X1 port map( A1 => n25184, A2 => n25462, B1 => n7476, B2 => 
                           n25174, ZN => n6443);
   U23409 : OAI22_X1 port map( A1 => n25185, A2 => n25465, B1 => n7474, B2 => 
                           n21273, ZN => n6444);
   U23410 : OAI22_X1 port map( A1 => n25185, A2 => n25468, B1 => n7472, B2 => 
                           n25174, ZN => n6445);
   U23411 : OAI22_X1 port map( A1 => n25185, A2 => n25471, B1 => n7470, B2 => 
                           n25175, ZN => n6446);
   U23412 : OAI22_X1 port map( A1 => n25185, A2 => n25474, B1 => n7468, B2 => 
                           n25176, ZN => n6447);
   U23413 : OAI22_X1 port map( A1 => n25185, A2 => n25477, B1 => n7466, B2 => 
                           n25174, ZN => n6448);
   U23414 : OAI22_X1 port map( A1 => n25186, A2 => n25480, B1 => n7464, B2 => 
                           n25174, ZN => n6449);
   U23415 : OAI22_X1 port map( A1 => n25186, A2 => n25483, B1 => n7462, B2 => 
                           n25175, ZN => n6450);
   U23416 : OAI22_X1 port map( A1 => n25186, A2 => n25486, B1 => n7460, B2 => 
                           n25176, ZN => n6451);
   U23417 : OAI22_X1 port map( A1 => n25186, A2 => n25489, B1 => n7458, B2 => 
                           n25174, ZN => n6452);
   U23418 : OAI22_X1 port map( A1 => n25186, A2 => n25492, B1 => n7456, B2 => 
                           n25174, ZN => n6453);
   U23419 : OAI22_X1 port map( A1 => n25187, A2 => n25495, B1 => n7454, B2 => 
                           n21273, ZN => n6454);
   U23420 : OAI22_X1 port map( A1 => n25187, A2 => n25498, B1 => n7452, B2 => 
                           n25174, ZN => n6455);
   U23421 : OAI22_X1 port map( A1 => n25187, A2 => n25501, B1 => n7450, B2 => 
                           n21273, ZN => n6456);
   U23422 : OAI22_X1 port map( A1 => n25187, A2 => n25504, B1 => n7448, B2 => 
                           n25174, ZN => n6457);
   U23423 : OAI22_X1 port map( A1 => n25187, A2 => n25507, B1 => n7446, B2 => 
                           n21273, ZN => n6458);
   U23424 : OAI22_X1 port map( A1 => n25188, A2 => n25510, B1 => n7444, B2 => 
                           n25174, ZN => n6459);
   U23425 : OAI22_X1 port map( A1 => n25188, A2 => n25513, B1 => n7442, B2 => 
                           n21273, ZN => n6460);
   U23426 : OAI22_X1 port map( A1 => n25188, A2 => n25516, B1 => n7440, B2 => 
                           n25174, ZN => n6461);
   U23427 : OAI22_X1 port map( A1 => n25188, A2 => n25519, B1 => n7438, B2 => 
                           n21273, ZN => n6462);
   U23428 : OAI22_X1 port map( A1 => n25188, A2 => n25522, B1 => n7436, B2 => 
                           n25174, ZN => n6463);
   U23429 : OAI22_X1 port map( A1 => n25045, A2 => n25418, B1 => n8813, B2 => 
                           n25039, ZN => n5916);
   U23430 : OAI22_X1 port map( A1 => n25046, A2 => n25421, B1 => n8811, B2 => 
                           n25040, ZN => n5917);
   U23431 : OAI22_X1 port map( A1 => n25046, A2 => n25424, B1 => n8809, B2 => 
                           n25038, ZN => n5918);
   U23432 : OAI22_X1 port map( A1 => n25046, A2 => n25427, B1 => n8807, B2 => 
                           n25039, ZN => n5919);
   U23433 : OAI22_X1 port map( A1 => n25046, A2 => n25430, B1 => n8805, B2 => 
                           n25040, ZN => n5920);
   U23434 : OAI22_X1 port map( A1 => n25046, A2 => n25433, B1 => n8803, B2 => 
                           n25038, ZN => n5921);
   U23435 : OAI22_X1 port map( A1 => n25047, A2 => n25436, B1 => n8801, B2 => 
                           n25039, ZN => n5922);
   U23436 : OAI22_X1 port map( A1 => n25047, A2 => n25439, B1 => n8799, B2 => 
                           n25040, ZN => n5923);
   U23437 : OAI22_X1 port map( A1 => n25047, A2 => n25442, B1 => n8797, B2 => 
                           n25038, ZN => n5924);
   U23438 : OAI22_X1 port map( A1 => n25047, A2 => n25445, B1 => n8795, B2 => 
                           n25039, ZN => n5925);
   U23439 : OAI22_X1 port map( A1 => n25047, A2 => n25448, B1 => n8793, B2 => 
                           n25040, ZN => n5926);
   U23440 : OAI22_X1 port map( A1 => n25048, A2 => n25451, B1 => n8791, B2 => 
                           n25038, ZN => n5927);
   U23441 : OAI22_X1 port map( A1 => n25048, A2 => n25454, B1 => n8789, B2 => 
                           n21282, ZN => n5928);
   U23442 : OAI22_X1 port map( A1 => n25048, A2 => n25457, B1 => n8787, B2 => 
                           n25038, ZN => n5929);
   U23443 : OAI22_X1 port map( A1 => n25048, A2 => n25460, B1 => n8785, B2 => 
                           n21282, ZN => n5930);
   U23444 : OAI22_X1 port map( A1 => n25048, A2 => n25463, B1 => n8783, B2 => 
                           n25038, ZN => n5931);
   U23445 : OAI22_X1 port map( A1 => n25049, A2 => n25466, B1 => n8781, B2 => 
                           n21282, ZN => n5932);
   U23446 : OAI22_X1 port map( A1 => n25049, A2 => n25469, B1 => n8779, B2 => 
                           n25038, ZN => n5933);
   U23447 : OAI22_X1 port map( A1 => n25049, A2 => n25472, B1 => n8777, B2 => 
                           n25039, ZN => n5934);
   U23448 : OAI22_X1 port map( A1 => n25049, A2 => n25475, B1 => n8775, B2 => 
                           n25040, ZN => n5935);
   U23449 : OAI22_X1 port map( A1 => n25049, A2 => n25478, B1 => n8773, B2 => 
                           n25038, ZN => n5936);
   U23450 : OAI22_X1 port map( A1 => n25050, A2 => n25481, B1 => n8771, B2 => 
                           n25038, ZN => n5937);
   U23451 : OAI22_X1 port map( A1 => n25050, A2 => n25484, B1 => n8769, B2 => 
                           n25039, ZN => n5938);
   U23452 : OAI22_X1 port map( A1 => n25050, A2 => n25487, B1 => n8767, B2 => 
                           n25040, ZN => n5939);
   U23453 : OAI22_X1 port map( A1 => n25050, A2 => n25490, B1 => n8765, B2 => 
                           n25038, ZN => n5940);
   U23454 : OAI22_X1 port map( A1 => n25050, A2 => n25493, B1 => n8763, B2 => 
                           n25038, ZN => n5941);
   U23455 : OAI22_X1 port map( A1 => n25051, A2 => n25496, B1 => n8761, B2 => 
                           n21282, ZN => n5942);
   U23456 : OAI22_X1 port map( A1 => n25051, A2 => n25499, B1 => n8759, B2 => 
                           n25038, ZN => n5943);
   U23457 : OAI22_X1 port map( A1 => n25051, A2 => n25502, B1 => n8757, B2 => 
                           n21282, ZN => n5944);
   U23458 : OAI22_X1 port map( A1 => n25051, A2 => n25505, B1 => n8755, B2 => 
                           n25038, ZN => n5945);
   U23459 : OAI22_X1 port map( A1 => n25051, A2 => n25508, B1 => n8753, B2 => 
                           n21282, ZN => n5946);
   U23460 : OAI22_X1 port map( A1 => n25052, A2 => n25511, B1 => n8751, B2 => 
                           n25038, ZN => n5947);
   U23461 : OAI22_X1 port map( A1 => n25052, A2 => n25514, B1 => n8749, B2 => 
                           n21282, ZN => n5948);
   U23462 : OAI22_X1 port map( A1 => n25052, A2 => n25517, B1 => n8747, B2 => 
                           n25038, ZN => n5949);
   U23463 : OAI22_X1 port map( A1 => n25052, A2 => n25520, B1 => n8745, B2 => 
                           n21282, ZN => n5950);
   U23464 : OAI22_X1 port map( A1 => n25052, A2 => n25523, B1 => n8743, B2 => 
                           n25038, ZN => n5951);
   U23465 : OAI22_X1 port map( A1 => n25028, A2 => n25418, B1 => n8941, B2 => 
                           n25022, ZN => n5852);
   U23466 : OAI22_X1 port map( A1 => n25029, A2 => n25421, B1 => n8939, B2 => 
                           n25023, ZN => n5853);
   U23467 : OAI22_X1 port map( A1 => n25029, A2 => n25424, B1 => n8937, B2 => 
                           n25021, ZN => n5854);
   U23468 : OAI22_X1 port map( A1 => n25029, A2 => n25427, B1 => n8935, B2 => 
                           n25022, ZN => n5855);
   U23469 : OAI22_X1 port map( A1 => n25029, A2 => n25430, B1 => n8933, B2 => 
                           n25023, ZN => n5856);
   U23470 : OAI22_X1 port map( A1 => n25029, A2 => n25433, B1 => n8931, B2 => 
                           n25021, ZN => n5857);
   U23471 : OAI22_X1 port map( A1 => n25030, A2 => n25436, B1 => n8929, B2 => 
                           n25022, ZN => n5858);
   U23472 : OAI22_X1 port map( A1 => n25030, A2 => n25439, B1 => n8927, B2 => 
                           n25023, ZN => n5859);
   U23473 : OAI22_X1 port map( A1 => n25030, A2 => n25442, B1 => n8925, B2 => 
                           n25021, ZN => n5860);
   U23474 : OAI22_X1 port map( A1 => n25030, A2 => n25445, B1 => n8923, B2 => 
                           n25022, ZN => n5861);
   U23475 : OAI22_X1 port map( A1 => n25030, A2 => n25448, B1 => n8921, B2 => 
                           n25023, ZN => n5862);
   U23476 : OAI22_X1 port map( A1 => n25031, A2 => n25451, B1 => n8919, B2 => 
                           n25021, ZN => n5863);
   U23477 : OAI22_X1 port map( A1 => n25031, A2 => n25454, B1 => n8917, B2 => 
                           n21283, ZN => n5864);
   U23478 : OAI22_X1 port map( A1 => n25031, A2 => n25457, B1 => n8915, B2 => 
                           n25021, ZN => n5865);
   U23479 : OAI22_X1 port map( A1 => n25031, A2 => n25460, B1 => n8913, B2 => 
                           n21283, ZN => n5866);
   U23480 : OAI22_X1 port map( A1 => n25031, A2 => n25463, B1 => n8911, B2 => 
                           n25021, ZN => n5867);
   U23481 : OAI22_X1 port map( A1 => n25032, A2 => n25466, B1 => n8909, B2 => 
                           n21283, ZN => n5868);
   U23482 : OAI22_X1 port map( A1 => n25032, A2 => n25469, B1 => n8907, B2 => 
                           n25021, ZN => n5869);
   U23483 : OAI22_X1 port map( A1 => n25032, A2 => n25472, B1 => n8905, B2 => 
                           n25022, ZN => n5870);
   U23484 : OAI22_X1 port map( A1 => n25032, A2 => n25475, B1 => n8903, B2 => 
                           n25023, ZN => n5871);
   U23485 : OAI22_X1 port map( A1 => n25032, A2 => n25478, B1 => n8901, B2 => 
                           n25021, ZN => n5872);
   U23486 : OAI22_X1 port map( A1 => n25033, A2 => n25481, B1 => n8899, B2 => 
                           n25021, ZN => n5873);
   U23487 : OAI22_X1 port map( A1 => n25033, A2 => n25484, B1 => n8897, B2 => 
                           n25022, ZN => n5874);
   U23488 : OAI22_X1 port map( A1 => n25033, A2 => n25487, B1 => n8895, B2 => 
                           n25023, ZN => n5875);
   U23489 : OAI22_X1 port map( A1 => n25033, A2 => n25490, B1 => n8893, B2 => 
                           n25021, ZN => n5876);
   U23490 : OAI22_X1 port map( A1 => n25033, A2 => n25493, B1 => n8891, B2 => 
                           n25021, ZN => n5877);
   U23491 : OAI22_X1 port map( A1 => n25034, A2 => n25496, B1 => n8889, B2 => 
                           n21283, ZN => n5878);
   U23492 : OAI22_X1 port map( A1 => n25034, A2 => n25499, B1 => n8887, B2 => 
                           n25021, ZN => n5879);
   U23493 : OAI22_X1 port map( A1 => n25034, A2 => n25502, B1 => n8885, B2 => 
                           n21283, ZN => n5880);
   U23494 : OAI22_X1 port map( A1 => n25034, A2 => n25505, B1 => n8883, B2 => 
                           n25021, ZN => n5881);
   U23495 : OAI22_X1 port map( A1 => n25034, A2 => n25508, B1 => n8881, B2 => 
                           n21283, ZN => n5882);
   U23496 : OAI22_X1 port map( A1 => n25035, A2 => n25511, B1 => n8879, B2 => 
                           n25021, ZN => n5883);
   U23497 : OAI22_X1 port map( A1 => n25035, A2 => n25514, B1 => n8877, B2 => 
                           n21283, ZN => n5884);
   U23498 : OAI22_X1 port map( A1 => n25035, A2 => n25517, B1 => n8875, B2 => 
                           n25021, ZN => n5885);
   U23499 : OAI22_X1 port map( A1 => n25035, A2 => n25520, B1 => n8873, B2 => 
                           n21283, ZN => n5886);
   U23500 : OAI22_X1 port map( A1 => n25035, A2 => n25523, B1 => n8871, B2 => 
                           n25021, ZN => n5887);
   U23501 : OAI22_X1 port map( A1 => n24858, A2 => n25419, B1 => n8940, B2 => 
                           n24852, ZN => n5212);
   U23502 : OAI22_X1 port map( A1 => n24859, A2 => n25422, B1 => n8938, B2 => 
                           n24853, ZN => n5213);
   U23503 : OAI22_X1 port map( A1 => n24859, A2 => n25425, B1 => n8936, B2 => 
                           n24851, ZN => n5214);
   U23504 : OAI22_X1 port map( A1 => n24859, A2 => n25428, B1 => n8934, B2 => 
                           n24852, ZN => n5215);
   U23505 : OAI22_X1 port map( A1 => n24859, A2 => n25431, B1 => n8932, B2 => 
                           n24853, ZN => n5216);
   U23506 : OAI22_X1 port map( A1 => n24859, A2 => n25434, B1 => n8930, B2 => 
                           n24851, ZN => n5217);
   U23507 : OAI22_X1 port map( A1 => n24860, A2 => n25437, B1 => n8928, B2 => 
                           n24852, ZN => n5218);
   U23508 : OAI22_X1 port map( A1 => n24860, A2 => n25440, B1 => n8926, B2 => 
                           n24853, ZN => n5219);
   U23509 : OAI22_X1 port map( A1 => n24860, A2 => n25443, B1 => n8924, B2 => 
                           n24851, ZN => n5220);
   U23510 : OAI22_X1 port map( A1 => n24860, A2 => n25446, B1 => n8922, B2 => 
                           n24852, ZN => n5221);
   U23511 : OAI22_X1 port map( A1 => n24860, A2 => n25449, B1 => n8920, B2 => 
                           n24853, ZN => n5222);
   U23512 : OAI22_X1 port map( A1 => n24861, A2 => n25452, B1 => n8918, B2 => 
                           n24851, ZN => n5223);
   U23513 : OAI22_X1 port map( A1 => n24861, A2 => n25455, B1 => n8916, B2 => 
                           n21294, ZN => n5224);
   U23514 : OAI22_X1 port map( A1 => n24861, A2 => n25458, B1 => n8914, B2 => 
                           n24851, ZN => n5225);
   U23515 : OAI22_X1 port map( A1 => n24861, A2 => n25461, B1 => n8912, B2 => 
                           n21294, ZN => n5226);
   U23516 : OAI22_X1 port map( A1 => n24861, A2 => n25464, B1 => n8910, B2 => 
                           n24851, ZN => n5227);
   U23517 : OAI22_X1 port map( A1 => n24862, A2 => n25467, B1 => n8908, B2 => 
                           n21294, ZN => n5228);
   U23518 : OAI22_X1 port map( A1 => n24862, A2 => n25470, B1 => n8906, B2 => 
                           n24851, ZN => n5229);
   U23519 : OAI22_X1 port map( A1 => n24862, A2 => n25473, B1 => n8904, B2 => 
                           n24852, ZN => n5230);
   U23520 : OAI22_X1 port map( A1 => n24862, A2 => n25476, B1 => n8902, B2 => 
                           n24853, ZN => n5231);
   U23521 : OAI22_X1 port map( A1 => n24862, A2 => n25479, B1 => n8900, B2 => 
                           n24851, ZN => n5232);
   U23522 : OAI22_X1 port map( A1 => n24863, A2 => n25482, B1 => n8898, B2 => 
                           n24851, ZN => n5233);
   U23523 : OAI22_X1 port map( A1 => n24863, A2 => n25485, B1 => n8896, B2 => 
                           n24852, ZN => n5234);
   U23524 : OAI22_X1 port map( A1 => n24863, A2 => n25488, B1 => n8894, B2 => 
                           n24853, ZN => n5235);
   U23525 : OAI22_X1 port map( A1 => n24863, A2 => n25491, B1 => n8892, B2 => 
                           n24851, ZN => n5236);
   U23526 : OAI22_X1 port map( A1 => n24863, A2 => n25494, B1 => n8890, B2 => 
                           n24851, ZN => n5237);
   U23527 : OAI22_X1 port map( A1 => n24864, A2 => n25497, B1 => n8888, B2 => 
                           n21294, ZN => n5238);
   U23528 : OAI22_X1 port map( A1 => n24864, A2 => n25500, B1 => n8886, B2 => 
                           n24851, ZN => n5239);
   U23529 : OAI22_X1 port map( A1 => n24864, A2 => n25503, B1 => n8884, B2 => 
                           n21294, ZN => n5240);
   U23530 : OAI22_X1 port map( A1 => n24864, A2 => n25506, B1 => n8882, B2 => 
                           n24851, ZN => n5241);
   U23531 : OAI22_X1 port map( A1 => n24864, A2 => n25509, B1 => n8880, B2 => 
                           n21294, ZN => n5242);
   U23532 : OAI22_X1 port map( A1 => n24865, A2 => n25512, B1 => n8878, B2 => 
                           n24851, ZN => n5243);
   U23533 : OAI22_X1 port map( A1 => n24865, A2 => n25515, B1 => n8876, B2 => 
                           n21294, ZN => n5244);
   U23534 : OAI22_X1 port map( A1 => n24865, A2 => n25518, B1 => n8874, B2 => 
                           n24851, ZN => n5245);
   U23535 : OAI22_X1 port map( A1 => n24865, A2 => n25521, B1 => n8872, B2 => 
                           n21294, ZN => n5246);
   U23536 : OAI22_X1 port map( A1 => n24865, A2 => n25524, B1 => n8870, B2 => 
                           n24851, ZN => n5247);
   U23537 : OAI22_X1 port map( A1 => n24926, A2 => n25419, B1 => n7379, B2 => 
                           n24920, ZN => n5468);
   U23538 : OAI22_X1 port map( A1 => n24927, A2 => n25422, B1 => n7377, B2 => 
                           n24921, ZN => n5469);
   U23539 : OAI22_X1 port map( A1 => n24927, A2 => n25425, B1 => n7375, B2 => 
                           n24919, ZN => n5470);
   U23540 : OAI22_X1 port map( A1 => n24927, A2 => n25428, B1 => n7373, B2 => 
                           n24920, ZN => n5471);
   U23541 : OAI22_X1 port map( A1 => n24927, A2 => n25431, B1 => n7371, B2 => 
                           n24921, ZN => n5472);
   U23542 : OAI22_X1 port map( A1 => n24927, A2 => n25434, B1 => n7369, B2 => 
                           n24919, ZN => n5473);
   U23543 : OAI22_X1 port map( A1 => n24928, A2 => n25437, B1 => n7367, B2 => 
                           n24920, ZN => n5474);
   U23544 : OAI22_X1 port map( A1 => n24928, A2 => n25440, B1 => n7365, B2 => 
                           n24921, ZN => n5475);
   U23545 : OAI22_X1 port map( A1 => n24928, A2 => n25443, B1 => n7363, B2 => 
                           n24919, ZN => n5476);
   U23546 : OAI22_X1 port map( A1 => n24928, A2 => n25446, B1 => n7361, B2 => 
                           n24920, ZN => n5477);
   U23547 : OAI22_X1 port map( A1 => n24928, A2 => n25449, B1 => n7359, B2 => 
                           n24921, ZN => n5478);
   U23548 : OAI22_X1 port map( A1 => n24929, A2 => n25452, B1 => n7357, B2 => 
                           n24919, ZN => n5479);
   U23549 : OAI22_X1 port map( A1 => n24929, A2 => n25455, B1 => n7355, B2 => 
                           n21290, ZN => n5480);
   U23550 : OAI22_X1 port map( A1 => n24929, A2 => n25458, B1 => n7353, B2 => 
                           n24919, ZN => n5481);
   U23551 : OAI22_X1 port map( A1 => n24929, A2 => n25461, B1 => n7351, B2 => 
                           n21290, ZN => n5482);
   U23552 : OAI22_X1 port map( A1 => n24929, A2 => n25464, B1 => n7349, B2 => 
                           n24919, ZN => n5483);
   U23553 : OAI22_X1 port map( A1 => n24930, A2 => n25467, B1 => n7347, B2 => 
                           n21290, ZN => n5484);
   U23554 : OAI22_X1 port map( A1 => n24930, A2 => n25470, B1 => n7345, B2 => 
                           n24919, ZN => n5485);
   U23555 : OAI22_X1 port map( A1 => n24930, A2 => n25473, B1 => n7343, B2 => 
                           n24920, ZN => n5486);
   U23556 : OAI22_X1 port map( A1 => n24930, A2 => n25476, B1 => n7341, B2 => 
                           n24921, ZN => n5487);
   U23557 : OAI22_X1 port map( A1 => n24930, A2 => n25479, B1 => n7339, B2 => 
                           n24919, ZN => n5488);
   U23558 : OAI22_X1 port map( A1 => n24931, A2 => n25482, B1 => n7337, B2 => 
                           n24919, ZN => n5489);
   U23559 : OAI22_X1 port map( A1 => n24931, A2 => n25485, B1 => n7335, B2 => 
                           n24920, ZN => n5490);
   U23560 : OAI22_X1 port map( A1 => n24931, A2 => n25488, B1 => n7333, B2 => 
                           n24921, ZN => n5491);
   U23561 : OAI22_X1 port map( A1 => n24931, A2 => n25491, B1 => n7331, B2 => 
                           n24919, ZN => n5492);
   U23562 : OAI22_X1 port map( A1 => n24931, A2 => n25494, B1 => n7329, B2 => 
                           n24919, ZN => n5493);
   U23563 : OAI22_X1 port map( A1 => n24932, A2 => n25497, B1 => n7327, B2 => 
                           n21290, ZN => n5494);
   U23564 : OAI22_X1 port map( A1 => n24932, A2 => n25500, B1 => n7325, B2 => 
                           n24919, ZN => n5495);
   U23565 : OAI22_X1 port map( A1 => n24932, A2 => n25503, B1 => n7323, B2 => 
                           n21290, ZN => n5496);
   U23566 : OAI22_X1 port map( A1 => n24932, A2 => n25506, B1 => n7321, B2 => 
                           n24919, ZN => n5497);
   U23567 : OAI22_X1 port map( A1 => n24932, A2 => n25509, B1 => n7319, B2 => 
                           n21290, ZN => n5498);
   U23568 : OAI22_X1 port map( A1 => n24933, A2 => n25512, B1 => n7317, B2 => 
                           n24919, ZN => n5499);
   U23569 : OAI22_X1 port map( A1 => n24933, A2 => n25515, B1 => n7315, B2 => 
                           n21290, ZN => n5500);
   U23570 : OAI22_X1 port map( A1 => n24933, A2 => n25518, B1 => n7313, B2 => 
                           n24919, ZN => n5501);
   U23571 : OAI22_X1 port map( A1 => n24933, A2 => n25521, B1 => n7311, B2 => 
                           n21290, ZN => n5502);
   U23572 : OAI22_X1 port map( A1 => n24933, A2 => n25524, B1 => n7309, B2 => 
                           n24919, ZN => n5503);
   U23573 : OAI22_X1 port map( A1 => n24960, A2 => n25418, B1 => n9197, B2 => 
                           n24954, ZN => n5596);
   U23574 : OAI22_X1 port map( A1 => n24961, A2 => n25421, B1 => n9195, B2 => 
                           n24955, ZN => n5597);
   U23575 : OAI22_X1 port map( A1 => n24961, A2 => n25424, B1 => n9193, B2 => 
                           n24953, ZN => n5598);
   U23576 : OAI22_X1 port map( A1 => n24961, A2 => n25427, B1 => n9191, B2 => 
                           n24954, ZN => n5599);
   U23577 : OAI22_X1 port map( A1 => n24961, A2 => n25430, B1 => n9189, B2 => 
                           n24955, ZN => n5600);
   U23578 : OAI22_X1 port map( A1 => n24961, A2 => n25433, B1 => n9187, B2 => 
                           n24953, ZN => n5601);
   U23579 : OAI22_X1 port map( A1 => n24962, A2 => n25436, B1 => n9185, B2 => 
                           n24954, ZN => n5602);
   U23580 : OAI22_X1 port map( A1 => n24962, A2 => n25439, B1 => n9183, B2 => 
                           n24955, ZN => n5603);
   U23581 : OAI22_X1 port map( A1 => n24962, A2 => n25442, B1 => n9181, B2 => 
                           n24953, ZN => n5604);
   U23582 : OAI22_X1 port map( A1 => n24962, A2 => n25445, B1 => n9179, B2 => 
                           n24954, ZN => n5605);
   U23583 : OAI22_X1 port map( A1 => n24962, A2 => n25448, B1 => n9177, B2 => 
                           n24955, ZN => n5606);
   U23584 : OAI22_X1 port map( A1 => n24963, A2 => n25451, B1 => n9175, B2 => 
                           n24953, ZN => n5607);
   U23585 : OAI22_X1 port map( A1 => n24963, A2 => n25454, B1 => n9173, B2 => 
                           n21287, ZN => n5608);
   U23586 : OAI22_X1 port map( A1 => n24963, A2 => n25457, B1 => n9171, B2 => 
                           n24953, ZN => n5609);
   U23587 : OAI22_X1 port map( A1 => n24963, A2 => n25460, B1 => n9169, B2 => 
                           n21287, ZN => n5610);
   U23588 : OAI22_X1 port map( A1 => n24963, A2 => n25463, B1 => n9167, B2 => 
                           n24953, ZN => n5611);
   U23589 : OAI22_X1 port map( A1 => n24964, A2 => n25466, B1 => n9165, B2 => 
                           n21287, ZN => n5612);
   U23590 : OAI22_X1 port map( A1 => n24964, A2 => n25469, B1 => n9163, B2 => 
                           n24953, ZN => n5613);
   U23591 : OAI22_X1 port map( A1 => n24964, A2 => n25472, B1 => n9161, B2 => 
                           n24954, ZN => n5614);
   U23592 : OAI22_X1 port map( A1 => n24964, A2 => n25475, B1 => n9159, B2 => 
                           n24955, ZN => n5615);
   U23593 : OAI22_X1 port map( A1 => n24964, A2 => n25478, B1 => n9157, B2 => 
                           n24953, ZN => n5616);
   U23594 : OAI22_X1 port map( A1 => n24965, A2 => n25481, B1 => n9155, B2 => 
                           n24953, ZN => n5617);
   U23595 : OAI22_X1 port map( A1 => n24965, A2 => n25484, B1 => n9153, B2 => 
                           n24954, ZN => n5618);
   U23596 : OAI22_X1 port map( A1 => n24965, A2 => n25487, B1 => n9151, B2 => 
                           n24955, ZN => n5619);
   U23597 : OAI22_X1 port map( A1 => n24965, A2 => n25490, B1 => n9149, B2 => 
                           n24953, ZN => n5620);
   U23598 : OAI22_X1 port map( A1 => n24965, A2 => n25493, B1 => n9147, B2 => 
                           n24953, ZN => n5621);
   U23599 : OAI22_X1 port map( A1 => n24966, A2 => n25496, B1 => n9145, B2 => 
                           n21287, ZN => n5622);
   U23600 : OAI22_X1 port map( A1 => n24966, A2 => n25499, B1 => n9143, B2 => 
                           n24953, ZN => n5623);
   U23601 : OAI22_X1 port map( A1 => n24966, A2 => n25502, B1 => n9141, B2 => 
                           n21287, ZN => n5624);
   U23602 : OAI22_X1 port map( A1 => n24966, A2 => n25505, B1 => n9139, B2 => 
                           n24953, ZN => n5625);
   U23603 : OAI22_X1 port map( A1 => n24966, A2 => n25508, B1 => n9137, B2 => 
                           n21287, ZN => n5626);
   U23604 : OAI22_X1 port map( A1 => n24967, A2 => n25511, B1 => n9135, B2 => 
                           n24953, ZN => n5627);
   U23605 : OAI22_X1 port map( A1 => n24967, A2 => n25514, B1 => n9133, B2 => 
                           n21287, ZN => n5628);
   U23606 : OAI22_X1 port map( A1 => n24967, A2 => n25517, B1 => n9131, B2 => 
                           n24953, ZN => n5629);
   U23607 : OAI22_X1 port map( A1 => n24967, A2 => n25520, B1 => n9129, B2 => 
                           n21287, ZN => n5630);
   U23608 : OAI22_X1 port map( A1 => n24967, A2 => n25523, B1 => n9127, B2 => 
                           n24953, ZN => n5631);
   U23609 : OAI22_X1 port map( A1 => n24977, A2 => n25418, B1 => n7507, B2 => 
                           n24971, ZN => n5660);
   U23610 : OAI22_X1 port map( A1 => n24978, A2 => n25421, B1 => n7505, B2 => 
                           n24972, ZN => n5661);
   U23611 : OAI22_X1 port map( A1 => n24978, A2 => n25424, B1 => n7503, B2 => 
                           n24970, ZN => n5662);
   U23612 : OAI22_X1 port map( A1 => n24978, A2 => n25427, B1 => n7501, B2 => 
                           n24971, ZN => n5663);
   U23613 : OAI22_X1 port map( A1 => n24978, A2 => n25430, B1 => n7499, B2 => 
                           n24972, ZN => n5664);
   U23614 : OAI22_X1 port map( A1 => n24978, A2 => n25433, B1 => n7497, B2 => 
                           n24970, ZN => n5665);
   U23615 : OAI22_X1 port map( A1 => n24979, A2 => n25436, B1 => n7495, B2 => 
                           n24971, ZN => n5666);
   U23616 : OAI22_X1 port map( A1 => n24979, A2 => n25439, B1 => n7493, B2 => 
                           n24972, ZN => n5667);
   U23617 : OAI22_X1 port map( A1 => n24979, A2 => n25442, B1 => n7491, B2 => 
                           n24970, ZN => n5668);
   U23618 : OAI22_X1 port map( A1 => n24979, A2 => n25445, B1 => n7489, B2 => 
                           n24971, ZN => n5669);
   U23619 : OAI22_X1 port map( A1 => n24979, A2 => n25448, B1 => n7487, B2 => 
                           n24972, ZN => n5670);
   U23620 : OAI22_X1 port map( A1 => n24980, A2 => n25451, B1 => n7485, B2 => 
                           n24970, ZN => n5671);
   U23621 : OAI22_X1 port map( A1 => n24980, A2 => n25454, B1 => n7483, B2 => 
                           n21286, ZN => n5672);
   U23622 : OAI22_X1 port map( A1 => n24980, A2 => n25457, B1 => n7481, B2 => 
                           n24970, ZN => n5673);
   U23623 : OAI22_X1 port map( A1 => n24980, A2 => n25460, B1 => n7479, B2 => 
                           n21286, ZN => n5674);
   U23624 : OAI22_X1 port map( A1 => n24980, A2 => n25463, B1 => n7477, B2 => 
                           n24970, ZN => n5675);
   U23625 : OAI22_X1 port map( A1 => n24981, A2 => n25466, B1 => n7475, B2 => 
                           n21286, ZN => n5676);
   U23626 : OAI22_X1 port map( A1 => n24981, A2 => n25469, B1 => n7473, B2 => 
                           n24970, ZN => n5677);
   U23627 : OAI22_X1 port map( A1 => n24981, A2 => n25472, B1 => n7471, B2 => 
                           n24971, ZN => n5678);
   U23628 : OAI22_X1 port map( A1 => n24981, A2 => n25475, B1 => n7469, B2 => 
                           n24972, ZN => n5679);
   U23629 : OAI22_X1 port map( A1 => n24981, A2 => n25478, B1 => n7467, B2 => 
                           n24970, ZN => n5680);
   U23630 : OAI22_X1 port map( A1 => n24982, A2 => n25481, B1 => n7465, B2 => 
                           n24970, ZN => n5681);
   U23631 : OAI22_X1 port map( A1 => n24982, A2 => n25484, B1 => n7463, B2 => 
                           n24971, ZN => n5682);
   U23632 : OAI22_X1 port map( A1 => n24982, A2 => n25487, B1 => n7461, B2 => 
                           n24972, ZN => n5683);
   U23633 : OAI22_X1 port map( A1 => n24982, A2 => n25490, B1 => n7459, B2 => 
                           n24970, ZN => n5684);
   U23634 : OAI22_X1 port map( A1 => n24982, A2 => n25493, B1 => n7457, B2 => 
                           n24970, ZN => n5685);
   U23635 : OAI22_X1 port map( A1 => n24983, A2 => n25496, B1 => n7455, B2 => 
                           n21286, ZN => n5686);
   U23636 : OAI22_X1 port map( A1 => n24983, A2 => n25499, B1 => n7453, B2 => 
                           n24970, ZN => n5687);
   U23637 : OAI22_X1 port map( A1 => n24983, A2 => n25502, B1 => n7451, B2 => 
                           n21286, ZN => n5688);
   U23638 : OAI22_X1 port map( A1 => n24983, A2 => n25505, B1 => n7449, B2 => 
                           n24970, ZN => n5689);
   U23639 : OAI22_X1 port map( A1 => n24983, A2 => n25508, B1 => n7447, B2 => 
                           n21286, ZN => n5690);
   U23640 : OAI22_X1 port map( A1 => n24984, A2 => n25511, B1 => n7445, B2 => 
                           n24970, ZN => n5691);
   U23641 : OAI22_X1 port map( A1 => n24984, A2 => n25514, B1 => n7443, B2 => 
                           n21286, ZN => n5692);
   U23642 : OAI22_X1 port map( A1 => n24984, A2 => n25517, B1 => n7441, B2 => 
                           n24970, ZN => n5693);
   U23643 : OAI22_X1 port map( A1 => n24984, A2 => n25520, B1 => n7439, B2 => 
                           n21286, ZN => n5694);
   U23644 : OAI22_X1 port map( A1 => n24984, A2 => n25523, B1 => n7437, B2 => 
                           n24970, ZN => n5695);
   U23645 : OAI22_X1 port map( A1 => n25113, A2 => n25418, B1 => n9068, B2 => 
                           n25107, ZN => n6172);
   U23646 : OAI22_X1 port map( A1 => n25114, A2 => n25421, B1 => n9066, B2 => 
                           n25108, ZN => n6173);
   U23647 : OAI22_X1 port map( A1 => n25114, A2 => n25424, B1 => n9064, B2 => 
                           n25106, ZN => n6174);
   U23648 : OAI22_X1 port map( A1 => n25114, A2 => n25427, B1 => n9062, B2 => 
                           n25107, ZN => n6175);
   U23649 : OAI22_X1 port map( A1 => n25114, A2 => n25430, B1 => n9060, B2 => 
                           n25108, ZN => n6176);
   U23650 : OAI22_X1 port map( A1 => n25114, A2 => n25433, B1 => n9058, B2 => 
                           n25106, ZN => n6177);
   U23651 : OAI22_X1 port map( A1 => n25115, A2 => n25436, B1 => n9056, B2 => 
                           n25107, ZN => n6178);
   U23652 : OAI22_X1 port map( A1 => n25115, A2 => n25439, B1 => n9054, B2 => 
                           n25108, ZN => n6179);
   U23653 : OAI22_X1 port map( A1 => n25115, A2 => n25442, B1 => n9052, B2 => 
                           n25106, ZN => n6180);
   U23654 : OAI22_X1 port map( A1 => n25115, A2 => n25445, B1 => n9050, B2 => 
                           n25107, ZN => n6181);
   U23655 : OAI22_X1 port map( A1 => n25115, A2 => n25448, B1 => n9048, B2 => 
                           n25108, ZN => n6182);
   U23656 : OAI22_X1 port map( A1 => n25116, A2 => n25451, B1 => n9046, B2 => 
                           n25106, ZN => n6183);
   U23657 : OAI22_X1 port map( A1 => n25116, A2 => n25454, B1 => n9044, B2 => 
                           n21277, ZN => n6184);
   U23658 : OAI22_X1 port map( A1 => n25116, A2 => n25457, B1 => n9042, B2 => 
                           n25106, ZN => n6185);
   U23659 : OAI22_X1 port map( A1 => n25116, A2 => n25460, B1 => n9040, B2 => 
                           n21277, ZN => n6186);
   U23660 : OAI22_X1 port map( A1 => n25116, A2 => n25463, B1 => n9038, B2 => 
                           n25106, ZN => n6187);
   U23661 : OAI22_X1 port map( A1 => n25117, A2 => n25466, B1 => n9036, B2 => 
                           n21277, ZN => n6188);
   U23662 : OAI22_X1 port map( A1 => n25117, A2 => n25469, B1 => n9034, B2 => 
                           n25106, ZN => n6189);
   U23663 : OAI22_X1 port map( A1 => n25117, A2 => n25472, B1 => n9032, B2 => 
                           n25107, ZN => n6190);
   U23664 : OAI22_X1 port map( A1 => n25117, A2 => n25475, B1 => n9030, B2 => 
                           n25108, ZN => n6191);
   U23665 : OAI22_X1 port map( A1 => n25117, A2 => n25478, B1 => n9028, B2 => 
                           n25106, ZN => n6192);
   U23666 : OAI22_X1 port map( A1 => n25118, A2 => n25481, B1 => n9026, B2 => 
                           n25106, ZN => n6193);
   U23667 : OAI22_X1 port map( A1 => n25118, A2 => n25484, B1 => n9024, B2 => 
                           n25107, ZN => n6194);
   U23668 : OAI22_X1 port map( A1 => n25118, A2 => n25487, B1 => n9022, B2 => 
                           n25108, ZN => n6195);
   U23669 : OAI22_X1 port map( A1 => n25118, A2 => n25490, B1 => n9020, B2 => 
                           n25106, ZN => n6196);
   U23670 : OAI22_X1 port map( A1 => n25118, A2 => n25493, B1 => n9018, B2 => 
                           n25106, ZN => n6197);
   U23671 : OAI22_X1 port map( A1 => n25119, A2 => n25496, B1 => n9016, B2 => 
                           n21277, ZN => n6198);
   U23672 : OAI22_X1 port map( A1 => n25119, A2 => n25499, B1 => n9014, B2 => 
                           n25106, ZN => n6199);
   U23673 : OAI22_X1 port map( A1 => n25119, A2 => n25502, B1 => n9012, B2 => 
                           n21277, ZN => n6200);
   U23674 : OAI22_X1 port map( A1 => n25119, A2 => n25505, B1 => n9010, B2 => 
                           n25106, ZN => n6201);
   U23675 : OAI22_X1 port map( A1 => n25119, A2 => n25508, B1 => n9008, B2 => 
                           n21277, ZN => n6202);
   U23676 : OAI22_X1 port map( A1 => n25120, A2 => n25511, B1 => n9006, B2 => 
                           n25106, ZN => n6203);
   U23677 : OAI22_X1 port map( A1 => n25120, A2 => n25514, B1 => n9004, B2 => 
                           n21277, ZN => n6204);
   U23678 : OAI22_X1 port map( A1 => n25120, A2 => n25517, B1 => n9002, B2 => 
                           n25106, ZN => n6205);
   U23679 : OAI22_X1 port map( A1 => n25120, A2 => n25520, B1 => n9000, B2 => 
                           n21277, ZN => n6206);
   U23680 : OAI22_X1 port map( A1 => n25120, A2 => n25523, B1 => n8998, B2 => 
                           n25106, ZN => n6207);
   U23681 : OAI22_X1 port map( A1 => n25130, A2 => n25418, B1 => n872, B2 => 
                           n25124, ZN => n6236);
   U23682 : OAI22_X1 port map( A1 => n25131, A2 => n25421, B1 => n871, B2 => 
                           n25125, ZN => n6237);
   U23683 : OAI22_X1 port map( A1 => n25131, A2 => n25424, B1 => n870, B2 => 
                           n25123, ZN => n6238);
   U23684 : OAI22_X1 port map( A1 => n25131, A2 => n25427, B1 => n869, B2 => 
                           n25124, ZN => n6239);
   U23685 : OAI22_X1 port map( A1 => n25131, A2 => n25430, B1 => n868, B2 => 
                           n25125, ZN => n6240);
   U23686 : OAI22_X1 port map( A1 => n25131, A2 => n25433, B1 => n867, B2 => 
                           n25123, ZN => n6241);
   U23687 : OAI22_X1 port map( A1 => n25132, A2 => n25436, B1 => n866, B2 => 
                           n25124, ZN => n6242);
   U23688 : OAI22_X1 port map( A1 => n25132, A2 => n25439, B1 => n865, B2 => 
                           n25125, ZN => n6243);
   U23689 : OAI22_X1 port map( A1 => n25132, A2 => n25442, B1 => n864, B2 => 
                           n25123, ZN => n6244);
   U23690 : OAI22_X1 port map( A1 => n25132, A2 => n25445, B1 => n863, B2 => 
                           n25124, ZN => n6245);
   U23691 : OAI22_X1 port map( A1 => n25132, A2 => n25448, B1 => n862, B2 => 
                           n25125, ZN => n6246);
   U23692 : OAI22_X1 port map( A1 => n25133, A2 => n25451, B1 => n861, B2 => 
                           n25123, ZN => n6247);
   U23693 : OAI22_X1 port map( A1 => n25133, A2 => n25454, B1 => n860, B2 => 
                           n21276, ZN => n6248);
   U23694 : OAI22_X1 port map( A1 => n25133, A2 => n25457, B1 => n859, B2 => 
                           n25123, ZN => n6249);
   U23695 : OAI22_X1 port map( A1 => n25133, A2 => n25460, B1 => n858, B2 => 
                           n21276, ZN => n6250);
   U23696 : OAI22_X1 port map( A1 => n25133, A2 => n25463, B1 => n857, B2 => 
                           n25123, ZN => n6251);
   U23697 : OAI22_X1 port map( A1 => n25134, A2 => n25466, B1 => n856, B2 => 
                           n21276, ZN => n6252);
   U23698 : OAI22_X1 port map( A1 => n25134, A2 => n25469, B1 => n855, B2 => 
                           n25123, ZN => n6253);
   U23699 : OAI22_X1 port map( A1 => n25134, A2 => n25472, B1 => n854, B2 => 
                           n25124, ZN => n6254);
   U23700 : OAI22_X1 port map( A1 => n25134, A2 => n25475, B1 => n853, B2 => 
                           n25125, ZN => n6255);
   U23701 : OAI22_X1 port map( A1 => n25134, A2 => n25478, B1 => n852, B2 => 
                           n25123, ZN => n6256);
   U23702 : OAI22_X1 port map( A1 => n25135, A2 => n25481, B1 => n851, B2 => 
                           n25123, ZN => n6257);
   U23703 : OAI22_X1 port map( A1 => n25135, A2 => n25484, B1 => n850, B2 => 
                           n25124, ZN => n6258);
   U23704 : OAI22_X1 port map( A1 => n25135, A2 => n25487, B1 => n849, B2 => 
                           n25125, ZN => n6259);
   U23705 : OAI22_X1 port map( A1 => n25135, A2 => n25490, B1 => n848, B2 => 
                           n25123, ZN => n6260);
   U23706 : OAI22_X1 port map( A1 => n25135, A2 => n25493, B1 => n847, B2 => 
                           n25123, ZN => n6261);
   U23707 : OAI22_X1 port map( A1 => n25136, A2 => n25496, B1 => n846, B2 => 
                           n21276, ZN => n6262);
   U23708 : OAI22_X1 port map( A1 => n25136, A2 => n25499, B1 => n845, B2 => 
                           n25123, ZN => n6263);
   U23709 : OAI22_X1 port map( A1 => n25136, A2 => n25502, B1 => n844, B2 => 
                           n21276, ZN => n6264);
   U23710 : OAI22_X1 port map( A1 => n25136, A2 => n25505, B1 => n843, B2 => 
                           n25123, ZN => n6265);
   U23711 : OAI22_X1 port map( A1 => n25136, A2 => n25508, B1 => n842, B2 => 
                           n21276, ZN => n6266);
   U23712 : OAI22_X1 port map( A1 => n25137, A2 => n25511, B1 => n841, B2 => 
                           n25123, ZN => n6267);
   U23713 : OAI22_X1 port map( A1 => n25137, A2 => n25514, B1 => n840, B2 => 
                           n21276, ZN => n6268);
   U23714 : OAI22_X1 port map( A1 => n25137, A2 => n25517, B1 => n839, B2 => 
                           n25123, ZN => n6269);
   U23715 : OAI22_X1 port map( A1 => n25137, A2 => n25520, B1 => n838, B2 => 
                           n21276, ZN => n6270);
   U23716 : OAI22_X1 port map( A1 => n25137, A2 => n25523, B1 => n837, B2 => 
                           n25123, ZN => n6271);
   U23717 : OAI22_X1 port map( A1 => n25164, A2 => n25417, B1 => n9196, B2 => 
                           n25158, ZN => n6364);
   U23718 : OAI22_X1 port map( A1 => n25165, A2 => n25420, B1 => n9194, B2 => 
                           n25159, ZN => n6365);
   U23719 : OAI22_X1 port map( A1 => n25165, A2 => n25423, B1 => n9192, B2 => 
                           n25157, ZN => n6366);
   U23720 : OAI22_X1 port map( A1 => n25165, A2 => n25426, B1 => n9190, B2 => 
                           n25158, ZN => n6367);
   U23721 : OAI22_X1 port map( A1 => n25165, A2 => n25429, B1 => n9188, B2 => 
                           n25159, ZN => n6368);
   U23722 : OAI22_X1 port map( A1 => n25165, A2 => n25432, B1 => n9186, B2 => 
                           n25157, ZN => n6369);
   U23723 : OAI22_X1 port map( A1 => n25166, A2 => n25435, B1 => n9184, B2 => 
                           n25158, ZN => n6370);
   U23724 : OAI22_X1 port map( A1 => n25166, A2 => n25438, B1 => n9182, B2 => 
                           n25159, ZN => n6371);
   U23725 : OAI22_X1 port map( A1 => n25166, A2 => n25441, B1 => n9180, B2 => 
                           n25157, ZN => n6372);
   U23726 : OAI22_X1 port map( A1 => n25166, A2 => n25444, B1 => n9178, B2 => 
                           n25158, ZN => n6373);
   U23727 : OAI22_X1 port map( A1 => n25166, A2 => n25447, B1 => n9176, B2 => 
                           n25159, ZN => n6374);
   U23728 : OAI22_X1 port map( A1 => n25167, A2 => n25450, B1 => n9174, B2 => 
                           n25157, ZN => n6375);
   U23729 : OAI22_X1 port map( A1 => n25167, A2 => n25453, B1 => n9172, B2 => 
                           n21274, ZN => n6376);
   U23730 : OAI22_X1 port map( A1 => n25167, A2 => n25456, B1 => n9170, B2 => 
                           n25157, ZN => n6377);
   U23731 : OAI22_X1 port map( A1 => n25167, A2 => n25459, B1 => n9168, B2 => 
                           n21274, ZN => n6378);
   U23732 : OAI22_X1 port map( A1 => n25167, A2 => n25462, B1 => n9166, B2 => 
                           n25157, ZN => n6379);
   U23733 : OAI22_X1 port map( A1 => n25168, A2 => n25465, B1 => n9164, B2 => 
                           n21274, ZN => n6380);
   U23734 : OAI22_X1 port map( A1 => n25168, A2 => n25468, B1 => n9162, B2 => 
                           n25157, ZN => n6381);
   U23735 : OAI22_X1 port map( A1 => n25168, A2 => n25471, B1 => n9160, B2 => 
                           n25158, ZN => n6382);
   U23736 : OAI22_X1 port map( A1 => n25168, A2 => n25474, B1 => n9158, B2 => 
                           n25159, ZN => n6383);
   U23737 : OAI22_X1 port map( A1 => n25168, A2 => n25477, B1 => n9156, B2 => 
                           n25157, ZN => n6384);
   U23738 : OAI22_X1 port map( A1 => n25169, A2 => n25480, B1 => n9154, B2 => 
                           n25157, ZN => n6385);
   U23739 : OAI22_X1 port map( A1 => n25169, A2 => n25483, B1 => n9152, B2 => 
                           n25158, ZN => n6386);
   U23740 : OAI22_X1 port map( A1 => n25169, A2 => n25486, B1 => n9150, B2 => 
                           n25159, ZN => n6387);
   U23741 : OAI22_X1 port map( A1 => n25169, A2 => n25489, B1 => n9148, B2 => 
                           n25157, ZN => n6388);
   U23742 : OAI22_X1 port map( A1 => n25169, A2 => n25492, B1 => n9146, B2 => 
                           n25157, ZN => n6389);
   U23743 : OAI22_X1 port map( A1 => n25170, A2 => n25495, B1 => n9144, B2 => 
                           n21274, ZN => n6390);
   U23744 : OAI22_X1 port map( A1 => n25170, A2 => n25498, B1 => n9142, B2 => 
                           n25157, ZN => n6391);
   U23745 : OAI22_X1 port map( A1 => n25170, A2 => n25501, B1 => n9140, B2 => 
                           n21274, ZN => n6392);
   U23746 : OAI22_X1 port map( A1 => n25170, A2 => n25504, B1 => n9138, B2 => 
                           n25157, ZN => n6393);
   U23747 : OAI22_X1 port map( A1 => n25170, A2 => n25507, B1 => n9136, B2 => 
                           n21274, ZN => n6394);
   U23748 : OAI22_X1 port map( A1 => n25171, A2 => n25510, B1 => n9134, B2 => 
                           n25157, ZN => n6395);
   U23749 : OAI22_X1 port map( A1 => n25171, A2 => n25513, B1 => n9132, B2 => 
                           n21274, ZN => n6396);
   U23750 : OAI22_X1 port map( A1 => n25171, A2 => n25516, B1 => n9130, B2 => 
                           n25157, ZN => n6397);
   U23751 : OAI22_X1 port map( A1 => n25171, A2 => n25519, B1 => n9128, B2 => 
                           n21274, ZN => n6398);
   U23752 : OAI22_X1 port map( A1 => n25171, A2 => n25522, B1 => n9126, B2 => 
                           n25157, ZN => n6399);
   U23753 : OAI22_X1 port map( A1 => n25274, A2 => n25525, B1 => n17230, B2 => 
                           n21263, ZN => n6784);
   U23754 : OAI22_X1 port map( A1 => n25274, A2 => n25528, B1 => n17227, B2 => 
                           n21263, ZN => n6785);
   U23755 : OAI22_X1 port map( A1 => n25274, A2 => n25531, B1 => n17224, B2 => 
                           n25259, ZN => n6786);
   U23756 : OAI22_X1 port map( A1 => n25274, A2 => n25551, B1 => n17221, B2 => 
                           n21263, ZN => n6787);
   U23757 : OAI22_X1 port map( A1 => n24968, A2 => n25526, B1 => n9125, B2 => 
                           n21287, ZN => n5632);
   U23758 : OAI22_X1 port map( A1 => n24968, A2 => n25529, B1 => n9123, B2 => 
                           n21287, ZN => n5633);
   U23759 : OAI22_X1 port map( A1 => n24968, A2 => n25532, B1 => n9121, B2 => 
                           n24953, ZN => n5634);
   U23760 : OAI22_X1 port map( A1 => n24968, A2 => n25552, B1 => n9119, B2 => 
                           n21287, ZN => n5635);
   U23761 : OAI22_X1 port map( A1 => n25036, A2 => n25526, B1 => n8869, B2 => 
                           n21283, ZN => n5888);
   U23762 : OAI22_X1 port map( A1 => n25036, A2 => n25529, B1 => n8867, B2 => 
                           n21283, ZN => n5889);
   U23763 : OAI22_X1 port map( A1 => n25036, A2 => n25532, B1 => n8865, B2 => 
                           n25021, ZN => n5890);
   U23764 : OAI22_X1 port map( A1 => n25036, A2 => n25552, B1 => n8863, B2 => 
                           n21283, ZN => n5891);
   U23765 : OAI22_X1 port map( A1 => n24866, A2 => n25527, B1 => n8868, B2 => 
                           n21294, ZN => n5248);
   U23766 : OAI22_X1 port map( A1 => n24866, A2 => n25530, B1 => n8866, B2 => 
                           n21294, ZN => n5249);
   U23767 : OAI22_X1 port map( A1 => n24866, A2 => n25533, B1 => n8864, B2 => 
                           n24851, ZN => n5250);
   U23768 : OAI22_X1 port map( A1 => n24866, A2 => n25553, B1 => n8862, B2 => 
                           n21294, ZN => n5251);
   U23769 : OAI22_X1 port map( A1 => n25172, A2 => n25525, B1 => n9124, B2 => 
                           n21274, ZN => n6400);
   U23770 : OAI22_X1 port map( A1 => n25172, A2 => n25528, B1 => n9122, B2 => 
                           n21274, ZN => n6401);
   U23771 : OAI22_X1 port map( A1 => n25172, A2 => n25531, B1 => n9120, B2 => 
                           n25157, ZN => n6402);
   U23772 : OAI22_X1 port map( A1 => n25172, A2 => n25551, B1 => n9118, B2 => 
                           n21274, ZN => n6403);
   U23773 : OAI22_X1 port map( A1 => n25189, A2 => n25525, B1 => n7434, B2 => 
                           n21273, ZN => n6464);
   U23774 : OAI22_X1 port map( A1 => n25189, A2 => n25528, B1 => n7432, B2 => 
                           n21273, ZN => n6465);
   U23775 : OAI22_X1 port map( A1 => n25189, A2 => n25531, B1 => n7430, B2 => 
                           n25174, ZN => n6466);
   U23776 : OAI22_X1 port map( A1 => n25189, A2 => n25551, B1 => n7428, B2 => 
                           n21273, ZN => n6467);
   U23777 : OAI22_X1 port map( A1 => n24934, A2 => n25527, B1 => n7307, B2 => 
                           n21290, ZN => n5504);
   U23778 : OAI22_X1 port map( A1 => n24934, A2 => n25530, B1 => n7305, B2 => 
                           n21290, ZN => n5505);
   U23779 : OAI22_X1 port map( A1 => n24934, A2 => n25533, B1 => n7303, B2 => 
                           n24919, ZN => n5506);
   U23780 : OAI22_X1 port map( A1 => n24934, A2 => n25553, B1 => n7301, B2 => 
                           n21290, ZN => n5507);
   U23781 : OAI22_X1 port map( A1 => n25138, A2 => n25526, B1 => n836, B2 => 
                           n21276, ZN => n6272);
   U23782 : OAI22_X1 port map( A1 => n25138, A2 => n25529, B1 => n835, B2 => 
                           n21276, ZN => n6273);
   U23783 : OAI22_X1 port map( A1 => n25138, A2 => n25532, B1 => n834, B2 => 
                           n25123, ZN => n6274);
   U23784 : OAI22_X1 port map( A1 => n25138, A2 => n25552, B1 => n833, B2 => 
                           n21276, ZN => n6275);
   U23785 : OAI22_X1 port map( A1 => n25053, A2 => n25526, B1 => n8741, B2 => 
                           n21282, ZN => n5952);
   U23786 : OAI22_X1 port map( A1 => n25053, A2 => n25529, B1 => n8739, B2 => 
                           n21282, ZN => n5953);
   U23787 : OAI22_X1 port map( A1 => n25053, A2 => n25532, B1 => n8737, B2 => 
                           n25038, ZN => n5954);
   U23788 : OAI22_X1 port map( A1 => n25053, A2 => n25552, B1 => n8735, B2 => 
                           n21282, ZN => n5955);
   U23789 : OAI22_X1 port map( A1 => n24985, A2 => n25526, B1 => n7435, B2 => 
                           n21286, ZN => n5696);
   U23790 : OAI22_X1 port map( A1 => n24985, A2 => n25529, B1 => n7433, B2 => 
                           n21286, ZN => n5697);
   U23791 : OAI22_X1 port map( A1 => n24985, A2 => n25532, B1 => n7431, B2 => 
                           n24970, ZN => n5698);
   U23792 : OAI22_X1 port map( A1 => n24985, A2 => n25552, B1 => n7429, B2 => 
                           n21286, ZN => n5699);
   U23793 : OAI22_X1 port map( A1 => n25121, A2 => n25526, B1 => n8996, B2 => 
                           n21277, ZN => n6208);
   U23794 : OAI22_X1 port map( A1 => n25121, A2 => n25529, B1 => n8994, B2 => 
                           n21277, ZN => n6209);
   U23795 : OAI22_X1 port map( A1 => n25121, A2 => n25532, B1 => n8992, B2 => 
                           n25106, ZN => n6210);
   U23796 : OAI22_X1 port map( A1 => n25121, A2 => n25552, B1 => n8990, B2 => 
                           n21277, ZN => n6211);
   U23797 : OAI22_X1 port map( A1 => n24900, A2 => n25527, B1 => n21292, B2 => 
                           n20530, ZN => n5376);
   U23798 : OAI22_X1 port map( A1 => n24900, A2 => n25530, B1 => n21292, B2 => 
                           n20529, ZN => n5377);
   U23799 : OAI22_X1 port map( A1 => n24900, A2 => n25533, B1 => n24885, B2 => 
                           n20528, ZN => n5378);
   U23800 : OAI22_X1 port map( A1 => n24900, A2 => n25553, B1 => n21292, B2 => 
                           n20527, ZN => n5379);
   U23801 : OAI221_X1 port map( B1 => n19207, B2 => n24809, C1 => n11843, C2 =>
                           n24798, A => n21389, ZN => n5056);
   U23802 : OAI21_X1 port map( B1 => n21390, B2 => n21391, A => n24797, ZN => 
                           n21389);
   U23803 : NAND4_X1 port map( A1 => n21400, A2 => n21401, A3 => n21402, A4 => 
                           n21403, ZN => n21390);
   U23804 : NAND4_X1 port map( A1 => n21392, A2 => n21393, A3 => n21394, A4 => 
                           n21395, ZN => n21391);
   U23805 : OAI221_X1 port map( B1 => n19206, B2 => n24809, C1 => n11844, C2 =>
                           n24798, A => n21370, ZN => n5057);
   U23806 : OAI21_X1 port map( B1 => n21371, B2 => n21372, A => n24797, ZN => 
                           n21370);
   U23807 : NAND4_X1 port map( A1 => n21381, A2 => n21382, A3 => n21383, A4 => 
                           n21384, ZN => n21371);
   U23808 : NAND4_X1 port map( A1 => n21373, A2 => n21374, A3 => n21375, A4 => 
                           n21376, ZN => n21372);
   U23809 : OAI221_X1 port map( B1 => n19205, B2 => n24809, C1 => n11845, C2 =>
                           n24798, A => n21351, ZN => n5058);
   U23810 : OAI21_X1 port map( B1 => n21352, B2 => n21353, A => n24797, ZN => 
                           n21351);
   U23811 : NAND4_X1 port map( A1 => n21362, A2 => n21363, A3 => n21364, A4 => 
                           n21365, ZN => n21352);
   U23812 : NAND4_X1 port map( A1 => n21354, A2 => n21355, A3 => n21356, A4 => 
                           n21357, ZN => n21353);
   U23813 : OAI221_X1 port map( B1 => n19204, B2 => n24809, C1 => n11846, C2 =>
                           n24800, A => n21299, ZN => n5059);
   U23814 : OAI21_X1 port map( B1 => n21300, B2 => n21301, A => n24797, ZN => 
                           n21299);
   U23815 : NAND4_X1 port map( A1 => n21327, A2 => n21328, A3 => n21329, A4 => 
                           n21330, ZN => n21300);
   U23816 : NAND4_X1 port map( A1 => n21303, A2 => n21304, A3 => n21305, A4 => 
                           n21306, ZN => n21301);
   U23817 : OAI221_X1 port map( B1 => n19267, B2 => n24804, C1 => n11783, C2 =>
                           n24803, A => n22529, ZN => n4996);
   U23818 : OAI21_X1 port map( B1 => n22530, B2 => n22531, A => n24792, ZN => 
                           n22529);
   U23819 : NAND4_X1 port map( A1 => n22548, A2 => n22549, A3 => n22550, A4 => 
                           n22551, ZN => n22530);
   U23820 : NAND4_X1 port map( A1 => n22532, A2 => n22533, A3 => n22534, A4 => 
                           n22535, ZN => n22531);
   U23821 : OAI221_X1 port map( B1 => n19266, B2 => n24804, C1 => n11784, C2 =>
                           n24803, A => n22510, ZN => n4997);
   U23822 : OAI21_X1 port map( B1 => n22511, B2 => n22512, A => n24792, ZN => 
                           n22510);
   U23823 : NAND4_X1 port map( A1 => n22521, A2 => n22522, A3 => n22523, A4 => 
                           n22524, ZN => n22511);
   U23824 : NAND4_X1 port map( A1 => n22513, A2 => n22514, A3 => n22515, A4 => 
                           n22516, ZN => n22512);
   U23825 : OAI221_X1 port map( B1 => n19265, B2 => n24804, C1 => n11785, C2 =>
                           n24803, A => n22491, ZN => n4998);
   U23826 : OAI21_X1 port map( B1 => n22492, B2 => n22493, A => n24792, ZN => 
                           n22491);
   U23827 : NAND4_X1 port map( A1 => n22502, A2 => n22503, A3 => n22504, A4 => 
                           n22505, ZN => n22492);
   U23828 : NAND4_X1 port map( A1 => n22494, A2 => n22495, A3 => n22496, A4 => 
                           n22497, ZN => n22493);
   U23829 : OAI221_X1 port map( B1 => n19264, B2 => n24804, C1 => n11786, C2 =>
                           n24803, A => n22472, ZN => n4999);
   U23830 : OAI21_X1 port map( B1 => n22473, B2 => n22474, A => n24792, ZN => 
                           n22472);
   U23831 : NAND4_X1 port map( A1 => n22483, A2 => n22484, A3 => n22485, A4 => 
                           n22486, ZN => n22473);
   U23832 : NAND4_X1 port map( A1 => n22475, A2 => n22476, A3 => n22477, A4 => 
                           n22478, ZN => n22474);
   U23833 : OAI221_X1 port map( B1 => n19263, B2 => n24804, C1 => n11787, C2 =>
                           n24802, A => n22453, ZN => n5000);
   U23834 : OAI21_X1 port map( B1 => n22454, B2 => n22455, A => n24792, ZN => 
                           n22453);
   U23835 : NAND4_X1 port map( A1 => n22464, A2 => n22465, A3 => n22466, A4 => 
                           n22467, ZN => n22454);
   U23836 : NAND4_X1 port map( A1 => n22456, A2 => n22457, A3 => n22458, A4 => 
                           n22459, ZN => n22455);
   U23837 : OAI221_X1 port map( B1 => n19262, B2 => n24804, C1 => n11788, C2 =>
                           n24802, A => n22434, ZN => n5001);
   U23838 : OAI21_X1 port map( B1 => n22435, B2 => n22436, A => n24792, ZN => 
                           n22434);
   U23839 : NAND4_X1 port map( A1 => n22445, A2 => n22446, A3 => n22447, A4 => 
                           n22448, ZN => n22435);
   U23840 : NAND4_X1 port map( A1 => n22437, A2 => n22438, A3 => n22439, A4 => 
                           n22440, ZN => n22436);
   U23841 : OAI221_X1 port map( B1 => n19261, B2 => n24804, C1 => n11789, C2 =>
                           n24802, A => n22415, ZN => n5002);
   U23842 : OAI21_X1 port map( B1 => n22416, B2 => n22417, A => n24792, ZN => 
                           n22415);
   U23843 : NAND4_X1 port map( A1 => n22426, A2 => n22427, A3 => n22428, A4 => 
                           n22429, ZN => n22416);
   U23844 : NAND4_X1 port map( A1 => n22418, A2 => n22419, A3 => n22420, A4 => 
                           n22421, ZN => n22417);
   U23845 : OAI221_X1 port map( B1 => n19260, B2 => n24804, C1 => n11790, C2 =>
                           n24802, A => n22396, ZN => n5003);
   U23846 : OAI21_X1 port map( B1 => n22397, B2 => n22398, A => n24792, ZN => 
                           n22396);
   U23847 : NAND4_X1 port map( A1 => n22407, A2 => n22408, A3 => n22409, A4 => 
                           n22410, ZN => n22397);
   U23848 : NAND4_X1 port map( A1 => n22399, A2 => n22400, A3 => n22401, A4 => 
                           n22402, ZN => n22398);
   U23849 : OAI221_X1 port map( B1 => n19259, B2 => n24804, C1 => n11791, C2 =>
                           n24802, A => n22377, ZN => n5004);
   U23850 : OAI21_X1 port map( B1 => n22378, B2 => n22379, A => n24792, ZN => 
                           n22377);
   U23851 : NAND4_X1 port map( A1 => n22388, A2 => n22389, A3 => n22390, A4 => 
                           n22391, ZN => n22378);
   U23852 : NAND4_X1 port map( A1 => n22380, A2 => n22381, A3 => n22382, A4 => 
                           n22383, ZN => n22379);
   U23853 : OAI221_X1 port map( B1 => n19258, B2 => n24804, C1 => n11792, C2 =>
                           n24802, A => n22358, ZN => n5005);
   U23854 : OAI21_X1 port map( B1 => n22359, B2 => n22360, A => n24792, ZN => 
                           n22358);
   U23855 : NAND4_X1 port map( A1 => n22369, A2 => n22370, A3 => n22371, A4 => 
                           n22372, ZN => n22359);
   U23856 : NAND4_X1 port map( A1 => n22361, A2 => n22362, A3 => n22363, A4 => 
                           n22364, ZN => n22360);
   U23857 : OAI221_X1 port map( B1 => n19257, B2 => n24804, C1 => n11793, C2 =>
                           n24802, A => n22339, ZN => n5006);
   U23858 : OAI21_X1 port map( B1 => n22340, B2 => n22341, A => n24792, ZN => 
                           n22339);
   U23859 : NAND4_X1 port map( A1 => n22350, A2 => n22351, A3 => n22352, A4 => 
                           n22353, ZN => n22340);
   U23860 : NAND4_X1 port map( A1 => n22342, A2 => n22343, A3 => n22344, A4 => 
                           n22345, ZN => n22341);
   U23861 : OAI221_X1 port map( B1 => n19256, B2 => n24804, C1 => n11794, C2 =>
                           n24802, A => n22320, ZN => n5007);
   U23862 : OAI21_X1 port map( B1 => n22321, B2 => n22322, A => n24792, ZN => 
                           n22320);
   U23863 : NAND4_X1 port map( A1 => n22331, A2 => n22332, A3 => n22333, A4 => 
                           n22334, ZN => n22321);
   U23864 : NAND4_X1 port map( A1 => n22323, A2 => n22324, A3 => n22325, A4 => 
                           n22326, ZN => n22322);
   U23865 : OAI221_X1 port map( B1 => n19255, B2 => n24805, C1 => n11795, C2 =>
                           n24802, A => n22301, ZN => n5008);
   U23866 : OAI21_X1 port map( B1 => n22302, B2 => n22303, A => n24793, ZN => 
                           n22301);
   U23867 : NAND4_X1 port map( A1 => n22312, A2 => n22313, A3 => n22314, A4 => 
                           n22315, ZN => n22302);
   U23868 : NAND4_X1 port map( A1 => n22304, A2 => n22305, A3 => n22306, A4 => 
                           n22307, ZN => n22303);
   U23869 : OAI221_X1 port map( B1 => n19254, B2 => n24805, C1 => n11796, C2 =>
                           n24802, A => n22282, ZN => n5009);
   U23870 : OAI21_X1 port map( B1 => n22283, B2 => n22284, A => n24793, ZN => 
                           n22282);
   U23871 : NAND4_X1 port map( A1 => n22293, A2 => n22294, A3 => n22295, A4 => 
                           n22296, ZN => n22283);
   U23872 : NAND4_X1 port map( A1 => n22285, A2 => n22286, A3 => n22287, A4 => 
                           n22288, ZN => n22284);
   U23873 : OAI221_X1 port map( B1 => n19253, B2 => n24805, C1 => n11797, C2 =>
                           n24802, A => n22263, ZN => n5010);
   U23874 : OAI21_X1 port map( B1 => n22264, B2 => n22265, A => n24793, ZN => 
                           n22263);
   U23875 : NAND4_X1 port map( A1 => n22274, A2 => n22275, A3 => n22276, A4 => 
                           n22277, ZN => n22264);
   U23876 : NAND4_X1 port map( A1 => n22266, A2 => n22267, A3 => n22268, A4 => 
                           n22269, ZN => n22265);
   U23877 : OAI221_X1 port map( B1 => n19252, B2 => n24805, C1 => n11798, C2 =>
                           n24802, A => n22244, ZN => n5011);
   U23878 : OAI21_X1 port map( B1 => n22245, B2 => n22246, A => n24793, ZN => 
                           n22244);
   U23879 : NAND4_X1 port map( A1 => n22255, A2 => n22256, A3 => n22257, A4 => 
                           n22258, ZN => n22245);
   U23880 : NAND4_X1 port map( A1 => n22247, A2 => n22248, A3 => n22249, A4 => 
                           n22250, ZN => n22246);
   U23881 : OAI221_X1 port map( B1 => n19251, B2 => n24805, C1 => n11799, C2 =>
                           n24801, A => n22225, ZN => n5012);
   U23882 : OAI21_X1 port map( B1 => n22226, B2 => n22227, A => n24793, ZN => 
                           n22225);
   U23883 : NAND4_X1 port map( A1 => n22236, A2 => n22237, A3 => n22238, A4 => 
                           n22239, ZN => n22226);
   U23884 : NAND4_X1 port map( A1 => n22228, A2 => n22229, A3 => n22230, A4 => 
                           n22231, ZN => n22227);
   U23885 : OAI221_X1 port map( B1 => n19250, B2 => n24805, C1 => n11800, C2 =>
                           n24801, A => n22206, ZN => n5013);
   U23886 : OAI21_X1 port map( B1 => n22207, B2 => n22208, A => n24793, ZN => 
                           n22206);
   U23887 : NAND4_X1 port map( A1 => n22217, A2 => n22218, A3 => n22219, A4 => 
                           n22220, ZN => n22207);
   U23888 : NAND4_X1 port map( A1 => n22209, A2 => n22210, A3 => n22211, A4 => 
                           n22212, ZN => n22208);
   U23889 : OAI221_X1 port map( B1 => n19249, B2 => n24805, C1 => n11801, C2 =>
                           n24801, A => n22187, ZN => n5014);
   U23890 : OAI21_X1 port map( B1 => n22188, B2 => n22189, A => n24793, ZN => 
                           n22187);
   U23891 : NAND4_X1 port map( A1 => n22198, A2 => n22199, A3 => n22200, A4 => 
                           n22201, ZN => n22188);
   U23892 : NAND4_X1 port map( A1 => n22190, A2 => n22191, A3 => n22192, A4 => 
                           n22193, ZN => n22189);
   U23893 : OAI221_X1 port map( B1 => n19248, B2 => n24805, C1 => n11802, C2 =>
                           n24801, A => n22168, ZN => n5015);
   U23894 : OAI21_X1 port map( B1 => n22169, B2 => n22170, A => n24793, ZN => 
                           n22168);
   U23895 : NAND4_X1 port map( A1 => n22179, A2 => n22180, A3 => n22181, A4 => 
                           n22182, ZN => n22169);
   U23896 : NAND4_X1 port map( A1 => n22171, A2 => n22172, A3 => n22173, A4 => 
                           n22174, ZN => n22170);
   U23897 : OAI221_X1 port map( B1 => n19247, B2 => n24805, C1 => n11803, C2 =>
                           n24801, A => n22149, ZN => n5016);
   U23898 : OAI21_X1 port map( B1 => n22150, B2 => n22151, A => n24793, ZN => 
                           n22149);
   U23899 : NAND4_X1 port map( A1 => n22160, A2 => n22161, A3 => n22162, A4 => 
                           n22163, ZN => n22150);
   U23900 : NAND4_X1 port map( A1 => n22152, A2 => n22153, A3 => n22154, A4 => 
                           n22155, ZN => n22151);
   U23901 : OAI221_X1 port map( B1 => n19246, B2 => n24805, C1 => n11804, C2 =>
                           n24801, A => n22130, ZN => n5017);
   U23902 : OAI21_X1 port map( B1 => n22131, B2 => n22132, A => n24793, ZN => 
                           n22130);
   U23903 : NAND4_X1 port map( A1 => n22141, A2 => n22142, A3 => n22143, A4 => 
                           n22144, ZN => n22131);
   U23904 : NAND4_X1 port map( A1 => n22133, A2 => n22134, A3 => n22135, A4 => 
                           n22136, ZN => n22132);
   U23905 : OAI221_X1 port map( B1 => n19245, B2 => n24805, C1 => n11805, C2 =>
                           n24801, A => n22111, ZN => n5018);
   U23906 : OAI21_X1 port map( B1 => n22112, B2 => n22113, A => n24793, ZN => 
                           n22111);
   U23907 : NAND4_X1 port map( A1 => n22122, A2 => n22123, A3 => n22124, A4 => 
                           n22125, ZN => n22112);
   U23908 : NAND4_X1 port map( A1 => n22114, A2 => n22115, A3 => n22116, A4 => 
                           n22117, ZN => n22113);
   U23909 : OAI221_X1 port map( B1 => n19244, B2 => n24805, C1 => n11806, C2 =>
                           n24801, A => n22092, ZN => n5019);
   U23910 : OAI21_X1 port map( B1 => n22093, B2 => n22094, A => n24793, ZN => 
                           n22092);
   U23911 : NAND4_X1 port map( A1 => n22103, A2 => n22104, A3 => n22105, A4 => 
                           n22106, ZN => n22093);
   U23912 : NAND4_X1 port map( A1 => n22095, A2 => n22096, A3 => n22097, A4 => 
                           n22098, ZN => n22094);
   U23913 : OAI221_X1 port map( B1 => n19243, B2 => n24806, C1 => n11807, C2 =>
                           n24801, A => n22073, ZN => n5020);
   U23914 : OAI21_X1 port map( B1 => n22074, B2 => n22075, A => n24794, ZN => 
                           n22073);
   U23915 : NAND4_X1 port map( A1 => n22084, A2 => n22085, A3 => n22086, A4 => 
                           n22087, ZN => n22074);
   U23916 : NAND4_X1 port map( A1 => n22076, A2 => n22077, A3 => n22078, A4 => 
                           n22079, ZN => n22075);
   U23917 : OAI221_X1 port map( B1 => n19242, B2 => n24806, C1 => n11808, C2 =>
                           n24801, A => n22054, ZN => n5021);
   U23918 : OAI21_X1 port map( B1 => n22055, B2 => n22056, A => n24794, ZN => 
                           n22054);
   U23919 : NAND4_X1 port map( A1 => n22065, A2 => n22066, A3 => n22067, A4 => 
                           n22068, ZN => n22055);
   U23920 : NAND4_X1 port map( A1 => n22057, A2 => n22058, A3 => n22059, A4 => 
                           n22060, ZN => n22056);
   U23921 : OAI221_X1 port map( B1 => n19241, B2 => n24806, C1 => n11809, C2 =>
                           n24801, A => n22035, ZN => n5022);
   U23922 : OAI21_X1 port map( B1 => n22036, B2 => n22037, A => n24794, ZN => 
                           n22035);
   U23923 : NAND4_X1 port map( A1 => n22046, A2 => n22047, A3 => n22048, A4 => 
                           n22049, ZN => n22036);
   U23924 : NAND4_X1 port map( A1 => n22038, A2 => n22039, A3 => n22040, A4 => 
                           n22041, ZN => n22037);
   U23925 : OAI221_X1 port map( B1 => n19240, B2 => n24806, C1 => n11810, C2 =>
                           n24801, A => n22016, ZN => n5023);
   U23926 : OAI21_X1 port map( B1 => n22017, B2 => n22018, A => n24794, ZN => 
                           n22016);
   U23927 : NAND4_X1 port map( A1 => n22027, A2 => n22028, A3 => n22029, A4 => 
                           n22030, ZN => n22017);
   U23928 : NAND4_X1 port map( A1 => n22019, A2 => n22020, A3 => n22021, A4 => 
                           n22022, ZN => n22018);
   U23929 : OAI221_X1 port map( B1 => n19239, B2 => n24806, C1 => n11811, C2 =>
                           n24800, A => n21997, ZN => n5024);
   U23930 : OAI21_X1 port map( B1 => n21998, B2 => n21999, A => n24794, ZN => 
                           n21997);
   U23931 : NAND4_X1 port map( A1 => n22008, A2 => n22009, A3 => n22010, A4 => 
                           n22011, ZN => n21998);
   U23932 : NAND4_X1 port map( A1 => n22000, A2 => n22001, A3 => n22002, A4 => 
                           n22003, ZN => n21999);
   U23933 : OAI221_X1 port map( B1 => n19238, B2 => n24806, C1 => n11812, C2 =>
                           n24800, A => n21978, ZN => n5025);
   U23934 : OAI21_X1 port map( B1 => n21979, B2 => n21980, A => n24794, ZN => 
                           n21978);
   U23935 : NAND4_X1 port map( A1 => n21989, A2 => n21990, A3 => n21991, A4 => 
                           n21992, ZN => n21979);
   U23936 : NAND4_X1 port map( A1 => n21981, A2 => n21982, A3 => n21983, A4 => 
                           n21984, ZN => n21980);
   U23937 : OAI221_X1 port map( B1 => n19237, B2 => n24806, C1 => n11813, C2 =>
                           n24800, A => n21959, ZN => n5026);
   U23938 : OAI21_X1 port map( B1 => n21960, B2 => n21961, A => n24794, ZN => 
                           n21959);
   U23939 : NAND4_X1 port map( A1 => n21970, A2 => n21971, A3 => n21972, A4 => 
                           n21973, ZN => n21960);
   U23940 : NAND4_X1 port map( A1 => n21962, A2 => n21963, A3 => n21964, A4 => 
                           n21965, ZN => n21961);
   U23941 : OAI221_X1 port map( B1 => n19236, B2 => n24806, C1 => n11814, C2 =>
                           n24800, A => n21940, ZN => n5027);
   U23942 : OAI21_X1 port map( B1 => n21941, B2 => n21942, A => n24794, ZN => 
                           n21940);
   U23943 : NAND4_X1 port map( A1 => n21951, A2 => n21952, A3 => n21953, A4 => 
                           n21954, ZN => n21941);
   U23944 : NAND4_X1 port map( A1 => n21943, A2 => n21944, A3 => n21945, A4 => 
                           n21946, ZN => n21942);
   U23945 : OAI221_X1 port map( B1 => n19235, B2 => n24806, C1 => n11815, C2 =>
                           n24800, A => n21921, ZN => n5028);
   U23946 : OAI21_X1 port map( B1 => n21922, B2 => n21923, A => n24794, ZN => 
                           n21921);
   U23947 : NAND4_X1 port map( A1 => n21932, A2 => n21933, A3 => n21934, A4 => 
                           n21935, ZN => n21922);
   U23948 : NAND4_X1 port map( A1 => n21924, A2 => n21925, A3 => n21926, A4 => 
                           n21927, ZN => n21923);
   U23949 : OAI221_X1 port map( B1 => n19234, B2 => n24806, C1 => n11816, C2 =>
                           n24800, A => n21902, ZN => n5029);
   U23950 : OAI21_X1 port map( B1 => n21903, B2 => n21904, A => n24794, ZN => 
                           n21902);
   U23951 : NAND4_X1 port map( A1 => n21913, A2 => n21914, A3 => n21915, A4 => 
                           n21916, ZN => n21903);
   U23952 : NAND4_X1 port map( A1 => n21905, A2 => n21906, A3 => n21907, A4 => 
                           n21908, ZN => n21904);
   U23953 : OAI221_X1 port map( B1 => n19233, B2 => n24806, C1 => n11817, C2 =>
                           n24800, A => n21883, ZN => n5030);
   U23954 : OAI21_X1 port map( B1 => n21884, B2 => n21885, A => n24794, ZN => 
                           n21883);
   U23955 : NAND4_X1 port map( A1 => n21894, A2 => n21895, A3 => n21896, A4 => 
                           n21897, ZN => n21884);
   U23956 : NAND4_X1 port map( A1 => n21886, A2 => n21887, A3 => n21888, A4 => 
                           n21889, ZN => n21885);
   U23957 : OAI221_X1 port map( B1 => n19232, B2 => n24806, C1 => n11818, C2 =>
                           n24800, A => n21864, ZN => n5031);
   U23958 : OAI21_X1 port map( B1 => n21865, B2 => n21866, A => n24794, ZN => 
                           n21864);
   U23959 : NAND4_X1 port map( A1 => n21875, A2 => n21876, A3 => n21877, A4 => 
                           n21878, ZN => n21865);
   U23960 : NAND4_X1 port map( A1 => n21867, A2 => n21868, A3 => n21869, A4 => 
                           n21870, ZN => n21866);
   U23961 : OAI221_X1 port map( B1 => n19231, B2 => n24807, C1 => n11819, C2 =>
                           n24800, A => n21845, ZN => n5032);
   U23962 : OAI21_X1 port map( B1 => n21846, B2 => n21847, A => n24795, ZN => 
                           n21845);
   U23963 : NAND4_X1 port map( A1 => n21856, A2 => n21857, A3 => n21858, A4 => 
                           n21859, ZN => n21846);
   U23964 : NAND4_X1 port map( A1 => n21848, A2 => n21849, A3 => n21850, A4 => 
                           n21851, ZN => n21847);
   U23965 : OAI221_X1 port map( B1 => n19230, B2 => n24807, C1 => n11820, C2 =>
                           n24800, A => n21826, ZN => n5033);
   U23966 : OAI21_X1 port map( B1 => n21827, B2 => n21828, A => n24795, ZN => 
                           n21826);
   U23967 : NAND4_X1 port map( A1 => n21837, A2 => n21838, A3 => n21839, A4 => 
                           n21840, ZN => n21827);
   U23968 : NAND4_X1 port map( A1 => n21829, A2 => n21830, A3 => n21831, A4 => 
                           n21832, ZN => n21828);
   U23969 : OAI221_X1 port map( B1 => n19229, B2 => n24807, C1 => n11821, C2 =>
                           n24800, A => n21807, ZN => n5034);
   U23970 : OAI21_X1 port map( B1 => n21808, B2 => n21809, A => n24795, ZN => 
                           n21807);
   U23971 : NAND4_X1 port map( A1 => n21818, A2 => n21819, A3 => n21820, A4 => 
                           n21821, ZN => n21808);
   U23972 : NAND4_X1 port map( A1 => n21810, A2 => n21811, A3 => n21812, A4 => 
                           n21813, ZN => n21809);
   U23973 : OAI221_X1 port map( B1 => n19228, B2 => n24807, C1 => n11822, C2 =>
                           n24799, A => n21788, ZN => n5035);
   U23974 : OAI21_X1 port map( B1 => n21789, B2 => n21790, A => n24795, ZN => 
                           n21788);
   U23975 : NAND4_X1 port map( A1 => n21799, A2 => n21800, A3 => n21801, A4 => 
                           n21802, ZN => n21789);
   U23976 : NAND4_X1 port map( A1 => n21791, A2 => n21792, A3 => n21793, A4 => 
                           n21794, ZN => n21790);
   U23977 : OAI221_X1 port map( B1 => n19227, B2 => n24807, C1 => n11823, C2 =>
                           n24799, A => n21769, ZN => n5036);
   U23978 : OAI21_X1 port map( B1 => n21770, B2 => n21771, A => n24795, ZN => 
                           n21769);
   U23979 : NAND4_X1 port map( A1 => n21780, A2 => n21781, A3 => n21782, A4 => 
                           n21783, ZN => n21770);
   U23980 : NAND4_X1 port map( A1 => n21772, A2 => n21773, A3 => n21774, A4 => 
                           n21775, ZN => n21771);
   U23981 : OAI221_X1 port map( B1 => n19226, B2 => n24807, C1 => n11824, C2 =>
                           n24799, A => n21750, ZN => n5037);
   U23982 : OAI21_X1 port map( B1 => n21751, B2 => n21752, A => n24795, ZN => 
                           n21750);
   U23983 : NAND4_X1 port map( A1 => n21761, A2 => n21762, A3 => n21763, A4 => 
                           n21764, ZN => n21751);
   U23984 : NAND4_X1 port map( A1 => n21753, A2 => n21754, A3 => n21755, A4 => 
                           n21756, ZN => n21752);
   U23985 : OAI221_X1 port map( B1 => n19225, B2 => n24807, C1 => n11825, C2 =>
                           n24799, A => n21731, ZN => n5038);
   U23986 : OAI21_X1 port map( B1 => n21732, B2 => n21733, A => n24795, ZN => 
                           n21731);
   U23987 : NAND4_X1 port map( A1 => n21742, A2 => n21743, A3 => n21744, A4 => 
                           n21745, ZN => n21732);
   U23988 : NAND4_X1 port map( A1 => n21734, A2 => n21735, A3 => n21736, A4 => 
                           n21737, ZN => n21733);
   U23989 : OAI221_X1 port map( B1 => n19224, B2 => n24807, C1 => n11826, C2 =>
                           n24799, A => n21712, ZN => n5039);
   U23990 : OAI21_X1 port map( B1 => n21713, B2 => n21714, A => n24795, ZN => 
                           n21712);
   U23991 : NAND4_X1 port map( A1 => n21723, A2 => n21724, A3 => n21725, A4 => 
                           n21726, ZN => n21713);
   U23992 : NAND4_X1 port map( A1 => n21715, A2 => n21716, A3 => n21717, A4 => 
                           n21718, ZN => n21714);
   U23993 : OAI221_X1 port map( B1 => n19223, B2 => n24807, C1 => n11827, C2 =>
                           n24799, A => n21693, ZN => n5040);
   U23994 : OAI21_X1 port map( B1 => n21694, B2 => n21695, A => n24795, ZN => 
                           n21693);
   U23995 : NAND4_X1 port map( A1 => n21704, A2 => n21705, A3 => n21706, A4 => 
                           n21707, ZN => n21694);
   U23996 : NAND4_X1 port map( A1 => n21696, A2 => n21697, A3 => n21698, A4 => 
                           n21699, ZN => n21695);
   U23997 : OAI221_X1 port map( B1 => n19222, B2 => n24807, C1 => n11828, C2 =>
                           n24799, A => n21674, ZN => n5041);
   U23998 : OAI21_X1 port map( B1 => n21675, B2 => n21676, A => n24795, ZN => 
                           n21674);
   U23999 : NAND4_X1 port map( A1 => n21685, A2 => n21686, A3 => n21687, A4 => 
                           n21688, ZN => n21675);
   U24000 : NAND4_X1 port map( A1 => n21677, A2 => n21678, A3 => n21679, A4 => 
                           n21680, ZN => n21676);
   U24001 : OAI221_X1 port map( B1 => n19221, B2 => n24807, C1 => n11829, C2 =>
                           n24799, A => n21655, ZN => n5042);
   U24002 : OAI21_X1 port map( B1 => n21656, B2 => n21657, A => n24795, ZN => 
                           n21655);
   U24003 : NAND4_X1 port map( A1 => n21666, A2 => n21667, A3 => n21668, A4 => 
                           n21669, ZN => n21656);
   U24004 : NAND4_X1 port map( A1 => n21658, A2 => n21659, A3 => n21660, A4 => 
                           n21661, ZN => n21657);
   U24005 : OAI221_X1 port map( B1 => n19220, B2 => n24807, C1 => n11830, C2 =>
                           n24799, A => n21636, ZN => n5043);
   U24006 : OAI21_X1 port map( B1 => n21637, B2 => n21638, A => n24795, ZN => 
                           n21636);
   U24007 : NAND4_X1 port map( A1 => n21647, A2 => n21648, A3 => n21649, A4 => 
                           n21650, ZN => n21637);
   U24008 : NAND4_X1 port map( A1 => n21639, A2 => n21640, A3 => n21641, A4 => 
                           n21642, ZN => n21638);
   U24009 : OAI221_X1 port map( B1 => n19219, B2 => n24808, C1 => n11831, C2 =>
                           n24799, A => n21617, ZN => n5044);
   U24010 : OAI21_X1 port map( B1 => n21618, B2 => n21619, A => n24796, ZN => 
                           n21617);
   U24011 : NAND4_X1 port map( A1 => n21628, A2 => n21629, A3 => n21630, A4 => 
                           n21631, ZN => n21618);
   U24012 : NAND4_X1 port map( A1 => n21620, A2 => n21621, A3 => n21622, A4 => 
                           n21623, ZN => n21619);
   U24013 : OAI221_X1 port map( B1 => n19218, B2 => n24808, C1 => n11832, C2 =>
                           n24799, A => n21598, ZN => n5045);
   U24014 : OAI21_X1 port map( B1 => n21599, B2 => n21600, A => n24796, ZN => 
                           n21598);
   U24015 : NAND4_X1 port map( A1 => n21609, A2 => n21610, A3 => n21611, A4 => 
                           n21612, ZN => n21599);
   U24016 : NAND4_X1 port map( A1 => n21601, A2 => n21602, A3 => n21603, A4 => 
                           n21604, ZN => n21600);
   U24017 : OAI221_X1 port map( B1 => n19217, B2 => n24808, C1 => n11833, C2 =>
                           n24799, A => n21579, ZN => n5046);
   U24018 : OAI21_X1 port map( B1 => n21580, B2 => n21581, A => n24796, ZN => 
                           n21579);
   U24019 : NAND4_X1 port map( A1 => n21590, A2 => n21591, A3 => n21592, A4 => 
                           n21593, ZN => n21580);
   U24020 : NAND4_X1 port map( A1 => n21582, A2 => n21583, A3 => n21584, A4 => 
                           n21585, ZN => n21581);
   U24021 : OAI221_X1 port map( B1 => n19216, B2 => n24808, C1 => n11834, C2 =>
                           n24798, A => n21560, ZN => n5047);
   U24022 : OAI21_X1 port map( B1 => n21561, B2 => n21562, A => n24796, ZN => 
                           n21560);
   U24023 : NAND4_X1 port map( A1 => n21571, A2 => n21572, A3 => n21573, A4 => 
                           n21574, ZN => n21561);
   U24024 : NAND4_X1 port map( A1 => n21563, A2 => n21564, A3 => n21565, A4 => 
                           n21566, ZN => n21562);
   U24025 : OAI221_X1 port map( B1 => n19215, B2 => n24808, C1 => n11835, C2 =>
                           n24798, A => n21541, ZN => n5048);
   U24026 : OAI21_X1 port map( B1 => n21542, B2 => n21543, A => n24796, ZN => 
                           n21541);
   U24027 : NAND4_X1 port map( A1 => n21552, A2 => n21553, A3 => n21554, A4 => 
                           n21555, ZN => n21542);
   U24028 : NAND4_X1 port map( A1 => n21544, A2 => n21545, A3 => n21546, A4 => 
                           n21547, ZN => n21543);
   U24029 : OAI221_X1 port map( B1 => n19214, B2 => n24808, C1 => n11836, C2 =>
                           n24798, A => n21522, ZN => n5049);
   U24030 : OAI21_X1 port map( B1 => n21523, B2 => n21524, A => n24796, ZN => 
                           n21522);
   U24031 : NAND4_X1 port map( A1 => n21533, A2 => n21534, A3 => n21535, A4 => 
                           n21536, ZN => n21523);
   U24032 : NAND4_X1 port map( A1 => n21525, A2 => n21526, A3 => n21527, A4 => 
                           n21528, ZN => n21524);
   U24033 : OAI221_X1 port map( B1 => n19213, B2 => n24808, C1 => n11837, C2 =>
                           n24798, A => n21503, ZN => n5050);
   U24034 : OAI21_X1 port map( B1 => n21504, B2 => n21505, A => n24796, ZN => 
                           n21503);
   U24035 : NAND4_X1 port map( A1 => n21514, A2 => n21515, A3 => n21516, A4 => 
                           n21517, ZN => n21504);
   U24036 : NAND4_X1 port map( A1 => n21506, A2 => n21507, A3 => n21508, A4 => 
                           n21509, ZN => n21505);
   U24037 : OAI221_X1 port map( B1 => n19212, B2 => n24808, C1 => n11838, C2 =>
                           n24798, A => n21484, ZN => n5051);
   U24038 : OAI21_X1 port map( B1 => n21485, B2 => n21486, A => n24796, ZN => 
                           n21484);
   U24039 : NAND4_X1 port map( A1 => n21495, A2 => n21496, A3 => n21497, A4 => 
                           n21498, ZN => n21485);
   U24040 : NAND4_X1 port map( A1 => n21487, A2 => n21488, A3 => n21489, A4 => 
                           n21490, ZN => n21486);
   U24041 : OAI221_X1 port map( B1 => n19211, B2 => n24808, C1 => n11839, C2 =>
                           n24798, A => n21465, ZN => n5052);
   U24042 : OAI21_X1 port map( B1 => n21466, B2 => n21467, A => n24796, ZN => 
                           n21465);
   U24043 : NAND4_X1 port map( A1 => n21476, A2 => n21477, A3 => n21478, A4 => 
                           n21479, ZN => n21466);
   U24044 : NAND4_X1 port map( A1 => n21468, A2 => n21469, A3 => n21470, A4 => 
                           n21471, ZN => n21467);
   U24045 : OAI221_X1 port map( B1 => n19210, B2 => n24808, C1 => n11840, C2 =>
                           n24798, A => n21446, ZN => n5053);
   U24046 : OAI21_X1 port map( B1 => n21447, B2 => n21448, A => n24796, ZN => 
                           n21446);
   U24047 : NAND4_X1 port map( A1 => n21457, A2 => n21458, A3 => n21459, A4 => 
                           n21460, ZN => n21447);
   U24048 : NAND4_X1 port map( A1 => n21449, A2 => n21450, A3 => n21451, A4 => 
                           n21452, ZN => n21448);
   U24049 : OAI221_X1 port map( B1 => n19209, B2 => n24808, C1 => n11841, C2 =>
                           n24798, A => n21427, ZN => n5054);
   U24050 : OAI21_X1 port map( B1 => n21428, B2 => n21429, A => n24796, ZN => 
                           n21427);
   U24051 : NAND4_X1 port map( A1 => n21438, A2 => n21439, A3 => n21440, A4 => 
                           n21441, ZN => n21428);
   U24052 : NAND4_X1 port map( A1 => n21430, A2 => n21431, A3 => n21432, A4 => 
                           n21433, ZN => n21429);
   U24053 : OAI221_X1 port map( B1 => n19208, B2 => n24808, C1 => n11842, C2 =>
                           n24798, A => n21408, ZN => n5055);
   U24054 : OAI21_X1 port map( B1 => n21409, B2 => n21410, A => n24796, ZN => 
                           n21408);
   U24055 : NAND4_X1 port map( A1 => n21419, A2 => n21420, A3 => n21421, A4 => 
                           n21422, ZN => n21409);
   U24056 : NAND4_X1 port map( A1 => n21411, A2 => n21412, A3 => n21413, A4 => 
                           n21414, ZN => n21410);
   U24057 : NAND4_X1 port map( A1 => n23008, A2 => n23009, A3 => n23010, A4 => 
                           n23011, ZN => n4972);
   U24058 : AOI221_X1 port map( B1 => n24441, B2 => n24332, C1 => n24435, C2 =>
                           n19877, A => n23024, ZN => n23009);
   U24059 : AOI221_X1 port map( B1 => n24417, B2 => n19483, C1 => n24410, C2 =>
                           OUT2_40_port, A => n23025, ZN => n23008);
   U24060 : NOR4_X1 port map( A1 => n23020, A2 => n23021, A3 => n23022, A4 => 
                           n23023, ZN => n23010);
   U24061 : NAND4_X1 port map( A1 => n22990, A2 => n22991, A3 => n22992, A4 => 
                           n22993, ZN => n4973);
   U24062 : AOI221_X1 port map( B1 => n24441, B2 => n24333, C1 => n24435, C2 =>
                           n19876, A => n23006, ZN => n22991);
   U24063 : AOI221_X1 port map( B1 => n24417, B2 => n19482, C1 => n24409, C2 =>
                           OUT2_41_port, A => n23007, ZN => n22990);
   U24064 : NOR4_X1 port map( A1 => n23002, A2 => n23003, A3 => n23004, A4 => 
                           n23005, ZN => n22992);
   U24065 : NAND4_X1 port map( A1 => n22972, A2 => n22973, A3 => n22974, A4 => 
                           n22975, ZN => n4974);
   U24066 : AOI221_X1 port map( B1 => n24441, B2 => n24334, C1 => n24435, C2 =>
                           n19875, A => n22988, ZN => n22973);
   U24067 : AOI221_X1 port map( B1 => n24417, B2 => n19481, C1 => n24409, C2 =>
                           OUT2_42_port, A => n22989, ZN => n22972);
   U24068 : NOR4_X1 port map( A1 => n22984, A2 => n22985, A3 => n22986, A4 => 
                           n22987, ZN => n22974);
   U24069 : NAND4_X1 port map( A1 => n22954, A2 => n22955, A3 => n22956, A4 => 
                           n22957, ZN => n4975);
   U24070 : AOI221_X1 port map( B1 => n24441, B2 => n24335, C1 => n24435, C2 =>
                           n19874, A => n22970, ZN => n22955);
   U24071 : AOI221_X1 port map( B1 => n24417, B2 => n19480, C1 => n24409, C2 =>
                           OUT2_43_port, A => n22971, ZN => n22954);
   U24072 : NOR4_X1 port map( A1 => n22966, A2 => n22967, A3 => n22968, A4 => 
                           n22969, ZN => n22956);
   U24073 : NAND4_X1 port map( A1 => n22936, A2 => n22937, A3 => n22938, A4 => 
                           n22939, ZN => n4976);
   U24074 : AOI221_X1 port map( B1 => n24441, B2 => n24336, C1 => n24435, C2 =>
                           n19873, A => n22952, ZN => n22937);
   U24075 : AOI221_X1 port map( B1 => n24417, B2 => n19479, C1 => n24409, C2 =>
                           OUT2_44_port, A => n22953, ZN => n22936);
   U24076 : NOR4_X1 port map( A1 => n22948, A2 => n22949, A3 => n22950, A4 => 
                           n22951, ZN => n22938);
   U24077 : NAND4_X1 port map( A1 => n22918, A2 => n22919, A3 => n22920, A4 => 
                           n22921, ZN => n4977);
   U24078 : AOI221_X1 port map( B1 => n24441, B2 => n24337, C1 => n24435, C2 =>
                           n19872, A => n22934, ZN => n22919);
   U24079 : AOI221_X1 port map( B1 => n24417, B2 => n19478, C1 => n24409, C2 =>
                           OUT2_45_port, A => n22935, ZN => n22918);
   U24080 : NOR4_X1 port map( A1 => n22930, A2 => n22931, A3 => n22932, A4 => 
                           n22933, ZN => n22920);
   U24081 : NAND4_X1 port map( A1 => n22900, A2 => n22901, A3 => n22902, A4 => 
                           n22903, ZN => n4978);
   U24082 : AOI221_X1 port map( B1 => n24441, B2 => n24338, C1 => n24435, C2 =>
                           n19871, A => n22916, ZN => n22901);
   U24083 : AOI221_X1 port map( B1 => n24417, B2 => n19477, C1 => n24409, C2 =>
                           OUT2_46_port, A => n22917, ZN => n22900);
   U24084 : NOR4_X1 port map( A1 => n22912, A2 => n22913, A3 => n22914, A4 => 
                           n22915, ZN => n22902);
   U24085 : NAND4_X1 port map( A1 => n22882, A2 => n22883, A3 => n22884, A4 => 
                           n22885, ZN => n4979);
   U24086 : AOI221_X1 port map( B1 => n24441, B2 => n24339, C1 => n24435, C2 =>
                           n19870, A => n22898, ZN => n22883);
   U24087 : AOI221_X1 port map( B1 => n24417, B2 => n19476, C1 => n24409, C2 =>
                           OUT2_47_port, A => n22899, ZN => n22882);
   U24088 : NOR4_X1 port map( A1 => n22894, A2 => n22895, A3 => n22896, A4 => 
                           n22897, ZN => n22884);
   U24089 : NAND4_X1 port map( A1 => n22864, A2 => n22865, A3 => n22866, A4 => 
                           n22867, ZN => n4980);
   U24090 : AOI221_X1 port map( B1 => n24442, B2 => n24340, C1 => n24436, C2 =>
                           n19869, A => n22880, ZN => n22865);
   U24091 : AOI221_X1 port map( B1 => n24418, B2 => n19475, C1 => n24409, C2 =>
                           OUT2_48_port, A => n22881, ZN => n22864);
   U24092 : NOR4_X1 port map( A1 => n22876, A2 => n22877, A3 => n22878, A4 => 
                           n22879, ZN => n22866);
   U24093 : NAND4_X1 port map( A1 => n22846, A2 => n22847, A3 => n22848, A4 => 
                           n22849, ZN => n4981);
   U24094 : AOI221_X1 port map( B1 => n24442, B2 => n24341, C1 => n24436, C2 =>
                           n19868, A => n22862, ZN => n22847);
   U24095 : AOI221_X1 port map( B1 => n24418, B2 => n19474, C1 => n24409, C2 =>
                           OUT2_49_port, A => n22863, ZN => n22846);
   U24096 : NOR4_X1 port map( A1 => n22858, A2 => n22859, A3 => n22860, A4 => 
                           n22861, ZN => n22848);
   U24097 : NAND4_X1 port map( A1 => n22828, A2 => n22829, A3 => n22830, A4 => 
                           n22831, ZN => n4982);
   U24098 : AOI221_X1 port map( B1 => n24442, B2 => n24342, C1 => n24436, C2 =>
                           n19867, A => n22844, ZN => n22829);
   U24099 : AOI221_X1 port map( B1 => n24418, B2 => n19473, C1 => n24409, C2 =>
                           OUT2_50_port, A => n22845, ZN => n22828);
   U24100 : NOR4_X1 port map( A1 => n22840, A2 => n22841, A3 => n22842, A4 => 
                           n22843, ZN => n22830);
   U24101 : NAND4_X1 port map( A1 => n22810, A2 => n22811, A3 => n22812, A4 => 
                           n22813, ZN => n4983);
   U24102 : AOI221_X1 port map( B1 => n24442, B2 => n24343, C1 => n24436, C2 =>
                           n19866, A => n22826, ZN => n22811);
   U24103 : AOI221_X1 port map( B1 => n24418, B2 => n19472, C1 => n24409, C2 =>
                           OUT2_51_port, A => n22827, ZN => n22810);
   U24104 : NOR4_X1 port map( A1 => n22822, A2 => n22823, A3 => n22824, A4 => 
                           n22825, ZN => n22812);
   U24105 : NAND4_X1 port map( A1 => n22792, A2 => n22793, A3 => n22794, A4 => 
                           n22795, ZN => n4984);
   U24106 : AOI221_X1 port map( B1 => n24442, B2 => n24344, C1 => n24436, C2 =>
                           n19865, A => n22808, ZN => n22793);
   U24107 : AOI221_X1 port map( B1 => n24418, B2 => n19471, C1 => n24409, C2 =>
                           OUT2_52_port, A => n22809, ZN => n22792);
   U24108 : NOR4_X1 port map( A1 => n22804, A2 => n22805, A3 => n22806, A4 => 
                           n22807, ZN => n22794);
   U24109 : NAND4_X1 port map( A1 => n22774, A2 => n22775, A3 => n22776, A4 => 
                           n22777, ZN => n4985);
   U24110 : AOI221_X1 port map( B1 => n24442, B2 => n24345, C1 => n24436, C2 =>
                           n19864, A => n22790, ZN => n22775);
   U24111 : AOI221_X1 port map( B1 => n24418, B2 => n19470, C1 => n24408, C2 =>
                           OUT2_53_port, A => n22791, ZN => n22774);
   U24112 : NOR4_X1 port map( A1 => n22786, A2 => n22787, A3 => n22788, A4 => 
                           n22789, ZN => n22776);
   U24113 : NAND4_X1 port map( A1 => n22756, A2 => n22757, A3 => n22758, A4 => 
                           n22759, ZN => n4986);
   U24114 : AOI221_X1 port map( B1 => n24442, B2 => n24346, C1 => n24436, C2 =>
                           n19863, A => n22772, ZN => n22757);
   U24115 : AOI221_X1 port map( B1 => n24418, B2 => n19469, C1 => n24408, C2 =>
                           OUT2_54_port, A => n22773, ZN => n22756);
   U24116 : NOR4_X1 port map( A1 => n22768, A2 => n22769, A3 => n22770, A4 => 
                           n22771, ZN => n22758);
   U24117 : NAND4_X1 port map( A1 => n22738, A2 => n22739, A3 => n22740, A4 => 
                           n22741, ZN => n4987);
   U24118 : AOI221_X1 port map( B1 => n24442, B2 => n24347, C1 => n24436, C2 =>
                           n19862, A => n22754, ZN => n22739);
   U24119 : AOI221_X1 port map( B1 => n24418, B2 => n19468, C1 => n24408, C2 =>
                           OUT2_55_port, A => n22755, ZN => n22738);
   U24120 : NOR4_X1 port map( A1 => n22750, A2 => n22751, A3 => n22752, A4 => 
                           n22753, ZN => n22740);
   U24121 : NAND4_X1 port map( A1 => n22720, A2 => n22721, A3 => n22722, A4 => 
                           n22723, ZN => n4988);
   U24122 : AOI221_X1 port map( B1 => n24442, B2 => n24348, C1 => n24436, C2 =>
                           n19861, A => n22736, ZN => n22721);
   U24123 : AOI221_X1 port map( B1 => n24418, B2 => n19467, C1 => n24408, C2 =>
                           OUT2_56_port, A => n22737, ZN => n22720);
   U24124 : NOR4_X1 port map( A1 => n22732, A2 => n22733, A3 => n22734, A4 => 
                           n22735, ZN => n22722);
   U24125 : NAND4_X1 port map( A1 => n22702, A2 => n22703, A3 => n22704, A4 => 
                           n22705, ZN => n4989);
   U24126 : AOI221_X1 port map( B1 => n24442, B2 => n24349, C1 => n24436, C2 =>
                           n19860, A => n22718, ZN => n22703);
   U24127 : AOI221_X1 port map( B1 => n24418, B2 => n19466, C1 => n24408, C2 =>
                           OUT2_57_port, A => n22719, ZN => n22702);
   U24128 : NOR4_X1 port map( A1 => n22714, A2 => n22715, A3 => n22716, A4 => 
                           n22717, ZN => n22704);
   U24129 : NAND4_X1 port map( A1 => n22684, A2 => n22685, A3 => n22686, A4 => 
                           n22687, ZN => n4990);
   U24130 : AOI221_X1 port map( B1 => n24442, B2 => n24350, C1 => n24436, C2 =>
                           n19859, A => n22700, ZN => n22685);
   U24131 : AOI221_X1 port map( B1 => n24418, B2 => n19465, C1 => n24408, C2 =>
                           OUT2_58_port, A => n22701, ZN => n22684);
   U24132 : NOR4_X1 port map( A1 => n22696, A2 => n22697, A3 => n22698, A4 => 
                           n22699, ZN => n22686);
   U24133 : NAND4_X1 port map( A1 => n22666, A2 => n22667, A3 => n22668, A4 => 
                           n22669, ZN => n4991);
   U24134 : AOI221_X1 port map( B1 => n24442, B2 => n24351, C1 => n24436, C2 =>
                           n19858, A => n22682, ZN => n22667);
   U24135 : AOI221_X1 port map( B1 => n24418, B2 => n19464, C1 => n24408, C2 =>
                           OUT2_59_port, A => n22683, ZN => n22666);
   U24136 : NOR4_X1 port map( A1 => n22678, A2 => n22679, A3 => n22680, A4 => 
                           n22681, ZN => n22668);
   U24137 : NAND4_X1 port map( A1 => n22648, A2 => n22649, A3 => n22650, A4 => 
                           n22651, ZN => n4992);
   U24138 : AOI221_X1 port map( B1 => n24443, B2 => n24352, C1 => n24437, C2 =>
                           n19809, A => n22664, ZN => n22649);
   U24139 : AOI221_X1 port map( B1 => n24419, B2 => n19463, C1 => n24408, C2 =>
                           OUT2_60_port, A => n22665, ZN => n22648);
   U24140 : NOR4_X1 port map( A1 => n22660, A2 => n22661, A3 => n22662, A4 => 
                           n22663, ZN => n22650);
   U24141 : NAND4_X1 port map( A1 => n22630, A2 => n22631, A3 => n22632, A4 => 
                           n22633, ZN => n4993);
   U24142 : AOI221_X1 port map( B1 => n24443, B2 => n24353, C1 => n24437, C2 =>
                           n19808, A => n22646, ZN => n22631);
   U24143 : AOI221_X1 port map( B1 => n24419, B2 => n19462, C1 => n24408, C2 =>
                           OUT2_61_port, A => n22647, ZN => n22630);
   U24144 : NOR4_X1 port map( A1 => n22642, A2 => n22643, A3 => n22644, A4 => 
                           n22645, ZN => n22632);
   U24145 : NAND4_X1 port map( A1 => n22612, A2 => n22613, A3 => n22614, A4 => 
                           n22615, ZN => n4994);
   U24146 : AOI221_X1 port map( B1 => n24443, B2 => n24354, C1 => n24437, C2 =>
                           n19807, A => n22628, ZN => n22613);
   U24147 : AOI221_X1 port map( B1 => n24419, B2 => n19461, C1 => n24408, C2 =>
                           OUT2_62_port, A => n22629, ZN => n22612);
   U24148 : NOR4_X1 port map( A1 => n22624, A2 => n22625, A3 => n22626, A4 => 
                           n22627, ZN => n22614);
   U24149 : NAND4_X1 port map( A1 => n22560, A2 => n22561, A3 => n22562, A4 => 
                           n22563, ZN => n4995);
   U24150 : AOI221_X1 port map( B1 => n24443, B2 => n24355, C1 => n24437, C2 =>
                           n19806, A => n22604, ZN => n22561);
   U24151 : AOI221_X1 port map( B1 => n24419, B2 => n19460, C1 => n24410, C2 =>
                           OUT2_63_port, A => n22609, ZN => n22560);
   U24152 : NOR4_X1 port map( A1 => n22589, A2 => n22590, A3 => n22591, A4 => 
                           n22592, ZN => n22562);
   U24153 : NAND4_X1 port map( A1 => n23728, A2 => n23729, A3 => n23730, A4 => 
                           n23731, ZN => n4932);
   U24154 : AOI221_X1 port map( B1 => n24438, B2 => n24356, C1 => n24432, C2 =>
                           n20049, A => n23762, ZN => n23729);
   U24155 : AOI221_X1 port map( B1 => n24414, B2 => n19523, C1 => n24408, C2 =>
                           OUT2_0_port, A => n23763, ZN => n23728);
   U24156 : NOR4_X1 port map( A1 => n23750, A2 => n23751, A3 => n23752, A4 => 
                           n23753, ZN => n23730);
   U24157 : NAND4_X1 port map( A1 => n23710, A2 => n23711, A3 => n23712, A4 => 
                           n23713, ZN => n4933);
   U24158 : AOI221_X1 port map( B1 => n24438, B2 => n24357, C1 => n24432, C2 =>
                           n20048, A => n23726, ZN => n23711);
   U24159 : AOI221_X1 port map( B1 => n24414, B2 => n19522, C1 => n24413, C2 =>
                           OUT2_1_port, A => n23727, ZN => n23710);
   U24160 : NOR4_X1 port map( A1 => n23722, A2 => n23723, A3 => n23724, A4 => 
                           n23725, ZN => n23712);
   U24161 : NAND4_X1 port map( A1 => n23692, A2 => n23693, A3 => n23694, A4 => 
                           n23695, ZN => n4934);
   U24162 : AOI221_X1 port map( B1 => n24438, B2 => n24358, C1 => n24432, C2 =>
                           n20047, A => n23708, ZN => n23693);
   U24163 : AOI221_X1 port map( B1 => n24414, B2 => n19521, C1 => n24413, C2 =>
                           OUT2_2_port, A => n23709, ZN => n23692);
   U24164 : NOR4_X1 port map( A1 => n23704, A2 => n23705, A3 => n23706, A4 => 
                           n23707, ZN => n23694);
   U24165 : NAND4_X1 port map( A1 => n23674, A2 => n23675, A3 => n23676, A4 => 
                           n23677, ZN => n4935);
   U24166 : AOI221_X1 port map( B1 => n24438, B2 => n24359, C1 => n24432, C2 =>
                           n20046, A => n23690, ZN => n23675);
   U24167 : AOI221_X1 port map( B1 => n24414, B2 => n19520, C1 => n24413, C2 =>
                           OUT2_3_port, A => n23691, ZN => n23674);
   U24168 : NOR4_X1 port map( A1 => n23686, A2 => n23687, A3 => n23688, A4 => 
                           n23689, ZN => n23676);
   U24169 : NAND4_X1 port map( A1 => n23656, A2 => n23657, A3 => n23658, A4 => 
                           n23659, ZN => n4936);
   U24170 : AOI221_X1 port map( B1 => n24438, B2 => n24360, C1 => n24432, C2 =>
                           n20045, A => n23672, ZN => n23657);
   U24171 : AOI221_X1 port map( B1 => n24414, B2 => n19519, C1 => n24413, C2 =>
                           OUT2_4_port, A => n23673, ZN => n23656);
   U24172 : NOR4_X1 port map( A1 => n23668, A2 => n23669, A3 => n23670, A4 => 
                           n23671, ZN => n23658);
   U24173 : NAND4_X1 port map( A1 => n23638, A2 => n23639, A3 => n23640, A4 => 
                           n23641, ZN => n4937);
   U24174 : AOI221_X1 port map( B1 => n24438, B2 => n24361, C1 => n24432, C2 =>
                           n20044, A => n23654, ZN => n23639);
   U24175 : AOI221_X1 port map( B1 => n24414, B2 => n19518, C1 => n24413, C2 =>
                           OUT2_5_port, A => n23655, ZN => n23638);
   U24176 : NOR4_X1 port map( A1 => n23650, A2 => n23651, A3 => n23652, A4 => 
                           n23653, ZN => n23640);
   U24177 : NAND4_X1 port map( A1 => n23620, A2 => n23621, A3 => n23622, A4 => 
                           n23623, ZN => n4938);
   U24178 : AOI221_X1 port map( B1 => n24438, B2 => n24362, C1 => n24432, C2 =>
                           n20043, A => n23636, ZN => n23621);
   U24179 : AOI221_X1 port map( B1 => n24414, B2 => n19517, C1 => n24412, C2 =>
                           OUT2_6_port, A => n23637, ZN => n23620);
   U24180 : NOR4_X1 port map( A1 => n23632, A2 => n23633, A3 => n23634, A4 => 
                           n23635, ZN => n23622);
   U24181 : NAND4_X1 port map( A1 => n23602, A2 => n23603, A3 => n23604, A4 => 
                           n23605, ZN => n4939);
   U24182 : AOI221_X1 port map( B1 => n24438, B2 => n24363, C1 => n24432, C2 =>
                           n20042, A => n23618, ZN => n23603);
   U24183 : AOI221_X1 port map( B1 => n24414, B2 => n19516, C1 => n24412, C2 =>
                           OUT2_7_port, A => n23619, ZN => n23602);
   U24184 : NOR4_X1 port map( A1 => n23614, A2 => n23615, A3 => n23616, A4 => 
                           n23617, ZN => n23604);
   U24185 : NAND4_X1 port map( A1 => n23584, A2 => n23585, A3 => n23586, A4 => 
                           n23587, ZN => n4940);
   U24186 : AOI221_X1 port map( B1 => n24438, B2 => n24364, C1 => n24432, C2 =>
                           n20041, A => n23600, ZN => n23585);
   U24187 : AOI221_X1 port map( B1 => n24414, B2 => n19515, C1 => n24412, C2 =>
                           OUT2_8_port, A => n23601, ZN => n23584);
   U24188 : NOR4_X1 port map( A1 => n23596, A2 => n23597, A3 => n23598, A4 => 
                           n23599, ZN => n23586);
   U24189 : NAND4_X1 port map( A1 => n23566, A2 => n23567, A3 => n23568, A4 => 
                           n23569, ZN => n4941);
   U24190 : AOI221_X1 port map( B1 => n24438, B2 => n24365, C1 => n24432, C2 =>
                           n20040, A => n23582, ZN => n23567);
   U24191 : AOI221_X1 port map( B1 => n24414, B2 => n19514, C1 => n24412, C2 =>
                           OUT2_9_port, A => n23583, ZN => n23566);
   U24192 : NOR4_X1 port map( A1 => n23578, A2 => n23579, A3 => n23580, A4 => 
                           n23581, ZN => n23568);
   U24193 : NAND4_X1 port map( A1 => n23548, A2 => n23549, A3 => n23550, A4 => 
                           n23551, ZN => n4942);
   U24194 : AOI221_X1 port map( B1 => n24438, B2 => n24366, C1 => n24432, C2 =>
                           n20039, A => n23564, ZN => n23549);
   U24195 : AOI221_X1 port map( B1 => n24414, B2 => n19513, C1 => n24412, C2 =>
                           OUT2_10_port, A => n23565, ZN => n23548);
   U24196 : NOR4_X1 port map( A1 => n23560, A2 => n23561, A3 => n23562, A4 => 
                           n23563, ZN => n23550);
   U24197 : NAND4_X1 port map( A1 => n23530, A2 => n23531, A3 => n23532, A4 => 
                           n23533, ZN => n4943);
   U24198 : AOI221_X1 port map( B1 => n24438, B2 => n24367, C1 => n24432, C2 =>
                           n20038, A => n23546, ZN => n23531);
   U24199 : AOI221_X1 port map( B1 => n24414, B2 => n19512, C1 => n24412, C2 =>
                           OUT2_11_port, A => n23547, ZN => n23530);
   U24200 : NOR4_X1 port map( A1 => n23542, A2 => n23543, A3 => n23544, A4 => 
                           n23545, ZN => n23532);
   U24201 : NAND4_X1 port map( A1 => n23512, A2 => n23513, A3 => n23514, A4 => 
                           n23515, ZN => n4944);
   U24202 : AOI221_X1 port map( B1 => n24439, B2 => n24368, C1 => n24433, C2 =>
                           n20037, A => n23528, ZN => n23513);
   U24203 : AOI221_X1 port map( B1 => n24415, B2 => n19511, C1 => n24412, C2 =>
                           OUT2_12_port, A => n23529, ZN => n23512);
   U24204 : NOR4_X1 port map( A1 => n23524, A2 => n23525, A3 => n23526, A4 => 
                           n23527, ZN => n23514);
   U24205 : NAND4_X1 port map( A1 => n23494, A2 => n23495, A3 => n23496, A4 => 
                           n23497, ZN => n4945);
   U24206 : AOI221_X1 port map( B1 => n24439, B2 => n24369, C1 => n24433, C2 =>
                           n20036, A => n23510, ZN => n23495);
   U24207 : AOI221_X1 port map( B1 => n24415, B2 => n19510, C1 => n24412, C2 =>
                           OUT2_13_port, A => n23511, ZN => n23494);
   U24208 : NOR4_X1 port map( A1 => n23506, A2 => n23507, A3 => n23508, A4 => 
                           n23509, ZN => n23496);
   U24209 : NAND4_X1 port map( A1 => n23476, A2 => n23477, A3 => n23478, A4 => 
                           n23479, ZN => n4946);
   U24210 : AOI221_X1 port map( B1 => n24439, B2 => n24370, C1 => n24433, C2 =>
                           n20035, A => n23492, ZN => n23477);
   U24211 : AOI221_X1 port map( B1 => n24415, B2 => n19509, C1 => n24412, C2 =>
                           OUT2_14_port, A => n23493, ZN => n23476);
   U24212 : NOR4_X1 port map( A1 => n23488, A2 => n23489, A3 => n23490, A4 => 
                           n23491, ZN => n23478);
   U24213 : NAND4_X1 port map( A1 => n23458, A2 => n23459, A3 => n23460, A4 => 
                           n23461, ZN => n4947);
   U24214 : AOI221_X1 port map( B1 => n24439, B2 => n24371, C1 => n24433, C2 =>
                           n20034, A => n23474, ZN => n23459);
   U24215 : AOI221_X1 port map( B1 => n24415, B2 => n19508, C1 => n24412, C2 =>
                           OUT2_15_port, A => n23475, ZN => n23458);
   U24216 : NOR4_X1 port map( A1 => n23470, A2 => n23471, A3 => n23472, A4 => 
                           n23473, ZN => n23460);
   U24217 : NAND4_X1 port map( A1 => n23440, A2 => n23441, A3 => n23442, A4 => 
                           n23443, ZN => n4948);
   U24218 : AOI221_X1 port map( B1 => n24439, B2 => n24372, C1 => n24433, C2 =>
                           n20033, A => n23456, ZN => n23441);
   U24219 : AOI221_X1 port map( B1 => n24415, B2 => n19507, C1 => n24412, C2 =>
                           OUT2_16_port, A => n23457, ZN => n23440);
   U24220 : NOR4_X1 port map( A1 => n23452, A2 => n23453, A3 => n23454, A4 => 
                           n23455, ZN => n23442);
   U24221 : NAND4_X1 port map( A1 => n23422, A2 => n23423, A3 => n23424, A4 => 
                           n23425, ZN => n4949);
   U24222 : AOI221_X1 port map( B1 => n24439, B2 => n24373, C1 => n24433, C2 =>
                           n20032, A => n23438, ZN => n23423);
   U24223 : AOI221_X1 port map( B1 => n24415, B2 => n19506, C1 => n24412, C2 =>
                           OUT2_17_port, A => n23439, ZN => n23422);
   U24224 : NOR4_X1 port map( A1 => n23434, A2 => n23435, A3 => n23436, A4 => 
                           n23437, ZN => n23424);
   U24225 : NAND4_X1 port map( A1 => n23404, A2 => n23405, A3 => n23406, A4 => 
                           n23407, ZN => n4950);
   U24226 : AOI221_X1 port map( B1 => n24439, B2 => n24374, C1 => n24433, C2 =>
                           n20031, A => n23420, ZN => n23405);
   U24227 : AOI221_X1 port map( B1 => n24415, B2 => n19505, C1 => n24411, C2 =>
                           OUT2_18_port, A => n23421, ZN => n23404);
   U24228 : NOR4_X1 port map( A1 => n23416, A2 => n23417, A3 => n23418, A4 => 
                           n23419, ZN => n23406);
   U24229 : NAND4_X1 port map( A1 => n23386, A2 => n23387, A3 => n23388, A4 => 
                           n23389, ZN => n4951);
   U24230 : AOI221_X1 port map( B1 => n24439, B2 => n24375, C1 => n24433, C2 =>
                           n20030, A => n23402, ZN => n23387);
   U24231 : AOI221_X1 port map( B1 => n24415, B2 => n19504, C1 => n24411, C2 =>
                           OUT2_19_port, A => n23403, ZN => n23386);
   U24232 : NOR4_X1 port map( A1 => n23398, A2 => n23399, A3 => n23400, A4 => 
                           n23401, ZN => n23388);
   U24233 : NAND4_X1 port map( A1 => n23368, A2 => n23369, A3 => n23370, A4 => 
                           n23371, ZN => n4952);
   U24234 : AOI221_X1 port map( B1 => n24439, B2 => n24376, C1 => n24433, C2 =>
                           n20029, A => n23384, ZN => n23369);
   U24235 : AOI221_X1 port map( B1 => n24415, B2 => n19503, C1 => n24411, C2 =>
                           OUT2_20_port, A => n23385, ZN => n23368);
   U24236 : NOR4_X1 port map( A1 => n23380, A2 => n23381, A3 => n23382, A4 => 
                           n23383, ZN => n23370);
   U24237 : NAND4_X1 port map( A1 => n23350, A2 => n23351, A3 => n23352, A4 => 
                           n23353, ZN => n4953);
   U24238 : AOI221_X1 port map( B1 => n24439, B2 => n24377, C1 => n24433, C2 =>
                           n20028, A => n23366, ZN => n23351);
   U24239 : AOI221_X1 port map( B1 => n24415, B2 => n19502, C1 => n24411, C2 =>
                           OUT2_21_port, A => n23367, ZN => n23350);
   U24240 : NOR4_X1 port map( A1 => n23362, A2 => n23363, A3 => n23364, A4 => 
                           n23365, ZN => n23352);
   U24241 : NAND4_X1 port map( A1 => n23332, A2 => n23333, A3 => n23334, A4 => 
                           n23335, ZN => n4954);
   U24242 : AOI221_X1 port map( B1 => n24439, B2 => n24378, C1 => n24433, C2 =>
                           n20027, A => n23348, ZN => n23333);
   U24243 : AOI221_X1 port map( B1 => n24415, B2 => n19501, C1 => n24411, C2 =>
                           OUT2_22_port, A => n23349, ZN => n23332);
   U24244 : NOR4_X1 port map( A1 => n23344, A2 => n23345, A3 => n23346, A4 => 
                           n23347, ZN => n23334);
   U24245 : NAND4_X1 port map( A1 => n23314, A2 => n23315, A3 => n23316, A4 => 
                           n23317, ZN => n4955);
   U24246 : AOI221_X1 port map( B1 => n24439, B2 => n24379, C1 => n24433, C2 =>
                           n20026, A => n23330, ZN => n23315);
   U24247 : AOI221_X1 port map( B1 => n24415, B2 => n19500, C1 => n24411, C2 =>
                           OUT2_23_port, A => n23331, ZN => n23314);
   U24248 : NOR4_X1 port map( A1 => n23326, A2 => n23327, A3 => n23328, A4 => 
                           n23329, ZN => n23316);
   U24249 : NAND4_X1 port map( A1 => n23296, A2 => n23297, A3 => n23298, A4 => 
                           n23299, ZN => n4956);
   U24250 : AOI221_X1 port map( B1 => n24440, B2 => n24380, C1 => n24434, C2 =>
                           n19893, A => n23312, ZN => n23297);
   U24251 : AOI221_X1 port map( B1 => n24416, B2 => n19499, C1 => n24411, C2 =>
                           OUT2_24_port, A => n23313, ZN => n23296);
   U24252 : NOR4_X1 port map( A1 => n23308, A2 => n23309, A3 => n23310, A4 => 
                           n23311, ZN => n23298);
   U24253 : NAND4_X1 port map( A1 => n23278, A2 => n23279, A3 => n23280, A4 => 
                           n23281, ZN => n4957);
   U24254 : AOI221_X1 port map( B1 => n24440, B2 => n24381, C1 => n24434, C2 =>
                           n19892, A => n23294, ZN => n23279);
   U24255 : AOI221_X1 port map( B1 => n24416, B2 => n19498, C1 => n24411, C2 =>
                           OUT2_25_port, A => n23295, ZN => n23278);
   U24256 : NOR4_X1 port map( A1 => n23290, A2 => n23291, A3 => n23292, A4 => 
                           n23293, ZN => n23280);
   U24257 : NAND4_X1 port map( A1 => n23260, A2 => n23261, A3 => n23262, A4 => 
                           n23263, ZN => n4958);
   U24258 : AOI221_X1 port map( B1 => n24440, B2 => n24382, C1 => n24434, C2 =>
                           n19891, A => n23276, ZN => n23261);
   U24259 : AOI221_X1 port map( B1 => n24416, B2 => n19497, C1 => n24411, C2 =>
                           OUT2_26_port, A => n23277, ZN => n23260);
   U24260 : NOR4_X1 port map( A1 => n23272, A2 => n23273, A3 => n23274, A4 => 
                           n23275, ZN => n23262);
   U24261 : NAND4_X1 port map( A1 => n23242, A2 => n23243, A3 => n23244, A4 => 
                           n23245, ZN => n4959);
   U24262 : AOI221_X1 port map( B1 => n24440, B2 => n24383, C1 => n24434, C2 =>
                           n19890, A => n23258, ZN => n23243);
   U24263 : AOI221_X1 port map( B1 => n24416, B2 => n19496, C1 => n24411, C2 =>
                           OUT2_27_port, A => n23259, ZN => n23242);
   U24264 : NOR4_X1 port map( A1 => n23254, A2 => n23255, A3 => n23256, A4 => 
                           n23257, ZN => n23244);
   U24265 : NAND4_X1 port map( A1 => n23224, A2 => n23225, A3 => n23226, A4 => 
                           n23227, ZN => n4960);
   U24266 : AOI221_X1 port map( B1 => n24440, B2 => n24384, C1 => n24434, C2 =>
                           n19889, A => n23240, ZN => n23225);
   U24267 : AOI221_X1 port map( B1 => n24416, B2 => n19495, C1 => n24411, C2 =>
                           OUT2_28_port, A => n23241, ZN => n23224);
   U24268 : NOR4_X1 port map( A1 => n23236, A2 => n23237, A3 => n23238, A4 => 
                           n23239, ZN => n23226);
   U24269 : NAND4_X1 port map( A1 => n23206, A2 => n23207, A3 => n23208, A4 => 
                           n23209, ZN => n4961);
   U24270 : AOI221_X1 port map( B1 => n24440, B2 => n24385, C1 => n24434, C2 =>
                           n19888, A => n23222, ZN => n23207);
   U24271 : AOI221_X1 port map( B1 => n24416, B2 => n19494, C1 => n24411, C2 =>
                           OUT2_29_port, A => n23223, ZN => n23206);
   U24272 : NOR4_X1 port map( A1 => n23218, A2 => n23219, A3 => n23220, A4 => 
                           n23221, ZN => n23208);
   U24273 : NAND4_X1 port map( A1 => n23188, A2 => n23189, A3 => n23190, A4 => 
                           n23191, ZN => n4962);
   U24274 : AOI221_X1 port map( B1 => n24440, B2 => n24386, C1 => n24434, C2 =>
                           n19887, A => n23204, ZN => n23189);
   U24275 : AOI221_X1 port map( B1 => n24416, B2 => n19493, C1 => n24410, C2 =>
                           OUT2_30_port, A => n23205, ZN => n23188);
   U24276 : NOR4_X1 port map( A1 => n23200, A2 => n23201, A3 => n23202, A4 => 
                           n23203, ZN => n23190);
   U24277 : NAND4_X1 port map( A1 => n23170, A2 => n23171, A3 => n23172, A4 => 
                           n23173, ZN => n4963);
   U24278 : AOI221_X1 port map( B1 => n24440, B2 => n24387, C1 => n24434, C2 =>
                           n19886, A => n23186, ZN => n23171);
   U24279 : AOI221_X1 port map( B1 => n24416, B2 => n19492, C1 => n24410, C2 =>
                           OUT2_31_port, A => n23187, ZN => n23170);
   U24280 : NOR4_X1 port map( A1 => n23182, A2 => n23183, A3 => n23184, A4 => 
                           n23185, ZN => n23172);
   U24281 : NAND4_X1 port map( A1 => n23152, A2 => n23153, A3 => n23154, A4 => 
                           n23155, ZN => n4964);
   U24282 : AOI221_X1 port map( B1 => n24440, B2 => n24388, C1 => n24434, C2 =>
                           n19885, A => n23168, ZN => n23153);
   U24283 : AOI221_X1 port map( B1 => n24416, B2 => n19491, C1 => n24410, C2 =>
                           OUT2_32_port, A => n23169, ZN => n23152);
   U24284 : NOR4_X1 port map( A1 => n23164, A2 => n23165, A3 => n23166, A4 => 
                           n23167, ZN => n23154);
   U24285 : NAND4_X1 port map( A1 => n23134, A2 => n23135, A3 => n23136, A4 => 
                           n23137, ZN => n4965);
   U24286 : AOI221_X1 port map( B1 => n24440, B2 => n24389, C1 => n24434, C2 =>
                           n19884, A => n23150, ZN => n23135);
   U24287 : AOI221_X1 port map( B1 => n24416, B2 => n19490, C1 => n24410, C2 =>
                           OUT2_33_port, A => n23151, ZN => n23134);
   U24288 : NOR4_X1 port map( A1 => n23146, A2 => n23147, A3 => n23148, A4 => 
                           n23149, ZN => n23136);
   U24289 : NAND4_X1 port map( A1 => n23116, A2 => n23117, A3 => n23118, A4 => 
                           n23119, ZN => n4966);
   U24290 : AOI221_X1 port map( B1 => n24440, B2 => n24390, C1 => n24434, C2 =>
                           n19883, A => n23132, ZN => n23117);
   U24291 : AOI221_X1 port map( B1 => n24416, B2 => n19489, C1 => n24410, C2 =>
                           OUT2_34_port, A => n23133, ZN => n23116);
   U24292 : NOR4_X1 port map( A1 => n23128, A2 => n23129, A3 => n23130, A4 => 
                           n23131, ZN => n23118);
   U24293 : NAND4_X1 port map( A1 => n23098, A2 => n23099, A3 => n23100, A4 => 
                           n23101, ZN => n4967);
   U24294 : AOI221_X1 port map( B1 => n24440, B2 => n24391, C1 => n24434, C2 =>
                           n19882, A => n23114, ZN => n23099);
   U24295 : AOI221_X1 port map( B1 => n24416, B2 => n19488, C1 => n24410, C2 =>
                           OUT2_35_port, A => n23115, ZN => n23098);
   U24296 : NOR4_X1 port map( A1 => n23110, A2 => n23111, A3 => n23112, A4 => 
                           n23113, ZN => n23100);
   U24297 : NAND4_X1 port map( A1 => n23080, A2 => n23081, A3 => n23082, A4 => 
                           n23083, ZN => n4968);
   U24298 : AOI221_X1 port map( B1 => n24441, B2 => n24392, C1 => n24435, C2 =>
                           n19881, A => n23096, ZN => n23081);
   U24299 : AOI221_X1 port map( B1 => n24417, B2 => n19487, C1 => n24410, C2 =>
                           OUT2_36_port, A => n23097, ZN => n23080);
   U24300 : NOR4_X1 port map( A1 => n23092, A2 => n23093, A3 => n23094, A4 => 
                           n23095, ZN => n23082);
   U24301 : NAND4_X1 port map( A1 => n23062, A2 => n23063, A3 => n23064, A4 => 
                           n23065, ZN => n4969);
   U24302 : AOI221_X1 port map( B1 => n24441, B2 => n24393, C1 => n24435, C2 =>
                           n19880, A => n23078, ZN => n23063);
   U24303 : AOI221_X1 port map( B1 => n24417, B2 => n19486, C1 => n24410, C2 =>
                           OUT2_37_port, A => n23079, ZN => n23062);
   U24304 : NOR4_X1 port map( A1 => n23074, A2 => n23075, A3 => n23076, A4 => 
                           n23077, ZN => n23064);
   U24305 : NAND4_X1 port map( A1 => n23044, A2 => n23045, A3 => n23046, A4 => 
                           n23047, ZN => n4970);
   U24306 : AOI221_X1 port map( B1 => n24441, B2 => n24394, C1 => n24435, C2 =>
                           n19879, A => n23060, ZN => n23045);
   U24307 : AOI221_X1 port map( B1 => n24417, B2 => n19485, C1 => n24410, C2 =>
                           OUT2_38_port, A => n23061, ZN => n23044);
   U24308 : NOR4_X1 port map( A1 => n23056, A2 => n23057, A3 => n23058, A4 => 
                           n23059, ZN => n23046);
   U24309 : NAND4_X1 port map( A1 => n23026, A2 => n23027, A3 => n23028, A4 => 
                           n23029, ZN => n4971);
   U24310 : AOI221_X1 port map( B1 => n24441, B2 => n24395, C1 => n24435, C2 =>
                           n19878, A => n23042, ZN => n23027);
   U24311 : AOI221_X1 port map( B1 => n24417, B2 => n19484, C1 => n24410, C2 =>
                           OUT2_39_port, A => n23043, ZN => n23026);
   U24312 : NOR4_X1 port map( A1 => n23038, A2 => n23039, A3 => n23040, A4 => 
                           n23041, ZN => n23028);
   U24313 : OAI22_X1 port map( A1 => n24888, A2 => n25347, B1 => n24886, B2 => 
                           n20906, ZN => n5316);
   U24314 : OAI22_X1 port map( A1 => n24888, A2 => n25350, B1 => n24886, B2 => 
                           n20905, ZN => n5317);
   U24315 : OAI22_X1 port map( A1 => n24888, A2 => n25353, B1 => n24886, B2 => 
                           n20904, ZN => n5318);
   U24316 : OAI22_X1 port map( A1 => n24888, A2 => n25356, B1 => n24886, B2 => 
                           n20903, ZN => n5319);
   U24317 : OAI22_X1 port map( A1 => n24888, A2 => n25359, B1 => n24886, B2 => 
                           n20902, ZN => n5320);
   U24318 : OAI22_X1 port map( A1 => n24889, A2 => n25362, B1 => n24886, B2 => 
                           n20901, ZN => n5321);
   U24319 : OAI22_X1 port map( A1 => n24889, A2 => n25365, B1 => n24886, B2 => 
                           n20900, ZN => n5322);
   U24320 : OAI22_X1 port map( A1 => n24889, A2 => n25368, B1 => n24886, B2 => 
                           n20899, ZN => n5323);
   U24321 : OAI22_X1 port map( A1 => n24889, A2 => n25371, B1 => n24886, B2 => 
                           n20898, ZN => n5324);
   U24322 : OAI22_X1 port map( A1 => n24889, A2 => n25374, B1 => n24886, B2 => 
                           n20897, ZN => n5325);
   U24323 : OAI22_X1 port map( A1 => n24890, A2 => n25377, B1 => n24886, B2 => 
                           n20896, ZN => n5326);
   U24324 : OAI22_X1 port map( A1 => n24890, A2 => n25380, B1 => n24886, B2 => 
                           n20895, ZN => n5327);
   U24325 : OAI22_X1 port map( A1 => n24890, A2 => n25383, B1 => n24887, B2 => 
                           n20894, ZN => n5328);
   U24326 : OAI22_X1 port map( A1 => n24890, A2 => n25386, B1 => n24887, B2 => 
                           n20893, ZN => n5329);
   U24327 : OAI22_X1 port map( A1 => n24890, A2 => n25389, B1 => n24887, B2 => 
                           n20892, ZN => n5330);
   U24328 : OAI22_X1 port map( A1 => n24891, A2 => n25392, B1 => n24887, B2 => 
                           n20891, ZN => n5331);
   U24329 : OAI22_X1 port map( A1 => n24891, A2 => n25395, B1 => n24887, B2 => 
                           n20890, ZN => n5332);
   U24330 : OAI22_X1 port map( A1 => n24891, A2 => n25398, B1 => n24887, B2 => 
                           n20889, ZN => n5333);
   U24331 : OAI22_X1 port map( A1 => n24891, A2 => n25401, B1 => n24887, B2 => 
                           n20888, ZN => n5334);
   U24332 : OAI22_X1 port map( A1 => n24891, A2 => n25404, B1 => n24887, B2 => 
                           n20887, ZN => n5335);
   U24333 : OAI22_X1 port map( A1 => n24892, A2 => n25407, B1 => n24887, B2 => 
                           n20886, ZN => n5336);
   U24334 : OAI22_X1 port map( A1 => n24892, A2 => n25410, B1 => n24887, B2 => 
                           n20885, ZN => n5337);
   U24335 : OAI22_X1 port map( A1 => n24892, A2 => n25413, B1 => n24887, B2 => 
                           n20884, ZN => n5338);
   U24336 : OAI22_X1 port map( A1 => n24892, A2 => n25416, B1 => n24887, B2 => 
                           n20883, ZN => n5339);
   U24337 : OAI22_X1 port map( A1 => n24892, A2 => n25419, B1 => n24886, B2 => 
                           n20882, ZN => n5340);
   U24338 : OAI22_X1 port map( A1 => n24893, A2 => n25422, B1 => n24887, B2 => 
                           n20881, ZN => n5341);
   U24339 : OAI22_X1 port map( A1 => n24893, A2 => n25425, B1 => n24885, B2 => 
                           n20880, ZN => n5342);
   U24340 : OAI22_X1 port map( A1 => n24893, A2 => n25428, B1 => n24886, B2 => 
                           n20879, ZN => n5343);
   U24341 : OAI22_X1 port map( A1 => n24893, A2 => n25431, B1 => n24887, B2 => 
                           n20878, ZN => n5344);
   U24342 : OAI22_X1 port map( A1 => n24893, A2 => n25434, B1 => n24885, B2 => 
                           n20877, ZN => n5345);
   U24343 : OAI22_X1 port map( A1 => n24894, A2 => n25437, B1 => n24886, B2 => 
                           n20876, ZN => n5346);
   U24344 : OAI22_X1 port map( A1 => n24894, A2 => n25440, B1 => n24887, B2 => 
                           n20875, ZN => n5347);
   U24345 : OAI22_X1 port map( A1 => n24894, A2 => n25443, B1 => n24885, B2 => 
                           n20874, ZN => n5348);
   U24346 : OAI22_X1 port map( A1 => n24894, A2 => n25446, B1 => n24886, B2 => 
                           n20873, ZN => n5349);
   U24347 : OAI22_X1 port map( A1 => n24894, A2 => n25449, B1 => n24887, B2 => 
                           n20872, ZN => n5350);
   U24348 : OAI22_X1 port map( A1 => n24895, A2 => n25452, B1 => n24885, B2 => 
                           n20871, ZN => n5351);
   U24349 : OAI22_X1 port map( A1 => n24895, A2 => n25455, B1 => n21292, B2 => 
                           n20870, ZN => n5352);
   U24350 : OAI22_X1 port map( A1 => n24895, A2 => n25458, B1 => n24885, B2 => 
                           n20869, ZN => n5353);
   U24351 : OAI22_X1 port map( A1 => n24895, A2 => n25461, B1 => n21292, B2 => 
                           n20868, ZN => n5354);
   U24352 : OAI22_X1 port map( A1 => n24895, A2 => n25464, B1 => n24885, B2 => 
                           n20867, ZN => n5355);
   U24353 : OAI22_X1 port map( A1 => n24896, A2 => n25467, B1 => n21292, B2 => 
                           n20866, ZN => n5356);
   U24354 : OAI22_X1 port map( A1 => n24896, A2 => n25470, B1 => n24885, B2 => 
                           n20865, ZN => n5357);
   U24355 : OAI22_X1 port map( A1 => n24896, A2 => n25473, B1 => n24886, B2 => 
                           n20864, ZN => n5358);
   U24356 : OAI22_X1 port map( A1 => n24896, A2 => n25476, B1 => n24887, B2 => 
                           n20863, ZN => n5359);
   U24357 : OAI22_X1 port map( A1 => n24896, A2 => n25479, B1 => n24885, B2 => 
                           n20862, ZN => n5360);
   U24358 : OAI22_X1 port map( A1 => n24897, A2 => n25482, B1 => n24885, B2 => 
                           n20861, ZN => n5361);
   U24359 : OAI22_X1 port map( A1 => n24897, A2 => n25485, B1 => n24886, B2 => 
                           n20860, ZN => n5362);
   U24360 : OAI22_X1 port map( A1 => n24897, A2 => n25488, B1 => n24887, B2 => 
                           n20859, ZN => n5363);
   U24361 : OAI22_X1 port map( A1 => n24897, A2 => n25491, B1 => n24885, B2 => 
                           n20858, ZN => n5364);
   U24362 : OAI22_X1 port map( A1 => n24897, A2 => n25494, B1 => n24885, B2 => 
                           n20857, ZN => n5365);
   U24363 : OAI22_X1 port map( A1 => n24898, A2 => n25497, B1 => n21292, B2 => 
                           n20856, ZN => n5366);
   U24364 : OAI22_X1 port map( A1 => n24898, A2 => n25500, B1 => n24885, B2 => 
                           n20855, ZN => n5367);
   U24365 : OAI22_X1 port map( A1 => n24898, A2 => n25503, B1 => n21292, B2 => 
                           n20854, ZN => n5368);
   U24366 : OAI22_X1 port map( A1 => n24898, A2 => n25506, B1 => n24885, B2 => 
                           n20853, ZN => n5369);
   U24367 : OAI22_X1 port map( A1 => n24898, A2 => n25509, B1 => n21292, B2 => 
                           n20852, ZN => n5370);
   U24368 : OAI22_X1 port map( A1 => n24899, A2 => n25512, B1 => n24885, B2 => 
                           n20851, ZN => n5371);
   U24369 : OAI22_X1 port map( A1 => n24899, A2 => n25515, B1 => n21292, B2 => 
                           n20850, ZN => n5372);
   U24370 : OAI22_X1 port map( A1 => n24899, A2 => n25518, B1 => n24885, B2 => 
                           n20849, ZN => n5373);
   U24371 : OAI22_X1 port map( A1 => n24899, A2 => n25521, B1 => n21292, B2 => 
                           n20848, ZN => n5374);
   U24372 : OAI22_X1 port map( A1 => n24899, A2 => n25524, B1 => n24885, B2 => 
                           n20847, ZN => n5375);
   U24373 : NOR3_X1 port map( A1 => n19199, A2 => ADD_RD2(0), A3 => n19200, ZN 
                           => n23748);
   U24374 : NOR3_X1 port map( A1 => n19199, A2 => ADD_RD2(3), A3 => n19203, ZN 
                           => n23745);
   U24375 : NOR3_X1 port map( A1 => n19203, A2 => ADD_RD2(4), A3 => n19200, ZN 
                           => n23742);
   U24376 : NOR3_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(4), A3 => n19196,
                           ZN => n22553);
   U24377 : NOR2_X1 port map( A1 => n19197, A2 => ADD_RD1(2), ZN => n22543);
   U24378 : NOR3_X1 port map( A1 => n19196, A2 => ADD_RD1(4), A3 => n19198, ZN 
                           => n22554);
   U24379 : NOR3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), A3 => 
                           ADD_RD1(0), ZN => n22558);
   U24380 : NOR3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), A3 => n19198,
                           ZN => n22557);
   U24381 : NOR3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(3), A3 => n19199,
                           ZN => n23738);
   U24382 : NOR3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(4), A3 => n19200,
                           ZN => n23741);
   U24383 : AND2_X1 port map( A1 => ADD_RD1(2), A2 => n19197, ZN => n22538);
   U24384 : NOR2_X1 port map( A1 => n24408, A2 => WR, ZN => n23761);
   U24385 : NOR2_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), ZN => n23757)
                           ;
   U24386 : NOR2_X1 port map( A1 => n19201, A2 => ADD_RD2(1), ZN => n23759);
   U24387 : NOR2_X1 port map( A1 => n19202, A2 => ADD_RD2(2), ZN => n23758);
   U24388 : AND2_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), ZN => n22540)
                           ;
   U24389 : NAND2_X1 port map( A1 => n24803, A2 => WR, ZN => n21297);
   U24390 : INV_X1 port map( A => ADD_RD2(3), ZN => n19200);
   U24391 : INV_X1 port map( A => ADD_RD2(4), ZN => n19199);
   U24392 : NAND2_X1 port map( A1 => RD2, A2 => ENABLE, ZN => n22608);
   U24393 : AND2_X1 port map( A1 => n23760, A2 => ADD_RD2(0), ZN => n23756);
   U24394 : AND3_X1 port map( A1 => n19198, A2 => n19196, A3 => ADD_RD1(4), ZN 
                           => n22545);
   U24395 : AND3_X1 port map( A1 => ADD_RD1(3), A2 => n19198, A3 => ADD_RD1(4),
                           ZN => n22537);
   U24396 : AND3_X1 port map( A1 => ADD_RD1(0), A2 => n19196, A3 => ADD_RD1(4),
                           ZN => n22546);
   U24397 : AND3_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(3), A3 => 
                           ADD_RD1(4), ZN => n22539);
   U24398 : INV_X1 port map( A => ADD_RD2(0), ZN => n19203);
   U24399 : NAND2_X1 port map( A1 => DATAIN(0), A2 => n25562, ZN => n21252);
   U24400 : NAND2_X1 port map( A1 => DATAIN(1), A2 => n25562, ZN => n21251);
   U24401 : NAND2_X1 port map( A1 => DATAIN(2), A2 => n25562, ZN => n21250);
   U24402 : NAND2_X1 port map( A1 => DATAIN(4), A2 => n25562, ZN => n21248);
   U24403 : NAND2_X1 port map( A1 => DATAIN(3), A2 => n25561, ZN => n21249);
   U24404 : NAND2_X1 port map( A1 => DATAIN(5), A2 => n25561, ZN => n21247);
   U24405 : NAND2_X1 port map( A1 => DATAIN(6), A2 => n25561, ZN => n21246);
   U24406 : NAND2_X1 port map( A1 => DATAIN(7), A2 => n25561, ZN => n21245);
   U24407 : NAND2_X1 port map( A1 => DATAIN(8), A2 => n25561, ZN => n21244);
   U24408 : NAND2_X1 port map( A1 => DATAIN(9), A2 => n25561, ZN => n21243);
   U24409 : NAND2_X1 port map( A1 => DATAIN(10), A2 => n25561, ZN => n21242);
   U24410 : NAND2_X1 port map( A1 => DATAIN(11), A2 => n25561, ZN => n21241);
   U24411 : NAND2_X1 port map( A1 => DATAIN(12), A2 => n25561, ZN => n21240);
   U24412 : NAND2_X1 port map( A1 => DATAIN(13), A2 => n25561, ZN => n21239);
   U24413 : NAND2_X1 port map( A1 => DATAIN(14), A2 => n25561, ZN => n21238);
   U24414 : NAND2_X1 port map( A1 => DATAIN(15), A2 => n25560, ZN => n21237);
   U24415 : NAND2_X1 port map( A1 => DATAIN(16), A2 => n25561, ZN => n21236);
   U24416 : NAND2_X1 port map( A1 => DATAIN(17), A2 => n25560, ZN => n21235);
   U24417 : NAND2_X1 port map( A1 => DATAIN(18), A2 => n25560, ZN => n21234);
   U24418 : NAND2_X1 port map( A1 => DATAIN(19), A2 => n25560, ZN => n21233);
   U24419 : NAND2_X1 port map( A1 => DATAIN(20), A2 => n25560, ZN => n21232);
   U24420 : NAND2_X1 port map( A1 => DATAIN(21), A2 => n25560, ZN => n21231);
   U24421 : NAND2_X1 port map( A1 => DATAIN(22), A2 => n25560, ZN => n21230);
   U24422 : NAND2_X1 port map( A1 => DATAIN(23), A2 => n25559, ZN => n21229);
   U24423 : NAND2_X1 port map( A1 => DATAIN(24), A2 => n25560, ZN => n21228);
   U24424 : NAND2_X1 port map( A1 => DATAIN(25), A2 => n25560, ZN => n21227);
   U24425 : NAND2_X1 port map( A1 => DATAIN(26), A2 => n25560, ZN => n21226);
   U24426 : NAND2_X1 port map( A1 => DATAIN(27), A2 => n25560, ZN => n21225);
   U24427 : NAND2_X1 port map( A1 => DATAIN(28), A2 => n25560, ZN => n21224);
   U24428 : NAND2_X1 port map( A1 => DATAIN(29), A2 => n25559, ZN => n21223);
   U24429 : NAND2_X1 port map( A1 => DATAIN(30), A2 => n25559, ZN => n21222);
   U24430 : NAND2_X1 port map( A1 => DATAIN(31), A2 => n25559, ZN => n21221);
   U24431 : NAND2_X1 port map( A1 => DATAIN(32), A2 => n25559, ZN => n21220);
   U24432 : NAND2_X1 port map( A1 => DATAIN(33), A2 => n25559, ZN => n21219);
   U24433 : NAND2_X1 port map( A1 => DATAIN(34), A2 => n25559, ZN => n21218);
   U24434 : NAND2_X1 port map( A1 => DATAIN(35), A2 => n25559, ZN => n21217);
   U24435 : NAND2_X1 port map( A1 => DATAIN(36), A2 => n25559, ZN => n21216);
   U24436 : NAND2_X1 port map( A1 => DATAIN(37), A2 => n25559, ZN => n21215);
   U24437 : NAND2_X1 port map( A1 => DATAIN(38), A2 => n25559, ZN => n21214);
   U24438 : NAND2_X1 port map( A1 => DATAIN(39), A2 => n25559, ZN => n21213);
   U24439 : NAND2_X1 port map( A1 => DATAIN(40), A2 => n25558, ZN => n21212);
   U24440 : NAND2_X1 port map( A1 => DATAIN(41), A2 => n25558, ZN => n21211);
   U24441 : NAND2_X1 port map( A1 => DATAIN(42), A2 => n25558, ZN => n21210);
   U24442 : NAND2_X1 port map( A1 => DATAIN(43), A2 => n25558, ZN => n21209);
   U24443 : NAND2_X1 port map( A1 => DATAIN(44), A2 => n25558, ZN => n21208);
   U24444 : NAND2_X1 port map( A1 => DATAIN(45), A2 => n25558, ZN => n21207);
   U24445 : NAND2_X1 port map( A1 => DATAIN(46), A2 => n25558, ZN => n21206);
   U24446 : NAND2_X1 port map( A1 => DATAIN(47), A2 => n25558, ZN => n21205);
   U24447 : NAND2_X1 port map( A1 => DATAIN(48), A2 => n25558, ZN => n21204);
   U24448 : NAND2_X1 port map( A1 => DATAIN(49), A2 => n25558, ZN => n21203);
   U24449 : NAND2_X1 port map( A1 => DATAIN(50), A2 => n25558, ZN => n21202);
   U24450 : NAND2_X1 port map( A1 => DATAIN(51), A2 => n25558, ZN => n21201);
   U24451 : NAND2_X1 port map( A1 => DATAIN(52), A2 => n25557, ZN => n21200);
   U24452 : NAND2_X1 port map( A1 => DATAIN(53), A2 => n25557, ZN => n21199);
   U24453 : NAND2_X1 port map( A1 => DATAIN(54), A2 => n25557, ZN => n21198);
   U24454 : NAND2_X1 port map( A1 => DATAIN(55), A2 => n25557, ZN => n21197);
   U24455 : NAND2_X1 port map( A1 => DATAIN(56), A2 => n25557, ZN => n21196);
   U24456 : NAND2_X1 port map( A1 => DATAIN(57), A2 => n25557, ZN => n21195);
   U24457 : NAND2_X1 port map( A1 => DATAIN(58), A2 => n25557, ZN => n21194);
   U24458 : NAND2_X1 port map( A1 => DATAIN(59), A2 => n25557, ZN => n21193);
   U24459 : NAND2_X1 port map( A1 => DATAIN(60), A2 => n25557, ZN => n21192);
   U24460 : NAND2_X1 port map( A1 => DATAIN(61), A2 => n25557, ZN => n21191);
   U24461 : NAND2_X1 port map( A1 => DATAIN(62), A2 => n25557, ZN => n21190);
   U24462 : NAND2_X1 port map( A1 => DATAIN(63), A2 => n25557, ZN => n21188);
   U24463 : AND2_X1 port map( A1 => RD1, A2 => ENABLE, ZN => n21298);
   U24464 : INV_X1 port map( A => ADD_RD1(0), ZN => n19198);
   U24465 : INV_X1 port map( A => ADD_RD1(3), ZN => n19196);
   U24466 : AND2_X1 port map( A1 => WR, A2 => ENABLE, ZN => n21269);
   U24467 : INV_X1 port map( A => ADD_WR(2), ZN => n19193);
   U24468 : INV_X1 port map( A => ADD_WR(0), ZN => n19195);
   U24469 : INV_X1 port map( A => ADD_WR(1), ZN => n19194);
   U24470 : INV_X1 port map( A => ADD_RD2(2), ZN => n19201);
   U24471 : INV_X1 port map( A => DATAIN(40), ZN => n19227);
   U24472 : INV_X1 port map( A => DATAIN(41), ZN => n19226);
   U24473 : INV_X1 port map( A => DATAIN(42), ZN => n19225);
   U24474 : INV_X1 port map( A => DATAIN(43), ZN => n19224);
   U24475 : INV_X1 port map( A => DATAIN(44), ZN => n19223);
   U24476 : INV_X1 port map( A => DATAIN(45), ZN => n19222);
   U24477 : INV_X1 port map( A => DATAIN(46), ZN => n19221);
   U24478 : INV_X1 port map( A => DATAIN(47), ZN => n19220);
   U24479 : INV_X1 port map( A => DATAIN(48), ZN => n19219);
   U24480 : INV_X1 port map( A => DATAIN(49), ZN => n19218);
   U24481 : INV_X1 port map( A => DATAIN(50), ZN => n19217);
   U24482 : INV_X1 port map( A => DATAIN(51), ZN => n19216);
   U24483 : INV_X1 port map( A => DATAIN(52), ZN => n19215);
   U24484 : INV_X1 port map( A => DATAIN(53), ZN => n19214);
   U24485 : INV_X1 port map( A => DATAIN(54), ZN => n19213);
   U24486 : INV_X1 port map( A => DATAIN(55), ZN => n19212);
   U24487 : INV_X1 port map( A => DATAIN(56), ZN => n19211);
   U24488 : INV_X1 port map( A => DATAIN(57), ZN => n19210);
   U24489 : INV_X1 port map( A => DATAIN(58), ZN => n19209);
   U24490 : INV_X1 port map( A => DATAIN(59), ZN => n19208);
   U24491 : INV_X1 port map( A => DATAIN(60), ZN => n19207);
   U24492 : INV_X1 port map( A => DATAIN(61), ZN => n19206);
   U24493 : INV_X1 port map( A => DATAIN(62), ZN => n19205);
   U24494 : INV_X1 port map( A => DATAIN(63), ZN => n19204);
   U24495 : INV_X1 port map( A => DATAIN(0), ZN => n19267);
   U24496 : INV_X1 port map( A => DATAIN(1), ZN => n19266);
   U24497 : INV_X1 port map( A => DATAIN(2), ZN => n19265);
   U24498 : INV_X1 port map( A => DATAIN(3), ZN => n19264);
   U24499 : INV_X1 port map( A => DATAIN(4), ZN => n19263);
   U24500 : INV_X1 port map( A => DATAIN(5), ZN => n19262);
   U24501 : INV_X1 port map( A => DATAIN(6), ZN => n19261);
   U24502 : INV_X1 port map( A => DATAIN(7), ZN => n19260);
   U24503 : INV_X1 port map( A => DATAIN(8), ZN => n19259);
   U24504 : INV_X1 port map( A => DATAIN(9), ZN => n19258);
   U24505 : INV_X1 port map( A => DATAIN(10), ZN => n19257);
   U24506 : INV_X1 port map( A => DATAIN(11), ZN => n19256);
   U24507 : INV_X1 port map( A => DATAIN(12), ZN => n19255);
   U24508 : INV_X1 port map( A => DATAIN(13), ZN => n19254);
   U24509 : INV_X1 port map( A => DATAIN(14), ZN => n19253);
   U24510 : INV_X1 port map( A => DATAIN(15), ZN => n19252);
   U24511 : INV_X1 port map( A => DATAIN(16), ZN => n19251);
   U24512 : INV_X1 port map( A => DATAIN(17), ZN => n19250);
   U24513 : INV_X1 port map( A => DATAIN(18), ZN => n19249);
   U24514 : INV_X1 port map( A => DATAIN(19), ZN => n19248);
   U24515 : INV_X1 port map( A => DATAIN(20), ZN => n19247);
   U24516 : INV_X1 port map( A => DATAIN(21), ZN => n19246);
   U24517 : INV_X1 port map( A => DATAIN(22), ZN => n19245);
   U24518 : INV_X1 port map( A => DATAIN(23), ZN => n19244);
   U24519 : INV_X1 port map( A => DATAIN(24), ZN => n19243);
   U24520 : INV_X1 port map( A => DATAIN(25), ZN => n19242);
   U24521 : INV_X1 port map( A => DATAIN(26), ZN => n19241);
   U24522 : INV_X1 port map( A => DATAIN(27), ZN => n19240);
   U24523 : INV_X1 port map( A => DATAIN(28), ZN => n19239);
   U24524 : INV_X1 port map( A => DATAIN(29), ZN => n19238);
   U24525 : INV_X1 port map( A => DATAIN(30), ZN => n19237);
   U24526 : INV_X1 port map( A => DATAIN(31), ZN => n19236);
   U24527 : INV_X1 port map( A => DATAIN(32), ZN => n19235);
   U24528 : INV_X1 port map( A => DATAIN(33), ZN => n19234);
   U24529 : INV_X1 port map( A => DATAIN(34), ZN => n19233);
   U24530 : INV_X1 port map( A => DATAIN(35), ZN => n19232);
   U24531 : INV_X1 port map( A => DATAIN(36), ZN => n19231);
   U24532 : INV_X1 port map( A => DATAIN(37), ZN => n19230);
   U24533 : INV_X1 port map( A => DATAIN(38), ZN => n19229);
   U24534 : INV_X1 port map( A => DATAIN(39), ZN => n19228);
   U24535 : INV_X1 port map( A => ADD_RD2(1), ZN => n19202);
   U24536 : INV_X1 port map( A => ADD_RD1(1), ZN => n19197);
   U24537 : INV_X1 port map( A => WR, ZN => n19190);
   U24538 : INV_X1 port map( A => ADD_WR(4), ZN => n19191);
   U24539 : INV_X1 port map( A => ADD_WR(3), ZN => n19192);
   U24540 : INV_X1 port map( A => RESET, ZN => n19189);
   U24541 : CLKBUF_X1 port map( A => n22611, Z => n24401);
   U24542 : CLKBUF_X1 port map( A => n22610, Z => n24407);
   U24543 : CLKBUF_X1 port map( A => n22608, Z => n24413);
   U24544 : CLKBUF_X1 port map( A => n22607, Z => n24419);
   U24545 : CLKBUF_X1 port map( A => n22606, Z => n24425);
   U24546 : CLKBUF_X1 port map( A => n22605, Z => n24431);
   U24547 : CLKBUF_X1 port map( A => n22603, Z => n24437);
   U24548 : CLKBUF_X1 port map( A => n22602, Z => n24443);
   U24549 : CLKBUF_X1 port map( A => n22601, Z => n24449);
   U24550 : CLKBUF_X1 port map( A => n22600, Z => n24455);
   U24551 : CLKBUF_X1 port map( A => n22599, Z => n24461);
   U24552 : CLKBUF_X1 port map( A => n22598, Z => n24467);
   U24553 : CLKBUF_X1 port map( A => n22597, Z => n24473);
   U24554 : CLKBUF_X1 port map( A => n22596, Z => n24479);
   U24555 : CLKBUF_X1 port map( A => n22595, Z => n24485);
   U24556 : CLKBUF_X1 port map( A => n22594, Z => n24491);
   U24557 : CLKBUF_X1 port map( A => n22593, Z => n24497);
   U24558 : CLKBUF_X1 port map( A => n22588, Z => n24503);
   U24559 : CLKBUF_X1 port map( A => n22587, Z => n24509);
   U24560 : CLKBUF_X1 port map( A => n22586, Z => n24515);
   U24561 : CLKBUF_X1 port map( A => n22584, Z => n24521);
   U24562 : CLKBUF_X1 port map( A => n22583, Z => n24527);
   U24563 : CLKBUF_X1 port map( A => n22582, Z => n24533);
   U24564 : CLKBUF_X1 port map( A => n22581, Z => n24539);
   U24565 : CLKBUF_X1 port map( A => n22579, Z => n24545);
   U24566 : CLKBUF_X1 port map( A => n22578, Z => n24551);
   U24567 : CLKBUF_X1 port map( A => n22577, Z => n24557);
   U24568 : CLKBUF_X1 port map( A => n22576, Z => n24563);
   U24569 : CLKBUF_X1 port map( A => n22574, Z => n24569);
   U24570 : CLKBUF_X1 port map( A => n22573, Z => n24575);
   U24571 : CLKBUF_X1 port map( A => n22572, Z => n24581);
   U24572 : CLKBUF_X1 port map( A => n22571, Z => n24587);
   U24573 : CLKBUF_X1 port map( A => n22569, Z => n24593);
   U24574 : CLKBUF_X1 port map( A => n22568, Z => n24599);
   U24575 : CLKBUF_X1 port map( A => n21350, Z => n24605);
   U24576 : CLKBUF_X1 port map( A => n21349, Z => n24611);
   U24577 : CLKBUF_X1 port map( A => n21347, Z => n24617);
   U24578 : CLKBUF_X1 port map( A => n21346, Z => n24623);
   U24579 : CLKBUF_X1 port map( A => n21345, Z => n24629);
   U24580 : CLKBUF_X1 port map( A => n21344, Z => n24635);
   U24581 : CLKBUF_X1 port map( A => n21342, Z => n24641);
   U24582 : CLKBUF_X1 port map( A => n21341, Z => n24647);
   U24583 : CLKBUF_X1 port map( A => n21340, Z => n24653);
   U24584 : CLKBUF_X1 port map( A => n21339, Z => n24659);
   U24585 : CLKBUF_X1 port map( A => n21337, Z => n24665);
   U24586 : CLKBUF_X1 port map( A => n21336, Z => n24671);
   U24587 : CLKBUF_X1 port map( A => n21335, Z => n24677);
   U24588 : CLKBUF_X1 port map( A => n21334, Z => n24683);
   U24589 : CLKBUF_X1 port map( A => n21332, Z => n24689);
   U24590 : CLKBUF_X1 port map( A => n21331, Z => n24695);
   U24591 : CLKBUF_X1 port map( A => n21326, Z => n24701);
   U24592 : CLKBUF_X1 port map( A => n21325, Z => n24707);
   U24593 : CLKBUF_X1 port map( A => n21323, Z => n24713);
   U24594 : CLKBUF_X1 port map( A => n21322, Z => n24719);
   U24595 : CLKBUF_X1 port map( A => n21321, Z => n24725);
   U24596 : CLKBUF_X1 port map( A => n21320, Z => n24731);
   U24597 : CLKBUF_X1 port map( A => n21318, Z => n24737);
   U24598 : CLKBUF_X1 port map( A => n21317, Z => n24743);
   U24599 : CLKBUF_X1 port map( A => n21316, Z => n24749);
   U24600 : CLKBUF_X1 port map( A => n21315, Z => n24755);
   U24601 : CLKBUF_X1 port map( A => n21313, Z => n24761);
   U24602 : CLKBUF_X1 port map( A => n21312, Z => n24767);
   U24603 : CLKBUF_X1 port map( A => n21311, Z => n24773);
   U24604 : CLKBUF_X1 port map( A => n21310, Z => n24779);
   U24605 : CLKBUF_X1 port map( A => n21308, Z => n24785);
   U24606 : CLKBUF_X1 port map( A => n21307, Z => n24791);
   U24607 : CLKBUF_X1 port map( A => n21302, Z => n24797);
   U24608 : CLKBUF_X1 port map( A => n21298, Z => n24803);
   U24609 : CLKBUF_X1 port map( A => n21297, Z => n24809);
   U24610 : CLKBUF_X1 port map( A => n19189, Z => n25554);
   U24611 : CLKBUF_X1 port map( A => n19189, Z => n25555);
   U24612 : CLKBUF_X1 port map( A => n19189, Z => n25556);

end SYN_beh;
