package constants is

  constant OP_CODE_SIZE : integer := 6;
  constant FUNC_SIZE : integer := 11;
  constant CW_SIZE : integer := 13;

end package constants;
