package constants is

  constant numBit : integer := 32;    -- Number of bits of the input operands
  constant radixN : integer := 3;     -- Number of the radix of the Booth's multiplier

end package constants;
