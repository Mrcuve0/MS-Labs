
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_registerFile_TLE is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_registerFile_TLE;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_registerFile_TLE.all;

entity 
   controlUnit_RF_N8_M8_F4_windowBlocks3_NData32_NAddr_Windowed5_DW01_incdec_0 
   is

   port( A : in std_logic_vector (31 downto 0);  INC_DEC : in std_logic;  SUM :
         out std_logic_vector (31 downto 0));

end controlUnit_RF_N8_M8_F4_windowBlocks3_NData32_NAddr_Windowed5_DW01_incdec_0
   ;

architecture SYN_rpl of 
   controlUnit_RF_N8_M8_F4_windowBlocks3_NData32_NAddr_Windowed5_DW01_incdec_0 
   is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port, n7, n8, n9, 
      n_1000, n_1001 : std_logic;

begin
   
   U1_31 : FA_X1 port map( A => A(31), B => INC_DEC, CI => carry_31_port, CO =>
                           n_1000, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => INC_DEC, CI => carry_30_port, CO =>
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => INC_DEC, CI => carry_29_port, CO =>
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => n8, CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => INC_DEC, CI => carry_27_port, CO =>
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => n8, CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => INC_DEC, CI => carry_25_port, CO =>
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => n8, CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => INC_DEC, CI => carry_23_port, CO =>
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => INC_DEC, CI => carry_22_port, CO =>
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => INC_DEC, CI => carry_21_port, CO =>
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => n8, CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => n8, CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => n8, CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => n8, CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => n8, CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => n8, CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => n8, CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => n8, CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => n8, CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => n7, CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => n7, CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => n7, CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => n7, CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => n7, CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => n7, CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => n7, CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => n7, CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => n7, CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => n7, CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => n7, CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => n7, CI => n9, CO => carry_1_port, S 
                           => n_1001);
   U1 : INV_X1 port map( A => n9, ZN => n7);
   U2 : INV_X1 port map( A => n9, ZN => n8);
   U3 : INV_X1 port map( A => INC_DEC, ZN => n9);
   U4 : INV_X1 port map( A => A(0), ZN => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_registerFile_TLE.all;

entity physical_RF_NData32_NRegs72_NAddr7 is

   port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (6 downto 0);  DATAIN : in 
         std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31
         downto 0));

end physical_RF_NData32_NRegs72_NAddr7;

architecture SYN_beh of physical_RF_NData32_NRegs72_NAddr7 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X4
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component TINV_X1
      port( I, EN : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
      n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, 
      n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, 
      n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, 
      n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, 
      n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, 
      n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, 
      n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, 
      n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, 
      n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, 
      n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, 
      n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, 
      n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, 
      n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, 
      n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, 
      n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, 
      n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, 
      n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, 
      n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, 
      n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, 
      n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, 
      n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, 
      n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, 
      n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, 
      n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, 
      n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, 
      n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, 
      n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, 
      n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, 
      n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, 
      n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, 
      n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, 
      n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, 
      n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, 
      n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, 
      n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, 
      n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, 
      n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, 
      n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, 
      n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, 
      n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, 
      n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, 
      n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, 
      n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, 
      n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, 
      n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, 
      n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, 
      n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, 
      n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, 
      n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, 
      n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, 
      n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, 
      n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, 
      n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, 
      n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, 
      n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, 
      n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, 
      n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, 
      n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, 
      n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, 
      n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, 
      n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, 
      n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, 
      n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, 
      n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, 
      n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, 
      n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, 
      n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, 
      n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, 
      n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, 
      n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, 
      n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, 
      n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, 
      n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, 
      n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, 
      n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, 
      n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, 
      n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, 
      n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, 
      n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, 
      n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, 
      n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, 
      n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, 
      n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, 
      n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, 
      n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, 
      n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, 
      n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, 
      n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, 
      n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, 
      n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, 
      n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, 
      n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, 
      n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, 
      n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, 
      n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, 
      n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, 
      n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, 
      n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, 
      n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, 
      n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, 
      n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, 
      n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, 
      n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, 
      n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, 
      n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, 
      n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, 
      n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, 
      n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, 
      n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, 
      n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, 
      n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, 
      n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, 
      n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, 
      n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, 
      n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, 
      n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, 
      n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, 
      n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, 
      n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, 
      n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, 
      n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, 
      n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, 
      n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, 
      n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, 
      n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, 
      n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, 
      n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, 
      n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, 
      n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, 
      n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, 
      n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, 
      n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, 
      n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, 
      n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, 
      n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, 
      n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, 
      n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, 
      n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, 
      n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, 
      n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, 
      n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, 
      n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, 
      n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, 
      n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, 
      n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, 
      n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, 
      n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, 
      n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, 
      n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, 
      n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, 
      n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, 
      n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, 
      n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, 
      n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, 
      n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, 
      n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, 
      n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, 
      n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, 
      n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, 
      n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, 
      n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, 
      n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, 
      n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, 
      n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, 
      n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, 
      n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, 
      n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, 
      n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, 
      n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, 
      n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, 
      n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, 
      n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, 
      n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, 
      n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, 
      n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, 
      n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, 
      n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, 
      n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, 
      n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, 
      n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, 
      n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, 
      n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, 
      n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, 
      n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, 
      n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, 
      n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, 
      n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, 
      n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, 
      n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, 
      n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, 
      n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, 
      n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, 
      n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, 
      n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, 
      n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, 
      n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, 
      n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, 
      n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, 
      n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, 
      n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, 
      n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, 
      n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, 
      n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, 
      n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, 
      n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, 
      n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, 
      n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, 
      n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, 
      n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, 
      n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, 
      n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, 
      n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, 
      n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, 
      n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, 
      n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, 
      n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, 
      n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, 
      n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, 
      n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, 
      n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, 
      n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, 
      n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, 
      n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, 
      n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, 
      n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, 
      n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, 
      n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, 
      n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, 
      n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, 
      n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, 
      n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, 
      n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, 
      n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, 
      n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, 
      n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, 
      n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, 
      n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, 
      n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, 
      n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, 
      n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, 
      n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, 
      n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, 
      n9976, n9977, n97, n98, n99, n578, n580, n582, n584, n586, n588, n590, 
      n592, n594, n596, n598, n600, n602, n604, n606, n608, n610, n612, n614, 
      n616, n622, n625, n628, n631, n634, n637, n640, n643, n646, n649, n652, 
      n653, n655, n656, n658, n659, n661, n662, n664, n665, n666, n667, n668, 
      n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, 
      n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, 
      n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, 
      n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n716, n717, 
      n719, n720, n722, n723, n725, n726, n728, n729, n731, n732, n734, n735, 
      n737, n738, n740, n741, n743, n744, n746, n747, n749, n750, n752, n753, 
      n755, n756, n758, n759, n761, n762, n764, n765, n767, n768, n770, n771, 
      n773, n774, n776, n777, n779, n780, n782, n783, n785, n786, n788, n789, 
      n791, n792, n794, n795, n797, n798, n800, n801, n803, n804, n806, n807, 
      n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, 
      n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, 
      n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, 
      n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, 
      n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, 
      n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, 
      n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, 
      n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, 
      n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, 
      n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, 
      n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, 
      n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, 
      n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, 
      n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, 
      n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, 
      n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1449, 
      n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, 
      n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, 
      n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, 
      n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, 
      n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, 
      n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, 
      n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, 
      n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, 
      n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, 
      n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, 
      n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, 
      n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, 
      n1570, n1571, n1572, n1573, n1574, n1575, n1576, n5383, n5385, n5387, 
      n5393, n5395, n5397, n5403, n5405, n5407, n5413, n5415, n5417, n5423, 
      n5425, n5427, n5433, n5435, n5437, n5443, n5445, n5447, n5452, n5453, 
      n5455, n5457, n5462, n5463, n5465, n5467, n5472, n5473, n5475, n5477, 
      n5482, n5483, n5485, n5487, n5492, n5493, n5495, n5497, n5502, n5503, 
      n5505, n5507, n5512, n5513, n5515, n5517, n5522, n5523, n5525, n5527, 
      n5532, n5533, n5535, n5537, n5542, n5543, n5545, n5547, n5552, n5553, 
      n5555, n5557, n5562, n5563, n5565, n5567, n5572, n5573, n5575, n5577, 
      n5582, n5583, n5585, n5587, n5592, n5593, n5595, n5597, n5602, n5603, 
      n5605, n5607, n5612, n5613, n5615, n5617, n5622, n5623, n5625, n5627, 
      n5632, n5633, n5635, n5637, n5642, n5643, n5645, n5647, n5652, n5653, 
      n5655, n5657, n5662, n5663, n5665, n5667, n5672, n5673, n5675, n5677, 
      n5682, n5683, n5685, n5687, n5692, n5693, n5695, n5697, n5699, n5701, 
      n5703, n5705, n5707, n5709, n5711, n5713, n5715, n5717, n5719, n5721, 
      n5723, n5725, n5727, n5729, n5731, n5733, n5735, n5737, n5739, n5741, 
      n5743, n5745, n5747, n5749, n5751, n5753, n5755, n5757, n5759, n5761, 
      n5763, n5765, n5767, n5769, n5771, n5773, n5775, n5776, n5777, n5778, 
      n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, 
      n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, 
      n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, 
      n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, 
      n5819, n5820, n5822, n5824, n5890, n5891, n5892, n5893, n5894, n5895, 
      n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, 
      n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, 
      n5916, n5917, n5918, n5919, n5920, n5921, n5954, n5955, n5956, n5957, 
      n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, 
      n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, 
      n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n6018, n6019, 
      n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, 
      n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, 
      n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, 
      n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, 
      n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, 
      n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, 
      n6080, n6081, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, 
      n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, 
      n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, 
      n6174, n6175, n6176, n6177, n6210, n6211, n6212, n6213, n6214, n6215, 
      n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, 
      n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, 
      n6236, n6237, n6238, n6239, n6240, n6241, n6659, n6661, n6663, n6665, 
      n6667, n6669, n6671, n6673, n6675, n6677, n6679, n6681, n6683, n6685, 
      n6687, n6689, n6691, n6693, n6695, n6697, n6699, n6701, n6703, n6705, 
      n6707, n6709, n6711, n6713, n6715, n6717, n6719, n6721, n6723, n6725, 
      n6727, n6729, n6731, n6733, n6735, n6737, n6739, n6741, n6743, n6745, 
      n6747, n6749, n6751, n6753, n6755, n6757, n6759, n6761, n6763, n6765, 
      n6767, n6769, n6771, n6773, n6775, n6777, n6779, n6781, n6783, n6785, 
      n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, 
      n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, 
      n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6830, n6831, 
      n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, 
      n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, 
      n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, 
      n6890, n6891, n6892, n6893, n6914, n6915, n6916, n6917, n6918, n6919, 
      n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, 
      n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, 
      n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, 
      n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, 
      n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, 
      n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, 
      n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, 
      n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, 
      n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, 
      n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, 
      n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, 
      n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, 
      n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, 
      n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, 
      n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, 
      n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, 
      n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, 
      n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, 
      n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, 
      n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, 
      n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, 
      n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, 
      n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, 
      n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, 
      n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, 
      n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, 
      n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, 
      n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, 
      n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, 
      n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, 
      n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, 
      n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, 
      n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, 
      n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n2832, n2833, 
      n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, 
      n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, 
      n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, 
      n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, 
      n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, 
      n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, 
      n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, 
      n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, 
      n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, 
      n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, 
      n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, 
      n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, 
      n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, 
      n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, 
      n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, 
      n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, 
      n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, 
      n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, 
      n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, 
      n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, 
      n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, 
      n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, 
      n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, 
      n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, 
      n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, 
      n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, 
      n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, 
      n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, 
      n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, 
      n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, 
      n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, 
      n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, 
      n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, 
      n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, 
      n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, 
      n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, 
      n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, 
      n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, 
      n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, 
      n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, 
      n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, 
      n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, 
      n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, 
      n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, 
      n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, 
      n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, 
      n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, 
      n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, 
      n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, 
      n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, 
      n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, 
      n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, 
      n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, 
      n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, 
      n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, 
      n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, 
      n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, 
      n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, 
      n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, 
      n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, 
      n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, 
      n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, 
      n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, 
      n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, 
      n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, 
      n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, 
      n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, 
      n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, 
      n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, 
      n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, 
      n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, 
      n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, 
      n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, 
      n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, 
      n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, 
      n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, 
      n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, 
      n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, 
      n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, 
      n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, 
      n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, 
      n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, 
      n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, 
      n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, 
      n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, 
      n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, 
      n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, 
      n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, 
      n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, 
      n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, 
      n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, 
      n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, 
      n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, 
      n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, 
      n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, 
      n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, 
      n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, 
      n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, 
      n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, 
      n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, 
      n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, 
      n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, 
      n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, 
      n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, 
      n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, 
      n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, 
      n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, 
      n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, 
      n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, 
      n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, 
      n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, 
      n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, 
      n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, 
      n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, 
      n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, 
      n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, 
      n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, 
      n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, 
      n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, 
      n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, 
      n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, 
      n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, 
      n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, 
      n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, 
      n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, 
      n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, 
      n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, 
      n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, 
      n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, 
      n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, 
      n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, 
      n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, 
      n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, 
      n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, 
      n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, 
      n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, 
      n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, 
      n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, 
      n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, 
      n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, 
      n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, 
      n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, 
      n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, 
      n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, 
      n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, 
      n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, 
      n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, 
      n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, 
      n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, 
      n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, 
      n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, 
      n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, 
      n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, 
      n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, 
      n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, 
      n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, 
      n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, 
      n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, 
      n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, 
      n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, 
      n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, 
      n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, 
      n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, 
      n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, 
      n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, 
      n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, 
      n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, 
      n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, 
      n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, 
      n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, 
      n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, 
      n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, 
      n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, 
      n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, 
      n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, 
      n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, 
      n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, 
      n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, 
      n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, 
      n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, 
      n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, 
      n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, 
      n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, 
      n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, 
      n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, 
      n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, 
      n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, 
      n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, 
      n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, 
      n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, 
      n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, 
      n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, 
      n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, 
      n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, 
      n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, 
      n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, 
      n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, 
      n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, 
      n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, 
      n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, 
      n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, 
      n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, 
      n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, 
      n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, 
      n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, 
      n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, 
      n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, 
      n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, 
      n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, 
      n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, 
      n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, 
      n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, 
      n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, 
      n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, 
      n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, 
      n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, 
      n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, 
      n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, 
      n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, 
      n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, 
      n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, 
      n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, 
      n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, 
      n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, 
      n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, 
      n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, 
      n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, 
      n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, 
      n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, 
      n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, 
      n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, 
      n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, 
      n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, 
      n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, 
      n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, 
      n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, 
      n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, 
      n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, 
      n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, 
      n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, 
      n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, 
      n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, 
      n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, 
      n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, 
      n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, 
      n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, 
      n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, 
      n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, 
      n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, 
      n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, 
      n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, 
      n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, 
      n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, 
      n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, 
      n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5384, 
      n5386, n5388, n5389, n5390, n5391, n5392, n5394, n5396, n5398, n5399, 
      n5400, n5401, n5402, n5404, n5406, n5408, n5409, n5410, n5411, n5412, 
      n5414, n5416, n5418, n5419, n5420, n5421, n5422, n5424, n5426, n5428, 
      n5429, n5430, n5431, n5432, n5434, n5436, n5438, n5439, n5440, n5441, 
      n5442, n5444, n5446, n5448, n5449, n5450, n5451, n5454, n5456, n5458, 
      n5459, n5460, n5461, n5464, n5466, n5468, n5469, n5470, n5471, n5474, 
      n5476, n5478, n5479, n5480, n5481, n5484, n5486, n5488, n5489, n5490, 
      n5491, n5494, n5496, n5498, n5499, n5500, n5501, n5504, n5506, n5508, 
      n5509, n5510, n5511, n5514, n5516, n5518, n5519, n5520, n5521, n5524, 
      n5526, n5528, n5529, n5530, n5531, n5534, n5536, n5538, n5539, n5540, 
      n5541, n5544, n5546, n5548, n5549, n5550, n5551, n5554, n5556, n5558, 
      n5559, n5560, n5561, n5564, n5566, n5568, n5569, n5570, n5571, n5574, 
      n5576, n5578, n5579, n5580, n5581, n5584, n5586, n5588, n5589, n5590, 
      n5591, n5594, n5596, n5598, n5599, n5600, n5601, n5604, n5606, n5608, 
      n5609, n5610, n5611, n5614, n5616, n5618, n5619, n5620, n5621, n5624, 
      n5626, n5628, n5629, n5630, n5631, n5634, n5636, n5638, n5639, n5640, 
      n5641, n5644, n5646, n5648, n5649, n5650, n5651, n5654, n5656, n5658, 
      n5659, n5660, n5661, n5664, n5666, n5668, n5669, n5670, n5671, n5674, 
      n5676, n5678, n5679, n5680, n5681, n5684, n5686, n5688, n5689, n5690, 
      n5691, n5694, n5696, n5698, n5700, n5702, n5704, n5706, n5708, n5710, 
      n5712, n5714, n5716, n5718, n5720, n5722, n5724, n5726, n5728, n5730, 
      n5732, n5734, n5736, n5738, n5740, n5742, n5744, n5746, n5748, n5750, 
      n5752, n5754, n12645, n12646, n12647, n12648, n12649, n12650, n12651, 
      n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660, 
      n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669, 
      n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678, 
      n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687, 
      n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696, 
      n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705, 
      n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714, 
      n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723, 
      n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732, 
      n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741, 
      n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750, 
      n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759, 
      n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768, 
      n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777, 
      n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786, 
      n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795, 
      n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804, 
      n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813, 
      n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822, 
      n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831, 
      n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840, 
      n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849, 
      n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858, 
      n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867, 
      n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876, 
      n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885, 
      n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894, 
      n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903, 
      n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912, 
      n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921, 
      n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930, 
      n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939, 
      n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948, 
      n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957, 
      n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966, 
      n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975, 
      n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984, 
      n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993, 
      n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002, 
      n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011, 
      n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020, 
      n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029, 
      n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038, 
      n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047, 
      n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056, 
      n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065, 
      n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074, 
      n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083, 
      n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092, 
      n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101, 
      n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110, 
      n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119, 
      n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128, 
      n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137, 
      n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146, 
      n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155, 
      n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164, 
      n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173, 
      n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182, 
      n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191, 
      n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200, 
      n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209, 
      n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218, 
      n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227, 
      n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236, 
      n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245, 
      n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254, 
      n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263, 
      n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272, 
      n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281, 
      n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290, 
      n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299, 
      n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308, 
      n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317, 
      n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326, 
      n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335, 
      n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344, 
      n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353, 
      n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362, 
      n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371, 
      n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380, 
      n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389, 
      n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398, 
      n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407, 
      n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416, 
      n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425, 
      n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434, 
      n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443, 
      n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452, 
      n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461, 
      n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470, 
      n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479, 
      n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488, 
      n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497, 
      n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506, 
      n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515, 
      n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524, 
      n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533, 
      n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542, 
      n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551, 
      n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560, 
      n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569, 
      n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578, 
      n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587, 
      n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596, 
      n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605, 
      n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614, 
      n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623, 
      n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632, 
      n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641, 
      n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650, 
      n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659, 
      n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668, 
      n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677, 
      n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686, 
      n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695, 
      n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704, 
      n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713, 
      n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722, 
      n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731, 
      n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740, 
      n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749, 
      n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758, 
      n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767, 
      n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776, 
      n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785, 
      n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794, 
      n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803, 
      n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812, 
      n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821, 
      n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829, n13830, 
      n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839, 
      n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848, 
      n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857, 
      n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866, 
      n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875, 
      n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884, 
      n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893, 
      n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901, n13902, 
      n13903, n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911, 
      n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920, 
      n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929, 
      n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938, 
      n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947, 
      n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956, 
      n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965, 
      n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973, n13974, 
      n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983, 
      n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992, 
      n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001, 
      n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010, 
      n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019, 
      n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028, 
      n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037, 
      n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046, 
      n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055, 
      n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064, 
      n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073, 
      n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082, 
      n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091, 
      n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100, 
      n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109, 
      n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118, 
      n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127, 
      n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136, 
      n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145, 
      n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154, 
      n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163, 
      n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172, 
      n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181, 
      n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190, 
      n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199, 
      n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208, 
      n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217, 
      n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226, 
      n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235, 
      n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244, 
      n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253, 
      n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262, 
      n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271, 
      n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280, 
      n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289, 
      n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298, 
      n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307, 
      n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316, 
      n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325, 
      n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334, 
      n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343, 
      n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352, 
      n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361, 
      n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370, 
      n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379, 
      n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388, 
      n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397, 
      n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406, 
      n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415, 
      n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424, 
      n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433, 
      n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442, 
      n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451, 
      n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460, 
      n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469, 
      n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478, 
      n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487, 
      n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496, 
      n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505, 
      n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514, 
      n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523, 
      n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532, 
      n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541, 
      n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550, 
      n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559, 
      n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568, 
      n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577, 
      n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586, 
      n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595, 
      n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604, 
      n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613, 
      n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622, 
      n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631, 
      n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640, 
      n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649, 
      n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658, 
      n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667, 
      n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676, 
      n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685, 
      n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694, 
      n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703, 
      n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712, 
      n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721, 
      n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730, 
      n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739, 
      n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748, 
      n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757, 
      n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766, 
      n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775, 
      n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784, 
      n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793, 
      n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802, 
      n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811, 
      n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820, 
      n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829, 
      n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838, 
      n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847, 
      n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856, 
      n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865, 
      n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874, 
      n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883, 
      n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892, 
      n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901, 
      n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910, 
      n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919, 
      n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928, 
      n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937, 
      n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946, 
      n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955, 
      n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964, 
      n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973, 
      n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982, 
      n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991, 
      n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000, 
      n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009, 
      n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018, 
      n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027, 
      n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036, 
      n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045, 
      n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054, 
      n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063, 
      n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072, 
      n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081, 
      n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090, 
      n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099, 
      n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108, 
      n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117, 
      n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126, 
      n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135, 
      n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144, 
      n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153, 
      n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162, 
      n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171, 
      n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179, n15180, 
      n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189, 
      n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198, 
      n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207, 
      n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216, 
      n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225, 
      n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234, 
      n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243, 
      n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252, 
      n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261, 
      n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270, 
      n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279, 
      n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288, 
      n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297, 
      n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306, 
      n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315, 
      n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324, 
      n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333, 
      n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342, 
      n15343, n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351, 
      n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360, 
      n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369, 
      n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378, 
      n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387, 
      n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396, 
      n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405, 
      n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414, 
      n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423, 
      n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432, 
      n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441, 
      n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450, 
      n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459, 
      n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468, 
      n15469, n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477, 
      n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15485, n15486, 
      n15487, n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495, 
      n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504, 
      n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513, 
      n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522, 
      n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531, 
      n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540, 
      n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549, 
      n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557, n15558, 
      n15559, n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567, 
      n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576, 
      n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585, 
      n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594, 
      n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603, 
      n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612, 
      n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621, 
      n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629, n15630, 
      n15631, n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639, 
      n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648, 
      n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657, 
      n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666, 
      n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674, n15675, 
      n15676, n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684, 
      n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693, 
      n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701, n15702, 
      n15703, n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711, 
      n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720, 
      n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729, 
      n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738, 
      n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746, n15747, 
      n15748, n15749, n15750, n15751, n15752, n15753, n15754, n15755, n15756, 
      n15757, n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765, 
      n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773, n15774, 
      n15775, n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783, 
      n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792, 
      n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801, 
      n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810, 
      n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818, n15819, 
      n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827, n15828, 
      n15829, n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837, 
      n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845, n15846, 
      n15847, n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855, 
      n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864, 
      n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873, 
      n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882, 
      n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890, n15891, 
      n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899, n15900, 
      n15901, n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909, 
      n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917, n15918, 
      n15919, n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927, 
      n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936, 
      n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945, 
      n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954, 
      n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962, n15963, 
      n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971, n15972, 
      n15973, n15974, n15975, n15976, n15977, n15978, n15979, n15980, n15981, 
      n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989, n15990, 
      n15991, n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999, 
      n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008, 
      n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017, 
      n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026, 
      n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034, n16035, 
      n16036, n16037, n16038, n16039, n16040, n16041, n16042, n16043, n16044, 
      n16045, n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053, 
      n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061, n16062, 
      n16063, n16064, n16065, n16066, n16067, n16068, n16069, n16070, n16071, 
      n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080, 
      n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089, 
      n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098, 
      n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106, n16107, 
      n_1002, n_1003, n_1004, n_1005, n_1006, n_1007, n_1008, n_1009, n_1010, 
      n_1011, n_1012, n_1013, n_1014, n_1015, n_1016, n_1017, n_1018, n_1019, 
      n_1020, n_1021, n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, n_1028, 
      n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, n_1037, 
      n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, n_1044, n_1045, n_1046, 
      n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, n_1055, 
      n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, 
      n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, 
      n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, 
      n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, 
      n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, 
      n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, 
      n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, 
      n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, n_1127, 
      n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, 
      n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, n_1145, 
      n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, 
      n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, 
      n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, 
      n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, 
      n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, 
      n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, 
      n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, 
      n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, 
      n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, 
      n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, 
      n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, 
      n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, 
      n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, 
      n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, 
      n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, 
      n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, 
      n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, 
      n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, 
      n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, 
      n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, 
      n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, 
      n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, 
      n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, 
      n_1353, n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, 
      n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, 
      n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, 
      n_1380, n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, 
      n_1389, n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, 
      n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, 
      n_1407, n_1408, n_1409, n_1410, n_1411, n_1412, n_1413, n_1414, n_1415, 
      n_1416, n_1417, n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, 
      n_1425, n_1426, n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, 
      n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, 
      n_1443, n_1444, n_1445, n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, 
      n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, 
      n_1461, n_1462, n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, 
      n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, 
      n_1479, n_1480, n_1481, n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, 
      n_1488, n_1489, n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, 
      n_1497, n_1498, n_1499, n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, 
      n_1506, n_1507, n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, 
      n_1515, n_1516, n_1517, n_1518, n_1519, n_1520, n_1521, n_1522, n_1523, 
      n_1524, n_1525, n_1526, n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, 
      n_1533, n_1534, n_1535, n_1536, n_1537, n_1538, n_1539, n_1540, n_1541, 
      n_1542, n_1543, n_1544, n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, 
      n_1551, n_1552, n_1553, n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, 
      n_1560, n_1561, n_1562, n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, 
      n_1569, n_1570, n_1571, n_1572, n_1573, n_1574, n_1575, n_1576, n_1577, 
      n_1578, n_1579, n_1580, n_1581, n_1582, n_1583, n_1584, n_1585, n_1586, 
      n_1587, n_1588, n_1589, n_1590, n_1591, n_1592, n_1593, n_1594, n_1595, 
      n_1596, n_1597, n_1598, n_1599, n_1600, n_1601, n_1602, n_1603, n_1604, 
      n_1605, n_1606, n_1607, n_1608, n_1609, n_1610, n_1611, n_1612, n_1613, 
      n_1614, n_1615, n_1616, n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, 
      n_1623, n_1624, n_1625, n_1626, n_1627, n_1628, n_1629, n_1630, n_1631, 
      n_1632, n_1633, n_1634, n_1635, n_1636, n_1637, n_1638, n_1639, n_1640, 
      n_1641, n_1642, n_1643, n_1644, n_1645, n_1646, n_1647, n_1648, n_1649, 
      n_1650, n_1651, n_1652, n_1653, n_1654, n_1655, n_1656, n_1657, n_1658, 
      n_1659, n_1660, n_1661, n_1662, n_1663, n_1664, n_1665, n_1666, n_1667, 
      n_1668, n_1669, n_1670, n_1671, n_1672, n_1673, n_1674, n_1675, n_1676, 
      n_1677, n_1678, n_1679, n_1680, n_1681, n_1682, n_1683, n_1684, n_1685, 
      n_1686, n_1687, n_1688, n_1689, n_1690, n_1691, n_1692, n_1693, n_1694, 
      n_1695, n_1696, n_1697, n_1698, n_1699, n_1700, n_1701, n_1702, n_1703, 
      n_1704, n_1705, n_1706, n_1707, n_1708, n_1709, n_1710, n_1711, n_1712, 
      n_1713, n_1714, n_1715, n_1716, n_1717, n_1718, n_1719, n_1720, n_1721, 
      n_1722, n_1723, n_1724, n_1725, n_1726, n_1727, n_1728, n_1729, n_1730, 
      n_1731, n_1732, n_1733, n_1734, n_1735, n_1736, n_1737, n_1738, n_1739, 
      n_1740, n_1741, n_1742, n_1743, n_1744, n_1745, n_1746, n_1747, n_1748, 
      n_1749, n_1750, n_1751, n_1752, n_1753, n_1754, n_1755, n_1756, n_1757, 
      n_1758, n_1759, n_1760, n_1761, n_1762, n_1763, n_1764, n_1765, n_1766, 
      n_1767, n_1768, n_1769, n_1770, n_1771, n_1772, n_1773, n_1774, n_1775, 
      n_1776, n_1777, n_1778, n_1779, n_1780, n_1781, n_1782, n_1783, n_1784, 
      n_1785, n_1786, n_1787, n_1788, n_1789, n_1790, n_1791, n_1792, n_1793, 
      n_1794, n_1795, n_1796, n_1797, n_1798, n_1799, n_1800, n_1801, n_1802, 
      n_1803, n_1804, n_1805, n_1806, n_1807, n_1808, n_1809, n_1810, n_1811, 
      n_1812, n_1813, n_1814, n_1815, n_1816, n_1817, n_1818, n_1819, n_1820, 
      n_1821, n_1822, n_1823, n_1824, n_1825, n_1826, n_1827, n_1828, n_1829, 
      n_1830, n_1831, n_1832, n_1833, n_1834, n_1835, n_1836, n_1837, n_1838, 
      n_1839, n_1840, n_1841, n_1842, n_1843, n_1844, n_1845, n_1846, n_1847, 
      n_1848, n_1849, n_1850, n_1851, n_1852, n_1853, n_1854, n_1855, n_1856, 
      n_1857, n_1858, n_1859, n_1860, n_1861, n_1862, n_1863, n_1864, n_1865, 
      n_1866, n_1867, n_1868, n_1869, n_1870, n_1871, n_1872, n_1873, n_1874, 
      n_1875, n_1876, n_1877, n_1878, n_1879, n_1880, n_1881, n_1882, n_1883, 
      n_1884, n_1885, n_1886, n_1887, n_1888, n_1889, n_1890, n_1891, n_1892, 
      n_1893, n_1894, n_1895, n_1896, n_1897, n_1898, n_1899, n_1900, n_1901, 
      n_1902, n_1903, n_1904, n_1905, n_1906, n_1907, n_1908, n_1909, n_1910, 
      n_1911, n_1912, n_1913, n_1914, n_1915, n_1916, n_1917, n_1918, n_1919, 
      n_1920, n_1921, n_1922, n_1923, n_1924, n_1925, n_1926, n_1927, n_1928, 
      n_1929, n_1930, n_1931, n_1932, n_1933, n_1934, n_1935, n_1936, n_1937, 
      n_1938, n_1939, n_1940, n_1941, n_1942, n_1943, n_1944, n_1945, n_1946, 
      n_1947, n_1948, n_1949, n_1950, n_1951, n_1952, n_1953, n_1954, n_1955, 
      n_1956, n_1957, n_1958, n_1959, n_1960, n_1961, n_1962, n_1963, n_1964, 
      n_1965, n_1966, n_1967, n_1968, n_1969, n_1970, n_1971, n_1972, n_1973, 
      n_1974, n_1975, n_1976, n_1977, n_1978, n_1979, n_1980, n_1981, n_1982, 
      n_1983, n_1984, n_1985, n_1986, n_1987, n_1988, n_1989, n_1990, n_1991, 
      n_1992, n_1993, n_1994, n_1995, n_1996, n_1997, n_1998, n_1999, n_2000, 
      n_2001, n_2002, n_2003, n_2004, n_2005, n_2006, n_2007, n_2008, n_2009, 
      n_2010, n_2011, n_2012, n_2013, n_2014, n_2015, n_2016, n_2017, n_2018, 
      n_2019, n_2020, n_2021, n_2022, n_2023, n_2024, n_2025, n_2026, n_2027, 
      n_2028, n_2029, n_2030, n_2031, n_2032, n_2033, n_2034, n_2035, n_2036, 
      n_2037, n_2038, n_2039, n_2040, n_2041, n_2042, n_2043, n_2044, n_2045, 
      n_2046, n_2047, n_2048, n_2049, n_2050, n_2051, n_2052, n_2053, n_2054, 
      n_2055, n_2056, n_2057, n_2058, n_2059, n_2060, n_2061, n_2062, n_2063, 
      n_2064, n_2065, n_2066, n_2067, n_2068, n_2069, n_2070, n_2071, n_2072, 
      n_2073, n_2074, n_2075, n_2076, n_2077, n_2078, n_2079, n_2080, n_2081, 
      n_2082, n_2083, n_2084, n_2085, n_2086, n_2087, n_2088, n_2089, n_2090, 
      n_2091, n_2092, n_2093, n_2094, n_2095, n_2096, n_2097, n_2098, n_2099, 
      n_2100, n_2101, n_2102, n_2103, n_2104, n_2105, n_2106, n_2107, n_2108, 
      n_2109, n_2110, n_2111, n_2112, n_2113, n_2114, n_2115, n_2116, n_2117, 
      n_2118, n_2119, n_2120, n_2121, n_2122, n_2123, n_2124, n_2125, n_2126, 
      n_2127, n_2128, n_2129, n_2130, n_2131, n_2132, n_2133, n_2134, n_2135, 
      n_2136, n_2137, n_2138, n_2139, n_2140, n_2141, n_2142, n_2143, n_2144, 
      n_2145, n_2146, n_2147, n_2148, n_2149, n_2150, n_2151, n_2152, n_2153, 
      n_2154, n_2155, n_2156, n_2157, n_2158, n_2159, n_2160, n_2161, n_2162, 
      n_2163, n_2164, n_2165, n_2166, n_2167, n_2168, n_2169, n_2170, n_2171, 
      n_2172, n_2173, n_2174, n_2175, n_2176, n_2177, n_2178, n_2179, n_2180, 
      n_2181, n_2182, n_2183, n_2184, n_2185, n_2186, n_2187, n_2188, n_2189, 
      n_2190, n_2191, n_2192, n_2193, n_2194, n_2195, n_2196, n_2197, n_2198, 
      n_2199, n_2200, n_2201, n_2202, n_2203, n_2204, n_2205, n_2206, n_2207, 
      n_2208, n_2209, n_2210, n_2211, n_2212, n_2213, n_2214, n_2215, n_2216, 
      n_2217 : std_logic;

begin
   
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n9913, CK => CLK, Q => n714,
                           QN => n12648);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n9912, CK => CLK, Q => n717,
                           QN => n12647);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n9911, CK => CLK, Q => n720,
                           QN => n12646);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n9910, CK => CLK, Q => n723,
                           QN => n12645);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n9909, CK => CLK, Q => n726,
                           QN => n12652);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n9908, CK => CLK, Q => n729,
                           QN => n12651);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n9907, CK => CLK, Q => n732,
                           QN => n12650);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n9906, CK => CLK, Q => n735,
                           QN => n12649);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n9905, CK => CLK, Q => n738,
                           QN => n12708);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n9904, CK => CLK, Q => n741,
                           QN => n12706);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n9903, CK => CLK, Q => n744,
                           QN => n12704);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n9902, CK => CLK, Q => n747,
                           QN => n12702);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n9901, CK => CLK, Q => n750,
                           QN => n12700);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n9900, CK => CLK, Q => n753,
                           QN => n12698);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n9899, CK => CLK, Q => n756,
                           QN => n12696);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n9898, CK => CLK, Q => n759,
                           QN => n12694);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n9897, CK => CLK, Q => n762,
                           QN => n12692);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n9896, CK => CLK, Q => n765,
                           QN => n12690);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n9895, CK => CLK, Q => n768,
                           QN => n12688);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n9894, CK => CLK, Q => n771,
                           QN => n12686);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n9893, CK => CLK, Q => n774,
                           QN => n12684);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n9892, CK => CLK, Q => n777,
                           QN => n12682);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n9891, CK => CLK, Q => n780, 
                           QN => n12680);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n9890, CK => CLK, Q => n783, 
                           QN => n12678);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n9889, CK => CLK, Q => n786, 
                           QN => n12676);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n9888, CK => CLK, Q => n789, 
                           QN => n12674);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n9887, CK => CLK, Q => n792, 
                           QN => n12672);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n9886, CK => CLK, Q => n795, 
                           QN => n12670);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n9885, CK => CLK, Q => n798, 
                           QN => n12668);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n9884, CK => CLK, Q => n801, 
                           QN => n12666);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n9883, CK => CLK, Q => n804, 
                           QN => n12664);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n9882, CK => CLK, Q => n807, 
                           QN => n12662);
   REGISTERS_reg_6_31_inst : DFF_X1 port map( D => n9785, CK => CLK, Q => 
                           n_1002, QN => n14108);
   REGISTERS_reg_6_30_inst : DFF_X1 port map( D => n9784, CK => CLK, Q => 
                           n_1003, QN => n14109);
   REGISTERS_reg_6_29_inst : DFF_X1 port map( D => n9783, CK => CLK, Q => 
                           n_1004, QN => n14110);
   REGISTERS_reg_6_28_inst : DFF_X1 port map( D => n9782, CK => CLK, Q => 
                           n_1005, QN => n14111);
   REGISTERS_reg_6_27_inst : DFF_X1 port map( D => n9781, CK => CLK, Q => 
                           n_1006, QN => n14112);
   REGISTERS_reg_6_26_inst : DFF_X1 port map( D => n9780, CK => CLK, Q => 
                           n_1007, QN => n14113);
   REGISTERS_reg_6_25_inst : DFF_X1 port map( D => n9779, CK => CLK, Q => 
                           n_1008, QN => n14114);
   REGISTERS_reg_6_24_inst : DFF_X1 port map( D => n9778, CK => CLK, Q => 
                           n_1009, QN => n14115);
   REGISTERS_reg_6_23_inst : DFF_X1 port map( D => n9777, CK => CLK, Q => 
                           n_1010, QN => n14116);
   REGISTERS_reg_6_22_inst : DFF_X1 port map( D => n9776, CK => CLK, Q => 
                           n_1011, QN => n14117);
   REGISTERS_reg_6_21_inst : DFF_X1 port map( D => n9775, CK => CLK, Q => 
                           n_1012, QN => n14118);
   REGISTERS_reg_6_20_inst : DFF_X1 port map( D => n9774, CK => CLK, Q => 
                           n_1013, QN => n14119);
   REGISTERS_reg_6_19_inst : DFF_X1 port map( D => n9773, CK => CLK, Q => 
                           n_1014, QN => n14120);
   REGISTERS_reg_6_18_inst : DFF_X1 port map( D => n9772, CK => CLK, Q => 
                           n_1015, QN => n14121);
   REGISTERS_reg_6_17_inst : DFF_X1 port map( D => n9771, CK => CLK, Q => 
                           n_1016, QN => n14122);
   REGISTERS_reg_6_16_inst : DFF_X1 port map( D => n9770, CK => CLK, Q => 
                           n_1017, QN => n14123);
   REGISTERS_reg_6_15_inst : DFF_X1 port map( D => n9769, CK => CLK, Q => 
                           n_1018, QN => n14124);
   REGISTERS_reg_6_14_inst : DFF_X1 port map( D => n9768, CK => CLK, Q => 
                           n_1019, QN => n14125);
   REGISTERS_reg_6_13_inst : DFF_X1 port map( D => n9767, CK => CLK, Q => 
                           n_1020, QN => n14126);
   REGISTERS_reg_6_12_inst : DFF_X1 port map( D => n9766, CK => CLK, Q => 
                           n_1021, QN => n14127);
   REGISTERS_reg_6_11_inst : DFF_X1 port map( D => n9765, CK => CLK, Q => 
                           n_1022, QN => n14128);
   REGISTERS_reg_6_10_inst : DFF_X1 port map( D => n9764, CK => CLK, Q => 
                           n_1023, QN => n14129);
   REGISTERS_reg_6_9_inst : DFF_X1 port map( D => n9763, CK => CLK, Q => n_1024
                           , QN => n14130);
   REGISTERS_reg_6_8_inst : DFF_X1 port map( D => n9762, CK => CLK, Q => n_1025
                           , QN => n14131);
   REGISTERS_reg_6_7_inst : DFF_X1 port map( D => n9761, CK => CLK, Q => n_1026
                           , QN => n14132);
   REGISTERS_reg_6_6_inst : DFF_X1 port map( D => n9760, CK => CLK, Q => n_1027
                           , QN => n14133);
   REGISTERS_reg_6_5_inst : DFF_X1 port map( D => n9759, CK => CLK, Q => n_1028
                           , QN => n14134);
   REGISTERS_reg_6_4_inst : DFF_X1 port map( D => n9758, CK => CLK, Q => n_1029
                           , QN => n14135);
   REGISTERS_reg_6_3_inst : DFF_X1 port map( D => n9757, CK => CLK, Q => n_1030
                           , QN => n14136);
   REGISTERS_reg_6_2_inst : DFF_X1 port map( D => n9756, CK => CLK, Q => n_1031
                           , QN => n14137);
   REGISTERS_reg_6_1_inst : DFF_X1 port map( D => n9755, CK => CLK, Q => n_1032
                           , QN => n14138);
   REGISTERS_reg_6_0_inst : DFF_X1 port map( D => n9754, CK => CLK, Q => n_1033
                           , QN => n14139);
   REGISTERS_reg_7_31_inst : DFF_X1 port map( D => n9753, CK => CLK, Q => 
                           n_1034, QN => n14140);
   REGISTERS_reg_7_30_inst : DFF_X1 port map( D => n9752, CK => CLK, Q => 
                           n_1035, QN => n14141);
   REGISTERS_reg_7_29_inst : DFF_X1 port map( D => n9751, CK => CLK, Q => 
                           n_1036, QN => n14142);
   REGISTERS_reg_7_28_inst : DFF_X1 port map( D => n9750, CK => CLK, Q => 
                           n_1037, QN => n14143);
   REGISTERS_reg_7_27_inst : DFF_X1 port map( D => n9749, CK => CLK, Q => 
                           n_1038, QN => n14144);
   REGISTERS_reg_7_26_inst : DFF_X1 port map( D => n9748, CK => CLK, Q => 
                           n_1039, QN => n14145);
   REGISTERS_reg_7_25_inst : DFF_X1 port map( D => n9747, CK => CLK, Q => 
                           n_1040, QN => n14146);
   REGISTERS_reg_7_24_inst : DFF_X1 port map( D => n9746, CK => CLK, Q => 
                           n_1041, QN => n14147);
   REGISTERS_reg_7_23_inst : DFF_X1 port map( D => n9745, CK => CLK, Q => 
                           n_1042, QN => n14148);
   REGISTERS_reg_7_22_inst : DFF_X1 port map( D => n9744, CK => CLK, Q => 
                           n_1043, QN => n14149);
   REGISTERS_reg_7_21_inst : DFF_X1 port map( D => n9743, CK => CLK, Q => 
                           n_1044, QN => n14150);
   REGISTERS_reg_7_20_inst : DFF_X1 port map( D => n9742, CK => CLK, Q => 
                           n_1045, QN => n14151);
   REGISTERS_reg_7_19_inst : DFF_X1 port map( D => n9741, CK => CLK, Q => 
                           n_1046, QN => n14152);
   REGISTERS_reg_7_18_inst : DFF_X1 port map( D => n9740, CK => CLK, Q => 
                           n_1047, QN => n14153);
   REGISTERS_reg_7_17_inst : DFF_X1 port map( D => n9739, CK => CLK, Q => 
                           n_1048, QN => n14154);
   REGISTERS_reg_7_16_inst : DFF_X1 port map( D => n9738, CK => CLK, Q => 
                           n_1049, QN => n14155);
   REGISTERS_reg_7_15_inst : DFF_X1 port map( D => n9737, CK => CLK, Q => 
                           n_1050, QN => n14156);
   REGISTERS_reg_7_14_inst : DFF_X1 port map( D => n9736, CK => CLK, Q => 
                           n_1051, QN => n14157);
   REGISTERS_reg_7_13_inst : DFF_X1 port map( D => n9735, CK => CLK, Q => 
                           n_1052, QN => n14158);
   REGISTERS_reg_7_12_inst : DFF_X1 port map( D => n9734, CK => CLK, Q => 
                           n_1053, QN => n14159);
   REGISTERS_reg_7_11_inst : DFF_X1 port map( D => n9733, CK => CLK, Q => 
                           n_1054, QN => n14160);
   REGISTERS_reg_7_10_inst : DFF_X1 port map( D => n9732, CK => CLK, Q => 
                           n_1055, QN => n14161);
   REGISTERS_reg_7_9_inst : DFF_X1 port map( D => n9731, CK => CLK, Q => n_1056
                           , QN => n14162);
   REGISTERS_reg_7_8_inst : DFF_X1 port map( D => n9730, CK => CLK, Q => n_1057
                           , QN => n14163);
   REGISTERS_reg_7_7_inst : DFF_X1 port map( D => n9729, CK => CLK, Q => n_1058
                           , QN => n14164);
   REGISTERS_reg_7_6_inst : DFF_X1 port map( D => n9728, CK => CLK, Q => n_1059
                           , QN => n14165);
   REGISTERS_reg_7_5_inst : DFF_X1 port map( D => n9727, CK => CLK, Q => n_1060
                           , QN => n14166);
   REGISTERS_reg_7_4_inst : DFF_X1 port map( D => n9726, CK => CLK, Q => n_1061
                           , QN => n14167);
   REGISTERS_reg_7_3_inst : DFF_X1 port map( D => n9725, CK => CLK, Q => n_1062
                           , QN => n14168);
   REGISTERS_reg_7_2_inst : DFF_X1 port map( D => n9724, CK => CLK, Q => n_1063
                           , QN => n14169);
   REGISTERS_reg_7_1_inst : DFF_X1 port map( D => n9723, CK => CLK, Q => n_1064
                           , QN => n14170);
   REGISTERS_reg_7_0_inst : DFF_X1 port map( D => n9722, CK => CLK, Q => n_1065
                           , QN => n14171);
   REGISTERS_reg_8_31_inst : DFF_X1 port map( D => n9721, CK => CLK, Q => 
                           n_1066, QN => n14172);
   REGISTERS_reg_8_30_inst : DFF_X1 port map( D => n9720, CK => CLK, Q => 
                           n_1067, QN => n14173);
   REGISTERS_reg_8_29_inst : DFF_X1 port map( D => n9719, CK => CLK, Q => 
                           n_1068, QN => n14174);
   REGISTERS_reg_8_28_inst : DFF_X1 port map( D => n9718, CK => CLK, Q => 
                           n_1069, QN => n14175);
   REGISTERS_reg_8_27_inst : DFF_X1 port map( D => n9717, CK => CLK, Q => 
                           n_1070, QN => n14176);
   REGISTERS_reg_8_26_inst : DFF_X1 port map( D => n9716, CK => CLK, Q => 
                           n_1071, QN => n14177);
   REGISTERS_reg_8_25_inst : DFF_X1 port map( D => n9715, CK => CLK, Q => 
                           n_1072, QN => n14178);
   REGISTERS_reg_8_24_inst : DFF_X1 port map( D => n9714, CK => CLK, Q => 
                           n_1073, QN => n14179);
   REGISTERS_reg_8_23_inst : DFF_X1 port map( D => n9713, CK => CLK, Q => 
                           n_1074, QN => n14180);
   REGISTERS_reg_8_22_inst : DFF_X1 port map( D => n9712, CK => CLK, Q => 
                           n_1075, QN => n14181);
   REGISTERS_reg_8_21_inst : DFF_X1 port map( D => n9711, CK => CLK, Q => 
                           n_1076, QN => n14182);
   REGISTERS_reg_8_20_inst : DFF_X1 port map( D => n9710, CK => CLK, Q => 
                           n_1077, QN => n14183);
   REGISTERS_reg_8_19_inst : DFF_X1 port map( D => n9709, CK => CLK, Q => 
                           n_1078, QN => n14184);
   REGISTERS_reg_8_18_inst : DFF_X1 port map( D => n9708, CK => CLK, Q => 
                           n_1079, QN => n14185);
   REGISTERS_reg_8_17_inst : DFF_X1 port map( D => n9707, CK => CLK, Q => 
                           n_1080, QN => n14186);
   REGISTERS_reg_8_16_inst : DFF_X1 port map( D => n9706, CK => CLK, Q => 
                           n_1081, QN => n14187);
   REGISTERS_reg_8_15_inst : DFF_X1 port map( D => n9705, CK => CLK, Q => 
                           n_1082, QN => n14188);
   REGISTERS_reg_8_14_inst : DFF_X1 port map( D => n9704, CK => CLK, Q => 
                           n_1083, QN => n14189);
   REGISTERS_reg_8_13_inst : DFF_X1 port map( D => n9703, CK => CLK, Q => 
                           n_1084, QN => n14190);
   REGISTERS_reg_8_12_inst : DFF_X1 port map( D => n9702, CK => CLK, Q => 
                           n_1085, QN => n14191);
   REGISTERS_reg_8_11_inst : DFF_X1 port map( D => n9701, CK => CLK, Q => 
                           n_1086, QN => n14192);
   REGISTERS_reg_8_10_inst : DFF_X1 port map( D => n9700, CK => CLK, Q => 
                           n_1087, QN => n14193);
   REGISTERS_reg_8_9_inst : DFF_X1 port map( D => n9699, CK => CLK, Q => n_1088
                           , QN => n14194);
   REGISTERS_reg_8_8_inst : DFF_X1 port map( D => n9698, CK => CLK, Q => n_1089
                           , QN => n14195);
   REGISTERS_reg_8_7_inst : DFF_X1 port map( D => n9697, CK => CLK, Q => n_1090
                           , QN => n14196);
   REGISTERS_reg_8_6_inst : DFF_X1 port map( D => n9696, CK => CLK, Q => n_1091
                           , QN => n14197);
   REGISTERS_reg_8_5_inst : DFF_X1 port map( D => n9695, CK => CLK, Q => n_1092
                           , QN => n14198);
   REGISTERS_reg_8_4_inst : DFF_X1 port map( D => n9694, CK => CLK, Q => n_1093
                           , QN => n14199);
   REGISTERS_reg_8_3_inst : DFF_X1 port map( D => n9693, CK => CLK, Q => n_1094
                           , QN => n14200);
   REGISTERS_reg_8_2_inst : DFF_X1 port map( D => n9692, CK => CLK, Q => n_1095
                           , QN => n14201);
   REGISTERS_reg_8_1_inst : DFF_X1 port map( D => n9691, CK => CLK, Q => n_1096
                           , QN => n14202);
   REGISTERS_reg_8_0_inst : DFF_X1 port map( D => n9690, CK => CLK, Q => n_1097
                           , QN => n14203);
   REGISTERS_reg_11_31_inst : DFF_X1 port map( D => n9625, CK => CLK, Q => n713
                           , QN => n12656);
   REGISTERS_reg_11_30_inst : DFF_X1 port map( D => n9624, CK => CLK, Q => n716
                           , QN => n12655);
   REGISTERS_reg_11_29_inst : DFF_X1 port map( D => n9623, CK => CLK, Q => n719
                           , QN => n12654);
   REGISTERS_reg_11_28_inst : DFF_X1 port map( D => n9622, CK => CLK, Q => n722
                           , QN => n12653);
   REGISTERS_reg_11_27_inst : DFF_X1 port map( D => n9621, CK => CLK, Q => n725
                           , QN => n12660);
   REGISTERS_reg_11_26_inst : DFF_X1 port map( D => n9620, CK => CLK, Q => n728
                           , QN => n12659);
   REGISTERS_reg_11_25_inst : DFF_X1 port map( D => n9619, CK => CLK, Q => n731
                           , QN => n12658);
   REGISTERS_reg_11_24_inst : DFF_X1 port map( D => n9618, CK => CLK, Q => n734
                           , QN => n12657);
   REGISTERS_reg_11_23_inst : DFF_X1 port map( D => n9617, CK => CLK, Q => n737
                           , QN => n12707);
   REGISTERS_reg_11_22_inst : DFF_X1 port map( D => n9616, CK => CLK, Q => n740
                           , QN => n12705);
   REGISTERS_reg_11_21_inst : DFF_X1 port map( D => n9615, CK => CLK, Q => n743
                           , QN => n12703);
   REGISTERS_reg_11_20_inst : DFF_X1 port map( D => n9614, CK => CLK, Q => n746
                           , QN => n12701);
   REGISTERS_reg_11_19_inst : DFF_X1 port map( D => n9613, CK => CLK, Q => n749
                           , QN => n12699);
   REGISTERS_reg_11_18_inst : DFF_X1 port map( D => n9612, CK => CLK, Q => n752
                           , QN => n12697);
   REGISTERS_reg_11_17_inst : DFF_X1 port map( D => n9611, CK => CLK, Q => n755
                           , QN => n12695);
   REGISTERS_reg_11_16_inst : DFF_X1 port map( D => n9610, CK => CLK, Q => n758
                           , QN => n12693);
   REGISTERS_reg_11_15_inst : DFF_X1 port map( D => n9609, CK => CLK, Q => n761
                           , QN => n12691);
   REGISTERS_reg_11_14_inst : DFF_X1 port map( D => n9608, CK => CLK, Q => n764
                           , QN => n12689);
   REGISTERS_reg_11_13_inst : DFF_X1 port map( D => n9607, CK => CLK, Q => n767
                           , QN => n12687);
   REGISTERS_reg_11_12_inst : DFF_X1 port map( D => n9606, CK => CLK, Q => n770
                           , QN => n12685);
   REGISTERS_reg_11_11_inst : DFF_X1 port map( D => n9605, CK => CLK, Q => n773
                           , QN => n12683);
   REGISTERS_reg_11_10_inst : DFF_X1 port map( D => n9604, CK => CLK, Q => n776
                           , QN => n12681);
   REGISTERS_reg_11_9_inst : DFF_X1 port map( D => n9603, CK => CLK, Q => n779,
                           QN => n12679);
   REGISTERS_reg_11_8_inst : DFF_X1 port map( D => n9602, CK => CLK, Q => n782,
                           QN => n12677);
   REGISTERS_reg_11_7_inst : DFF_X1 port map( D => n9601, CK => CLK, Q => n785,
                           QN => n12675);
   REGISTERS_reg_11_6_inst : DFF_X1 port map( D => n9600, CK => CLK, Q => n788,
                           QN => n12673);
   REGISTERS_reg_11_5_inst : DFF_X1 port map( D => n9599, CK => CLK, Q => n791,
                           QN => n12671);
   REGISTERS_reg_11_4_inst : DFF_X1 port map( D => n9598, CK => CLK, Q => n794,
                           QN => n12669);
   REGISTERS_reg_11_3_inst : DFF_X1 port map( D => n9597, CK => CLK, Q => n797,
                           QN => n12667);
   REGISTERS_reg_11_2_inst : DFF_X1 port map( D => n9596, CK => CLK, Q => n800,
                           QN => n12665);
   REGISTERS_reg_11_1_inst : DFF_X1 port map( D => n9595, CK => CLK, Q => n803,
                           QN => n12663);
   REGISTERS_reg_11_0_inst : DFF_X1 port map( D => n9594, CK => CLK, Q => n806,
                           QN => n12661);
   REGISTERS_reg_15_31_inst : DFF_X1 port map( D => n9497, CK => CLK, Q => 
                           n_1098, QN => n14280);
   REGISTERS_reg_15_30_inst : DFF_X1 port map( D => n9496, CK => CLK, Q => 
                           n_1099, QN => n14281);
   REGISTERS_reg_15_29_inst : DFF_X1 port map( D => n9495, CK => CLK, Q => 
                           n_1100, QN => n14282);
   REGISTERS_reg_15_28_inst : DFF_X1 port map( D => n9494, CK => CLK, Q => 
                           n_1101, QN => n14283);
   REGISTERS_reg_15_27_inst : DFF_X1 port map( D => n9493, CK => CLK, Q => 
                           n_1102, QN => n14284);
   REGISTERS_reg_15_26_inst : DFF_X1 port map( D => n9492, CK => CLK, Q => 
                           n_1103, QN => n14285);
   REGISTERS_reg_15_25_inst : DFF_X1 port map( D => n9491, CK => CLK, Q => 
                           n_1104, QN => n14286);
   REGISTERS_reg_15_24_inst : DFF_X1 port map( D => n9490, CK => CLK, Q => 
                           n_1105, QN => n14287);
   REGISTERS_reg_15_23_inst : DFF_X1 port map( D => n9489, CK => CLK, Q => 
                           n_1106, QN => n14288);
   REGISTERS_reg_15_22_inst : DFF_X1 port map( D => n9488, CK => CLK, Q => 
                           n_1107, QN => n14289);
   REGISTERS_reg_15_21_inst : DFF_X1 port map( D => n9487, CK => CLK, Q => 
                           n_1108, QN => n14290);
   REGISTERS_reg_15_20_inst : DFF_X1 port map( D => n9486, CK => CLK, Q => 
                           n_1109, QN => n14291);
   REGISTERS_reg_15_19_inst : DFF_X1 port map( D => n9485, CK => CLK, Q => 
                           n_1110, QN => n14292);
   REGISTERS_reg_15_18_inst : DFF_X1 port map( D => n9484, CK => CLK, Q => 
                           n_1111, QN => n14293);
   REGISTERS_reg_15_17_inst : DFF_X1 port map( D => n9483, CK => CLK, Q => 
                           n_1112, QN => n14294);
   REGISTERS_reg_15_16_inst : DFF_X1 port map( D => n9482, CK => CLK, Q => 
                           n_1113, QN => n14295);
   REGISTERS_reg_15_15_inst : DFF_X1 port map( D => n9481, CK => CLK, Q => 
                           n_1114, QN => n14296);
   REGISTERS_reg_15_14_inst : DFF_X1 port map( D => n9480, CK => CLK, Q => 
                           n_1115, QN => n14297);
   REGISTERS_reg_15_13_inst : DFF_X1 port map( D => n9479, CK => CLK, Q => 
                           n_1116, QN => n14298);
   REGISTERS_reg_15_12_inst : DFF_X1 port map( D => n9478, CK => CLK, Q => 
                           n_1117, QN => n14299);
   REGISTERS_reg_15_11_inst : DFF_X1 port map( D => n9477, CK => CLK, Q => 
                           n_1118, QN => n14300);
   REGISTERS_reg_15_10_inst : DFF_X1 port map( D => n9476, CK => CLK, Q => 
                           n_1119, QN => n14301);
   REGISTERS_reg_15_9_inst : DFF_X1 port map( D => n9475, CK => CLK, Q => 
                           n_1120, QN => n14302);
   REGISTERS_reg_15_8_inst : DFF_X1 port map( D => n9474, CK => CLK, Q => 
                           n_1121, QN => n14303);
   REGISTERS_reg_15_7_inst : DFF_X1 port map( D => n9473, CK => CLK, Q => 
                           n_1122, QN => n14304);
   REGISTERS_reg_15_6_inst : DFF_X1 port map( D => n9472, CK => CLK, Q => 
                           n_1123, QN => n14305);
   REGISTERS_reg_15_5_inst : DFF_X1 port map( D => n9471, CK => CLK, Q => 
                           n_1124, QN => n14306);
   REGISTERS_reg_15_4_inst : DFF_X1 port map( D => n9470, CK => CLK, Q => 
                           n_1125, QN => n14307);
   REGISTERS_reg_15_3_inst : DFF_X1 port map( D => n9469, CK => CLK, Q => 
                           n_1126, QN => n14308);
   REGISTERS_reg_15_2_inst : DFF_X1 port map( D => n9468, CK => CLK, Q => 
                           n_1127, QN => n14309);
   REGISTERS_reg_15_1_inst : DFF_X1 port map( D => n9467, CK => CLK, Q => 
                           n_1128, QN => n14310);
   REGISTERS_reg_15_0_inst : DFF_X1 port map( D => n9466, CK => CLK, Q => 
                           n_1129, QN => n14311);
   REGISTERS_reg_16_31_inst : DFF_X1 port map( D => n9465, CK => CLK, Q => 
                           n_1130, QN => n14312);
   REGISTERS_reg_16_30_inst : DFF_X1 port map( D => n9464, CK => CLK, Q => 
                           n_1131, QN => n14313);
   REGISTERS_reg_16_29_inst : DFF_X1 port map( D => n9463, CK => CLK, Q => 
                           n_1132, QN => n14314);
   REGISTERS_reg_16_28_inst : DFF_X1 port map( D => n9462, CK => CLK, Q => 
                           n_1133, QN => n14315);
   REGISTERS_reg_16_27_inst : DFF_X1 port map( D => n9461, CK => CLK, Q => 
                           n_1134, QN => n14316);
   REGISTERS_reg_16_26_inst : DFF_X1 port map( D => n9460, CK => CLK, Q => 
                           n_1135, QN => n14317);
   REGISTERS_reg_16_25_inst : DFF_X1 port map( D => n9459, CK => CLK, Q => 
                           n_1136, QN => n14318);
   REGISTERS_reg_16_24_inst : DFF_X1 port map( D => n9458, CK => CLK, Q => 
                           n_1137, QN => n14319);
   REGISTERS_reg_16_23_inst : DFF_X1 port map( D => n9457, CK => CLK, Q => 
                           n_1138, QN => n14320);
   REGISTERS_reg_16_22_inst : DFF_X1 port map( D => n9456, CK => CLK, Q => 
                           n_1139, QN => n14321);
   REGISTERS_reg_16_21_inst : DFF_X1 port map( D => n9455, CK => CLK, Q => 
                           n_1140, QN => n14322);
   REGISTERS_reg_16_20_inst : DFF_X1 port map( D => n9454, CK => CLK, Q => 
                           n_1141, QN => n14323);
   REGISTERS_reg_16_19_inst : DFF_X1 port map( D => n9453, CK => CLK, Q => 
                           n_1142, QN => n14324);
   REGISTERS_reg_16_18_inst : DFF_X1 port map( D => n9452, CK => CLK, Q => 
                           n_1143, QN => n14325);
   REGISTERS_reg_16_17_inst : DFF_X1 port map( D => n9451, CK => CLK, Q => 
                           n_1144, QN => n14326);
   REGISTERS_reg_16_16_inst : DFF_X1 port map( D => n9450, CK => CLK, Q => 
                           n_1145, QN => n14327);
   REGISTERS_reg_16_15_inst : DFF_X1 port map( D => n9449, CK => CLK, Q => 
                           n_1146, QN => n14328);
   REGISTERS_reg_16_14_inst : DFF_X1 port map( D => n9448, CK => CLK, Q => 
                           n_1147, QN => n14329);
   REGISTERS_reg_16_13_inst : DFF_X1 port map( D => n9447, CK => CLK, Q => 
                           n_1148, QN => n14330);
   REGISTERS_reg_16_12_inst : DFF_X1 port map( D => n9446, CK => CLK, Q => 
                           n_1149, QN => n14331);
   REGISTERS_reg_16_11_inst : DFF_X1 port map( D => n9445, CK => CLK, Q => 
                           n_1150, QN => n14332);
   REGISTERS_reg_16_10_inst : DFF_X1 port map( D => n9444, CK => CLK, Q => 
                           n_1151, QN => n14333);
   REGISTERS_reg_16_9_inst : DFF_X1 port map( D => n9443, CK => CLK, Q => 
                           n_1152, QN => n14334);
   REGISTERS_reg_16_8_inst : DFF_X1 port map( D => n9442, CK => CLK, Q => 
                           n_1153, QN => n14335);
   REGISTERS_reg_16_7_inst : DFF_X1 port map( D => n9441, CK => CLK, Q => 
                           n_1154, QN => n14336);
   REGISTERS_reg_16_6_inst : DFF_X1 port map( D => n9440, CK => CLK, Q => 
                           n_1155, QN => n14337);
   REGISTERS_reg_16_5_inst : DFF_X1 port map( D => n9439, CK => CLK, Q => 
                           n_1156, QN => n14338);
   REGISTERS_reg_16_4_inst : DFF_X1 port map( D => n9438, CK => CLK, Q => 
                           n_1157, QN => n14339);
   REGISTERS_reg_16_3_inst : DFF_X1 port map( D => n9437, CK => CLK, Q => 
                           n_1158, QN => n14340);
   REGISTERS_reg_16_2_inst : DFF_X1 port map( D => n9436, CK => CLK, Q => 
                           n_1159, QN => n14341);
   REGISTERS_reg_16_1_inst : DFF_X1 port map( D => n9435, CK => CLK, Q => 
                           n_1160, QN => n14342);
   REGISTERS_reg_16_0_inst : DFF_X1 port map( D => n9434, CK => CLK, Q => 
                           n_1161, QN => n14343);
   REGISTERS_reg_17_31_inst : DFF_X1 port map( D => n9433, CK => CLK, Q => 
                           n_1162, QN => n14344);
   REGISTERS_reg_17_30_inst : DFF_X1 port map( D => n9432, CK => CLK, Q => 
                           n_1163, QN => n14345);
   REGISTERS_reg_17_29_inst : DFF_X1 port map( D => n9431, CK => CLK, Q => 
                           n_1164, QN => n14346);
   REGISTERS_reg_17_28_inst : DFF_X1 port map( D => n9430, CK => CLK, Q => 
                           n_1165, QN => n14347);
   REGISTERS_reg_17_27_inst : DFF_X1 port map( D => n9429, CK => CLK, Q => 
                           n_1166, QN => n14348);
   REGISTERS_reg_17_26_inst : DFF_X1 port map( D => n9428, CK => CLK, Q => 
                           n_1167, QN => n14349);
   REGISTERS_reg_17_25_inst : DFF_X1 port map( D => n9427, CK => CLK, Q => 
                           n_1168, QN => n14350);
   REGISTERS_reg_17_24_inst : DFF_X1 port map( D => n9426, CK => CLK, Q => 
                           n_1169, QN => n14351);
   REGISTERS_reg_17_23_inst : DFF_X1 port map( D => n9425, CK => CLK, Q => 
                           n_1170, QN => n14352);
   REGISTERS_reg_17_22_inst : DFF_X1 port map( D => n9424, CK => CLK, Q => 
                           n_1171, QN => n14353);
   REGISTERS_reg_17_21_inst : DFF_X1 port map( D => n9423, CK => CLK, Q => 
                           n_1172, QN => n14354);
   REGISTERS_reg_17_20_inst : DFF_X1 port map( D => n9422, CK => CLK, Q => 
                           n_1173, QN => n14355);
   REGISTERS_reg_17_19_inst : DFF_X1 port map( D => n9421, CK => CLK, Q => 
                           n_1174, QN => n14356);
   REGISTERS_reg_17_18_inst : DFF_X1 port map( D => n9420, CK => CLK, Q => 
                           n_1175, QN => n14357);
   REGISTERS_reg_17_17_inst : DFF_X1 port map( D => n9419, CK => CLK, Q => 
                           n_1176, QN => n14358);
   REGISTERS_reg_17_16_inst : DFF_X1 port map( D => n9418, CK => CLK, Q => 
                           n_1177, QN => n14359);
   REGISTERS_reg_17_15_inst : DFF_X1 port map( D => n9417, CK => CLK, Q => 
                           n_1178, QN => n14360);
   REGISTERS_reg_17_14_inst : DFF_X1 port map( D => n9416, CK => CLK, Q => 
                           n_1179, QN => n14361);
   REGISTERS_reg_17_13_inst : DFF_X1 port map( D => n9415, CK => CLK, Q => 
                           n_1180, QN => n14362);
   REGISTERS_reg_17_12_inst : DFF_X1 port map( D => n9414, CK => CLK, Q => 
                           n_1181, QN => n14363);
   REGISTERS_reg_17_11_inst : DFF_X1 port map( D => n9413, CK => CLK, Q => 
                           n_1182, QN => n14364);
   REGISTERS_reg_17_10_inst : DFF_X1 port map( D => n9412, CK => CLK, Q => 
                           n_1183, QN => n14365);
   REGISTERS_reg_17_9_inst : DFF_X1 port map( D => n9411, CK => CLK, Q => 
                           n_1184, QN => n14366);
   REGISTERS_reg_17_8_inst : DFF_X1 port map( D => n9410, CK => CLK, Q => 
                           n_1185, QN => n14367);
   REGISTERS_reg_17_7_inst : DFF_X1 port map( D => n9409, CK => CLK, Q => 
                           n_1186, QN => n14368);
   REGISTERS_reg_17_6_inst : DFF_X1 port map( D => n9408, CK => CLK, Q => 
                           n_1187, QN => n14369);
   REGISTERS_reg_17_5_inst : DFF_X1 port map( D => n9407, CK => CLK, Q => 
                           n_1188, QN => n14370);
   REGISTERS_reg_17_4_inst : DFF_X1 port map( D => n9406, CK => CLK, Q => 
                           n_1189, QN => n14371);
   REGISTERS_reg_17_3_inst : DFF_X1 port map( D => n9405, CK => CLK, Q => 
                           n_1190, QN => n14372);
   REGISTERS_reg_17_2_inst : DFF_X1 port map( D => n9404, CK => CLK, Q => 
                           n_1191, QN => n14373);
   REGISTERS_reg_17_1_inst : DFF_X1 port map( D => n9403, CK => CLK, Q => 
                           n_1192, QN => n14374);
   REGISTERS_reg_17_0_inst : DFF_X1 port map( D => n9402, CK => CLK, Q => 
                           n_1193, QN => n14375);
   REGISTERS_reg_18_31_inst : DFF_X1 port map( D => n9401, CK => CLK, Q => 
                           n_1194, QN => n14376);
   REGISTERS_reg_18_30_inst : DFF_X1 port map( D => n9400, CK => CLK, Q => 
                           n_1195, QN => n14377);
   REGISTERS_reg_18_29_inst : DFF_X1 port map( D => n9399, CK => CLK, Q => 
                           n_1196, QN => n14378);
   REGISTERS_reg_18_28_inst : DFF_X1 port map( D => n9398, CK => CLK, Q => 
                           n_1197, QN => n14379);
   REGISTERS_reg_18_27_inst : DFF_X1 port map( D => n9397, CK => CLK, Q => 
                           n_1198, QN => n14380);
   REGISTERS_reg_18_26_inst : DFF_X1 port map( D => n9396, CK => CLK, Q => 
                           n_1199, QN => n14381);
   REGISTERS_reg_18_25_inst : DFF_X1 port map( D => n9395, CK => CLK, Q => 
                           n_1200, QN => n14382);
   REGISTERS_reg_18_24_inst : DFF_X1 port map( D => n9394, CK => CLK, Q => 
                           n_1201, QN => n14383);
   REGISTERS_reg_18_23_inst : DFF_X1 port map( D => n9393, CK => CLK, Q => 
                           n_1202, QN => n14384);
   REGISTERS_reg_18_22_inst : DFF_X1 port map( D => n9392, CK => CLK, Q => 
                           n_1203, QN => n14385);
   REGISTERS_reg_18_21_inst : DFF_X1 port map( D => n9391, CK => CLK, Q => 
                           n_1204, QN => n14386);
   REGISTERS_reg_18_20_inst : DFF_X1 port map( D => n9390, CK => CLK, Q => 
                           n_1205, QN => n14387);
   REGISTERS_reg_18_19_inst : DFF_X1 port map( D => n9389, CK => CLK, Q => 
                           n_1206, QN => n14388);
   REGISTERS_reg_18_18_inst : DFF_X1 port map( D => n9388, CK => CLK, Q => 
                           n_1207, QN => n14389);
   REGISTERS_reg_18_17_inst : DFF_X1 port map( D => n9387, CK => CLK, Q => 
                           n_1208, QN => n14390);
   REGISTERS_reg_18_16_inst : DFF_X1 port map( D => n9386, CK => CLK, Q => 
                           n_1209, QN => n14391);
   REGISTERS_reg_18_15_inst : DFF_X1 port map( D => n9385, CK => CLK, Q => 
                           n_1210, QN => n14392);
   REGISTERS_reg_18_14_inst : DFF_X1 port map( D => n9384, CK => CLK, Q => 
                           n_1211, QN => n14393);
   REGISTERS_reg_18_13_inst : DFF_X1 port map( D => n9383, CK => CLK, Q => 
                           n_1212, QN => n14394);
   REGISTERS_reg_18_12_inst : DFF_X1 port map( D => n9382, CK => CLK, Q => 
                           n_1213, QN => n14395);
   REGISTERS_reg_18_11_inst : DFF_X1 port map( D => n9381, CK => CLK, Q => 
                           n_1214, QN => n14396);
   REGISTERS_reg_18_10_inst : DFF_X1 port map( D => n9380, CK => CLK, Q => 
                           n_1215, QN => n14397);
   REGISTERS_reg_18_9_inst : DFF_X1 port map( D => n9379, CK => CLK, Q => 
                           n_1216, QN => n14398);
   REGISTERS_reg_18_8_inst : DFF_X1 port map( D => n9378, CK => CLK, Q => 
                           n_1217, QN => n14399);
   REGISTERS_reg_18_7_inst : DFF_X1 port map( D => n9377, CK => CLK, Q => 
                           n_1218, QN => n14400);
   REGISTERS_reg_18_6_inst : DFF_X1 port map( D => n9376, CK => CLK, Q => 
                           n_1219, QN => n14401);
   REGISTERS_reg_18_5_inst : DFF_X1 port map( D => n9375, CK => CLK, Q => 
                           n_1220, QN => n14402);
   REGISTERS_reg_18_4_inst : DFF_X1 port map( D => n9374, CK => CLK, Q => 
                           n_1221, QN => n14403);
   REGISTERS_reg_18_3_inst : DFF_X1 port map( D => n9373, CK => CLK, Q => 
                           n_1222, QN => n14404);
   REGISTERS_reg_18_2_inst : DFF_X1 port map( D => n9372, CK => CLK, Q => 
                           n_1223, QN => n14405);
   REGISTERS_reg_18_1_inst : DFF_X1 port map( D => n9371, CK => CLK, Q => 
                           n_1224, QN => n14406);
   REGISTERS_reg_18_0_inst : DFF_X1 port map( D => n9370, CK => CLK, Q => 
                           n_1225, QN => n14407);
   REGISTERS_reg_19_31_inst : DFF_X1 port map( D => n9369, CK => CLK, Q => 
                           n_1226, QN => n14408);
   REGISTERS_reg_19_30_inst : DFF_X1 port map( D => n9368, CK => CLK, Q => 
                           n_1227, QN => n14409);
   REGISTERS_reg_19_29_inst : DFF_X1 port map( D => n9367, CK => CLK, Q => 
                           n_1228, QN => n14410);
   REGISTERS_reg_19_28_inst : DFF_X1 port map( D => n9366, CK => CLK, Q => 
                           n_1229, QN => n14411);
   REGISTERS_reg_19_27_inst : DFF_X1 port map( D => n9365, CK => CLK, Q => 
                           n_1230, QN => n14412);
   REGISTERS_reg_19_26_inst : DFF_X1 port map( D => n9364, CK => CLK, Q => 
                           n_1231, QN => n14413);
   REGISTERS_reg_19_25_inst : DFF_X1 port map( D => n9363, CK => CLK, Q => 
                           n_1232, QN => n14414);
   REGISTERS_reg_19_24_inst : DFF_X1 port map( D => n9362, CK => CLK, Q => 
                           n_1233, QN => n14415);
   REGISTERS_reg_19_23_inst : DFF_X1 port map( D => n9361, CK => CLK, Q => 
                           n_1234, QN => n14416);
   REGISTERS_reg_19_22_inst : DFF_X1 port map( D => n9360, CK => CLK, Q => 
                           n_1235, QN => n14417);
   REGISTERS_reg_19_21_inst : DFF_X1 port map( D => n9359, CK => CLK, Q => 
                           n_1236, QN => n14418);
   REGISTERS_reg_19_20_inst : DFF_X1 port map( D => n9358, CK => CLK, Q => 
                           n_1237, QN => n14419);
   REGISTERS_reg_19_19_inst : DFF_X1 port map( D => n9357, CK => CLK, Q => 
                           n_1238, QN => n14420);
   REGISTERS_reg_19_18_inst : DFF_X1 port map( D => n9356, CK => CLK, Q => 
                           n_1239, QN => n14421);
   REGISTERS_reg_19_17_inst : DFF_X1 port map( D => n9355, CK => CLK, Q => 
                           n_1240, QN => n14422);
   REGISTERS_reg_19_16_inst : DFF_X1 port map( D => n9354, CK => CLK, Q => 
                           n_1241, QN => n14423);
   REGISTERS_reg_19_15_inst : DFF_X1 port map( D => n9353, CK => CLK, Q => 
                           n_1242, QN => n14424);
   REGISTERS_reg_19_14_inst : DFF_X1 port map( D => n9352, CK => CLK, Q => 
                           n_1243, QN => n14425);
   REGISTERS_reg_19_13_inst : DFF_X1 port map( D => n9351, CK => CLK, Q => 
                           n_1244, QN => n14426);
   REGISTERS_reg_19_12_inst : DFF_X1 port map( D => n9350, CK => CLK, Q => 
                           n_1245, QN => n14427);
   REGISTERS_reg_19_11_inst : DFF_X1 port map( D => n9349, CK => CLK, Q => 
                           n_1246, QN => n14428);
   REGISTERS_reg_19_10_inst : DFF_X1 port map( D => n9348, CK => CLK, Q => 
                           n_1247, QN => n14429);
   REGISTERS_reg_19_9_inst : DFF_X1 port map( D => n9347, CK => CLK, Q => 
                           n_1248, QN => n14430);
   REGISTERS_reg_19_8_inst : DFF_X1 port map( D => n9346, CK => CLK, Q => 
                           n_1249, QN => n14431);
   REGISTERS_reg_19_7_inst : DFF_X1 port map( D => n9345, CK => CLK, Q => 
                           n_1250, QN => n14432);
   REGISTERS_reg_19_6_inst : DFF_X1 port map( D => n9344, CK => CLK, Q => 
                           n_1251, QN => n14433);
   REGISTERS_reg_19_5_inst : DFF_X1 port map( D => n9343, CK => CLK, Q => 
                           n_1252, QN => n14434);
   REGISTERS_reg_19_4_inst : DFF_X1 port map( D => n9342, CK => CLK, Q => 
                           n_1253, QN => n14435);
   REGISTERS_reg_19_3_inst : DFF_X1 port map( D => n9341, CK => CLK, Q => 
                           n_1254, QN => n14436);
   REGISTERS_reg_19_2_inst : DFF_X1 port map( D => n9340, CK => CLK, Q => 
                           n_1255, QN => n14437);
   REGISTERS_reg_19_1_inst : DFF_X1 port map( D => n9339, CK => CLK, Q => 
                           n_1256, QN => n14438);
   REGISTERS_reg_19_0_inst : DFF_X1 port map( D => n9338, CK => CLK, Q => 
                           n_1257, QN => n14439);
   REGISTERS_reg_21_31_inst : DFF_X1 port map( D => n9305, CK => CLK, Q => n97,
                           QN => n14459);
   REGISTERS_reg_21_30_inst : DFF_X1 port map( D => n9304, CK => CLK, Q => n99,
                           QN => n14460);
   REGISTERS_reg_24_31_inst : DFF_X1 port map( D => n9209, CK => CLK, Q => 
                           n_1258, QN => n14493);
   REGISTERS_reg_24_30_inst : DFF_X1 port map( D => n9208, CK => CLK, Q => 
                           n_1259, QN => n14494);
   REGISTERS_reg_24_29_inst : DFF_X1 port map( D => n9207, CK => CLK, Q => 
                           n_1260, QN => n14495);
   REGISTERS_reg_24_28_inst : DFF_X1 port map( D => n9206, CK => CLK, Q => 
                           n_1261, QN => n14496);
   REGISTERS_reg_24_27_inst : DFF_X1 port map( D => n9205, CK => CLK, Q => 
                           n_1262, QN => n14497);
   REGISTERS_reg_24_26_inst : DFF_X1 port map( D => n9204, CK => CLK, Q => 
                           n_1263, QN => n14498);
   REGISTERS_reg_24_25_inst : DFF_X1 port map( D => n9203, CK => CLK, Q => 
                           n_1264, QN => n14499);
   REGISTERS_reg_24_24_inst : DFF_X1 port map( D => n9202, CK => CLK, Q => 
                           n_1265, QN => n14500);
   REGISTERS_reg_24_23_inst : DFF_X1 port map( D => n9201, CK => CLK, Q => 
                           n_1266, QN => n14501);
   REGISTERS_reg_24_22_inst : DFF_X1 port map( D => n9200, CK => CLK, Q => 
                           n_1267, QN => n14502);
   REGISTERS_reg_24_21_inst : DFF_X1 port map( D => n9199, CK => CLK, Q => 
                           n_1268, QN => n14503);
   REGISTERS_reg_24_20_inst : DFF_X1 port map( D => n9198, CK => CLK, Q => 
                           n_1269, QN => n14504);
   REGISTERS_reg_24_19_inst : DFF_X1 port map( D => n9197, CK => CLK, Q => 
                           n_1270, QN => n14505);
   REGISTERS_reg_24_18_inst : DFF_X1 port map( D => n9196, CK => CLK, Q => 
                           n_1271, QN => n14506);
   REGISTERS_reg_24_17_inst : DFF_X1 port map( D => n9195, CK => CLK, Q => 
                           n_1272, QN => n14507);
   REGISTERS_reg_24_16_inst : DFF_X1 port map( D => n9194, CK => CLK, Q => 
                           n_1273, QN => n14508);
   REGISTERS_reg_24_15_inst : DFF_X1 port map( D => n9193, CK => CLK, Q => 
                           n_1274, QN => n14509);
   REGISTERS_reg_24_14_inst : DFF_X1 port map( D => n9192, CK => CLK, Q => 
                           n_1275, QN => n14510);
   REGISTERS_reg_24_13_inst : DFF_X1 port map( D => n9191, CK => CLK, Q => 
                           n_1276, QN => n14511);
   REGISTERS_reg_24_12_inst : DFF_X1 port map( D => n9190, CK => CLK, Q => 
                           n_1277, QN => n14512);
   REGISTERS_reg_24_11_inst : DFF_X1 port map( D => n9189, CK => CLK, Q => 
                           n_1278, QN => n14513);
   REGISTERS_reg_24_10_inst : DFF_X1 port map( D => n9188, CK => CLK, Q => 
                           n_1279, QN => n14514);
   REGISTERS_reg_24_9_inst : DFF_X1 port map( D => n9187, CK => CLK, Q => 
                           n_1280, QN => n14515);
   REGISTERS_reg_24_8_inst : DFF_X1 port map( D => n9186, CK => CLK, Q => 
                           n_1281, QN => n14516);
   REGISTERS_reg_24_7_inst : DFF_X1 port map( D => n9185, CK => CLK, Q => 
                           n_1282, QN => n14517);
   REGISTERS_reg_24_6_inst : DFF_X1 port map( D => n9184, CK => CLK, Q => 
                           n_1283, QN => n14518);
   REGISTERS_reg_24_5_inst : DFF_X1 port map( D => n9183, CK => CLK, Q => 
                           n_1284, QN => n14519);
   REGISTERS_reg_24_4_inst : DFF_X1 port map( D => n9182, CK => CLK, Q => 
                           n_1285, QN => n14520);
   REGISTERS_reg_24_3_inst : DFF_X1 port map( D => n9181, CK => CLK, Q => 
                           n_1286, QN => n14521);
   REGISTERS_reg_24_2_inst : DFF_X1 port map( D => n9180, CK => CLK, Q => 
                           n_1287, QN => n14522);
   REGISTERS_reg_24_1_inst : DFF_X1 port map( D => n9179, CK => CLK, Q => 
                           n_1288, QN => n14523);
   REGISTERS_reg_24_0_inst : DFF_X1 port map( D => n9178, CK => CLK, Q => 
                           n_1289, QN => n14524);
   REGISTERS_reg_25_31_inst : DFF_X1 port map( D => n9177, CK => CLK, Q => 
                           n_1290, QN => n14525);
   REGISTERS_reg_25_30_inst : DFF_X1 port map( D => n9176, CK => CLK, Q => 
                           n_1291, QN => n14526);
   REGISTERS_reg_25_29_inst : DFF_X1 port map( D => n9175, CK => CLK, Q => 
                           n_1292, QN => n14527);
   REGISTERS_reg_25_28_inst : DFF_X1 port map( D => n9174, CK => CLK, Q => 
                           n_1293, QN => n14528);
   REGISTERS_reg_25_27_inst : DFF_X1 port map( D => n9173, CK => CLK, Q => 
                           n_1294, QN => n14529);
   REGISTERS_reg_25_26_inst : DFF_X1 port map( D => n9172, CK => CLK, Q => 
                           n_1295, QN => n14530);
   REGISTERS_reg_25_25_inst : DFF_X1 port map( D => n9171, CK => CLK, Q => 
                           n_1296, QN => n14531);
   REGISTERS_reg_25_24_inst : DFF_X1 port map( D => n9170, CK => CLK, Q => 
                           n_1297, QN => n14532);
   REGISTERS_reg_25_23_inst : DFF_X1 port map( D => n9169, CK => CLK, Q => 
                           n_1298, QN => n14533);
   REGISTERS_reg_25_22_inst : DFF_X1 port map( D => n9168, CK => CLK, Q => 
                           n_1299, QN => n14534);
   REGISTERS_reg_25_21_inst : DFF_X1 port map( D => n9167, CK => CLK, Q => 
                           n_1300, QN => n14535);
   REGISTERS_reg_25_20_inst : DFF_X1 port map( D => n9166, CK => CLK, Q => 
                           n_1301, QN => n14536);
   REGISTERS_reg_25_19_inst : DFF_X1 port map( D => n9165, CK => CLK, Q => 
                           n_1302, QN => n14537);
   REGISTERS_reg_25_18_inst : DFF_X1 port map( D => n9164, CK => CLK, Q => 
                           n_1303, QN => n14538);
   REGISTERS_reg_25_17_inst : DFF_X1 port map( D => n9163, CK => CLK, Q => 
                           n_1304, QN => n14539);
   REGISTERS_reg_25_16_inst : DFF_X1 port map( D => n9162, CK => CLK, Q => 
                           n_1305, QN => n14540);
   REGISTERS_reg_25_15_inst : DFF_X1 port map( D => n9161, CK => CLK, Q => 
                           n_1306, QN => n14541);
   REGISTERS_reg_25_14_inst : DFF_X1 port map( D => n9160, CK => CLK, Q => 
                           n_1307, QN => n14542);
   REGISTERS_reg_25_13_inst : DFF_X1 port map( D => n9159, CK => CLK, Q => 
                           n_1308, QN => n14543);
   REGISTERS_reg_25_12_inst : DFF_X1 port map( D => n9158, CK => CLK, Q => 
                           n_1309, QN => n14544);
   REGISTERS_reg_25_11_inst : DFF_X1 port map( D => n9157, CK => CLK, Q => 
                           n_1310, QN => n14545);
   REGISTERS_reg_25_10_inst : DFF_X1 port map( D => n9156, CK => CLK, Q => 
                           n_1311, QN => n14546);
   REGISTERS_reg_25_9_inst : DFF_X1 port map( D => n9155, CK => CLK, Q => 
                           n_1312, QN => n14547);
   REGISTERS_reg_25_8_inst : DFF_X1 port map( D => n9154, CK => CLK, Q => 
                           n_1313, QN => n14548);
   REGISTERS_reg_25_7_inst : DFF_X1 port map( D => n9153, CK => CLK, Q => 
                           n_1314, QN => n14549);
   REGISTERS_reg_25_6_inst : DFF_X1 port map( D => n9152, CK => CLK, Q => 
                           n_1315, QN => n14550);
   REGISTERS_reg_25_5_inst : DFF_X1 port map( D => n9151, CK => CLK, Q => 
                           n_1316, QN => n14551);
   REGISTERS_reg_25_4_inst : DFF_X1 port map( D => n9150, CK => CLK, Q => 
                           n_1317, QN => n14552);
   REGISTERS_reg_25_3_inst : DFF_X1 port map( D => n9149, CK => CLK, Q => 
                           n_1318, QN => n14553);
   REGISTERS_reg_25_2_inst : DFF_X1 port map( D => n9148, CK => CLK, Q => 
                           n_1319, QN => n14554);
   REGISTERS_reg_25_1_inst : DFF_X1 port map( D => n9147, CK => CLK, Q => 
                           n_1320, QN => n14555);
   REGISTERS_reg_25_0_inst : DFF_X1 port map( D => n9146, CK => CLK, Q => 
                           n_1321, QN => n14556);
   REGISTERS_reg_26_31_inst : DFF_X1 port map( D => n9145, CK => CLK, Q => 
                           n_1322, QN => n14557);
   REGISTERS_reg_26_30_inst : DFF_X1 port map( D => n9144, CK => CLK, Q => 
                           n_1323, QN => n14558);
   REGISTERS_reg_26_29_inst : DFF_X1 port map( D => n9143, CK => CLK, Q => 
                           n_1324, QN => n14559);
   REGISTERS_reg_26_28_inst : DFF_X1 port map( D => n9142, CK => CLK, Q => 
                           n_1325, QN => n14560);
   REGISTERS_reg_26_27_inst : DFF_X1 port map( D => n9141, CK => CLK, Q => 
                           n_1326, QN => n14561);
   REGISTERS_reg_26_26_inst : DFF_X1 port map( D => n9140, CK => CLK, Q => 
                           n_1327, QN => n14562);
   REGISTERS_reg_26_25_inst : DFF_X1 port map( D => n9139, CK => CLK, Q => 
                           n_1328, QN => n14563);
   REGISTERS_reg_26_24_inst : DFF_X1 port map( D => n9138, CK => CLK, Q => 
                           n_1329, QN => n14564);
   REGISTERS_reg_26_23_inst : DFF_X1 port map( D => n9137, CK => CLK, Q => 
                           n_1330, QN => n14565);
   REGISTERS_reg_26_22_inst : DFF_X1 port map( D => n9136, CK => CLK, Q => 
                           n_1331, QN => n14566);
   REGISTERS_reg_26_21_inst : DFF_X1 port map( D => n9135, CK => CLK, Q => 
                           n_1332, QN => n14567);
   REGISTERS_reg_26_20_inst : DFF_X1 port map( D => n9134, CK => CLK, Q => 
                           n_1333, QN => n14568);
   REGISTERS_reg_26_19_inst : DFF_X1 port map( D => n9133, CK => CLK, Q => 
                           n_1334, QN => n14569);
   REGISTERS_reg_26_18_inst : DFF_X1 port map( D => n9132, CK => CLK, Q => 
                           n_1335, QN => n14570);
   REGISTERS_reg_26_17_inst : DFF_X1 port map( D => n9131, CK => CLK, Q => 
                           n_1336, QN => n14571);
   REGISTERS_reg_26_16_inst : DFF_X1 port map( D => n9130, CK => CLK, Q => 
                           n_1337, QN => n14572);
   REGISTERS_reg_26_15_inst : DFF_X1 port map( D => n9129, CK => CLK, Q => 
                           n_1338, QN => n14573);
   REGISTERS_reg_26_14_inst : DFF_X1 port map( D => n9128, CK => CLK, Q => 
                           n_1339, QN => n14574);
   REGISTERS_reg_26_13_inst : DFF_X1 port map( D => n9127, CK => CLK, Q => 
                           n_1340, QN => n14575);
   REGISTERS_reg_26_12_inst : DFF_X1 port map( D => n9126, CK => CLK, Q => 
                           n_1341, QN => n14576);
   REGISTERS_reg_26_11_inst : DFF_X1 port map( D => n9125, CK => CLK, Q => 
                           n_1342, QN => n14577);
   REGISTERS_reg_26_10_inst : DFF_X1 port map( D => n9124, CK => CLK, Q => 
                           n_1343, QN => n14578);
   REGISTERS_reg_26_9_inst : DFF_X1 port map( D => n9123, CK => CLK, Q => 
                           n_1344, QN => n14579);
   REGISTERS_reg_26_8_inst : DFF_X1 port map( D => n9122, CK => CLK, Q => 
                           n_1345, QN => n14580);
   REGISTERS_reg_26_7_inst : DFF_X1 port map( D => n9121, CK => CLK, Q => 
                           n_1346, QN => n14581);
   REGISTERS_reg_26_6_inst : DFF_X1 port map( D => n9120, CK => CLK, Q => 
                           n_1347, QN => n14582);
   REGISTERS_reg_26_5_inst : DFF_X1 port map( D => n9119, CK => CLK, Q => 
                           n_1348, QN => n14583);
   REGISTERS_reg_26_4_inst : DFF_X1 port map( D => n9118, CK => CLK, Q => 
                           n_1349, QN => n14584);
   REGISTERS_reg_26_3_inst : DFF_X1 port map( D => n9117, CK => CLK, Q => 
                           n_1350, QN => n14585);
   REGISTERS_reg_26_2_inst : DFF_X1 port map( D => n9116, CK => CLK, Q => 
                           n_1351, QN => n14586);
   REGISTERS_reg_26_1_inst : DFF_X1 port map( D => n9115, CK => CLK, Q => 
                           n_1352, QN => n14587);
   REGISTERS_reg_26_0_inst : DFF_X1 port map( D => n9114, CK => CLK, Q => 
                           n_1353, QN => n14588);
   REGISTERS_reg_27_31_inst : DFF_X1 port map( D => n9113, CK => CLK, Q => 
                           n_1354, QN => n14589);
   REGISTERS_reg_27_30_inst : DFF_X1 port map( D => n9112, CK => CLK, Q => 
                           n_1355, QN => n14590);
   REGISTERS_reg_27_29_inst : DFF_X1 port map( D => n9111, CK => CLK, Q => 
                           n_1356, QN => n14591);
   REGISTERS_reg_27_28_inst : DFF_X1 port map( D => n9110, CK => CLK, Q => 
                           n_1357, QN => n14592);
   REGISTERS_reg_27_27_inst : DFF_X1 port map( D => n9109, CK => CLK, Q => 
                           n_1358, QN => n14593);
   REGISTERS_reg_27_26_inst : DFF_X1 port map( D => n9108, CK => CLK, Q => 
                           n_1359, QN => n14594);
   REGISTERS_reg_27_25_inst : DFF_X1 port map( D => n9107, CK => CLK, Q => 
                           n_1360, QN => n14595);
   REGISTERS_reg_27_24_inst : DFF_X1 port map( D => n9106, CK => CLK, Q => 
                           n_1361, QN => n14596);
   REGISTERS_reg_27_23_inst : DFF_X1 port map( D => n9105, CK => CLK, Q => 
                           n_1362, QN => n14597);
   REGISTERS_reg_27_22_inst : DFF_X1 port map( D => n9104, CK => CLK, Q => 
                           n_1363, QN => n14598);
   REGISTERS_reg_27_21_inst : DFF_X1 port map( D => n9103, CK => CLK, Q => 
                           n_1364, QN => n14599);
   REGISTERS_reg_27_20_inst : DFF_X1 port map( D => n9102, CK => CLK, Q => 
                           n_1365, QN => n14600);
   REGISTERS_reg_27_19_inst : DFF_X1 port map( D => n9101, CK => CLK, Q => 
                           n_1366, QN => n14601);
   REGISTERS_reg_27_18_inst : DFF_X1 port map( D => n9100, CK => CLK, Q => 
                           n_1367, QN => n14602);
   REGISTERS_reg_27_17_inst : DFF_X1 port map( D => n9099, CK => CLK, Q => 
                           n_1368, QN => n14603);
   REGISTERS_reg_27_16_inst : DFF_X1 port map( D => n9098, CK => CLK, Q => 
                           n_1369, QN => n14604);
   REGISTERS_reg_27_15_inst : DFF_X1 port map( D => n9097, CK => CLK, Q => 
                           n_1370, QN => n14605);
   REGISTERS_reg_27_14_inst : DFF_X1 port map( D => n9096, CK => CLK, Q => 
                           n_1371, QN => n14606);
   REGISTERS_reg_27_13_inst : DFF_X1 port map( D => n9095, CK => CLK, Q => 
                           n_1372, QN => n14607);
   REGISTERS_reg_27_12_inst : DFF_X1 port map( D => n9094, CK => CLK, Q => 
                           n_1373, QN => n14608);
   REGISTERS_reg_27_11_inst : DFF_X1 port map( D => n9093, CK => CLK, Q => 
                           n_1374, QN => n14609);
   REGISTERS_reg_27_10_inst : DFF_X1 port map( D => n9092, CK => CLK, Q => 
                           n_1375, QN => n14610);
   REGISTERS_reg_27_9_inst : DFF_X1 port map( D => n9091, CK => CLK, Q => 
                           n_1376, QN => n14611);
   REGISTERS_reg_27_8_inst : DFF_X1 port map( D => n9090, CK => CLK, Q => 
                           n_1377, QN => n14612);
   REGISTERS_reg_27_7_inst : DFF_X1 port map( D => n9089, CK => CLK, Q => 
                           n_1378, QN => n14613);
   REGISTERS_reg_27_6_inst : DFF_X1 port map( D => n9088, CK => CLK, Q => 
                           n_1379, QN => n14614);
   REGISTERS_reg_27_5_inst : DFF_X1 port map( D => n9087, CK => CLK, Q => 
                           n_1380, QN => n14615);
   REGISTERS_reg_27_4_inst : DFF_X1 port map( D => n9086, CK => CLK, Q => 
                           n_1381, QN => n14616);
   REGISTERS_reg_27_3_inst : DFF_X1 port map( D => n9085, CK => CLK, Q => 
                           n_1382, QN => n14617);
   REGISTERS_reg_27_2_inst : DFF_X1 port map( D => n9084, CK => CLK, Q => 
                           n_1383, QN => n14618);
   REGISTERS_reg_27_1_inst : DFF_X1 port map( D => n9083, CK => CLK, Q => 
                           n_1384, QN => n14619);
   REGISTERS_reg_27_0_inst : DFF_X1 port map( D => n9082, CK => CLK, Q => 
                           n_1385, QN => n14620);
   REGISTERS_reg_28_31_inst : DFF_X1 port map( D => n9081, CK => CLK, Q => 
                           n_1386, QN => n14621);
   REGISTERS_reg_28_30_inst : DFF_X1 port map( D => n9080, CK => CLK, Q => 
                           n_1387, QN => n14622);
   REGISTERS_reg_28_29_inst : DFF_X1 port map( D => n9079, CK => CLK, Q => 
                           n_1388, QN => n14623);
   REGISTERS_reg_28_28_inst : DFF_X1 port map( D => n9078, CK => CLK, Q => 
                           n_1389, QN => n14624);
   REGISTERS_reg_28_27_inst : DFF_X1 port map( D => n9077, CK => CLK, Q => 
                           n_1390, QN => n14625);
   REGISTERS_reg_28_26_inst : DFF_X1 port map( D => n9076, CK => CLK, Q => 
                           n_1391, QN => n14626);
   REGISTERS_reg_28_25_inst : DFF_X1 port map( D => n9075, CK => CLK, Q => 
                           n_1392, QN => n14627);
   REGISTERS_reg_28_24_inst : DFF_X1 port map( D => n9074, CK => CLK, Q => 
                           n_1393, QN => n14628);
   REGISTERS_reg_28_23_inst : DFF_X1 port map( D => n9073, CK => CLK, Q => 
                           n_1394, QN => n14629);
   REGISTERS_reg_28_22_inst : DFF_X1 port map( D => n9072, CK => CLK, Q => 
                           n_1395, QN => n14630);
   REGISTERS_reg_28_21_inst : DFF_X1 port map( D => n9071, CK => CLK, Q => 
                           n_1396, QN => n14631);
   REGISTERS_reg_28_20_inst : DFF_X1 port map( D => n9070, CK => CLK, Q => 
                           n_1397, QN => n14632);
   REGISTERS_reg_28_19_inst : DFF_X1 port map( D => n9069, CK => CLK, Q => 
                           n_1398, QN => n14633);
   REGISTERS_reg_28_18_inst : DFF_X1 port map( D => n9068, CK => CLK, Q => 
                           n_1399, QN => n14634);
   REGISTERS_reg_28_17_inst : DFF_X1 port map( D => n9067, CK => CLK, Q => 
                           n_1400, QN => n14635);
   REGISTERS_reg_28_16_inst : DFF_X1 port map( D => n9066, CK => CLK, Q => 
                           n_1401, QN => n14636);
   REGISTERS_reg_28_15_inst : DFF_X1 port map( D => n9065, CK => CLK, Q => 
                           n_1402, QN => n14637);
   REGISTERS_reg_28_14_inst : DFF_X1 port map( D => n9064, CK => CLK, Q => 
                           n_1403, QN => n14638);
   REGISTERS_reg_28_13_inst : DFF_X1 port map( D => n9063, CK => CLK, Q => 
                           n_1404, QN => n14639);
   REGISTERS_reg_28_12_inst : DFF_X1 port map( D => n9062, CK => CLK, Q => 
                           n_1405, QN => n14640);
   REGISTERS_reg_28_11_inst : DFF_X1 port map( D => n9061, CK => CLK, Q => 
                           n_1406, QN => n14641);
   REGISTERS_reg_28_10_inst : DFF_X1 port map( D => n9060, CK => CLK, Q => 
                           n_1407, QN => n14642);
   REGISTERS_reg_28_9_inst : DFF_X1 port map( D => n9059, CK => CLK, Q => 
                           n_1408, QN => n14643);
   REGISTERS_reg_28_8_inst : DFF_X1 port map( D => n9058, CK => CLK, Q => 
                           n_1409, QN => n14644);
   REGISTERS_reg_28_7_inst : DFF_X1 port map( D => n9057, CK => CLK, Q => 
                           n_1410, QN => n14645);
   REGISTERS_reg_28_6_inst : DFF_X1 port map( D => n9056, CK => CLK, Q => 
                           n_1411, QN => n14646);
   REGISTERS_reg_28_5_inst : DFF_X1 port map( D => n9055, CK => CLK, Q => 
                           n_1412, QN => n14647);
   REGISTERS_reg_28_4_inst : DFF_X1 port map( D => n9054, CK => CLK, Q => 
                           n_1413, QN => n14648);
   REGISTERS_reg_28_3_inst : DFF_X1 port map( D => n9053, CK => CLK, Q => 
                           n_1414, QN => n14649);
   REGISTERS_reg_28_2_inst : DFF_X1 port map( D => n9052, CK => CLK, Q => 
                           n_1415, QN => n14650);
   REGISTERS_reg_28_1_inst : DFF_X1 port map( D => n9051, CK => CLK, Q => 
                           n_1416, QN => n14651);
   REGISTERS_reg_28_0_inst : DFF_X1 port map( D => n9050, CK => CLK, Q => 
                           n_1417, QN => n14652);
   REGISTERS_reg_33_31_inst : DFF_X1 port map( D => n8921, CK => CLK, Q => 
                           n_1418, QN => n14692);
   REGISTERS_reg_33_30_inst : DFF_X1 port map( D => n8920, CK => CLK, Q => 
                           n_1419, QN => n14693);
   REGISTERS_reg_33_29_inst : DFF_X1 port map( D => n8919, CK => CLK, Q => 
                           n_1420, QN => n14694);
   REGISTERS_reg_33_28_inst : DFF_X1 port map( D => n8918, CK => CLK, Q => 
                           n_1421, QN => n14695);
   REGISTERS_reg_33_27_inst : DFF_X1 port map( D => n8917, CK => CLK, Q => 
                           n_1422, QN => n14696);
   REGISTERS_reg_33_26_inst : DFF_X1 port map( D => n8916, CK => CLK, Q => 
                           n_1423, QN => n14697);
   REGISTERS_reg_33_25_inst : DFF_X1 port map( D => n8915, CK => CLK, Q => 
                           n_1424, QN => n14698);
   REGISTERS_reg_33_24_inst : DFF_X1 port map( D => n8914, CK => CLK, Q => 
                           n_1425, QN => n14699);
   REGISTERS_reg_33_23_inst : DFF_X1 port map( D => n8913, CK => CLK, Q => 
                           n_1426, QN => n14700);
   REGISTERS_reg_33_22_inst : DFF_X1 port map( D => n8912, CK => CLK, Q => 
                           n_1427, QN => n14701);
   REGISTERS_reg_33_21_inst : DFF_X1 port map( D => n8911, CK => CLK, Q => 
                           n_1428, QN => n14702);
   REGISTERS_reg_33_20_inst : DFF_X1 port map( D => n8910, CK => CLK, Q => 
                           n_1429, QN => n14703);
   REGISTERS_reg_33_19_inst : DFF_X1 port map( D => n8909, CK => CLK, Q => 
                           n_1430, QN => n14704);
   REGISTERS_reg_33_18_inst : DFF_X1 port map( D => n8908, CK => CLK, Q => 
                           n_1431, QN => n14705);
   REGISTERS_reg_33_17_inst : DFF_X1 port map( D => n8907, CK => CLK, Q => 
                           n_1432, QN => n14706);
   REGISTERS_reg_33_16_inst : DFF_X1 port map( D => n8906, CK => CLK, Q => 
                           n_1433, QN => n14707);
   REGISTERS_reg_33_15_inst : DFF_X1 port map( D => n8905, CK => CLK, Q => 
                           n_1434, QN => n14708);
   REGISTERS_reg_33_14_inst : DFF_X1 port map( D => n8904, CK => CLK, Q => 
                           n_1435, QN => n14709);
   REGISTERS_reg_33_13_inst : DFF_X1 port map( D => n8903, CK => CLK, Q => 
                           n_1436, QN => n14710);
   REGISTERS_reg_33_12_inst : DFF_X1 port map( D => n8902, CK => CLK, Q => 
                           n_1437, QN => n14711);
   REGISTERS_reg_33_11_inst : DFF_X1 port map( D => n8901, CK => CLK, Q => 
                           n_1438, QN => n14712);
   REGISTERS_reg_33_10_inst : DFF_X1 port map( D => n8900, CK => CLK, Q => 
                           n_1439, QN => n14713);
   REGISTERS_reg_33_9_inst : DFF_X1 port map( D => n8899, CK => CLK, Q => 
                           n_1440, QN => n14714);
   REGISTERS_reg_33_8_inst : DFF_X1 port map( D => n8898, CK => CLK, Q => 
                           n_1441, QN => n14715);
   REGISTERS_reg_33_7_inst : DFF_X1 port map( D => n8897, CK => CLK, Q => 
                           n_1442, QN => n14716);
   REGISTERS_reg_33_6_inst : DFF_X1 port map( D => n8896, CK => CLK, Q => 
                           n_1443, QN => n14717);
   REGISTERS_reg_33_5_inst : DFF_X1 port map( D => n8895, CK => CLK, Q => 
                           n_1444, QN => n14718);
   REGISTERS_reg_33_4_inst : DFF_X1 port map( D => n8894, CK => CLK, Q => 
                           n_1445, QN => n14719);
   REGISTERS_reg_33_3_inst : DFF_X1 port map( D => n8893, CK => CLK, Q => 
                           n_1446, QN => n14720);
   REGISTERS_reg_33_2_inst : DFF_X1 port map( D => n8892, CK => CLK, Q => 
                           n_1447, QN => n14721);
   REGISTERS_reg_33_1_inst : DFF_X1 port map( D => n8891, CK => CLK, Q => 
                           n_1448, QN => n14722);
   REGISTERS_reg_33_0_inst : DFF_X1 port map( D => n8890, CK => CLK, Q => 
                           n_1449, QN => n14723);
   REGISTERS_reg_34_31_inst : DFF_X1 port map( D => n8889, CK => CLK, Q => 
                           n_1450, QN => n14724);
   REGISTERS_reg_34_30_inst : DFF_X1 port map( D => n8888, CK => CLK, Q => 
                           n_1451, QN => n14725);
   REGISTERS_reg_34_29_inst : DFF_X1 port map( D => n8887, CK => CLK, Q => 
                           n_1452, QN => n14726);
   REGISTERS_reg_34_28_inst : DFF_X1 port map( D => n8886, CK => CLK, Q => 
                           n_1453, QN => n14727);
   REGISTERS_reg_34_27_inst : DFF_X1 port map( D => n8885, CK => CLK, Q => 
                           n_1454, QN => n14728);
   REGISTERS_reg_34_26_inst : DFF_X1 port map( D => n8884, CK => CLK, Q => 
                           n_1455, QN => n14729);
   REGISTERS_reg_34_25_inst : DFF_X1 port map( D => n8883, CK => CLK, Q => 
                           n_1456, QN => n14730);
   REGISTERS_reg_34_24_inst : DFF_X1 port map( D => n8882, CK => CLK, Q => 
                           n_1457, QN => n14731);
   REGISTERS_reg_34_23_inst : DFF_X1 port map( D => n8881, CK => CLK, Q => 
                           n_1458, QN => n14732);
   REGISTERS_reg_34_22_inst : DFF_X1 port map( D => n8880, CK => CLK, Q => 
                           n_1459, QN => n14733);
   REGISTERS_reg_34_21_inst : DFF_X1 port map( D => n8879, CK => CLK, Q => 
                           n_1460, QN => n14734);
   REGISTERS_reg_34_20_inst : DFF_X1 port map( D => n8878, CK => CLK, Q => 
                           n_1461, QN => n14735);
   REGISTERS_reg_34_19_inst : DFF_X1 port map( D => n8877, CK => CLK, Q => 
                           n_1462, QN => n14736);
   REGISTERS_reg_34_18_inst : DFF_X1 port map( D => n8876, CK => CLK, Q => 
                           n_1463, QN => n14737);
   REGISTERS_reg_34_17_inst : DFF_X1 port map( D => n8875, CK => CLK, Q => 
                           n_1464, QN => n14738);
   REGISTERS_reg_34_16_inst : DFF_X1 port map( D => n8874, CK => CLK, Q => 
                           n_1465, QN => n14739);
   REGISTERS_reg_34_15_inst : DFF_X1 port map( D => n8873, CK => CLK, Q => 
                           n_1466, QN => n14740);
   REGISTERS_reg_34_14_inst : DFF_X1 port map( D => n8872, CK => CLK, Q => 
                           n_1467, QN => n14741);
   REGISTERS_reg_34_13_inst : DFF_X1 port map( D => n8871, CK => CLK, Q => 
                           n_1468, QN => n14742);
   REGISTERS_reg_34_12_inst : DFF_X1 port map( D => n8870, CK => CLK, Q => 
                           n_1469, QN => n14743);
   REGISTERS_reg_34_11_inst : DFF_X1 port map( D => n8869, CK => CLK, Q => 
                           n_1470, QN => n14744);
   REGISTERS_reg_34_10_inst : DFF_X1 port map( D => n8868, CK => CLK, Q => 
                           n_1471, QN => n14745);
   REGISTERS_reg_34_9_inst : DFF_X1 port map( D => n8867, CK => CLK, Q => 
                           n_1472, QN => n14746);
   REGISTERS_reg_34_8_inst : DFF_X1 port map( D => n8866, CK => CLK, Q => 
                           n_1473, QN => n14747);
   REGISTERS_reg_34_7_inst : DFF_X1 port map( D => n8865, CK => CLK, Q => 
                           n_1474, QN => n14748);
   REGISTERS_reg_34_6_inst : DFF_X1 port map( D => n8864, CK => CLK, Q => 
                           n_1475, QN => n14749);
   REGISTERS_reg_34_5_inst : DFF_X1 port map( D => n8863, CK => CLK, Q => 
                           n_1476, QN => n14750);
   REGISTERS_reg_34_4_inst : DFF_X1 port map( D => n8862, CK => CLK, Q => 
                           n_1477, QN => n14751);
   REGISTERS_reg_34_3_inst : DFF_X1 port map( D => n8861, CK => CLK, Q => 
                           n_1478, QN => n14752);
   REGISTERS_reg_34_2_inst : DFF_X1 port map( D => n8860, CK => CLK, Q => 
                           n_1479, QN => n14753);
   REGISTERS_reg_34_1_inst : DFF_X1 port map( D => n8859, CK => CLK, Q => 
                           n_1480, QN => n14754);
   REGISTERS_reg_34_0_inst : DFF_X1 port map( D => n8858, CK => CLK, Q => 
                           n_1481, QN => n14755);
   REGISTERS_reg_35_31_inst : DFF_X1 port map( D => n8857, CK => CLK, Q => 
                           n_1482, QN => n14756);
   REGISTERS_reg_35_30_inst : DFF_X1 port map( D => n8856, CK => CLK, Q => 
                           n_1483, QN => n14757);
   REGISTERS_reg_35_29_inst : DFF_X1 port map( D => n8855, CK => CLK, Q => 
                           n_1484, QN => n14758);
   REGISTERS_reg_35_28_inst : DFF_X1 port map( D => n8854, CK => CLK, Q => 
                           n_1485, QN => n14759);
   REGISTERS_reg_35_27_inst : DFF_X1 port map( D => n8853, CK => CLK, Q => 
                           n_1486, QN => n14760);
   REGISTERS_reg_35_26_inst : DFF_X1 port map( D => n8852, CK => CLK, Q => 
                           n_1487, QN => n14761);
   REGISTERS_reg_35_25_inst : DFF_X1 port map( D => n8851, CK => CLK, Q => 
                           n_1488, QN => n14762);
   REGISTERS_reg_35_24_inst : DFF_X1 port map( D => n8850, CK => CLK, Q => 
                           n_1489, QN => n14763);
   REGISTERS_reg_35_23_inst : DFF_X1 port map( D => n8849, CK => CLK, Q => 
                           n_1490, QN => n14764);
   REGISTERS_reg_35_22_inst : DFF_X1 port map( D => n8848, CK => CLK, Q => 
                           n_1491, QN => n14765);
   REGISTERS_reg_35_21_inst : DFF_X1 port map( D => n8847, CK => CLK, Q => 
                           n_1492, QN => n14766);
   REGISTERS_reg_35_20_inst : DFF_X1 port map( D => n8846, CK => CLK, Q => 
                           n_1493, QN => n14767);
   REGISTERS_reg_35_19_inst : DFF_X1 port map( D => n8845, CK => CLK, Q => 
                           n_1494, QN => n14768);
   REGISTERS_reg_35_18_inst : DFF_X1 port map( D => n8844, CK => CLK, Q => 
                           n_1495, QN => n14769);
   REGISTERS_reg_35_17_inst : DFF_X1 port map( D => n8843, CK => CLK, Q => 
                           n_1496, QN => n14770);
   REGISTERS_reg_35_16_inst : DFF_X1 port map( D => n8842, CK => CLK, Q => 
                           n_1497, QN => n14771);
   REGISTERS_reg_35_15_inst : DFF_X1 port map( D => n8841, CK => CLK, Q => 
                           n_1498, QN => n14772);
   REGISTERS_reg_35_14_inst : DFF_X1 port map( D => n8840, CK => CLK, Q => 
                           n_1499, QN => n14773);
   REGISTERS_reg_35_13_inst : DFF_X1 port map( D => n8839, CK => CLK, Q => 
                           n_1500, QN => n14774);
   REGISTERS_reg_35_12_inst : DFF_X1 port map( D => n8838, CK => CLK, Q => 
                           n_1501, QN => n14775);
   REGISTERS_reg_35_11_inst : DFF_X1 port map( D => n8837, CK => CLK, Q => 
                           n_1502, QN => n14776);
   REGISTERS_reg_35_10_inst : DFF_X1 port map( D => n8836, CK => CLK, Q => 
                           n_1503, QN => n14777);
   REGISTERS_reg_35_9_inst : DFF_X1 port map( D => n8835, CK => CLK, Q => 
                           n_1504, QN => n14778);
   REGISTERS_reg_35_8_inst : DFF_X1 port map( D => n8834, CK => CLK, Q => 
                           n_1505, QN => n14779);
   REGISTERS_reg_35_7_inst : DFF_X1 port map( D => n8833, CK => CLK, Q => 
                           n_1506, QN => n14780);
   REGISTERS_reg_35_6_inst : DFF_X1 port map( D => n8832, CK => CLK, Q => 
                           n_1507, QN => n14781);
   REGISTERS_reg_35_5_inst : DFF_X1 port map( D => n8831, CK => CLK, Q => 
                           n_1508, QN => n14782);
   REGISTERS_reg_35_4_inst : DFF_X1 port map( D => n8830, CK => CLK, Q => 
                           n_1509, QN => n14783);
   REGISTERS_reg_35_3_inst : DFF_X1 port map( D => n8829, CK => CLK, Q => 
                           n_1510, QN => n14784);
   REGISTERS_reg_35_2_inst : DFF_X1 port map( D => n8828, CK => CLK, Q => 
                           n_1511, QN => n14785);
   REGISTERS_reg_35_1_inst : DFF_X1 port map( D => n8827, CK => CLK, Q => 
                           n_1512, QN => n14786);
   REGISTERS_reg_35_0_inst : DFF_X1 port map( D => n8826, CK => CLK, Q => 
                           n_1513, QN => n14787);
   REGISTERS_reg_36_31_inst : DFF_X1 port map( D => n8825, CK => CLK, Q => 
                           n_1514, QN => n14788);
   REGISTERS_reg_36_30_inst : DFF_X1 port map( D => n8824, CK => CLK, Q => 
                           n_1515, QN => n14789);
   REGISTERS_reg_36_29_inst : DFF_X1 port map( D => n8823, CK => CLK, Q => 
                           n_1516, QN => n14790);
   REGISTERS_reg_36_28_inst : DFF_X1 port map( D => n8822, CK => CLK, Q => 
                           n_1517, QN => n14791);
   REGISTERS_reg_36_27_inst : DFF_X1 port map( D => n8821, CK => CLK, Q => 
                           n_1518, QN => n14792);
   REGISTERS_reg_36_26_inst : DFF_X1 port map( D => n8820, CK => CLK, Q => 
                           n_1519, QN => n14793);
   REGISTERS_reg_36_25_inst : DFF_X1 port map( D => n8819, CK => CLK, Q => 
                           n_1520, QN => n14794);
   REGISTERS_reg_36_24_inst : DFF_X1 port map( D => n8818, CK => CLK, Q => 
                           n_1521, QN => n14795);
   REGISTERS_reg_36_23_inst : DFF_X1 port map( D => n8817, CK => CLK, Q => 
                           n_1522, QN => n14796);
   REGISTERS_reg_36_22_inst : DFF_X1 port map( D => n8816, CK => CLK, Q => 
                           n_1523, QN => n14797);
   REGISTERS_reg_36_21_inst : DFF_X1 port map( D => n8815, CK => CLK, Q => 
                           n_1524, QN => n14798);
   REGISTERS_reg_36_20_inst : DFF_X1 port map( D => n8814, CK => CLK, Q => 
                           n_1525, QN => n14799);
   REGISTERS_reg_36_19_inst : DFF_X1 port map( D => n8813, CK => CLK, Q => 
                           n_1526, QN => n14800);
   REGISTERS_reg_36_18_inst : DFF_X1 port map( D => n8812, CK => CLK, Q => 
                           n_1527, QN => n14801);
   REGISTERS_reg_36_17_inst : DFF_X1 port map( D => n8811, CK => CLK, Q => 
                           n_1528, QN => n14802);
   REGISTERS_reg_36_16_inst : DFF_X1 port map( D => n8810, CK => CLK, Q => 
                           n_1529, QN => n14803);
   REGISTERS_reg_36_15_inst : DFF_X1 port map( D => n8809, CK => CLK, Q => 
                           n_1530, QN => n14804);
   REGISTERS_reg_36_14_inst : DFF_X1 port map( D => n8808, CK => CLK, Q => 
                           n_1531, QN => n14805);
   REGISTERS_reg_36_13_inst : DFF_X1 port map( D => n8807, CK => CLK, Q => 
                           n_1532, QN => n14806);
   REGISTERS_reg_36_12_inst : DFF_X1 port map( D => n8806, CK => CLK, Q => 
                           n_1533, QN => n14807);
   REGISTERS_reg_36_11_inst : DFF_X1 port map( D => n8805, CK => CLK, Q => 
                           n_1534, QN => n14808);
   REGISTERS_reg_36_10_inst : DFF_X1 port map( D => n8804, CK => CLK, Q => 
                           n_1535, QN => n14809);
   REGISTERS_reg_36_9_inst : DFF_X1 port map( D => n8803, CK => CLK, Q => 
                           n_1536, QN => n14810);
   REGISTERS_reg_36_8_inst : DFF_X1 port map( D => n8802, CK => CLK, Q => 
                           n_1537, QN => n14811);
   REGISTERS_reg_36_7_inst : DFF_X1 port map( D => n8801, CK => CLK, Q => 
                           n_1538, QN => n14812);
   REGISTERS_reg_36_6_inst : DFF_X1 port map( D => n8800, CK => CLK, Q => 
                           n_1539, QN => n14813);
   REGISTERS_reg_36_5_inst : DFF_X1 port map( D => n8799, CK => CLK, Q => 
                           n_1540, QN => n14814);
   REGISTERS_reg_36_4_inst : DFF_X1 port map( D => n8798, CK => CLK, Q => 
                           n_1541, QN => n14815);
   REGISTERS_reg_36_3_inst : DFF_X1 port map( D => n8797, CK => CLK, Q => 
                           n_1542, QN => n14816);
   REGISTERS_reg_36_2_inst : DFF_X1 port map( D => n8796, CK => CLK, Q => 
                           n_1543, QN => n14817);
   REGISTERS_reg_36_1_inst : DFF_X1 port map( D => n8795, CK => CLK, Q => 
                           n_1544, QN => n14818);
   REGISTERS_reg_36_0_inst : DFF_X1 port map( D => n8794, CK => CLK, Q => 
                           n_1545, QN => n14819);
   REGISTERS_reg_37_31_inst : DFF_X1 port map( D => n8793, CK => CLK, Q => 
                           n_1546, QN => n14820);
   REGISTERS_reg_37_30_inst : DFF_X1 port map( D => n8792, CK => CLK, Q => 
                           n_1547, QN => n14821);
   REGISTERS_reg_37_29_inst : DFF_X1 port map( D => n8791, CK => CLK, Q => 
                           n_1548, QN => n14822);
   REGISTERS_reg_37_28_inst : DFF_X1 port map( D => n8790, CK => CLK, Q => 
                           n_1549, QN => n14823);
   REGISTERS_reg_37_27_inst : DFF_X1 port map( D => n8789, CK => CLK, Q => 
                           n_1550, QN => n14824);
   REGISTERS_reg_37_26_inst : DFF_X1 port map( D => n8788, CK => CLK, Q => 
                           n_1551, QN => n14825);
   REGISTERS_reg_37_25_inst : DFF_X1 port map( D => n8787, CK => CLK, Q => 
                           n_1552, QN => n14826);
   REGISTERS_reg_37_24_inst : DFF_X1 port map( D => n8786, CK => CLK, Q => 
                           n_1553, QN => n14827);
   REGISTERS_reg_37_23_inst : DFF_X1 port map( D => n8785, CK => CLK, Q => 
                           n_1554, QN => n14828);
   REGISTERS_reg_37_22_inst : DFF_X1 port map( D => n8784, CK => CLK, Q => 
                           n_1555, QN => n14829);
   REGISTERS_reg_37_21_inst : DFF_X1 port map( D => n8783, CK => CLK, Q => 
                           n_1556, QN => n14830);
   REGISTERS_reg_37_20_inst : DFF_X1 port map( D => n8782, CK => CLK, Q => 
                           n_1557, QN => n14831);
   REGISTERS_reg_37_19_inst : DFF_X1 port map( D => n8781, CK => CLK, Q => 
                           n_1558, QN => n14832);
   REGISTERS_reg_37_18_inst : DFF_X1 port map( D => n8780, CK => CLK, Q => 
                           n_1559, QN => n14833);
   REGISTERS_reg_37_17_inst : DFF_X1 port map( D => n8779, CK => CLK, Q => 
                           n_1560, QN => n14834);
   REGISTERS_reg_37_16_inst : DFF_X1 port map( D => n8778, CK => CLK, Q => 
                           n_1561, QN => n14835);
   REGISTERS_reg_37_15_inst : DFF_X1 port map( D => n8777, CK => CLK, Q => 
                           n_1562, QN => n14836);
   REGISTERS_reg_37_14_inst : DFF_X1 port map( D => n8776, CK => CLK, Q => 
                           n_1563, QN => n14837);
   REGISTERS_reg_37_13_inst : DFF_X1 port map( D => n8775, CK => CLK, Q => 
                           n_1564, QN => n14838);
   REGISTERS_reg_37_12_inst : DFF_X1 port map( D => n8774, CK => CLK, Q => 
                           n_1565, QN => n14839);
   REGISTERS_reg_37_11_inst : DFF_X1 port map( D => n8773, CK => CLK, Q => 
                           n_1566, QN => n14840);
   REGISTERS_reg_37_10_inst : DFF_X1 port map( D => n8772, CK => CLK, Q => 
                           n_1567, QN => n14841);
   REGISTERS_reg_37_9_inst : DFF_X1 port map( D => n8771, CK => CLK, Q => 
                           n_1568, QN => n14842);
   REGISTERS_reg_37_8_inst : DFF_X1 port map( D => n8770, CK => CLK, Q => 
                           n_1569, QN => n14843);
   REGISTERS_reg_37_7_inst : DFF_X1 port map( D => n8769, CK => CLK, Q => 
                           n_1570, QN => n14844);
   REGISTERS_reg_37_6_inst : DFF_X1 port map( D => n8768, CK => CLK, Q => 
                           n_1571, QN => n14845);
   REGISTERS_reg_37_5_inst : DFF_X1 port map( D => n8767, CK => CLK, Q => 
                           n_1572, QN => n14846);
   REGISTERS_reg_37_4_inst : DFF_X1 port map( D => n8766, CK => CLK, Q => 
                           n_1573, QN => n14847);
   REGISTERS_reg_37_3_inst : DFF_X1 port map( D => n8765, CK => CLK, Q => 
                           n_1574, QN => n14848);
   REGISTERS_reg_37_2_inst : DFF_X1 port map( D => n8764, CK => CLK, Q => 
                           n_1575, QN => n14849);
   REGISTERS_reg_37_1_inst : DFF_X1 port map( D => n8763, CK => CLK, Q => 
                           n_1576, QN => n14850);
   REGISTERS_reg_37_0_inst : DFF_X1 port map( D => n8762, CK => CLK, Q => 
                           n_1577, QN => n14851);
   REGISTERS_reg_38_19_inst : DFF_X1 port map( D => n8749, CK => CLK, Q => n578
                           , QN => n12921);
   REGISTERS_reg_38_18_inst : DFF_X1 port map( D => n8748, CK => CLK, Q => n580
                           , QN => n12920);
   REGISTERS_reg_38_17_inst : DFF_X1 port map( D => n8747, CK => CLK, Q => n582
                           , QN => n12919);
   REGISTERS_reg_38_16_inst : DFF_X1 port map( D => n8746, CK => CLK, Q => n584
                           , QN => n12918);
   REGISTERS_reg_38_15_inst : DFF_X1 port map( D => n8745, CK => CLK, Q => n586
                           , QN => n12917);
   REGISTERS_reg_38_14_inst : DFF_X1 port map( D => n8744, CK => CLK, Q => n588
                           , QN => n12916);
   REGISTERS_reg_38_13_inst : DFF_X1 port map( D => n8743, CK => CLK, Q => n590
                           , QN => n12915);
   REGISTERS_reg_38_12_inst : DFF_X1 port map( D => n8742, CK => CLK, Q => n592
                           , QN => n12914);
   REGISTERS_reg_38_11_inst : DFF_X1 port map( D => n8741, CK => CLK, Q => n594
                           , QN => n12913);
   REGISTERS_reg_38_10_inst : DFF_X1 port map( D => n8740, CK => CLK, Q => n596
                           , QN => n12912);
   REGISTERS_reg_38_9_inst : DFF_X1 port map( D => n8739, CK => CLK, Q => n598,
                           QN => n12911);
   REGISTERS_reg_38_8_inst : DFF_X1 port map( D => n8738, CK => CLK, Q => n600,
                           QN => n12910);
   REGISTERS_reg_38_7_inst : DFF_X1 port map( D => n8737, CK => CLK, Q => n602,
                           QN => n12909);
   REGISTERS_reg_38_6_inst : DFF_X1 port map( D => n8736, CK => CLK, Q => n604,
                           QN => n12908);
   REGISTERS_reg_38_5_inst : DFF_X1 port map( D => n8735, CK => CLK, Q => n606,
                           QN => n12907);
   REGISTERS_reg_38_4_inst : DFF_X1 port map( D => n8734, CK => CLK, Q => n608,
                           QN => n12906);
   REGISTERS_reg_38_3_inst : DFF_X1 port map( D => n8733, CK => CLK, Q => n610,
                           QN => n12905);
   REGISTERS_reg_38_2_inst : DFF_X1 port map( D => n8732, CK => CLK, Q => n612,
                           QN => n12904);
   REGISTERS_reg_38_1_inst : DFF_X1 port map( D => n8731, CK => CLK, Q => n614,
                           QN => n12903);
   REGISTERS_reg_38_0_inst : DFF_X1 port map( D => n8730, CK => CLK, Q => n616,
                           QN => n12902);
   REGISTERS_reg_39_31_inst : DFF_X1 port map( D => n8729, CK => CLK, Q => n98,
                           QN => n12709);
   REGISTERS_reg_41_31_inst : DFF_X1 port map( D => n8665, CK => CLK, Q => 
                           n6241, QN => n12901);
   REGISTERS_reg_41_30_inst : DFF_X1 port map( D => n8664, CK => CLK, Q => 
                           n6240, QN => n12900);
   REGISTERS_reg_41_29_inst : DFF_X1 port map( D => n8663, CK => CLK, Q => 
                           n6239, QN => n12899);
   REGISTERS_reg_41_28_inst : DFF_X1 port map( D => n8662, CK => CLK, Q => 
                           n6238, QN => n12898);
   REGISTERS_reg_41_27_inst : DFF_X1 port map( D => n8661, CK => CLK, Q => 
                           n6237, QN => n12897);
   REGISTERS_reg_41_26_inst : DFF_X1 port map( D => n8660, CK => CLK, Q => 
                           n6236, QN => n12896);
   REGISTERS_reg_41_25_inst : DFF_X1 port map( D => n8659, CK => CLK, Q => 
                           n6235, QN => n12895);
   REGISTERS_reg_41_24_inst : DFF_X1 port map( D => n8658, CK => CLK, Q => 
                           n6234, QN => n12894);
   REGISTERS_reg_41_23_inst : DFF_X1 port map( D => n8657, CK => CLK, Q => 
                           n6233, QN => n12893);
   REGISTERS_reg_41_22_inst : DFF_X1 port map( D => n8656, CK => CLK, Q => 
                           n6232, QN => n12892);
   REGISTERS_reg_41_21_inst : DFF_X1 port map( D => n8655, CK => CLK, Q => 
                           n6231, QN => n12891);
   REGISTERS_reg_41_20_inst : DFF_X1 port map( D => n8654, CK => CLK, Q => 
                           n6230, QN => n12890);
   REGISTERS_reg_41_19_inst : DFF_X1 port map( D => n8653, CK => CLK, Q => 
                           n6229, QN => n12889);
   REGISTERS_reg_41_18_inst : DFF_X1 port map( D => n8652, CK => CLK, Q => 
                           n6228, QN => n12888);
   REGISTERS_reg_41_17_inst : DFF_X1 port map( D => n8651, CK => CLK, Q => 
                           n6227, QN => n12887);
   REGISTERS_reg_41_16_inst : DFF_X1 port map( D => n8650, CK => CLK, Q => 
                           n6226, QN => n12886);
   REGISTERS_reg_41_15_inst : DFF_X1 port map( D => n8649, CK => CLK, Q => 
                           n6225, QN => n12885);
   REGISTERS_reg_41_14_inst : DFF_X1 port map( D => n8648, CK => CLK, Q => 
                           n6224, QN => n12884);
   REGISTERS_reg_41_13_inst : DFF_X1 port map( D => n8647, CK => CLK, Q => 
                           n6223, QN => n12883);
   REGISTERS_reg_41_12_inst : DFF_X1 port map( D => n8646, CK => CLK, Q => 
                           n6222, QN => n12882);
   REGISTERS_reg_41_11_inst : DFF_X1 port map( D => n8645, CK => CLK, Q => 
                           n6221, QN => n12881);
   REGISTERS_reg_41_10_inst : DFF_X1 port map( D => n8644, CK => CLK, Q => 
                           n6220, QN => n12880);
   REGISTERS_reg_41_9_inst : DFF_X1 port map( D => n8643, CK => CLK, Q => n6219
                           , QN => n12879);
   REGISTERS_reg_41_8_inst : DFF_X1 port map( D => n8642, CK => CLK, Q => n6218
                           , QN => n12878);
   REGISTERS_reg_41_7_inst : DFF_X1 port map( D => n8641, CK => CLK, Q => n6217
                           , QN => n12877);
   REGISTERS_reg_41_6_inst : DFF_X1 port map( D => n8640, CK => CLK, Q => n6216
                           , QN => n12876);
   REGISTERS_reg_41_5_inst : DFF_X1 port map( D => n8639, CK => CLK, Q => n6215
                           , QN => n12875);
   REGISTERS_reg_41_4_inst : DFF_X1 port map( D => n8638, CK => CLK, Q => n6214
                           , QN => n12874);
   REGISTERS_reg_41_3_inst : DFF_X1 port map( D => n8637, CK => CLK, Q => n6213
                           , QN => n12873);
   REGISTERS_reg_41_2_inst : DFF_X1 port map( D => n8636, CK => CLK, Q => n6212
                           , QN => n12872);
   REGISTERS_reg_41_1_inst : DFF_X1 port map( D => n8635, CK => CLK, Q => n6211
                           , QN => n12871);
   REGISTERS_reg_41_0_inst : DFF_X1 port map( D => n8634, CK => CLK, Q => n6210
                           , QN => n12870);
   REGISTERS_reg_42_31_inst : DFF_X1 port map( D => n8633, CK => CLK, Q => 
                           n_1578, QN => n14852);
   REGISTERS_reg_42_30_inst : DFF_X1 port map( D => n8632, CK => CLK, Q => 
                           n_1579, QN => n14853);
   REGISTERS_reg_42_29_inst : DFF_X1 port map( D => n8631, CK => CLK, Q => 
                           n_1580, QN => n14854);
   REGISTERS_reg_42_28_inst : DFF_X1 port map( D => n8630, CK => CLK, Q => 
                           n_1581, QN => n14855);
   REGISTERS_reg_42_27_inst : DFF_X1 port map( D => n8629, CK => CLK, Q => 
                           n_1582, QN => n14856);
   REGISTERS_reg_42_26_inst : DFF_X1 port map( D => n8628, CK => CLK, Q => 
                           n_1583, QN => n14857);
   REGISTERS_reg_42_25_inst : DFF_X1 port map( D => n8627, CK => CLK, Q => 
                           n_1584, QN => n14858);
   REGISTERS_reg_42_24_inst : DFF_X1 port map( D => n8626, CK => CLK, Q => 
                           n_1585, QN => n14859);
   REGISTERS_reg_42_23_inst : DFF_X1 port map( D => n8625, CK => CLK, Q => 
                           n_1586, QN => n14860);
   REGISTERS_reg_42_22_inst : DFF_X1 port map( D => n8624, CK => CLK, Q => 
                           n_1587, QN => n14861);
   REGISTERS_reg_42_21_inst : DFF_X1 port map( D => n8623, CK => CLK, Q => 
                           n_1588, QN => n14862);
   REGISTERS_reg_42_20_inst : DFF_X1 port map( D => n8622, CK => CLK, Q => 
                           n_1589, QN => n14863);
   REGISTERS_reg_42_19_inst : DFF_X1 port map( D => n8621, CK => CLK, Q => 
                           n_1590, QN => n14864);
   REGISTERS_reg_42_18_inst : DFF_X1 port map( D => n8620, CK => CLK, Q => 
                           n_1591, QN => n14865);
   REGISTERS_reg_42_17_inst : DFF_X1 port map( D => n8619, CK => CLK, Q => 
                           n_1592, QN => n14866);
   REGISTERS_reg_42_16_inst : DFF_X1 port map( D => n8618, CK => CLK, Q => 
                           n_1593, QN => n14867);
   REGISTERS_reg_42_15_inst : DFF_X1 port map( D => n8617, CK => CLK, Q => 
                           n_1594, QN => n14868);
   REGISTERS_reg_42_14_inst : DFF_X1 port map( D => n8616, CK => CLK, Q => 
                           n_1595, QN => n14869);
   REGISTERS_reg_42_13_inst : DFF_X1 port map( D => n8615, CK => CLK, Q => 
                           n_1596, QN => n14870);
   REGISTERS_reg_42_12_inst : DFF_X1 port map( D => n8614, CK => CLK, Q => 
                           n_1597, QN => n14871);
   REGISTERS_reg_42_11_inst : DFF_X1 port map( D => n8613, CK => CLK, Q => 
                           n_1598, QN => n14872);
   REGISTERS_reg_42_10_inst : DFF_X1 port map( D => n8612, CK => CLK, Q => 
                           n_1599, QN => n14873);
   REGISTERS_reg_42_9_inst : DFF_X1 port map( D => n8611, CK => CLK, Q => 
                           n_1600, QN => n14874);
   REGISTERS_reg_42_8_inst : DFF_X1 port map( D => n8610, CK => CLK, Q => 
                           n_1601, QN => n14875);
   REGISTERS_reg_42_7_inst : DFF_X1 port map( D => n8609, CK => CLK, Q => 
                           n_1602, QN => n14876);
   REGISTERS_reg_42_6_inst : DFF_X1 port map( D => n8608, CK => CLK, Q => 
                           n_1603, QN => n14877);
   REGISTERS_reg_42_5_inst : DFF_X1 port map( D => n8607, CK => CLK, Q => 
                           n_1604, QN => n14878);
   REGISTERS_reg_42_4_inst : DFF_X1 port map( D => n8606, CK => CLK, Q => 
                           n_1605, QN => n14879);
   REGISTERS_reg_42_3_inst : DFF_X1 port map( D => n8605, CK => CLK, Q => 
                           n_1606, QN => n14880);
   REGISTERS_reg_42_2_inst : DFF_X1 port map( D => n8604, CK => CLK, Q => 
                           n_1607, QN => n14881);
   REGISTERS_reg_42_1_inst : DFF_X1 port map( D => n8603, CK => CLK, Q => 
                           n_1608, QN => n14882);
   REGISTERS_reg_42_0_inst : DFF_X1 port map( D => n8602, CK => CLK, Q => 
                           n_1609, QN => n14883);
   REGISTERS_reg_43_31_inst : DFF_X1 port map( D => n8601, CK => CLK, Q => 
                           n_1610, QN => n14884);
   REGISTERS_reg_43_30_inst : DFF_X1 port map( D => n8600, CK => CLK, Q => 
                           n_1611, QN => n14885);
   REGISTERS_reg_43_29_inst : DFF_X1 port map( D => n8599, CK => CLK, Q => 
                           n_1612, QN => n14886);
   REGISTERS_reg_43_28_inst : DFF_X1 port map( D => n8598, CK => CLK, Q => 
                           n_1613, QN => n14887);
   REGISTERS_reg_43_27_inst : DFF_X1 port map( D => n8597, CK => CLK, Q => 
                           n_1614, QN => n14888);
   REGISTERS_reg_43_26_inst : DFF_X1 port map( D => n8596, CK => CLK, Q => 
                           n_1615, QN => n14889);
   REGISTERS_reg_43_25_inst : DFF_X1 port map( D => n8595, CK => CLK, Q => 
                           n_1616, QN => n14890);
   REGISTERS_reg_43_24_inst : DFF_X1 port map( D => n8594, CK => CLK, Q => 
                           n_1617, QN => n14891);
   REGISTERS_reg_43_23_inst : DFF_X1 port map( D => n8593, CK => CLK, Q => 
                           n_1618, QN => n14892);
   REGISTERS_reg_43_22_inst : DFF_X1 port map( D => n8592, CK => CLK, Q => 
                           n_1619, QN => n14893);
   REGISTERS_reg_43_21_inst : DFF_X1 port map( D => n8591, CK => CLK, Q => 
                           n_1620, QN => n14894);
   REGISTERS_reg_43_20_inst : DFF_X1 port map( D => n8590, CK => CLK, Q => 
                           n_1621, QN => n14895);
   REGISTERS_reg_43_19_inst : DFF_X1 port map( D => n8589, CK => CLK, Q => 
                           n_1622, QN => n14896);
   REGISTERS_reg_43_18_inst : DFF_X1 port map( D => n8588, CK => CLK, Q => 
                           n_1623, QN => n14897);
   REGISTERS_reg_43_17_inst : DFF_X1 port map( D => n8587, CK => CLK, Q => 
                           n_1624, QN => n14898);
   REGISTERS_reg_43_16_inst : DFF_X1 port map( D => n8586, CK => CLK, Q => 
                           n_1625, QN => n14899);
   REGISTERS_reg_43_15_inst : DFF_X1 port map( D => n8585, CK => CLK, Q => 
                           n_1626, QN => n14900);
   REGISTERS_reg_43_14_inst : DFF_X1 port map( D => n8584, CK => CLK, Q => 
                           n_1627, QN => n14901);
   REGISTERS_reg_43_13_inst : DFF_X1 port map( D => n8583, CK => CLK, Q => 
                           n_1628, QN => n14902);
   REGISTERS_reg_43_12_inst : DFF_X1 port map( D => n8582, CK => CLK, Q => 
                           n_1629, QN => n14903);
   REGISTERS_reg_43_11_inst : DFF_X1 port map( D => n8581, CK => CLK, Q => 
                           n_1630, QN => n14904);
   REGISTERS_reg_43_10_inst : DFF_X1 port map( D => n8580, CK => CLK, Q => 
                           n_1631, QN => n14905);
   REGISTERS_reg_43_9_inst : DFF_X1 port map( D => n8579, CK => CLK, Q => 
                           n_1632, QN => n14906);
   REGISTERS_reg_43_8_inst : DFF_X1 port map( D => n8578, CK => CLK, Q => 
                           n_1633, QN => n14907);
   REGISTERS_reg_43_7_inst : DFF_X1 port map( D => n8577, CK => CLK, Q => 
                           n_1634, QN => n14908);
   REGISTERS_reg_43_6_inst : DFF_X1 port map( D => n8576, CK => CLK, Q => 
                           n_1635, QN => n14909);
   REGISTERS_reg_43_5_inst : DFF_X1 port map( D => n8575, CK => CLK, Q => 
                           n_1636, QN => n14910);
   REGISTERS_reg_43_4_inst : DFF_X1 port map( D => n8574, CK => CLK, Q => 
                           n_1637, QN => n14911);
   REGISTERS_reg_43_3_inst : DFF_X1 port map( D => n8573, CK => CLK, Q => 
                           n_1638, QN => n14912);
   REGISTERS_reg_43_2_inst : DFF_X1 port map( D => n8572, CK => CLK, Q => 
                           n_1639, QN => n14913);
   REGISTERS_reg_43_1_inst : DFF_X1 port map( D => n8571, CK => CLK, Q => 
                           n_1640, QN => n14914);
   REGISTERS_reg_43_0_inst : DFF_X1 port map( D => n8570, CK => CLK, Q => 
                           n_1641, QN => n14915);
   REGISTERS_reg_44_31_inst : DFF_X1 port map( D => n8569, CK => CLK, Q => 
                           n_1642, QN => n14916);
   REGISTERS_reg_44_30_inst : DFF_X1 port map( D => n8568, CK => CLK, Q => 
                           n_1643, QN => n14917);
   REGISTERS_reg_44_29_inst : DFF_X1 port map( D => n8567, CK => CLK, Q => 
                           n_1644, QN => n14918);
   REGISTERS_reg_44_28_inst : DFF_X1 port map( D => n8566, CK => CLK, Q => 
                           n_1645, QN => n14919);
   REGISTERS_reg_44_27_inst : DFF_X1 port map( D => n8565, CK => CLK, Q => 
                           n_1646, QN => n14920);
   REGISTERS_reg_44_26_inst : DFF_X1 port map( D => n8564, CK => CLK, Q => 
                           n_1647, QN => n14921);
   REGISTERS_reg_44_25_inst : DFF_X1 port map( D => n8563, CK => CLK, Q => 
                           n_1648, QN => n14922);
   REGISTERS_reg_44_24_inst : DFF_X1 port map( D => n8562, CK => CLK, Q => 
                           n_1649, QN => n14923);
   REGISTERS_reg_44_23_inst : DFF_X1 port map( D => n8561, CK => CLK, Q => 
                           n_1650, QN => n14924);
   REGISTERS_reg_44_22_inst : DFF_X1 port map( D => n8560, CK => CLK, Q => 
                           n_1651, QN => n14925);
   REGISTERS_reg_44_21_inst : DFF_X1 port map( D => n8559, CK => CLK, Q => 
                           n_1652, QN => n14926);
   REGISTERS_reg_44_20_inst : DFF_X1 port map( D => n8558, CK => CLK, Q => 
                           n_1653, QN => n14927);
   REGISTERS_reg_44_19_inst : DFF_X1 port map( D => n8557, CK => CLK, Q => 
                           n_1654, QN => n14928);
   REGISTERS_reg_44_18_inst : DFF_X1 port map( D => n8556, CK => CLK, Q => 
                           n_1655, QN => n14929);
   REGISTERS_reg_44_17_inst : DFF_X1 port map( D => n8555, CK => CLK, Q => 
                           n_1656, QN => n14930);
   REGISTERS_reg_44_16_inst : DFF_X1 port map( D => n8554, CK => CLK, Q => 
                           n_1657, QN => n14931);
   REGISTERS_reg_44_15_inst : DFF_X1 port map( D => n8553, CK => CLK, Q => 
                           n_1658, QN => n14932);
   REGISTERS_reg_44_14_inst : DFF_X1 port map( D => n8552, CK => CLK, Q => 
                           n_1659, QN => n14933);
   REGISTERS_reg_44_13_inst : DFF_X1 port map( D => n8551, CK => CLK, Q => 
                           n_1660, QN => n14934);
   REGISTERS_reg_44_12_inst : DFF_X1 port map( D => n8550, CK => CLK, Q => 
                           n_1661, QN => n14935);
   REGISTERS_reg_44_11_inst : DFF_X1 port map( D => n8549, CK => CLK, Q => 
                           n_1662, QN => n14936);
   REGISTERS_reg_44_10_inst : DFF_X1 port map( D => n8548, CK => CLK, Q => 
                           n_1663, QN => n14937);
   REGISTERS_reg_44_9_inst : DFF_X1 port map( D => n8547, CK => CLK, Q => 
                           n_1664, QN => n14938);
   REGISTERS_reg_44_8_inst : DFF_X1 port map( D => n8546, CK => CLK, Q => 
                           n_1665, QN => n14939);
   REGISTERS_reg_44_7_inst : DFF_X1 port map( D => n8545, CK => CLK, Q => 
                           n_1666, QN => n14940);
   REGISTERS_reg_44_6_inst : DFF_X1 port map( D => n8544, CK => CLK, Q => 
                           n_1667, QN => n14941);
   REGISTERS_reg_44_5_inst : DFF_X1 port map( D => n8543, CK => CLK, Q => 
                           n_1668, QN => n14942);
   REGISTERS_reg_44_4_inst : DFF_X1 port map( D => n8542, CK => CLK, Q => 
                           n_1669, QN => n14943);
   REGISTERS_reg_44_3_inst : DFF_X1 port map( D => n8541, CK => CLK, Q => 
                           n_1670, QN => n14944);
   REGISTERS_reg_44_2_inst : DFF_X1 port map( D => n8540, CK => CLK, Q => 
                           n_1671, QN => n14945);
   REGISTERS_reg_44_1_inst : DFF_X1 port map( D => n8539, CK => CLK, Q => 
                           n_1672, QN => n14946);
   REGISTERS_reg_44_0_inst : DFF_X1 port map( D => n8538, CK => CLK, Q => 
                           n_1673, QN => n14947);
   REGISTERS_reg_46_31_inst : DFF_X1 port map( D => n8505, CK => CLK, Q => 
                           n6177, QN => n12869);
   REGISTERS_reg_46_30_inst : DFF_X1 port map( D => n8504, CK => CLK, Q => 
                           n6176, QN => n12868);
   REGISTERS_reg_46_29_inst : DFF_X1 port map( D => n8503, CK => CLK, Q => 
                           n6175, QN => n12867);
   REGISTERS_reg_46_28_inst : DFF_X1 port map( D => n8502, CK => CLK, Q => 
                           n6174, QN => n12866);
   REGISTERS_reg_46_27_inst : DFF_X1 port map( D => n8501, CK => CLK, Q => 
                           n6173, QN => n12865);
   REGISTERS_reg_46_26_inst : DFF_X1 port map( D => n8500, CK => CLK, Q => 
                           n6172, QN => n12864);
   REGISTERS_reg_46_25_inst : DFF_X1 port map( D => n8499, CK => CLK, Q => 
                           n6171, QN => n12863);
   REGISTERS_reg_46_24_inst : DFF_X1 port map( D => n8498, CK => CLK, Q => 
                           n6170, QN => n12862);
   REGISTERS_reg_46_23_inst : DFF_X1 port map( D => n8497, CK => CLK, Q => 
                           n6169, QN => n12861);
   REGISTERS_reg_46_22_inst : DFF_X1 port map( D => n8496, CK => CLK, Q => 
                           n6168, QN => n12860);
   REGISTERS_reg_46_21_inst : DFF_X1 port map( D => n8495, CK => CLK, Q => 
                           n6167, QN => n12859);
   REGISTERS_reg_46_20_inst : DFF_X1 port map( D => n8494, CK => CLK, Q => 
                           n6166, QN => n12858);
   REGISTERS_reg_46_19_inst : DFF_X1 port map( D => n8493, CK => CLK, Q => 
                           n6165, QN => n12857);
   REGISTERS_reg_46_18_inst : DFF_X1 port map( D => n8492, CK => CLK, Q => 
                           n6164, QN => n12856);
   REGISTERS_reg_46_17_inst : DFF_X1 port map( D => n8491, CK => CLK, Q => 
                           n6163, QN => n12855);
   REGISTERS_reg_46_16_inst : DFF_X1 port map( D => n8490, CK => CLK, Q => 
                           n6162, QN => n12854);
   REGISTERS_reg_46_15_inst : DFF_X1 port map( D => n8489, CK => CLK, Q => 
                           n6161, QN => n12853);
   REGISTERS_reg_46_14_inst : DFF_X1 port map( D => n8488, CK => CLK, Q => 
                           n6160, QN => n12852);
   REGISTERS_reg_46_13_inst : DFF_X1 port map( D => n8487, CK => CLK, Q => 
                           n6159, QN => n12851);
   REGISTERS_reg_46_12_inst : DFF_X1 port map( D => n8486, CK => CLK, Q => 
                           n6158, QN => n12850);
   REGISTERS_reg_46_11_inst : DFF_X1 port map( D => n8485, CK => CLK, Q => 
                           n6157, QN => n12849);
   REGISTERS_reg_46_10_inst : DFF_X1 port map( D => n8484, CK => CLK, Q => 
                           n6156, QN => n12848);
   REGISTERS_reg_46_9_inst : DFF_X1 port map( D => n8483, CK => CLK, Q => n6155
                           , QN => n12847);
   REGISTERS_reg_46_8_inst : DFF_X1 port map( D => n8482, CK => CLK, Q => n6154
                           , QN => n12846);
   REGISTERS_reg_46_7_inst : DFF_X1 port map( D => n8481, CK => CLK, Q => n6153
                           , QN => n12845);
   REGISTERS_reg_46_6_inst : DFF_X1 port map( D => n8480, CK => CLK, Q => n6152
                           , QN => n12844);
   REGISTERS_reg_46_5_inst : DFF_X1 port map( D => n8479, CK => CLK, Q => n6151
                           , QN => n12843);
   REGISTERS_reg_46_4_inst : DFF_X1 port map( D => n8478, CK => CLK, Q => n6150
                           , QN => n12842);
   REGISTERS_reg_46_3_inst : DFF_X1 port map( D => n8477, CK => CLK, Q => n6149
                           , QN => n12841);
   REGISTERS_reg_46_2_inst : DFF_X1 port map( D => n8476, CK => CLK, Q => n6148
                           , QN => n12840);
   REGISTERS_reg_46_1_inst : DFF_X1 port map( D => n8475, CK => CLK, Q => n6147
                           , QN => n12839);
   REGISTERS_reg_46_0_inst : DFF_X1 port map( D => n8474, CK => CLK, Q => n6146
                           , QN => n12838);
   REGISTERS_reg_47_31_inst : DFF_X1 port map( D => n8473, CK => CLK, Q => 
                           n_1674, QN => n14949);
   REGISTERS_reg_47_30_inst : DFF_X1 port map( D => n8472, CK => CLK, Q => 
                           n_1675, QN => n14950);
   REGISTERS_reg_47_29_inst : DFF_X1 port map( D => n8471, CK => CLK, Q => 
                           n_1676, QN => n14951);
   REGISTERS_reg_47_28_inst : DFF_X1 port map( D => n8470, CK => CLK, Q => 
                           n_1677, QN => n14952);
   REGISTERS_reg_47_27_inst : DFF_X1 port map( D => n8469, CK => CLK, Q => 
                           n_1678, QN => n14953);
   REGISTERS_reg_47_26_inst : DFF_X1 port map( D => n8468, CK => CLK, Q => 
                           n_1679, QN => n14954);
   REGISTERS_reg_47_25_inst : DFF_X1 port map( D => n8467, CK => CLK, Q => 
                           n_1680, QN => n14955);
   REGISTERS_reg_47_24_inst : DFF_X1 port map( D => n8466, CK => CLK, Q => 
                           n_1681, QN => n14956);
   REGISTERS_reg_47_23_inst : DFF_X1 port map( D => n8465, CK => CLK, Q => 
                           n_1682, QN => n14957);
   REGISTERS_reg_47_22_inst : DFF_X1 port map( D => n8464, CK => CLK, Q => 
                           n_1683, QN => n14958);
   REGISTERS_reg_47_21_inst : DFF_X1 port map( D => n8463, CK => CLK, Q => 
                           n_1684, QN => n14959);
   REGISTERS_reg_47_20_inst : DFF_X1 port map( D => n8462, CK => CLK, Q => 
                           n_1685, QN => n14960);
   REGISTERS_reg_47_19_inst : DFF_X1 port map( D => n8461, CK => CLK, Q => 
                           n_1686, QN => n14961);
   REGISTERS_reg_47_18_inst : DFF_X1 port map( D => n8460, CK => CLK, Q => 
                           n_1687, QN => n14962);
   REGISTERS_reg_47_17_inst : DFF_X1 port map( D => n8459, CK => CLK, Q => 
                           n_1688, QN => n14963);
   REGISTERS_reg_47_16_inst : DFF_X1 port map( D => n8458, CK => CLK, Q => 
                           n_1689, QN => n14964);
   REGISTERS_reg_47_15_inst : DFF_X1 port map( D => n8457, CK => CLK, Q => 
                           n_1690, QN => n14965);
   REGISTERS_reg_47_14_inst : DFF_X1 port map( D => n8456, CK => CLK, Q => 
                           n_1691, QN => n14966);
   REGISTERS_reg_47_13_inst : DFF_X1 port map( D => n8455, CK => CLK, Q => 
                           n_1692, QN => n14967);
   REGISTERS_reg_47_12_inst : DFF_X1 port map( D => n8454, CK => CLK, Q => 
                           n_1693, QN => n14968);
   REGISTERS_reg_47_11_inst : DFF_X1 port map( D => n8453, CK => CLK, Q => 
                           n_1694, QN => n14969);
   REGISTERS_reg_47_10_inst : DFF_X1 port map( D => n8452, CK => CLK, Q => 
                           n_1695, QN => n14970);
   REGISTERS_reg_47_9_inst : DFF_X1 port map( D => n8451, CK => CLK, Q => 
                           n_1696, QN => n14971);
   REGISTERS_reg_47_8_inst : DFF_X1 port map( D => n8450, CK => CLK, Q => 
                           n_1697, QN => n14972);
   REGISTERS_reg_47_7_inst : DFF_X1 port map( D => n8449, CK => CLK, Q => 
                           n_1698, QN => n14973);
   REGISTERS_reg_47_6_inst : DFF_X1 port map( D => n8448, CK => CLK, Q => 
                           n_1699, QN => n14974);
   REGISTERS_reg_47_5_inst : DFF_X1 port map( D => n8447, CK => CLK, Q => 
                           n_1700, QN => n14975);
   REGISTERS_reg_47_4_inst : DFF_X1 port map( D => n8446, CK => CLK, Q => 
                           n_1701, QN => n14976);
   REGISTERS_reg_47_3_inst : DFF_X1 port map( D => n8445, CK => CLK, Q => 
                           n_1702, QN => n14977);
   REGISTERS_reg_47_2_inst : DFF_X1 port map( D => n8444, CK => CLK, Q => 
                           n_1703, QN => n14978);
   REGISTERS_reg_47_1_inst : DFF_X1 port map( D => n8443, CK => CLK, Q => 
                           n_1704, QN => n14979);
   REGISTERS_reg_47_0_inst : DFF_X1 port map( D => n8442, CK => CLK, Q => 
                           n_1705, QN => n14980);
   REGISTERS_reg_51_31_inst : DFF_X1 port map( D => n8345, CK => CLK, Q => 
                           n_1706, QN => n15014);
   REGISTERS_reg_51_30_inst : DFF_X1 port map( D => n8344, CK => CLK, Q => 
                           n_1707, QN => n15015);
   REGISTERS_reg_51_29_inst : DFF_X1 port map( D => n8343, CK => CLK, Q => 
                           n_1708, QN => n15016);
   REGISTERS_reg_51_28_inst : DFF_X1 port map( D => n8342, CK => CLK, Q => 
                           n_1709, QN => n15017);
   REGISTERS_reg_51_27_inst : DFF_X1 port map( D => n8341, CK => CLK, Q => 
                           n_1710, QN => n15018);
   REGISTERS_reg_51_26_inst : DFF_X1 port map( D => n8340, CK => CLK, Q => 
                           n_1711, QN => n15019);
   REGISTERS_reg_51_25_inst : DFF_X1 port map( D => n8339, CK => CLK, Q => 
                           n_1712, QN => n15020);
   REGISTERS_reg_51_24_inst : DFF_X1 port map( D => n8338, CK => CLK, Q => 
                           n_1713, QN => n15021);
   REGISTERS_reg_51_23_inst : DFF_X1 port map( D => n8337, CK => CLK, Q => 
                           n_1714, QN => n15022);
   REGISTERS_reg_51_22_inst : DFF_X1 port map( D => n8336, CK => CLK, Q => 
                           n_1715, QN => n15023);
   REGISTERS_reg_51_21_inst : DFF_X1 port map( D => n8335, CK => CLK, Q => 
                           n_1716, QN => n15024);
   REGISTERS_reg_51_20_inst : DFF_X1 port map( D => n8334, CK => CLK, Q => 
                           n_1717, QN => n15025);
   REGISTERS_reg_51_19_inst : DFF_X1 port map( D => n8333, CK => CLK, Q => 
                           n_1718, QN => n15026);
   REGISTERS_reg_51_18_inst : DFF_X1 port map( D => n8332, CK => CLK, Q => 
                           n_1719, QN => n15027);
   REGISTERS_reg_51_17_inst : DFF_X1 port map( D => n8331, CK => CLK, Q => 
                           n_1720, QN => n15028);
   REGISTERS_reg_51_16_inst : DFF_X1 port map( D => n8330, CK => CLK, Q => 
                           n_1721, QN => n15029);
   REGISTERS_reg_51_15_inst : DFF_X1 port map( D => n8329, CK => CLK, Q => 
                           n_1722, QN => n15030);
   REGISTERS_reg_51_14_inst : DFF_X1 port map( D => n8328, CK => CLK, Q => 
                           n_1723, QN => n15031);
   REGISTERS_reg_51_13_inst : DFF_X1 port map( D => n8327, CK => CLK, Q => 
                           n_1724, QN => n15032);
   REGISTERS_reg_51_12_inst : DFF_X1 port map( D => n8326, CK => CLK, Q => 
                           n_1725, QN => n15033);
   REGISTERS_reg_51_11_inst : DFF_X1 port map( D => n8325, CK => CLK, Q => 
                           n_1726, QN => n15034);
   REGISTERS_reg_51_10_inst : DFF_X1 port map( D => n8324, CK => CLK, Q => 
                           n_1727, QN => n15035);
   REGISTERS_reg_51_9_inst : DFF_X1 port map( D => n8323, CK => CLK, Q => 
                           n_1728, QN => n15036);
   REGISTERS_reg_51_8_inst : DFF_X1 port map( D => n8322, CK => CLK, Q => 
                           n_1729, QN => n15037);
   REGISTERS_reg_51_7_inst : DFF_X1 port map( D => n8321, CK => CLK, Q => 
                           n_1730, QN => n15038);
   REGISTERS_reg_51_6_inst : DFF_X1 port map( D => n8320, CK => CLK, Q => 
                           n_1731, QN => n15039);
   REGISTERS_reg_51_5_inst : DFF_X1 port map( D => n8319, CK => CLK, Q => 
                           n_1732, QN => n15040);
   REGISTERS_reg_51_4_inst : DFF_X1 port map( D => n8318, CK => CLK, Q => 
                           n_1733, QN => n15041);
   REGISTERS_reg_51_3_inst : DFF_X1 port map( D => n8317, CK => CLK, Q => 
                           n_1734, QN => n15042);
   REGISTERS_reg_51_2_inst : DFF_X1 port map( D => n8316, CK => CLK, Q => 
                           n_1735, QN => n15043);
   REGISTERS_reg_51_1_inst : DFF_X1 port map( D => n8315, CK => CLK, Q => 
                           n_1736, QN => n15044);
   REGISTERS_reg_51_0_inst : DFF_X1 port map( D => n8314, CK => CLK, Q => 
                           n_1737, QN => n15045);
   REGISTERS_reg_52_31_inst : DFF_X1 port map( D => n8313, CK => CLK, Q => 
                           n_1738, QN => n15046);
   REGISTERS_reg_52_30_inst : DFF_X1 port map( D => n8312, CK => CLK, Q => 
                           n_1739, QN => n15047);
   REGISTERS_reg_52_29_inst : DFF_X1 port map( D => n8311, CK => CLK, Q => 
                           n_1740, QN => n15048);
   REGISTERS_reg_52_28_inst : DFF_X1 port map( D => n8310, CK => CLK, Q => 
                           n_1741, QN => n15049);
   REGISTERS_reg_52_27_inst : DFF_X1 port map( D => n8309, CK => CLK, Q => 
                           n_1742, QN => n15050);
   REGISTERS_reg_52_26_inst : DFF_X1 port map( D => n8308, CK => CLK, Q => 
                           n_1743, QN => n15051);
   REGISTERS_reg_52_25_inst : DFF_X1 port map( D => n8307, CK => CLK, Q => 
                           n_1744, QN => n15052);
   REGISTERS_reg_52_24_inst : DFF_X1 port map( D => n8306, CK => CLK, Q => 
                           n_1745, QN => n15053);
   REGISTERS_reg_52_23_inst : DFF_X1 port map( D => n8305, CK => CLK, Q => 
                           n_1746, QN => n15054);
   REGISTERS_reg_52_22_inst : DFF_X1 port map( D => n8304, CK => CLK, Q => 
                           n_1747, QN => n15055);
   REGISTERS_reg_52_21_inst : DFF_X1 port map( D => n8303, CK => CLK, Q => 
                           n_1748, QN => n15056);
   REGISTERS_reg_52_20_inst : DFF_X1 port map( D => n8302, CK => CLK, Q => 
                           n_1749, QN => n15057);
   REGISTERS_reg_52_19_inst : DFF_X1 port map( D => n8301, CK => CLK, Q => 
                           n_1750, QN => n15058);
   REGISTERS_reg_52_18_inst : DFF_X1 port map( D => n8300, CK => CLK, Q => 
                           n_1751, QN => n15059);
   REGISTERS_reg_52_17_inst : DFF_X1 port map( D => n8299, CK => CLK, Q => 
                           n_1752, QN => n15060);
   REGISTERS_reg_52_16_inst : DFF_X1 port map( D => n8298, CK => CLK, Q => 
                           n_1753, QN => n15061);
   REGISTERS_reg_52_15_inst : DFF_X1 port map( D => n8297, CK => CLK, Q => 
                           n_1754, QN => n15062);
   REGISTERS_reg_52_14_inst : DFF_X1 port map( D => n8296, CK => CLK, Q => 
                           n_1755, QN => n15063);
   REGISTERS_reg_52_13_inst : DFF_X1 port map( D => n8295, CK => CLK, Q => 
                           n_1756, QN => n15064);
   REGISTERS_reg_52_12_inst : DFF_X1 port map( D => n8294, CK => CLK, Q => 
                           n_1757, QN => n15065);
   REGISTERS_reg_52_11_inst : DFF_X1 port map( D => n8293, CK => CLK, Q => 
                           n_1758, QN => n15066);
   REGISTERS_reg_52_10_inst : DFF_X1 port map( D => n8292, CK => CLK, Q => 
                           n_1759, QN => n15067);
   REGISTERS_reg_52_9_inst : DFF_X1 port map( D => n8291, CK => CLK, Q => 
                           n_1760, QN => n15068);
   REGISTERS_reg_52_8_inst : DFF_X1 port map( D => n8290, CK => CLK, Q => 
                           n_1761, QN => n15069);
   REGISTERS_reg_52_7_inst : DFF_X1 port map( D => n8289, CK => CLK, Q => 
                           n_1762, QN => n15070);
   REGISTERS_reg_52_6_inst : DFF_X1 port map( D => n8288, CK => CLK, Q => 
                           n_1763, QN => n15071);
   REGISTERS_reg_52_5_inst : DFF_X1 port map( D => n8287, CK => CLK, Q => 
                           n_1764, QN => n15072);
   REGISTERS_reg_52_4_inst : DFF_X1 port map( D => n8286, CK => CLK, Q => 
                           n_1765, QN => n15073);
   REGISTERS_reg_52_3_inst : DFF_X1 port map( D => n8285, CK => CLK, Q => 
                           n_1766, QN => n15074);
   REGISTERS_reg_52_2_inst : DFF_X1 port map( D => n8284, CK => CLK, Q => 
                           n_1767, QN => n15075);
   REGISTERS_reg_52_1_inst : DFF_X1 port map( D => n8283, CK => CLK, Q => 
                           n_1768, QN => n15076);
   REGISTERS_reg_52_0_inst : DFF_X1 port map( D => n8282, CK => CLK, Q => 
                           n_1769, QN => n15077);
   REGISTERS_reg_53_31_inst : DFF_X1 port map( D => n8281, CK => CLK, Q => 
                           n_1770, QN => n15078);
   REGISTERS_reg_53_30_inst : DFF_X1 port map( D => n8280, CK => CLK, Q => 
                           n_1771, QN => n15079);
   REGISTERS_reg_53_29_inst : DFF_X1 port map( D => n8279, CK => CLK, Q => 
                           n_1772, QN => n15080);
   REGISTERS_reg_53_28_inst : DFF_X1 port map( D => n8278, CK => CLK, Q => 
                           n_1773, QN => n15081);
   REGISTERS_reg_53_27_inst : DFF_X1 port map( D => n8277, CK => CLK, Q => 
                           n_1774, QN => n15082);
   REGISTERS_reg_53_26_inst : DFF_X1 port map( D => n8276, CK => CLK, Q => 
                           n_1775, QN => n15083);
   REGISTERS_reg_53_25_inst : DFF_X1 port map( D => n8275, CK => CLK, Q => 
                           n_1776, QN => n15084);
   REGISTERS_reg_53_24_inst : DFF_X1 port map( D => n8274, CK => CLK, Q => 
                           n_1777, QN => n15085);
   REGISTERS_reg_53_23_inst : DFF_X1 port map( D => n8273, CK => CLK, Q => 
                           n_1778, QN => n15086);
   REGISTERS_reg_53_22_inst : DFF_X1 port map( D => n8272, CK => CLK, Q => 
                           n_1779, QN => n15087);
   REGISTERS_reg_53_21_inst : DFF_X1 port map( D => n8271, CK => CLK, Q => 
                           n_1780, QN => n15088);
   REGISTERS_reg_53_20_inst : DFF_X1 port map( D => n8270, CK => CLK, Q => 
                           n_1781, QN => n15089);
   REGISTERS_reg_53_19_inst : DFF_X1 port map( D => n8269, CK => CLK, Q => 
                           n_1782, QN => n15090);
   REGISTERS_reg_53_18_inst : DFF_X1 port map( D => n8268, CK => CLK, Q => 
                           n_1783, QN => n15091);
   REGISTERS_reg_53_17_inst : DFF_X1 port map( D => n8267, CK => CLK, Q => 
                           n_1784, QN => n15092);
   REGISTERS_reg_53_16_inst : DFF_X1 port map( D => n8266, CK => CLK, Q => 
                           n_1785, QN => n15093);
   REGISTERS_reg_53_15_inst : DFF_X1 port map( D => n8265, CK => CLK, Q => 
                           n_1786, QN => n15094);
   REGISTERS_reg_53_14_inst : DFF_X1 port map( D => n8264, CK => CLK, Q => 
                           n_1787, QN => n15095);
   REGISTERS_reg_53_13_inst : DFF_X1 port map( D => n8263, CK => CLK, Q => 
                           n_1788, QN => n15096);
   REGISTERS_reg_53_12_inst : DFF_X1 port map( D => n8262, CK => CLK, Q => 
                           n_1789, QN => n15097);
   REGISTERS_reg_53_11_inst : DFF_X1 port map( D => n8261, CK => CLK, Q => 
                           n_1790, QN => n15098);
   REGISTERS_reg_53_10_inst : DFF_X1 port map( D => n8260, CK => CLK, Q => 
                           n_1791, QN => n15099);
   REGISTERS_reg_53_9_inst : DFF_X1 port map( D => n8259, CK => CLK, Q => 
                           n_1792, QN => n15100);
   REGISTERS_reg_53_8_inst : DFF_X1 port map( D => n8258, CK => CLK, Q => 
                           n_1793, QN => n15101);
   REGISTERS_reg_53_7_inst : DFF_X1 port map( D => n8257, CK => CLK, Q => 
                           n_1794, QN => n15102);
   REGISTERS_reg_53_6_inst : DFF_X1 port map( D => n8256, CK => CLK, Q => 
                           n_1795, QN => n15103);
   REGISTERS_reg_53_5_inst : DFF_X1 port map( D => n8255, CK => CLK, Q => 
                           n_1796, QN => n15104);
   REGISTERS_reg_53_4_inst : DFF_X1 port map( D => n8254, CK => CLK, Q => 
                           n_1797, QN => n15105);
   REGISTERS_reg_53_3_inst : DFF_X1 port map( D => n8253, CK => CLK, Q => 
                           n_1798, QN => n15106);
   REGISTERS_reg_53_2_inst : DFF_X1 port map( D => n8252, CK => CLK, Q => 
                           n_1799, QN => n15107);
   REGISTERS_reg_53_1_inst : DFF_X1 port map( D => n8251, CK => CLK, Q => 
                           n_1800, QN => n15108);
   REGISTERS_reg_53_0_inst : DFF_X1 port map( D => n8250, CK => CLK, Q => 
                           n_1801, QN => n15109);
   REGISTERS_reg_54_31_inst : DFF_X1 port map( D => n8249, CK => CLK, Q => 
                           n_1802, QN => n15110);
   REGISTERS_reg_54_30_inst : DFF_X1 port map( D => n8248, CK => CLK, Q => 
                           n_1803, QN => n15111);
   REGISTERS_reg_54_29_inst : DFF_X1 port map( D => n8247, CK => CLK, Q => 
                           n_1804, QN => n15112);
   REGISTERS_reg_54_28_inst : DFF_X1 port map( D => n8246, CK => CLK, Q => 
                           n_1805, QN => n15113);
   REGISTERS_reg_54_27_inst : DFF_X1 port map( D => n8245, CK => CLK, Q => 
                           n_1806, QN => n15114);
   REGISTERS_reg_54_26_inst : DFF_X1 port map( D => n8244, CK => CLK, Q => 
                           n_1807, QN => n15115);
   REGISTERS_reg_54_25_inst : DFF_X1 port map( D => n8243, CK => CLK, Q => 
                           n_1808, QN => n15116);
   REGISTERS_reg_54_24_inst : DFF_X1 port map( D => n8242, CK => CLK, Q => 
                           n_1809, QN => n15117);
   REGISTERS_reg_54_23_inst : DFF_X1 port map( D => n8241, CK => CLK, Q => 
                           n_1810, QN => n15118);
   REGISTERS_reg_54_22_inst : DFF_X1 port map( D => n8240, CK => CLK, Q => 
                           n_1811, QN => n15119);
   REGISTERS_reg_54_21_inst : DFF_X1 port map( D => n8239, CK => CLK, Q => 
                           n_1812, QN => n15120);
   REGISTERS_reg_54_20_inst : DFF_X1 port map( D => n8238, CK => CLK, Q => 
                           n_1813, QN => n15121);
   REGISTERS_reg_54_19_inst : DFF_X1 port map( D => n8237, CK => CLK, Q => 
                           n_1814, QN => n15122);
   REGISTERS_reg_54_18_inst : DFF_X1 port map( D => n8236, CK => CLK, Q => 
                           n_1815, QN => n15123);
   REGISTERS_reg_54_17_inst : DFF_X1 port map( D => n8235, CK => CLK, Q => 
                           n_1816, QN => n15124);
   REGISTERS_reg_54_16_inst : DFF_X1 port map( D => n8234, CK => CLK, Q => 
                           n_1817, QN => n15125);
   REGISTERS_reg_54_15_inst : DFF_X1 port map( D => n8233, CK => CLK, Q => 
                           n_1818, QN => n15126);
   REGISTERS_reg_54_14_inst : DFF_X1 port map( D => n8232, CK => CLK, Q => 
                           n_1819, QN => n15127);
   REGISTERS_reg_54_13_inst : DFF_X1 port map( D => n8231, CK => CLK, Q => 
                           n_1820, QN => n15128);
   REGISTERS_reg_54_12_inst : DFF_X1 port map( D => n8230, CK => CLK, Q => 
                           n_1821, QN => n15129);
   REGISTERS_reg_54_11_inst : DFF_X1 port map( D => n8229, CK => CLK, Q => 
                           n_1822, QN => n15130);
   REGISTERS_reg_54_10_inst : DFF_X1 port map( D => n8228, CK => CLK, Q => 
                           n_1823, QN => n15131);
   REGISTERS_reg_54_9_inst : DFF_X1 port map( D => n8227, CK => CLK, Q => 
                           n_1824, QN => n15132);
   REGISTERS_reg_54_8_inst : DFF_X1 port map( D => n8226, CK => CLK, Q => 
                           n_1825, QN => n15133);
   REGISTERS_reg_54_7_inst : DFF_X1 port map( D => n8225, CK => CLK, Q => 
                           n_1826, QN => n15134);
   REGISTERS_reg_54_6_inst : DFF_X1 port map( D => n8224, CK => CLK, Q => 
                           n_1827, QN => n15135);
   REGISTERS_reg_54_5_inst : DFF_X1 port map( D => n8223, CK => CLK, Q => 
                           n_1828, QN => n15136);
   REGISTERS_reg_54_4_inst : DFF_X1 port map( D => n8222, CK => CLK, Q => 
                           n_1829, QN => n15137);
   REGISTERS_reg_54_3_inst : DFF_X1 port map( D => n8221, CK => CLK, Q => 
                           n_1830, QN => n15138);
   REGISTERS_reg_54_2_inst : DFF_X1 port map( D => n8220, CK => CLK, Q => 
                           n_1831, QN => n15139);
   REGISTERS_reg_54_1_inst : DFF_X1 port map( D => n8219, CK => CLK, Q => 
                           n_1832, QN => n15140);
   REGISTERS_reg_54_0_inst : DFF_X1 port map( D => n8218, CK => CLK, Q => 
                           n_1833, QN => n15141);
   REGISTERS_reg_55_31_inst : DFF_X1 port map( D => n8217, CK => CLK, Q => 
                           n_1834, QN => n15142);
   REGISTERS_reg_55_30_inst : DFF_X1 port map( D => n8216, CK => CLK, Q => 
                           n_1835, QN => n15143);
   REGISTERS_reg_55_29_inst : DFF_X1 port map( D => n8215, CK => CLK, Q => 
                           n_1836, QN => n15144);
   REGISTERS_reg_55_28_inst : DFF_X1 port map( D => n8214, CK => CLK, Q => 
                           n_1837, QN => n15145);
   REGISTERS_reg_55_27_inst : DFF_X1 port map( D => n8213, CK => CLK, Q => 
                           n_1838, QN => n15146);
   REGISTERS_reg_55_26_inst : DFF_X1 port map( D => n8212, CK => CLK, Q => 
                           n_1839, QN => n15147);
   REGISTERS_reg_55_25_inst : DFF_X1 port map( D => n8211, CK => CLK, Q => 
                           n_1840, QN => n15148);
   REGISTERS_reg_55_24_inst : DFF_X1 port map( D => n8210, CK => CLK, Q => 
                           n_1841, QN => n15149);
   REGISTERS_reg_55_23_inst : DFF_X1 port map( D => n8209, CK => CLK, Q => 
                           n_1842, QN => n15150);
   REGISTERS_reg_55_22_inst : DFF_X1 port map( D => n8208, CK => CLK, Q => 
                           n_1843, QN => n15151);
   REGISTERS_reg_55_21_inst : DFF_X1 port map( D => n8207, CK => CLK, Q => 
                           n_1844, QN => n15152);
   REGISTERS_reg_55_20_inst : DFF_X1 port map( D => n8206, CK => CLK, Q => 
                           n_1845, QN => n15153);
   REGISTERS_reg_55_19_inst : DFF_X1 port map( D => n8205, CK => CLK, Q => 
                           n_1846, QN => n15154);
   REGISTERS_reg_55_18_inst : DFF_X1 port map( D => n8204, CK => CLK, Q => 
                           n_1847, QN => n15155);
   REGISTERS_reg_55_17_inst : DFF_X1 port map( D => n8203, CK => CLK, Q => 
                           n_1848, QN => n15156);
   REGISTERS_reg_55_16_inst : DFF_X1 port map( D => n8202, CK => CLK, Q => 
                           n_1849, QN => n15157);
   REGISTERS_reg_55_15_inst : DFF_X1 port map( D => n8201, CK => CLK, Q => 
                           n_1850, QN => n15158);
   REGISTERS_reg_55_14_inst : DFF_X1 port map( D => n8200, CK => CLK, Q => 
                           n_1851, QN => n15159);
   REGISTERS_reg_55_13_inst : DFF_X1 port map( D => n8199, CK => CLK, Q => 
                           n_1852, QN => n15160);
   REGISTERS_reg_55_12_inst : DFF_X1 port map( D => n8198, CK => CLK, Q => 
                           n_1853, QN => n15161);
   REGISTERS_reg_55_11_inst : DFF_X1 port map( D => n8197, CK => CLK, Q => 
                           n_1854, QN => n15162);
   REGISTERS_reg_55_10_inst : DFF_X1 port map( D => n8196, CK => CLK, Q => 
                           n_1855, QN => n15163);
   REGISTERS_reg_55_9_inst : DFF_X1 port map( D => n8195, CK => CLK, Q => 
                           n_1856, QN => n15164);
   REGISTERS_reg_55_8_inst : DFF_X1 port map( D => n8194, CK => CLK, Q => 
                           n_1857, QN => n15165);
   REGISTERS_reg_55_7_inst : DFF_X1 port map( D => n8193, CK => CLK, Q => 
                           n_1858, QN => n15166);
   REGISTERS_reg_55_6_inst : DFF_X1 port map( D => n8192, CK => CLK, Q => 
                           n_1859, QN => n15167);
   REGISTERS_reg_55_5_inst : DFF_X1 port map( D => n8191, CK => CLK, Q => 
                           n_1860, QN => n15168);
   REGISTERS_reg_55_4_inst : DFF_X1 port map( D => n8190, CK => CLK, Q => 
                           n_1861, QN => n15169);
   REGISTERS_reg_55_3_inst : DFF_X1 port map( D => n8189, CK => CLK, Q => 
                           n_1862, QN => n15170);
   REGISTERS_reg_55_2_inst : DFF_X1 port map( D => n8188, CK => CLK, Q => 
                           n_1863, QN => n15171);
   REGISTERS_reg_55_1_inst : DFF_X1 port map( D => n8187, CK => CLK, Q => 
                           n_1864, QN => n15172);
   REGISTERS_reg_55_0_inst : DFF_X1 port map( D => n8186, CK => CLK, Q => 
                           n_1865, QN => n15173);
   REGISTERS_reg_56_31_inst : DFF_X1 port map( D => n8185, CK => CLK, Q => 
                           n6081, QN => n12725);
   REGISTERS_reg_56_30_inst : DFF_X1 port map( D => n8184, CK => CLK, Q => 
                           n6080, QN => n12724);
   REGISTERS_reg_56_29_inst : DFF_X1 port map( D => n8183, CK => CLK, Q => 
                           n6079, QN => n12723);
   REGISTERS_reg_56_28_inst : DFF_X1 port map( D => n8182, CK => CLK, Q => 
                           n6078, QN => n12722);
   REGISTERS_reg_56_27_inst : DFF_X1 port map( D => n8181, CK => CLK, Q => 
                           n6077, QN => n12721);
   REGISTERS_reg_56_26_inst : DFF_X1 port map( D => n8180, CK => CLK, Q => 
                           n6076, QN => n12720);
   REGISTERS_reg_56_25_inst : DFF_X1 port map( D => n8179, CK => CLK, Q => 
                           n6075, QN => n12719);
   REGISTERS_reg_56_24_inst : DFF_X1 port map( D => n8178, CK => CLK, Q => 
                           n6074, QN => n12718);
   REGISTERS_reg_56_23_inst : DFF_X1 port map( D => n8177, CK => CLK, Q => 
                           n6073, QN => n12773);
   REGISTERS_reg_56_22_inst : DFF_X1 port map( D => n8176, CK => CLK, Q => 
                           n6072, QN => n12772);
   REGISTERS_reg_56_21_inst : DFF_X1 port map( D => n8175, CK => CLK, Q => 
                           n6071, QN => n12771);
   REGISTERS_reg_56_20_inst : DFF_X1 port map( D => n8174, CK => CLK, Q => 
                           n6070, QN => n12770);
   REGISTERS_reg_56_19_inst : DFF_X1 port map( D => n8173, CK => CLK, Q => 
                           n6069, QN => n12769);
   REGISTERS_reg_56_18_inst : DFF_X1 port map( D => n8172, CK => CLK, Q => 
                           n6068, QN => n12768);
   REGISTERS_reg_56_17_inst : DFF_X1 port map( D => n8171, CK => CLK, Q => 
                           n6067, QN => n12767);
   REGISTERS_reg_56_16_inst : DFF_X1 port map( D => n8170, CK => CLK, Q => 
                           n6066, QN => n12766);
   REGISTERS_reg_56_15_inst : DFF_X1 port map( D => n8169, CK => CLK, Q => 
                           n6065, QN => n12765);
   REGISTERS_reg_56_14_inst : DFF_X1 port map( D => n8168, CK => CLK, Q => 
                           n6064, QN => n12764);
   REGISTERS_reg_56_13_inst : DFF_X1 port map( D => n8167, CK => CLK, Q => 
                           n6063, QN => n12763);
   REGISTERS_reg_56_12_inst : DFF_X1 port map( D => n8166, CK => CLK, Q => 
                           n6062, QN => n12762);
   REGISTERS_reg_56_11_inst : DFF_X1 port map( D => n8165, CK => CLK, Q => 
                           n6061, QN => n12761);
   REGISTERS_reg_56_10_inst : DFF_X1 port map( D => n8164, CK => CLK, Q => 
                           n6060, QN => n12760);
   REGISTERS_reg_56_9_inst : DFF_X1 port map( D => n8163, CK => CLK, Q => n6059
                           , QN => n12759);
   REGISTERS_reg_56_8_inst : DFF_X1 port map( D => n8162, CK => CLK, Q => n6058
                           , QN => n12758);
   REGISTERS_reg_56_7_inst : DFF_X1 port map( D => n8161, CK => CLK, Q => n6057
                           , QN => n12757);
   REGISTERS_reg_56_6_inst : DFF_X1 port map( D => n8160, CK => CLK, Q => n6056
                           , QN => n12756);
   REGISTERS_reg_56_5_inst : DFF_X1 port map( D => n8159, CK => CLK, Q => n6055
                           , QN => n12755);
   REGISTERS_reg_56_4_inst : DFF_X1 port map( D => n8158, CK => CLK, Q => n6054
                           , QN => n12754);
   REGISTERS_reg_56_3_inst : DFF_X1 port map( D => n8157, CK => CLK, Q => n6053
                           , QN => n12753);
   REGISTERS_reg_56_2_inst : DFF_X1 port map( D => n8156, CK => CLK, Q => n6052
                           , QN => n12752);
   REGISTERS_reg_56_1_inst : DFF_X1 port map( D => n8155, CK => CLK, Q => n6051
                           , QN => n12751);
   REGISTERS_reg_56_0_inst : DFF_X1 port map( D => n8154, CK => CLK, Q => n6050
                           , QN => n12750);
   REGISTERS_reg_57_31_inst : DFF_X1 port map( D => n8153, CK => CLK, Q => 
                           n6049, QN => n12717);
   REGISTERS_reg_57_30_inst : DFF_X1 port map( D => n8152, CK => CLK, Q => 
                           n6048, QN => n12716);
   REGISTERS_reg_57_29_inst : DFF_X1 port map( D => n8151, CK => CLK, Q => 
                           n6047, QN => n12715);
   REGISTERS_reg_57_28_inst : DFF_X1 port map( D => n8150, CK => CLK, Q => 
                           n6046, QN => n12714);
   REGISTERS_reg_57_27_inst : DFF_X1 port map( D => n8149, CK => CLK, Q => 
                           n6045, QN => n12713);
   REGISTERS_reg_57_26_inst : DFF_X1 port map( D => n8148, CK => CLK, Q => 
                           n6044, QN => n12712);
   REGISTERS_reg_57_25_inst : DFF_X1 port map( D => n8147, CK => CLK, Q => 
                           n6043, QN => n12711);
   REGISTERS_reg_57_24_inst : DFF_X1 port map( D => n8146, CK => CLK, Q => 
                           n6042, QN => n12710);
   REGISTERS_reg_57_23_inst : DFF_X1 port map( D => n8145, CK => CLK, Q => 
                           n6041, QN => n12749);
   REGISTERS_reg_57_22_inst : DFF_X1 port map( D => n8144, CK => CLK, Q => 
                           n6040, QN => n12748);
   REGISTERS_reg_57_21_inst : DFF_X1 port map( D => n8143, CK => CLK, Q => 
                           n6039, QN => n12747);
   REGISTERS_reg_57_20_inst : DFF_X1 port map( D => n8142, CK => CLK, Q => 
                           n6038, QN => n12746);
   REGISTERS_reg_57_19_inst : DFF_X1 port map( D => n8141, CK => CLK, Q => 
                           n6037, QN => n12745);
   REGISTERS_reg_57_18_inst : DFF_X1 port map( D => n8140, CK => CLK, Q => 
                           n6036, QN => n12744);
   REGISTERS_reg_57_17_inst : DFF_X1 port map( D => n8139, CK => CLK, Q => 
                           n6035, QN => n12743);
   REGISTERS_reg_57_16_inst : DFF_X1 port map( D => n8138, CK => CLK, Q => 
                           n6034, QN => n12742);
   REGISTERS_reg_57_15_inst : DFF_X1 port map( D => n8137, CK => CLK, Q => 
                           n6033, QN => n12741);
   REGISTERS_reg_57_14_inst : DFF_X1 port map( D => n8136, CK => CLK, Q => 
                           n6032, QN => n12740);
   REGISTERS_reg_57_13_inst : DFF_X1 port map( D => n8135, CK => CLK, Q => 
                           n6031, QN => n12739);
   REGISTERS_reg_57_12_inst : DFF_X1 port map( D => n8134, CK => CLK, Q => 
                           n6030, QN => n12738);
   REGISTERS_reg_57_11_inst : DFF_X1 port map( D => n8133, CK => CLK, Q => 
                           n6029, QN => n12737);
   REGISTERS_reg_57_10_inst : DFF_X1 port map( D => n8132, CK => CLK, Q => 
                           n6028, QN => n12736);
   REGISTERS_reg_57_9_inst : DFF_X1 port map( D => n8131, CK => CLK, Q => n6027
                           , QN => n12735);
   REGISTERS_reg_57_8_inst : DFF_X1 port map( D => n8130, CK => CLK, Q => n6026
                           , QN => n12734);
   REGISTERS_reg_57_7_inst : DFF_X1 port map( D => n8129, CK => CLK, Q => n6025
                           , QN => n12733);
   REGISTERS_reg_57_6_inst : DFF_X1 port map( D => n8128, CK => CLK, Q => n6024
                           , QN => n12732);
   REGISTERS_reg_57_5_inst : DFF_X1 port map( D => n8127, CK => CLK, Q => n6023
                           , QN => n12731);
   REGISTERS_reg_57_4_inst : DFF_X1 port map( D => n8126, CK => CLK, Q => n6022
                           , QN => n12730);
   REGISTERS_reg_57_3_inst : DFF_X1 port map( D => n8125, CK => CLK, Q => n6021
                           , QN => n12729);
   REGISTERS_reg_57_2_inst : DFF_X1 port map( D => n8124, CK => CLK, Q => n6020
                           , QN => n12728);
   REGISTERS_reg_57_1_inst : DFF_X1 port map( D => n8123, CK => CLK, Q => n6019
                           , QN => n12727);
   REGISTERS_reg_57_0_inst : DFF_X1 port map( D => n8122, CK => CLK, Q => n6018
                           , QN => n12726);
   REGISTERS_reg_59_31_inst : DFF_X1 port map( D => n8089, CK => CLK, Q => 
                           n5985, QN => n12837);
   REGISTERS_reg_59_30_inst : DFF_X1 port map( D => n8088, CK => CLK, Q => 
                           n5984, QN => n12836);
   REGISTERS_reg_59_29_inst : DFF_X1 port map( D => n8087, CK => CLK, Q => 
                           n5983, QN => n12835);
   REGISTERS_reg_59_28_inst : DFF_X1 port map( D => n8086, CK => CLK, Q => 
                           n5982, QN => n12834);
   REGISTERS_reg_59_27_inst : DFF_X1 port map( D => n8085, CK => CLK, Q => 
                           n5981, QN => n12833);
   REGISTERS_reg_59_26_inst : DFF_X1 port map( D => n8084, CK => CLK, Q => 
                           n5980, QN => n12832);
   REGISTERS_reg_59_25_inst : DFF_X1 port map( D => n8083, CK => CLK, Q => 
                           n5979, QN => n12831);
   REGISTERS_reg_59_24_inst : DFF_X1 port map( D => n8082, CK => CLK, Q => 
                           n5978, QN => n12830);
   REGISTERS_reg_59_23_inst : DFF_X1 port map( D => n8081, CK => CLK, Q => 
                           n5977, QN => n12829);
   REGISTERS_reg_59_22_inst : DFF_X1 port map( D => n8080, CK => CLK, Q => 
                           n5976, QN => n12828);
   REGISTERS_reg_59_21_inst : DFF_X1 port map( D => n8079, CK => CLK, Q => 
                           n5975, QN => n12827);
   REGISTERS_reg_59_20_inst : DFF_X1 port map( D => n8078, CK => CLK, Q => 
                           n5974, QN => n12826);
   REGISTERS_reg_59_19_inst : DFF_X1 port map( D => n8077, CK => CLK, Q => 
                           n5973, QN => n12825);
   REGISTERS_reg_59_18_inst : DFF_X1 port map( D => n8076, CK => CLK, Q => 
                           n5972, QN => n12824);
   REGISTERS_reg_59_17_inst : DFF_X1 port map( D => n8075, CK => CLK, Q => 
                           n5971, QN => n12823);
   REGISTERS_reg_59_16_inst : DFF_X1 port map( D => n8074, CK => CLK, Q => 
                           n5970, QN => n12822);
   REGISTERS_reg_59_15_inst : DFF_X1 port map( D => n8073, CK => CLK, Q => 
                           n5969, QN => n12821);
   REGISTERS_reg_59_14_inst : DFF_X1 port map( D => n8072, CK => CLK, Q => 
                           n5968, QN => n12820);
   REGISTERS_reg_59_13_inst : DFF_X1 port map( D => n8071, CK => CLK, Q => 
                           n5967, QN => n12819);
   REGISTERS_reg_59_12_inst : DFF_X1 port map( D => n8070, CK => CLK, Q => 
                           n5966, QN => n12818);
   REGISTERS_reg_59_11_inst : DFF_X1 port map( D => n8069, CK => CLK, Q => 
                           n5965, QN => n12817);
   REGISTERS_reg_59_10_inst : DFF_X1 port map( D => n8068, CK => CLK, Q => 
                           n5964, QN => n12816);
   REGISTERS_reg_59_9_inst : DFF_X1 port map( D => n8067, CK => CLK, Q => n5963
                           , QN => n12815);
   REGISTERS_reg_59_8_inst : DFF_X1 port map( D => n8066, CK => CLK, Q => n5962
                           , QN => n12814);
   REGISTERS_reg_59_7_inst : DFF_X1 port map( D => n8065, CK => CLK, Q => n5961
                           , QN => n12813);
   REGISTERS_reg_59_6_inst : DFF_X1 port map( D => n8064, CK => CLK, Q => n5960
                           , QN => n12812);
   REGISTERS_reg_59_5_inst : DFF_X1 port map( D => n8063, CK => CLK, Q => n5959
                           , QN => n12811);
   REGISTERS_reg_59_4_inst : DFF_X1 port map( D => n8062, CK => CLK, Q => n5958
                           , QN => n12810);
   REGISTERS_reg_59_3_inst : DFF_X1 port map( D => n8061, CK => CLK, Q => n5957
                           , QN => n12809);
   REGISTERS_reg_59_2_inst : DFF_X1 port map( D => n8060, CK => CLK, Q => n5956
                           , QN => n12808);
   REGISTERS_reg_59_1_inst : DFF_X1 port map( D => n8059, CK => CLK, Q => n5955
                           , QN => n12807);
   REGISTERS_reg_59_0_inst : DFF_X1 port map( D => n8058, CK => CLK, Q => n5954
                           , QN => n12806);
   REGISTERS_reg_60_31_inst : DFF_X1 port map( D => n8057, CK => CLK, Q => 
                           n_1866, QN => n15206);
   REGISTERS_reg_60_30_inst : DFF_X1 port map( D => n8056, CK => CLK, Q => 
                           n_1867, QN => n15207);
   REGISTERS_reg_60_29_inst : DFF_X1 port map( D => n8055, CK => CLK, Q => 
                           n_1868, QN => n15208);
   REGISTERS_reg_60_28_inst : DFF_X1 port map( D => n8054, CK => CLK, Q => 
                           n_1869, QN => n15209);
   REGISTERS_reg_60_27_inst : DFF_X1 port map( D => n8053, CK => CLK, Q => 
                           n_1870, QN => n15210);
   REGISTERS_reg_60_26_inst : DFF_X1 port map( D => n8052, CK => CLK, Q => 
                           n_1871, QN => n15211);
   REGISTERS_reg_60_25_inst : DFF_X1 port map( D => n8051, CK => CLK, Q => 
                           n_1872, QN => n15212);
   REGISTERS_reg_60_24_inst : DFF_X1 port map( D => n8050, CK => CLK, Q => 
                           n_1873, QN => n15213);
   REGISTERS_reg_60_23_inst : DFF_X1 port map( D => n8049, CK => CLK, Q => 
                           n_1874, QN => n15214);
   REGISTERS_reg_60_22_inst : DFF_X1 port map( D => n8048, CK => CLK, Q => 
                           n_1875, QN => n15215);
   REGISTERS_reg_60_21_inst : DFF_X1 port map( D => n8047, CK => CLK, Q => 
                           n_1876, QN => n15216);
   REGISTERS_reg_60_20_inst : DFF_X1 port map( D => n8046, CK => CLK, Q => 
                           n_1877, QN => n15217);
   REGISTERS_reg_60_19_inst : DFF_X1 port map( D => n8045, CK => CLK, Q => 
                           n_1878, QN => n15218);
   REGISTERS_reg_60_18_inst : DFF_X1 port map( D => n8044, CK => CLK, Q => 
                           n_1879, QN => n15219);
   REGISTERS_reg_60_17_inst : DFF_X1 port map( D => n8043, CK => CLK, Q => 
                           n_1880, QN => n15220);
   REGISTERS_reg_60_16_inst : DFF_X1 port map( D => n8042, CK => CLK, Q => 
                           n_1881, QN => n15221);
   REGISTERS_reg_60_15_inst : DFF_X1 port map( D => n8041, CK => CLK, Q => 
                           n_1882, QN => n15222);
   REGISTERS_reg_60_14_inst : DFF_X1 port map( D => n8040, CK => CLK, Q => 
                           n_1883, QN => n15223);
   REGISTERS_reg_60_13_inst : DFF_X1 port map( D => n8039, CK => CLK, Q => 
                           n_1884, QN => n15224);
   REGISTERS_reg_60_12_inst : DFF_X1 port map( D => n8038, CK => CLK, Q => 
                           n_1885, QN => n15225);
   REGISTERS_reg_60_11_inst : DFF_X1 port map( D => n8037, CK => CLK, Q => 
                           n_1886, QN => n15226);
   REGISTERS_reg_60_10_inst : DFF_X1 port map( D => n8036, CK => CLK, Q => 
                           n_1887, QN => n15227);
   REGISTERS_reg_60_9_inst : DFF_X1 port map( D => n8035, CK => CLK, Q => 
                           n_1888, QN => n15228);
   REGISTERS_reg_60_8_inst : DFF_X1 port map( D => n8034, CK => CLK, Q => 
                           n_1889, QN => n15229);
   REGISTERS_reg_60_7_inst : DFF_X1 port map( D => n8033, CK => CLK, Q => 
                           n_1890, QN => n15230);
   REGISTERS_reg_60_6_inst : DFF_X1 port map( D => n8032, CK => CLK, Q => 
                           n_1891, QN => n15231);
   REGISTERS_reg_60_5_inst : DFF_X1 port map( D => n8031, CK => CLK, Q => 
                           n_1892, QN => n15232);
   REGISTERS_reg_60_4_inst : DFF_X1 port map( D => n8030, CK => CLK, Q => 
                           n_1893, QN => n15233);
   REGISTERS_reg_60_3_inst : DFF_X1 port map( D => n8029, CK => CLK, Q => 
                           n_1894, QN => n15234);
   REGISTERS_reg_60_2_inst : DFF_X1 port map( D => n8028, CK => CLK, Q => 
                           n_1895, QN => n15235);
   REGISTERS_reg_60_1_inst : DFF_X1 port map( D => n8027, CK => CLK, Q => 
                           n_1896, QN => n15236);
   REGISTERS_reg_60_0_inst : DFF_X1 port map( D => n8026, CK => CLK, Q => 
                           n_1897, QN => n15237);
   REGISTERS_reg_61_31_inst : DFF_X1 port map( D => n8025, CK => CLK, Q => 
                           n_1898, QN => n15238);
   REGISTERS_reg_61_30_inst : DFF_X1 port map( D => n8024, CK => CLK, Q => 
                           n_1899, QN => n15239);
   REGISTERS_reg_61_29_inst : DFF_X1 port map( D => n8023, CK => CLK, Q => 
                           n_1900, QN => n15240);
   REGISTERS_reg_61_28_inst : DFF_X1 port map( D => n8022, CK => CLK, Q => 
                           n_1901, QN => n15241);
   REGISTERS_reg_61_27_inst : DFF_X1 port map( D => n8021, CK => CLK, Q => 
                           n_1902, QN => n15242);
   REGISTERS_reg_61_26_inst : DFF_X1 port map( D => n8020, CK => CLK, Q => 
                           n_1903, QN => n15243);
   REGISTERS_reg_61_25_inst : DFF_X1 port map( D => n8019, CK => CLK, Q => 
                           n_1904, QN => n15244);
   REGISTERS_reg_61_24_inst : DFF_X1 port map( D => n8018, CK => CLK, Q => 
                           n_1905, QN => n15245);
   REGISTERS_reg_61_23_inst : DFF_X1 port map( D => n8017, CK => CLK, Q => 
                           n_1906, QN => n15246);
   REGISTERS_reg_61_22_inst : DFF_X1 port map( D => n8016, CK => CLK, Q => 
                           n_1907, QN => n15247);
   REGISTERS_reg_61_21_inst : DFF_X1 port map( D => n8015, CK => CLK, Q => 
                           n_1908, QN => n15248);
   REGISTERS_reg_61_20_inst : DFF_X1 port map( D => n8014, CK => CLK, Q => 
                           n_1909, QN => n15249);
   REGISTERS_reg_61_19_inst : DFF_X1 port map( D => n8013, CK => CLK, Q => 
                           n_1910, QN => n15250);
   REGISTERS_reg_61_18_inst : DFF_X1 port map( D => n8012, CK => CLK, Q => 
                           n_1911, QN => n15251);
   REGISTERS_reg_61_17_inst : DFF_X1 port map( D => n8011, CK => CLK, Q => 
                           n_1912, QN => n15252);
   REGISTERS_reg_61_16_inst : DFF_X1 port map( D => n8010, CK => CLK, Q => 
                           n_1913, QN => n15253);
   REGISTERS_reg_61_15_inst : DFF_X1 port map( D => n8009, CK => CLK, Q => 
                           n_1914, QN => n15254);
   REGISTERS_reg_61_14_inst : DFF_X1 port map( D => n8008, CK => CLK, Q => 
                           n_1915, QN => n15255);
   REGISTERS_reg_61_13_inst : DFF_X1 port map( D => n8007, CK => CLK, Q => 
                           n_1916, QN => n15256);
   REGISTERS_reg_61_12_inst : DFF_X1 port map( D => n8006, CK => CLK, Q => 
                           n_1917, QN => n15257);
   REGISTERS_reg_61_11_inst : DFF_X1 port map( D => n8005, CK => CLK, Q => 
                           n_1918, QN => n15258);
   REGISTERS_reg_61_10_inst : DFF_X1 port map( D => n8004, CK => CLK, Q => 
                           n_1919, QN => n15259);
   REGISTERS_reg_61_9_inst : DFF_X1 port map( D => n8003, CK => CLK, Q => 
                           n_1920, QN => n15260);
   REGISTERS_reg_61_8_inst : DFF_X1 port map( D => n8002, CK => CLK, Q => 
                           n_1921, QN => n15261);
   REGISTERS_reg_61_7_inst : DFF_X1 port map( D => n8001, CK => CLK, Q => 
                           n_1922, QN => n15262);
   REGISTERS_reg_61_6_inst : DFF_X1 port map( D => n8000, CK => CLK, Q => 
                           n_1923, QN => n15263);
   REGISTERS_reg_61_5_inst : DFF_X1 port map( D => n7999, CK => CLK, Q => 
                           n_1924, QN => n15264);
   REGISTERS_reg_61_4_inst : DFF_X1 port map( D => n7998, CK => CLK, Q => 
                           n_1925, QN => n15265);
   REGISTERS_reg_61_3_inst : DFF_X1 port map( D => n7997, CK => CLK, Q => 
                           n_1926, QN => n15266);
   REGISTERS_reg_61_2_inst : DFF_X1 port map( D => n7996, CK => CLK, Q => 
                           n_1927, QN => n15267);
   REGISTERS_reg_61_1_inst : DFF_X1 port map( D => n7995, CK => CLK, Q => 
                           n_1928, QN => n15268);
   REGISTERS_reg_61_0_inst : DFF_X1 port map( D => n7994, CK => CLK, Q => 
                           n_1929, QN => n15269);
   REGISTERS_reg_62_31_inst : DFF_X1 port map( D => n7993, CK => CLK, Q => 
                           n_1930, QN => n15270);
   REGISTERS_reg_62_30_inst : DFF_X1 port map( D => n7992, CK => CLK, Q => 
                           n_1931, QN => n15271);
   REGISTERS_reg_62_29_inst : DFF_X1 port map( D => n7991, CK => CLK, Q => 
                           n_1932, QN => n15272);
   REGISTERS_reg_62_28_inst : DFF_X1 port map( D => n7990, CK => CLK, Q => 
                           n_1933, QN => n15273);
   REGISTERS_reg_62_27_inst : DFF_X1 port map( D => n7989, CK => CLK, Q => 
                           n_1934, QN => n15274);
   REGISTERS_reg_62_26_inst : DFF_X1 port map( D => n7988, CK => CLK, Q => 
                           n_1935, QN => n15275);
   REGISTERS_reg_62_25_inst : DFF_X1 port map( D => n7987, CK => CLK, Q => 
                           n_1936, QN => n15276);
   REGISTERS_reg_62_24_inst : DFF_X1 port map( D => n7986, CK => CLK, Q => 
                           n_1937, QN => n15277);
   REGISTERS_reg_62_23_inst : DFF_X1 port map( D => n7985, CK => CLK, Q => 
                           n_1938, QN => n15278);
   REGISTERS_reg_62_22_inst : DFF_X1 port map( D => n7984, CK => CLK, Q => 
                           n_1939, QN => n15279);
   REGISTERS_reg_62_21_inst : DFF_X1 port map( D => n7983, CK => CLK, Q => 
                           n_1940, QN => n15280);
   REGISTERS_reg_62_20_inst : DFF_X1 port map( D => n7982, CK => CLK, Q => 
                           n_1941, QN => n15281);
   REGISTERS_reg_62_19_inst : DFF_X1 port map( D => n7981, CK => CLK, Q => 
                           n_1942, QN => n15282);
   REGISTERS_reg_62_18_inst : DFF_X1 port map( D => n7980, CK => CLK, Q => 
                           n_1943, QN => n15283);
   REGISTERS_reg_62_17_inst : DFF_X1 port map( D => n7979, CK => CLK, Q => 
                           n_1944, QN => n15284);
   REGISTERS_reg_62_16_inst : DFF_X1 port map( D => n7978, CK => CLK, Q => 
                           n_1945, QN => n15285);
   REGISTERS_reg_62_15_inst : DFF_X1 port map( D => n7977, CK => CLK, Q => 
                           n_1946, QN => n15286);
   REGISTERS_reg_62_14_inst : DFF_X1 port map( D => n7976, CK => CLK, Q => 
                           n_1947, QN => n15287);
   REGISTERS_reg_62_13_inst : DFF_X1 port map( D => n7975, CK => CLK, Q => 
                           n_1948, QN => n15288);
   REGISTERS_reg_62_12_inst : DFF_X1 port map( D => n7974, CK => CLK, Q => 
                           n_1949, QN => n15289);
   REGISTERS_reg_62_11_inst : DFF_X1 port map( D => n7973, CK => CLK, Q => 
                           n_1950, QN => n15290);
   REGISTERS_reg_62_10_inst : DFF_X1 port map( D => n7972, CK => CLK, Q => 
                           n_1951, QN => n15291);
   REGISTERS_reg_62_9_inst : DFF_X1 port map( D => n7971, CK => CLK, Q => 
                           n_1952, QN => n15292);
   REGISTERS_reg_62_8_inst : DFF_X1 port map( D => n7970, CK => CLK, Q => 
                           n_1953, QN => n15293);
   REGISTERS_reg_62_7_inst : DFF_X1 port map( D => n7969, CK => CLK, Q => 
                           n_1954, QN => n15294);
   REGISTERS_reg_62_6_inst : DFF_X1 port map( D => n7968, CK => CLK, Q => 
                           n_1955, QN => n15295);
   REGISTERS_reg_62_5_inst : DFF_X1 port map( D => n7967, CK => CLK, Q => 
                           n_1956, QN => n15296);
   REGISTERS_reg_62_4_inst : DFF_X1 port map( D => n7966, CK => CLK, Q => 
                           n_1957, QN => n15297);
   REGISTERS_reg_62_3_inst : DFF_X1 port map( D => n7965, CK => CLK, Q => 
                           n_1958, QN => n15298);
   REGISTERS_reg_62_2_inst : DFF_X1 port map( D => n7964, CK => CLK, Q => 
                           n_1959, QN => n15299);
   REGISTERS_reg_62_1_inst : DFF_X1 port map( D => n7963, CK => CLK, Q => 
                           n_1960, QN => n15300);
   REGISTERS_reg_62_0_inst : DFF_X1 port map( D => n7962, CK => CLK, Q => 
                           n_1961, QN => n15301);
   REGISTERS_reg_64_31_inst : DFF_X1 port map( D => n7929, CK => CLK, Q => 
                           n5921, QN => n12805);
   REGISTERS_reg_64_30_inst : DFF_X1 port map( D => n7928, CK => CLK, Q => 
                           n5920, QN => n12804);
   REGISTERS_reg_64_29_inst : DFF_X1 port map( D => n7927, CK => CLK, Q => 
                           n5919, QN => n12803);
   REGISTERS_reg_64_28_inst : DFF_X1 port map( D => n7926, CK => CLK, Q => 
                           n5918, QN => n12802);
   REGISTERS_reg_64_27_inst : DFF_X1 port map( D => n7925, CK => CLK, Q => 
                           n5917, QN => n12801);
   REGISTERS_reg_64_26_inst : DFF_X1 port map( D => n7924, CK => CLK, Q => 
                           n5916, QN => n12800);
   REGISTERS_reg_64_25_inst : DFF_X1 port map( D => n7923, CK => CLK, Q => 
                           n5915, QN => n12799);
   REGISTERS_reg_64_24_inst : DFF_X1 port map( D => n7922, CK => CLK, Q => 
                           n5914, QN => n12798);
   REGISTERS_reg_64_23_inst : DFF_X1 port map( D => n7921, CK => CLK, Q => 
                           n5913, QN => n12797);
   REGISTERS_reg_64_22_inst : DFF_X1 port map( D => n7920, CK => CLK, Q => 
                           n5912, QN => n12796);
   REGISTERS_reg_64_21_inst : DFF_X1 port map( D => n7919, CK => CLK, Q => 
                           n5911, QN => n12795);
   REGISTERS_reg_64_20_inst : DFF_X1 port map( D => n7918, CK => CLK, Q => 
                           n5910, QN => n12794);
   REGISTERS_reg_64_19_inst : DFF_X1 port map( D => n7917, CK => CLK, Q => 
                           n5909, QN => n12793);
   REGISTERS_reg_64_18_inst : DFF_X1 port map( D => n7916, CK => CLK, Q => 
                           n5908, QN => n12792);
   REGISTERS_reg_64_17_inst : DFF_X1 port map( D => n7915, CK => CLK, Q => 
                           n5907, QN => n12791);
   REGISTERS_reg_64_16_inst : DFF_X1 port map( D => n7914, CK => CLK, Q => 
                           n5906, QN => n12790);
   REGISTERS_reg_64_15_inst : DFF_X1 port map( D => n7913, CK => CLK, Q => 
                           n5905, QN => n12789);
   REGISTERS_reg_64_14_inst : DFF_X1 port map( D => n7912, CK => CLK, Q => 
                           n5904, QN => n12788);
   REGISTERS_reg_64_13_inst : DFF_X1 port map( D => n7911, CK => CLK, Q => 
                           n5903, QN => n12787);
   REGISTERS_reg_64_12_inst : DFF_X1 port map( D => n7910, CK => CLK, Q => 
                           n5902, QN => n12786);
   REGISTERS_reg_64_11_inst : DFF_X1 port map( D => n7909, CK => CLK, Q => 
                           n5901, QN => n12785);
   REGISTERS_reg_64_10_inst : DFF_X1 port map( D => n7908, CK => CLK, Q => 
                           n5900, QN => n12784);
   REGISTERS_reg_64_9_inst : DFF_X1 port map( D => n7907, CK => CLK, Q => n5899
                           , QN => n12783);
   REGISTERS_reg_64_8_inst : DFF_X1 port map( D => n7906, CK => CLK, Q => n5898
                           , QN => n12782);
   REGISTERS_reg_64_7_inst : DFF_X1 port map( D => n7905, CK => CLK, Q => n5897
                           , QN => n12781);
   REGISTERS_reg_64_6_inst : DFF_X1 port map( D => n7904, CK => CLK, Q => n5896
                           , QN => n12780);
   REGISTERS_reg_64_5_inst : DFF_X1 port map( D => n7903, CK => CLK, Q => n5895
                           , QN => n12779);
   REGISTERS_reg_64_4_inst : DFF_X1 port map( D => n7902, CK => CLK, Q => n5894
                           , QN => n12778);
   REGISTERS_reg_64_3_inst : DFF_X1 port map( D => n7901, CK => CLK, Q => n5893
                           , QN => n12777);
   REGISTERS_reg_64_2_inst : DFF_X1 port map( D => n7900, CK => CLK, Q => n5892
                           , QN => n12776);
   REGISTERS_reg_64_1_inst : DFF_X1 port map( D => n7899, CK => CLK, Q => n5891
                           , QN => n12775);
   REGISTERS_reg_64_0_inst : DFF_X1 port map( D => n7898, CK => CLK, Q => n5890
                           , QN => n12774);
   REGISTERS_reg_65_31_inst : DFF_X1 port map( D => n7897, CK => CLK, Q => 
                           n_1962, QN => n15334);
   REGISTERS_reg_65_30_inst : DFF_X1 port map( D => n7896, CK => CLK, Q => 
                           n_1963, QN => n15335);
   REGISTERS_reg_65_29_inst : DFF_X1 port map( D => n7895, CK => CLK, Q => 
                           n_1964, QN => n15336);
   REGISTERS_reg_65_28_inst : DFF_X1 port map( D => n7894, CK => CLK, Q => 
                           n_1965, QN => n15337);
   REGISTERS_reg_65_27_inst : DFF_X1 port map( D => n7893, CK => CLK, Q => 
                           n_1966, QN => n15338);
   REGISTERS_reg_65_26_inst : DFF_X1 port map( D => n7892, CK => CLK, Q => 
                           n_1967, QN => n15339);
   REGISTERS_reg_65_25_inst : DFF_X1 port map( D => n7891, CK => CLK, Q => 
                           n_1968, QN => n15340);
   REGISTERS_reg_65_24_inst : DFF_X1 port map( D => n7890, CK => CLK, Q => 
                           n_1969, QN => n15341);
   REGISTERS_reg_65_23_inst : DFF_X1 port map( D => n7889, CK => CLK, Q => 
                           n_1970, QN => n15342);
   REGISTERS_reg_65_22_inst : DFF_X1 port map( D => n7888, CK => CLK, Q => 
                           n_1971, QN => n15343);
   REGISTERS_reg_65_21_inst : DFF_X1 port map( D => n7887, CK => CLK, Q => 
                           n_1972, QN => n15344);
   REGISTERS_reg_65_20_inst : DFF_X1 port map( D => n7886, CK => CLK, Q => 
                           n_1973, QN => n15345);
   REGISTERS_reg_65_19_inst : DFF_X1 port map( D => n7885, CK => CLK, Q => 
                           n_1974, QN => n15346);
   REGISTERS_reg_65_18_inst : DFF_X1 port map( D => n7884, CK => CLK, Q => 
                           n_1975, QN => n15347);
   REGISTERS_reg_65_17_inst : DFF_X1 port map( D => n7883, CK => CLK, Q => 
                           n_1976, QN => n15348);
   REGISTERS_reg_65_16_inst : DFF_X1 port map( D => n7882, CK => CLK, Q => 
                           n_1977, QN => n15349);
   REGISTERS_reg_65_15_inst : DFF_X1 port map( D => n7881, CK => CLK, Q => 
                           n_1978, QN => n15350);
   REGISTERS_reg_65_14_inst : DFF_X1 port map( D => n7880, CK => CLK, Q => 
                           n_1979, QN => n15351);
   REGISTERS_reg_65_13_inst : DFF_X1 port map( D => n7879, CK => CLK, Q => 
                           n_1980, QN => n15352);
   REGISTERS_reg_65_12_inst : DFF_X1 port map( D => n7878, CK => CLK, Q => 
                           n_1981, QN => n15353);
   REGISTERS_reg_65_11_inst : DFF_X1 port map( D => n7877, CK => CLK, Q => 
                           n_1982, QN => n15354);
   REGISTERS_reg_65_10_inst : DFF_X1 port map( D => n7876, CK => CLK, Q => 
                           n_1983, QN => n15355);
   REGISTERS_reg_65_9_inst : DFF_X1 port map( D => n7875, CK => CLK, Q => 
                           n_1984, QN => n15356);
   REGISTERS_reg_65_8_inst : DFF_X1 port map( D => n7874, CK => CLK, Q => 
                           n_1985, QN => n15357);
   REGISTERS_reg_65_7_inst : DFF_X1 port map( D => n7873, CK => CLK, Q => 
                           n_1986, QN => n15358);
   REGISTERS_reg_65_6_inst : DFF_X1 port map( D => n7872, CK => CLK, Q => 
                           n_1987, QN => n15359);
   REGISTERS_reg_65_5_inst : DFF_X1 port map( D => n7871, CK => CLK, Q => 
                           n_1988, QN => n15360);
   REGISTERS_reg_65_4_inst : DFF_X1 port map( D => n7870, CK => CLK, Q => 
                           n_1989, QN => n15361);
   REGISTERS_reg_65_3_inst : DFF_X1 port map( D => n7869, CK => CLK, Q => 
                           n_1990, QN => n15362);
   REGISTERS_reg_65_2_inst : DFF_X1 port map( D => n7868, CK => CLK, Q => 
                           n_1991, QN => n15363);
   REGISTERS_reg_65_1_inst : DFF_X1 port map( D => n7867, CK => CLK, Q => 
                           n_1992, QN => n15364);
   REGISTERS_reg_65_0_inst : DFF_X1 port map( D => n7866, CK => CLK, Q => 
                           n_1993, QN => n15365);
   REGISTERS_reg_66_31_inst : DFF_X1 port map( D => n7865, CK => CLK, Q => 
                           n_1994, QN => n15366);
   REGISTERS_reg_66_30_inst : DFF_X1 port map( D => n7864, CK => CLK, Q => 
                           n_1995, QN => n15367);
   REGISTERS_reg_66_29_inst : DFF_X1 port map( D => n7863, CK => CLK, Q => 
                           n_1996, QN => n15368);
   REGISTERS_reg_66_28_inst : DFF_X1 port map( D => n7862, CK => CLK, Q => 
                           n_1997, QN => n15369);
   REGISTERS_reg_66_27_inst : DFF_X1 port map( D => n7861, CK => CLK, Q => 
                           n_1998, QN => n15370);
   REGISTERS_reg_66_26_inst : DFF_X1 port map( D => n7860, CK => CLK, Q => 
                           n_1999, QN => n15371);
   REGISTERS_reg_66_25_inst : DFF_X1 port map( D => n7859, CK => CLK, Q => 
                           n_2000, QN => n15372);
   REGISTERS_reg_66_24_inst : DFF_X1 port map( D => n7858, CK => CLK, Q => 
                           n_2001, QN => n15373);
   REGISTERS_reg_66_23_inst : DFF_X1 port map( D => n7857, CK => CLK, Q => 
                           n_2002, QN => n15374);
   REGISTERS_reg_66_22_inst : DFF_X1 port map( D => n7856, CK => CLK, Q => 
                           n_2003, QN => n15375);
   REGISTERS_reg_66_21_inst : DFF_X1 port map( D => n7855, CK => CLK, Q => 
                           n_2004, QN => n15376);
   REGISTERS_reg_66_20_inst : DFF_X1 port map( D => n7854, CK => CLK, Q => 
                           n_2005, QN => n15377);
   REGISTERS_reg_66_19_inst : DFF_X1 port map( D => n7853, CK => CLK, Q => 
                           n_2006, QN => n15378);
   REGISTERS_reg_66_18_inst : DFF_X1 port map( D => n7852, CK => CLK, Q => 
                           n_2007, QN => n15379);
   REGISTERS_reg_66_17_inst : DFF_X1 port map( D => n7851, CK => CLK, Q => 
                           n_2008, QN => n15380);
   REGISTERS_reg_66_16_inst : DFF_X1 port map( D => n7850, CK => CLK, Q => 
                           n_2009, QN => n15381);
   REGISTERS_reg_66_15_inst : DFF_X1 port map( D => n7849, CK => CLK, Q => 
                           n_2010, QN => n15382);
   REGISTERS_reg_66_14_inst : DFF_X1 port map( D => n7848, CK => CLK, Q => 
                           n_2011, QN => n15383);
   REGISTERS_reg_66_13_inst : DFF_X1 port map( D => n7847, CK => CLK, Q => 
                           n_2012, QN => n15384);
   REGISTERS_reg_66_12_inst : DFF_X1 port map( D => n7846, CK => CLK, Q => 
                           n_2013, QN => n15385);
   REGISTERS_reg_66_11_inst : DFF_X1 port map( D => n7845, CK => CLK, Q => 
                           n_2014, QN => n15386);
   REGISTERS_reg_66_10_inst : DFF_X1 port map( D => n7844, CK => CLK, Q => 
                           n_2015, QN => n15387);
   REGISTERS_reg_66_9_inst : DFF_X1 port map( D => n7843, CK => CLK, Q => 
                           n_2016, QN => n15388);
   REGISTERS_reg_66_8_inst : DFF_X1 port map( D => n7842, CK => CLK, Q => 
                           n_2017, QN => n15389);
   REGISTERS_reg_66_7_inst : DFF_X1 port map( D => n7841, CK => CLK, Q => 
                           n_2018, QN => n15390);
   REGISTERS_reg_66_6_inst : DFF_X1 port map( D => n7840, CK => CLK, Q => 
                           n_2019, QN => n15391);
   REGISTERS_reg_66_5_inst : DFF_X1 port map( D => n7839, CK => CLK, Q => 
                           n_2020, QN => n15392);
   REGISTERS_reg_66_4_inst : DFF_X1 port map( D => n7838, CK => CLK, Q => 
                           n_2021, QN => n15393);
   REGISTERS_reg_66_3_inst : DFF_X1 port map( D => n7837, CK => CLK, Q => 
                           n_2022, QN => n15394);
   REGISTERS_reg_66_2_inst : DFF_X1 port map( D => n7836, CK => CLK, Q => 
                           n_2023, QN => n15395);
   REGISTERS_reg_66_1_inst : DFF_X1 port map( D => n7835, CK => CLK, Q => 
                           n_2024, QN => n15396);
   REGISTERS_reg_66_0_inst : DFF_X1 port map( D => n7834, CK => CLK, Q => 
                           n_2025, QN => n15397);
   REGISTERS_reg_69_31_inst : DFF_X1 port map( D => n7769, CK => CLK, Q => 
                           n_2026, QN => n15462);
   REGISTERS_reg_69_30_inst : DFF_X1 port map( D => n7768, CK => CLK, Q => 
                           n_2027, QN => n15463);
   REGISTERS_reg_69_29_inst : DFF_X1 port map( D => n7767, CK => CLK, Q => 
                           n_2028, QN => n15464);
   REGISTERS_reg_69_28_inst : DFF_X1 port map( D => n7766, CK => CLK, Q => 
                           n_2029, QN => n15465);
   REGISTERS_reg_69_27_inst : DFF_X1 port map( D => n7765, CK => CLK, Q => 
                           n_2030, QN => n15466);
   REGISTERS_reg_69_26_inst : DFF_X1 port map( D => n7764, CK => CLK, Q => 
                           n_2031, QN => n15467);
   REGISTERS_reg_69_25_inst : DFF_X1 port map( D => n7763, CK => CLK, Q => 
                           n_2032, QN => n15468);
   REGISTERS_reg_69_24_inst : DFF_X1 port map( D => n7762, CK => CLK, Q => 
                           n_2033, QN => n15469);
   REGISTERS_reg_69_23_inst : DFF_X1 port map( D => n7761, CK => CLK, Q => 
                           n_2034, QN => n15470);
   REGISTERS_reg_69_22_inst : DFF_X1 port map( D => n7760, CK => CLK, Q => 
                           n_2035, QN => n15471);
   REGISTERS_reg_69_21_inst : DFF_X1 port map( D => n7759, CK => CLK, Q => 
                           n_2036, QN => n15472);
   REGISTERS_reg_69_20_inst : DFF_X1 port map( D => n7758, CK => CLK, Q => 
                           n_2037, QN => n15473);
   REGISTERS_reg_69_19_inst : DFF_X1 port map( D => n7757, CK => CLK, Q => 
                           n_2038, QN => n15474);
   REGISTERS_reg_69_18_inst : DFF_X1 port map( D => n7756, CK => CLK, Q => 
                           n_2039, QN => n15475);
   REGISTERS_reg_69_17_inst : DFF_X1 port map( D => n7755, CK => CLK, Q => 
                           n_2040, QN => n15476);
   REGISTERS_reg_69_16_inst : DFF_X1 port map( D => n7754, CK => CLK, Q => 
                           n_2041, QN => n15477);
   REGISTERS_reg_69_15_inst : DFF_X1 port map( D => n7753, CK => CLK, Q => 
                           n_2042, QN => n15478);
   REGISTERS_reg_69_14_inst : DFF_X1 port map( D => n7752, CK => CLK, Q => 
                           n_2043, QN => n15479);
   REGISTERS_reg_69_13_inst : DFF_X1 port map( D => n7751, CK => CLK, Q => 
                           n_2044, QN => n15480);
   REGISTERS_reg_69_12_inst : DFF_X1 port map( D => n7750, CK => CLK, Q => 
                           n_2045, QN => n15481);
   REGISTERS_reg_69_11_inst : DFF_X1 port map( D => n7749, CK => CLK, Q => 
                           n_2046, QN => n15482);
   REGISTERS_reg_69_10_inst : DFF_X1 port map( D => n7748, CK => CLK, Q => 
                           n_2047, QN => n15483);
   REGISTERS_reg_69_9_inst : DFF_X1 port map( D => n7747, CK => CLK, Q => 
                           n_2048, QN => n15484);
   REGISTERS_reg_69_8_inst : DFF_X1 port map( D => n7746, CK => CLK, Q => 
                           n_2049, QN => n15485);
   REGISTERS_reg_69_7_inst : DFF_X1 port map( D => n7745, CK => CLK, Q => 
                           n_2050, QN => n15486);
   REGISTERS_reg_69_6_inst : DFF_X1 port map( D => n7744, CK => CLK, Q => 
                           n_2051, QN => n15487);
   REGISTERS_reg_69_5_inst : DFF_X1 port map( D => n7743, CK => CLK, Q => 
                           n_2052, QN => n15488);
   REGISTERS_reg_69_4_inst : DFF_X1 port map( D => n7742, CK => CLK, Q => 
                           n_2053, QN => n15489);
   REGISTERS_reg_69_3_inst : DFF_X1 port map( D => n7741, CK => CLK, Q => 
                           n_2054, QN => n15490);
   REGISTERS_reg_69_2_inst : DFF_X1 port map( D => n7740, CK => CLK, Q => 
                           n_2055, QN => n15491);
   REGISTERS_reg_69_1_inst : DFF_X1 port map( D => n7739, CK => CLK, Q => 
                           n_2056, QN => n15492);
   REGISTERS_reg_69_0_inst : DFF_X1 port map( D => n7738, CK => CLK, Q => 
                           n_2057, QN => n15493);
   REGISTERS_reg_70_31_inst : DFF_X1 port map( D => n7737, CK => CLK, Q => 
                           n_2058, QN => n15494);
   REGISTERS_reg_70_30_inst : DFF_X1 port map( D => n7736, CK => CLK, Q => 
                           n_2059, QN => n15495);
   REGISTERS_reg_70_29_inst : DFF_X1 port map( D => n7735, CK => CLK, Q => 
                           n_2060, QN => n15496);
   REGISTERS_reg_70_28_inst : DFF_X1 port map( D => n7734, CK => CLK, Q => 
                           n_2061, QN => n15497);
   REGISTERS_reg_70_27_inst : DFF_X1 port map( D => n7733, CK => CLK, Q => 
                           n_2062, QN => n15498);
   REGISTERS_reg_70_26_inst : DFF_X1 port map( D => n7732, CK => CLK, Q => 
                           n_2063, QN => n15499);
   REGISTERS_reg_70_25_inst : DFF_X1 port map( D => n7731, CK => CLK, Q => 
                           n_2064, QN => n15500);
   REGISTERS_reg_70_24_inst : DFF_X1 port map( D => n7730, CK => CLK, Q => 
                           n_2065, QN => n15501);
   REGISTERS_reg_70_23_inst : DFF_X1 port map( D => n7729, CK => CLK, Q => 
                           n_2066, QN => n15502);
   REGISTERS_reg_70_22_inst : DFF_X1 port map( D => n7728, CK => CLK, Q => 
                           n_2067, QN => n15503);
   REGISTERS_reg_70_21_inst : DFF_X1 port map( D => n7727, CK => CLK, Q => 
                           n_2068, QN => n15504);
   REGISTERS_reg_70_20_inst : DFF_X1 port map( D => n7726, CK => CLK, Q => 
                           n_2069, QN => n15505);
   REGISTERS_reg_70_19_inst : DFF_X1 port map( D => n7725, CK => CLK, Q => 
                           n_2070, QN => n15506);
   REGISTERS_reg_70_18_inst : DFF_X1 port map( D => n7724, CK => CLK, Q => 
                           n_2071, QN => n15507);
   REGISTERS_reg_70_17_inst : DFF_X1 port map( D => n7723, CK => CLK, Q => 
                           n_2072, QN => n15508);
   REGISTERS_reg_70_16_inst : DFF_X1 port map( D => n7722, CK => CLK, Q => 
                           n_2073, QN => n15509);
   REGISTERS_reg_70_15_inst : DFF_X1 port map( D => n7721, CK => CLK, Q => 
                           n_2074, QN => n15510);
   REGISTERS_reg_70_14_inst : DFF_X1 port map( D => n7720, CK => CLK, Q => 
                           n_2075, QN => n15511);
   REGISTERS_reg_70_13_inst : DFF_X1 port map( D => n7719, CK => CLK, Q => 
                           n_2076, QN => n15512);
   REGISTERS_reg_70_12_inst : DFF_X1 port map( D => n7718, CK => CLK, Q => 
                           n_2077, QN => n15513);
   REGISTERS_reg_70_11_inst : DFF_X1 port map( D => n7717, CK => CLK, Q => 
                           n_2078, QN => n15514);
   REGISTERS_reg_70_10_inst : DFF_X1 port map( D => n7716, CK => CLK, Q => 
                           n_2079, QN => n15515);
   REGISTERS_reg_70_9_inst : DFF_X1 port map( D => n7715, CK => CLK, Q => 
                           n_2080, QN => n15516);
   REGISTERS_reg_70_8_inst : DFF_X1 port map( D => n7714, CK => CLK, Q => 
                           n_2081, QN => n15517);
   REGISTERS_reg_70_7_inst : DFF_X1 port map( D => n7713, CK => CLK, Q => 
                           n_2082, QN => n15518);
   REGISTERS_reg_70_6_inst : DFF_X1 port map( D => n7712, CK => CLK, Q => 
                           n_2083, QN => n15519);
   REGISTERS_reg_70_5_inst : DFF_X1 port map( D => n7711, CK => CLK, Q => 
                           n_2084, QN => n15520);
   REGISTERS_reg_70_4_inst : DFF_X1 port map( D => n7710, CK => CLK, Q => 
                           n_2085, QN => n15521);
   REGISTERS_reg_70_3_inst : DFF_X1 port map( D => n7709, CK => CLK, Q => 
                           n_2086, QN => n15522);
   REGISTERS_reg_70_2_inst : DFF_X1 port map( D => n7708, CK => CLK, Q => 
                           n_2087, QN => n15523);
   REGISTERS_reg_70_1_inst : DFF_X1 port map( D => n7707, CK => CLK, Q => 
                           n_2088, QN => n15524);
   REGISTERS_reg_70_0_inst : DFF_X1 port map( D => n7706, CK => CLK, Q => 
                           n_2089, QN => n15525);
   REGISTERS_reg_71_31_inst : DFF_X1 port map( D => n7705, CK => CLK, Q => 
                           n_2090, QN => n15526);
   REGISTERS_reg_71_30_inst : DFF_X1 port map( D => n7704, CK => CLK, Q => 
                           n_2091, QN => n15527);
   REGISTERS_reg_71_29_inst : DFF_X1 port map( D => n7703, CK => CLK, Q => 
                           n_2092, QN => n15528);
   REGISTERS_reg_71_28_inst : DFF_X1 port map( D => n7702, CK => CLK, Q => 
                           n_2093, QN => n15529);
   REGISTERS_reg_71_27_inst : DFF_X1 port map( D => n7701, CK => CLK, Q => 
                           n_2094, QN => n15530);
   REGISTERS_reg_71_26_inst : DFF_X1 port map( D => n7700, CK => CLK, Q => 
                           n_2095, QN => n15531);
   REGISTERS_reg_71_25_inst : DFF_X1 port map( D => n7699, CK => CLK, Q => 
                           n_2096, QN => n15532);
   REGISTERS_reg_71_24_inst : DFF_X1 port map( D => n7698, CK => CLK, Q => 
                           n_2097, QN => n15533);
   REGISTERS_reg_71_23_inst : DFF_X1 port map( D => n7697, CK => CLK, Q => 
                           n_2098, QN => n15534);
   REGISTERS_reg_71_22_inst : DFF_X1 port map( D => n7696, CK => CLK, Q => 
                           n_2099, QN => n15535);
   REGISTERS_reg_71_21_inst : DFF_X1 port map( D => n7695, CK => CLK, Q => 
                           n_2100, QN => n15536);
   REGISTERS_reg_71_20_inst : DFF_X1 port map( D => n7694, CK => CLK, Q => 
                           n_2101, QN => n15537);
   REGISTERS_reg_71_19_inst : DFF_X1 port map( D => n7693, CK => CLK, Q => 
                           n_2102, QN => n15538);
   REGISTERS_reg_71_18_inst : DFF_X1 port map( D => n7692, CK => CLK, Q => 
                           n_2103, QN => n15539);
   REGISTERS_reg_71_17_inst : DFF_X1 port map( D => n7691, CK => CLK, Q => 
                           n_2104, QN => n15540);
   REGISTERS_reg_71_16_inst : DFF_X1 port map( D => n7690, CK => CLK, Q => 
                           n_2105, QN => n15541);
   REGISTERS_reg_71_15_inst : DFF_X1 port map( D => n7689, CK => CLK, Q => 
                           n_2106, QN => n15542);
   REGISTERS_reg_71_14_inst : DFF_X1 port map( D => n7688, CK => CLK, Q => 
                           n_2107, QN => n15543);
   REGISTERS_reg_71_13_inst : DFF_X1 port map( D => n7687, CK => CLK, Q => 
                           n_2108, QN => n15544);
   REGISTERS_reg_71_12_inst : DFF_X1 port map( D => n7686, CK => CLK, Q => 
                           n_2109, QN => n15545);
   REGISTERS_reg_71_11_inst : DFF_X1 port map( D => n7685, CK => CLK, Q => 
                           n_2110, QN => n15546);
   REGISTERS_reg_71_10_inst : DFF_X1 port map( D => n7684, CK => CLK, Q => 
                           n_2111, QN => n15547);
   REGISTERS_reg_71_9_inst : DFF_X1 port map( D => n7683, CK => CLK, Q => 
                           n_2112, QN => n15548);
   REGISTERS_reg_71_8_inst : DFF_X1 port map( D => n7682, CK => CLK, Q => 
                           n_2113, QN => n15549);
   REGISTERS_reg_71_7_inst : DFF_X1 port map( D => n7681, CK => CLK, Q => 
                           n_2114, QN => n15550);
   REGISTERS_reg_71_6_inst : DFF_X1 port map( D => n7680, CK => CLK, Q => 
                           n_2115, QN => n15551);
   REGISTERS_reg_71_5_inst : DFF_X1 port map( D => n7679, CK => CLK, Q => 
                           n_2116, QN => n15552);
   REGISTERS_reg_71_4_inst : DFF_X1 port map( D => n7678, CK => CLK, Q => 
                           n_2117, QN => n15553);
   REGISTERS_reg_71_3_inst : DFF_X1 port map( D => n7677, CK => CLK, Q => 
                           n_2118, QN => n15554);
   REGISTERS_reg_71_2_inst : DFF_X1 port map( D => n7676, CK => CLK, Q => 
                           n_2119, QN => n15555);
   REGISTERS_reg_71_1_inst : DFF_X1 port map( D => n7675, CK => CLK, Q => 
                           n_2120, QN => n15556);
   REGISTERS_reg_71_0_inst : DFF_X1 port map( D => n7674, CK => CLK, Q => 
                           n_2121, QN => n15557);
   OUT1_tri_enable_reg_31_inst : DFF_X1 port map( D => n7672, CK => CLK, Q => 
                           n6659, QN => n1513);
   OUT1_tri_enable_reg_30_inst : DFF_X1 port map( D => n7670, CK => CLK, Q => 
                           n6661, QN => n1514);
   OUT1_tri_enable_reg_29_inst : DFF_X1 port map( D => n7668, CK => CLK, Q => 
                           n6663, QN => n1515);
   OUT1_tri_enable_reg_28_inst : DFF_X1 port map( D => n7666, CK => CLK, Q => 
                           n6665, QN => n1516);
   OUT1_tri_enable_reg_27_inst : DFF_X1 port map( D => n7664, CK => CLK, Q => 
                           n6667, QN => n1517);
   OUT1_tri_enable_reg_26_inst : DFF_X1 port map( D => n7662, CK => CLK, Q => 
                           n6669, QN => n1518);
   OUT1_tri_enable_reg_25_inst : DFF_X1 port map( D => n7660, CK => CLK, Q => 
                           n6671, QN => n1519);
   OUT1_tri_enable_reg_24_inst : DFF_X1 port map( D => n7658, CK => CLK, Q => 
                           n6673, QN => n1520);
   OUT1_reg_23_inst : DFF_X1 port map( D => n7657, CK => CLK, Q => n_2122, QN 
                           => n1457);
   OUT1_tri_enable_reg_23_inst : DFF_X1 port map( D => n7656, CK => CLK, Q => 
                           n6675, QN => n1521);
   OUT1_reg_22_inst : DFF_X1 port map( D => n7655, CK => CLK, Q => n_2123, QN 
                           => n1458);
   OUT1_tri_enable_reg_22_inst : DFF_X1 port map( D => n7654, CK => CLK, Q => 
                           n6677, QN => n1522);
   OUT1_reg_21_inst : DFF_X1 port map( D => n7653, CK => CLK, Q => n_2124, QN 
                           => n1459);
   OUT1_tri_enable_reg_21_inst : DFF_X1 port map( D => n7652, CK => CLK, Q => 
                           n6679, QN => n1523);
   OUT1_reg_20_inst : DFF_X1 port map( D => n7651, CK => CLK, Q => n_2125, QN 
                           => n1460);
   OUT1_tri_enable_reg_20_inst : DFF_X1 port map( D => n7650, CK => CLK, Q => 
                           n6681, QN => n1524);
   OUT1_reg_19_inst : DFF_X1 port map( D => n7649, CK => CLK, Q => n_2126, QN 
                           => n1461);
   OUT1_tri_enable_reg_19_inst : DFF_X1 port map( D => n7648, CK => CLK, Q => 
                           n6683, QN => n1525);
   OUT1_reg_18_inst : DFF_X1 port map( D => n7647, CK => CLK, Q => n_2127, QN 
                           => n1462);
   OUT1_tri_enable_reg_18_inst : DFF_X1 port map( D => n7646, CK => CLK, Q => 
                           n6685, QN => n1526);
   OUT1_reg_17_inst : DFF_X1 port map( D => n7645, CK => CLK, Q => n_2128, QN 
                           => n1463);
   OUT1_tri_enable_reg_17_inst : DFF_X1 port map( D => n7644, CK => CLK, Q => 
                           n6687, QN => n1527);
   OUT1_reg_16_inst : DFF_X1 port map( D => n7643, CK => CLK, Q => n_2129, QN 
                           => n1464);
   OUT1_tri_enable_reg_16_inst : DFF_X1 port map( D => n7642, CK => CLK, Q => 
                           n6689, QN => n1528);
   OUT1_reg_15_inst : DFF_X1 port map( D => n7641, CK => CLK, Q => n_2130, QN 
                           => n1465);
   OUT1_tri_enable_reg_15_inst : DFF_X1 port map( D => n7640, CK => CLK, Q => 
                           n6691, QN => n1529);
   OUT1_reg_14_inst : DFF_X1 port map( D => n7639, CK => CLK, Q => n_2131, QN 
                           => n1466);
   OUT1_tri_enable_reg_14_inst : DFF_X1 port map( D => n7638, CK => CLK, Q => 
                           n6693, QN => n1530);
   OUT1_reg_13_inst : DFF_X1 port map( D => n7637, CK => CLK, Q => n_2132, QN 
                           => n1467);
   OUT1_tri_enable_reg_13_inst : DFF_X1 port map( D => n7636, CK => CLK, Q => 
                           n6695, QN => n1531);
   OUT1_reg_12_inst : DFF_X1 port map( D => n7635, CK => CLK, Q => n_2133, QN 
                           => n1468);
   OUT1_tri_enable_reg_12_inst : DFF_X1 port map( D => n7634, CK => CLK, Q => 
                           n6697, QN => n1532);
   OUT1_reg_11_inst : DFF_X1 port map( D => n7633, CK => CLK, Q => n_2134, QN 
                           => n1469);
   OUT1_tri_enable_reg_11_inst : DFF_X1 port map( D => n7632, CK => CLK, Q => 
                           n6699, QN => n1533);
   OUT1_reg_10_inst : DFF_X1 port map( D => n7631, CK => CLK, Q => n_2135, QN 
                           => n1470);
   OUT1_tri_enable_reg_10_inst : DFF_X1 port map( D => n7630, CK => CLK, Q => 
                           n6701, QN => n1534);
   OUT1_reg_9_inst : DFF_X1 port map( D => n7629, CK => CLK, Q => n_2136, QN =>
                           n1471);
   OUT1_tri_enable_reg_9_inst : DFF_X1 port map( D => n7628, CK => CLK, Q => 
                           n6703, QN => n1535);
   OUT1_reg_8_inst : DFF_X1 port map( D => n7627, CK => CLK, Q => n_2137, QN =>
                           n1472);
   OUT1_tri_enable_reg_8_inst : DFF_X1 port map( D => n7626, CK => CLK, Q => 
                           n6705, QN => n1536);
   OUT1_reg_7_inst : DFF_X1 port map( D => n7625, CK => CLK, Q => n_2138, QN =>
                           n1473);
   OUT1_tri_enable_reg_7_inst : DFF_X1 port map( D => n7624, CK => CLK, Q => 
                           n6707, QN => n1537);
   OUT1_reg_6_inst : DFF_X1 port map( D => n7623, CK => CLK, Q => n_2139, QN =>
                           n1474);
   OUT1_tri_enable_reg_6_inst : DFF_X1 port map( D => n7622, CK => CLK, Q => 
                           n6709, QN => n1538);
   OUT1_reg_5_inst : DFF_X1 port map( D => n7621, CK => CLK, Q => n_2140, QN =>
                           n1475);
   OUT1_tri_enable_reg_5_inst : DFF_X1 port map( D => n7620, CK => CLK, Q => 
                           n6711, QN => n1539);
   OUT1_reg_4_inst : DFF_X1 port map( D => n7619, CK => CLK, Q => n_2141, QN =>
                           n1476);
   OUT1_tri_enable_reg_4_inst : DFF_X1 port map( D => n7618, CK => CLK, Q => 
                           n6713, QN => n1540);
   OUT1_reg_3_inst : DFF_X1 port map( D => n7617, CK => CLK, Q => n_2142, QN =>
                           n1477);
   OUT1_tri_enable_reg_3_inst : DFF_X1 port map( D => n7616, CK => CLK, Q => 
                           n6715, QN => n1541);
   OUT1_reg_2_inst : DFF_X1 port map( D => n7615, CK => CLK, Q => n_2143, QN =>
                           n1478);
   OUT1_tri_enable_reg_2_inst : DFF_X1 port map( D => n7614, CK => CLK, Q => 
                           n6717, QN => n1542);
   OUT1_reg_1_inst : DFF_X1 port map( D => n7613, CK => CLK, Q => n_2144, QN =>
                           n1479);
   OUT1_tri_enable_reg_1_inst : DFF_X1 port map( D => n7612, CK => CLK, Q => 
                           n6719, QN => n1543);
   OUT1_reg_0_inst : DFF_X1 port map( D => n7611, CK => CLK, Q => n_2145, QN =>
                           n1480);
   OUT1_tri_enable_reg_0_inst : DFF_X1 port map( D => n7610, CK => CLK, Q => 
                           n6721, QN => n1544);
   OUT2_tri_enable_reg_31_inst : DFF_X1 port map( D => n7608, CK => CLK, Q => 
                           n6723, QN => n1545);
   OUT2_tri_enable_reg_30_inst : DFF_X1 port map( D => n7606, CK => CLK, Q => 
                           n6725, QN => n1546);
   OUT2_tri_enable_reg_29_inst : DFF_X1 port map( D => n7604, CK => CLK, Q => 
                           n6727, QN => n1547);
   OUT2_tri_enable_reg_28_inst : DFF_X1 port map( D => n7602, CK => CLK, Q => 
                           n6729, QN => n1548);
   OUT2_tri_enable_reg_27_inst : DFF_X1 port map( D => n7600, CK => CLK, Q => 
                           n6731, QN => n1549);
   OUT2_tri_enable_reg_26_inst : DFF_X1 port map( D => n7598, CK => CLK, Q => 
                           n6733, QN => n1550);
   OUT2_tri_enable_reg_25_inst : DFF_X1 port map( D => n7596, CK => CLK, Q => 
                           n6735, QN => n1551);
   OUT2_tri_enable_reg_24_inst : DFF_X1 port map( D => n7594, CK => CLK, Q => 
                           n6737, QN => n1552);
   OUT2_reg_23_inst : DFF_X1 port map( D => n7593, CK => CLK, Q => n_2146, QN 
                           => n1489);
   OUT2_tri_enable_reg_23_inst : DFF_X1 port map( D => n7592, CK => CLK, Q => 
                           n6739, QN => n1553);
   OUT2_reg_22_inst : DFF_X1 port map( D => n7591, CK => CLK, Q => n_2147, QN 
                           => n1490);
   OUT2_tri_enable_reg_22_inst : DFF_X1 port map( D => n7590, CK => CLK, Q => 
                           n6741, QN => n1554);
   OUT2_reg_21_inst : DFF_X1 port map( D => n7589, CK => CLK, Q => n_2148, QN 
                           => n1491);
   OUT2_tri_enable_reg_21_inst : DFF_X1 port map( D => n7588, CK => CLK, Q => 
                           n6743, QN => n1555);
   OUT2_reg_20_inst : DFF_X1 port map( D => n7587, CK => CLK, Q => n_2149, QN 
                           => n1492);
   OUT2_tri_enable_reg_20_inst : DFF_X1 port map( D => n7586, CK => CLK, Q => 
                           n6745, QN => n1556);
   OUT2_reg_19_inst : DFF_X1 port map( D => n7585, CK => CLK, Q => n_2150, QN 
                           => n1493);
   OUT2_tri_enable_reg_19_inst : DFF_X1 port map( D => n7584, CK => CLK, Q => 
                           n6747, QN => n1557);
   OUT2_reg_18_inst : DFF_X1 port map( D => n7583, CK => CLK, Q => n_2151, QN 
                           => n1494);
   OUT2_tri_enable_reg_18_inst : DFF_X1 port map( D => n7582, CK => CLK, Q => 
                           n6749, QN => n1558);
   OUT2_reg_17_inst : DFF_X1 port map( D => n7581, CK => CLK, Q => n_2152, QN 
                           => n1495);
   OUT2_tri_enable_reg_17_inst : DFF_X1 port map( D => n7580, CK => CLK, Q => 
                           n6751, QN => n1559);
   OUT2_reg_16_inst : DFF_X1 port map( D => n7579, CK => CLK, Q => n_2153, QN 
                           => n1496);
   OUT2_tri_enable_reg_16_inst : DFF_X1 port map( D => n7578, CK => CLK, Q => 
                           n6753, QN => n1560);
   OUT2_reg_15_inst : DFF_X1 port map( D => n7577, CK => CLK, Q => n_2154, QN 
                           => n1497);
   OUT2_tri_enable_reg_15_inst : DFF_X1 port map( D => n7576, CK => CLK, Q => 
                           n6755, QN => n1561);
   OUT2_reg_14_inst : DFF_X1 port map( D => n7575, CK => CLK, Q => n_2155, QN 
                           => n1498);
   OUT2_tri_enable_reg_14_inst : DFF_X1 port map( D => n7574, CK => CLK, Q => 
                           n6757, QN => n1562);
   OUT2_reg_13_inst : DFF_X1 port map( D => n7573, CK => CLK, Q => n_2156, QN 
                           => n1499);
   OUT2_tri_enable_reg_13_inst : DFF_X1 port map( D => n7572, CK => CLK, Q => 
                           n6759, QN => n1563);
   OUT2_reg_12_inst : DFF_X1 port map( D => n7571, CK => CLK, Q => n_2157, QN 
                           => n1500);
   OUT2_tri_enable_reg_12_inst : DFF_X1 port map( D => n7570, CK => CLK, Q => 
                           n6761, QN => n1564);
   OUT2_reg_11_inst : DFF_X1 port map( D => n7569, CK => CLK, Q => n_2158, QN 
                           => n1501);
   OUT2_tri_enable_reg_11_inst : DFF_X1 port map( D => n7568, CK => CLK, Q => 
                           n6763, QN => n1565);
   OUT2_reg_10_inst : DFF_X1 port map( D => n7567, CK => CLK, Q => n_2159, QN 
                           => n1502);
   OUT2_tri_enable_reg_10_inst : DFF_X1 port map( D => n7566, CK => CLK, Q => 
                           n6765, QN => n1566);
   OUT2_reg_9_inst : DFF_X1 port map( D => n7565, CK => CLK, Q => n_2160, QN =>
                           n1503);
   OUT2_tri_enable_reg_9_inst : DFF_X1 port map( D => n7564, CK => CLK, Q => 
                           n6767, QN => n1567);
   OUT2_reg_8_inst : DFF_X1 port map( D => n7563, CK => CLK, Q => n_2161, QN =>
                           n1504);
   OUT2_tri_enable_reg_8_inst : DFF_X1 port map( D => n7562, CK => CLK, Q => 
                           n6769, QN => n1568);
   OUT2_reg_7_inst : DFF_X1 port map( D => n7561, CK => CLK, Q => n_2162, QN =>
                           n1505);
   OUT2_tri_enable_reg_7_inst : DFF_X1 port map( D => n7560, CK => CLK, Q => 
                           n6771, QN => n1569);
   OUT2_reg_6_inst : DFF_X1 port map( D => n7559, CK => CLK, Q => n_2163, QN =>
                           n1506);
   OUT2_tri_enable_reg_6_inst : DFF_X1 port map( D => n7558, CK => CLK, Q => 
                           n6773, QN => n1570);
   OUT2_reg_5_inst : DFF_X1 port map( D => n7557, CK => CLK, Q => n_2164, QN =>
                           n1507);
   OUT2_tri_enable_reg_5_inst : DFF_X1 port map( D => n7556, CK => CLK, Q => 
                           n6775, QN => n1571);
   OUT2_reg_4_inst : DFF_X1 port map( D => n7555, CK => CLK, Q => n_2165, QN =>
                           n1508);
   OUT2_tri_enable_reg_4_inst : DFF_X1 port map( D => n7554, CK => CLK, Q => 
                           n6777, QN => n1572);
   OUT2_reg_3_inst : DFF_X1 port map( D => n7553, CK => CLK, Q => n_2166, QN =>
                           n1509);
   OUT2_tri_enable_reg_3_inst : DFF_X1 port map( D => n7552, CK => CLK, Q => 
                           n6779, QN => n1573);
   OUT2_reg_2_inst : DFF_X1 port map( D => n7551, CK => CLK, Q => n_2167, QN =>
                           n1510);
   OUT2_tri_enable_reg_2_inst : DFF_X1 port map( D => n7550, CK => CLK, Q => 
                           n6781, QN => n1574);
   OUT2_reg_1_inst : DFF_X1 port map( D => n7549, CK => CLK, Q => n_2168, QN =>
                           n1511);
   OUT2_tri_enable_reg_1_inst : DFF_X1 port map( D => n7548, CK => CLK, Q => 
                           n6783, QN => n1575);
   OUT2_reg_0_inst : DFF_X1 port map( D => n7547, CK => CLK, Q => n_2169, QN =>
                           n1512);
   OUT2_tri_enable_reg_0_inst : DFF_X1 port map( D => n7546, CK => CLK, Q => 
                           n6785, QN => n1576);
   REGISTERS_reg_48_31_inst : DFF_X1 port map( D => n8441, CK => CLK, Q => 
                           n_2170, QN => n15923);
   REGISTERS_reg_48_30_inst : DFF_X1 port map( D => n8440, CK => CLK, Q => 
                           n_2171, QN => n15924);
   REGISTERS_reg_48_29_inst : DFF_X1 port map( D => n8439, CK => CLK, Q => 
                           n_2172, QN => n15925);
   REGISTERS_reg_48_28_inst : DFF_X1 port map( D => n8438, CK => CLK, Q => 
                           n_2173, QN => n15926);
   REGISTERS_reg_48_27_inst : DFF_X1 port map( D => n8437, CK => CLK, Q => 
                           n_2174, QN => n15927);
   REGISTERS_reg_48_26_inst : DFF_X1 port map( D => n8436, CK => CLK, Q => 
                           n_2175, QN => n15928);
   REGISTERS_reg_48_25_inst : DFF_X1 port map( D => n8435, CK => CLK, Q => 
                           n_2176, QN => n15929);
   REGISTERS_reg_48_24_inst : DFF_X1 port map( D => n8434, CK => CLK, Q => 
                           n_2177, QN => n15930);
   REGISTERS_reg_48_23_inst : DFF_X1 port map( D => n8433, CK => CLK, Q => 
                           n_2178, QN => n15947);
   REGISTERS_reg_48_22_inst : DFF_X1 port map( D => n8432, CK => CLK, Q => 
                           n_2179, QN => n15948);
   REGISTERS_reg_48_21_inst : DFF_X1 port map( D => n8431, CK => CLK, Q => 
                           n_2180, QN => n15949);
   REGISTERS_reg_48_20_inst : DFF_X1 port map( D => n8430, CK => CLK, Q => 
                           n_2181, QN => n15950);
   REGISTERS_reg_48_19_inst : DFF_X1 port map( D => n8429, CK => CLK, Q => 
                           n_2182, QN => n15951);
   REGISTERS_reg_48_18_inst : DFF_X1 port map( D => n8428, CK => CLK, Q => 
                           n_2183, QN => n15952);
   REGISTERS_reg_48_17_inst : DFF_X1 port map( D => n8427, CK => CLK, Q => 
                           n_2184, QN => n15953);
   REGISTERS_reg_48_16_inst : DFF_X1 port map( D => n8426, CK => CLK, Q => 
                           n_2185, QN => n15954);
   REGISTERS_reg_48_15_inst : DFF_X1 port map( D => n8425, CK => CLK, Q => 
                           n_2186, QN => n15955);
   REGISTERS_reg_48_14_inst : DFF_X1 port map( D => n8424, CK => CLK, Q => 
                           n_2187, QN => n15956);
   REGISTERS_reg_48_13_inst : DFF_X1 port map( D => n8423, CK => CLK, Q => 
                           n_2188, QN => n15957);
   REGISTERS_reg_48_12_inst : DFF_X1 port map( D => n8422, CK => CLK, Q => 
                           n_2189, QN => n15958);
   REGISTERS_reg_48_11_inst : DFF_X1 port map( D => n8421, CK => CLK, Q => 
                           n_2190, QN => n15959);
   REGISTERS_reg_48_10_inst : DFF_X1 port map( D => n8420, CK => CLK, Q => 
                           n_2191, QN => n15960);
   REGISTERS_reg_48_9_inst : DFF_X1 port map( D => n8419, CK => CLK, Q => 
                           n_2192, QN => n15961);
   REGISTERS_reg_48_8_inst : DFF_X1 port map( D => n8418, CK => CLK, Q => 
                           n_2193, QN => n15962);
   REGISTERS_reg_48_7_inst : DFF_X1 port map( D => n8417, CK => CLK, Q => 
                           n_2194, QN => n15963);
   REGISTERS_reg_48_6_inst : DFF_X1 port map( D => n8416, CK => CLK, Q => 
                           n_2195, QN => n15964);
   REGISTERS_reg_48_5_inst : DFF_X1 port map( D => n8415, CK => CLK, Q => 
                           n_2196, QN => n15965);
   REGISTERS_reg_48_4_inst : DFF_X1 port map( D => n8414, CK => CLK, Q => 
                           n_2197, QN => n15966);
   REGISTERS_reg_48_3_inst : DFF_X1 port map( D => n8413, CK => CLK, Q => 
                           n_2198, QN => n15967);
   REGISTERS_reg_48_2_inst : DFF_X1 port map( D => n8412, CK => CLK, Q => 
                           n_2199, QN => n15968);
   REGISTERS_reg_48_1_inst : DFF_X1 port map( D => n8411, CK => CLK, Q => 
                           n_2200, QN => n15969);
   REGISTERS_reg_48_0_inst : DFF_X1 port map( D => n8410, CK => CLK, Q => 
                           n_2201, QN => n15970);
   U5 : TINV_X1 port map( I => n1449, EN => n6659, ZN => OUT1(31));
   U6 : TINV_X1 port map( I => n1450, EN => n6661, ZN => OUT1(30));
   U7 : TINV_X1 port map( I => n1451, EN => n6663, ZN => OUT1(29));
   U8 : TINV_X1 port map( I => n1452, EN => n6665, ZN => OUT1(28));
   U9 : TINV_X1 port map( I => n1453, EN => n6667, ZN => OUT1(27));
   U10 : TINV_X1 port map( I => n1454, EN => n6669, ZN => OUT1(26));
   U11 : TINV_X1 port map( I => n1455, EN => n6671, ZN => OUT1(25));
   U12 : TINV_X1 port map( I => n1456, EN => n6673, ZN => OUT1(24));
   U13 : TINV_X1 port map( I => n1457, EN => n6675, ZN => OUT1(23));
   U14 : TINV_X1 port map( I => n1458, EN => n6677, ZN => OUT1(22));
   U15 : TINV_X1 port map( I => n1459, EN => n6679, ZN => OUT1(21));
   U16 : TINV_X1 port map( I => n1460, EN => n6681, ZN => OUT1(20));
   U17 : TINV_X1 port map( I => n1461, EN => n6683, ZN => OUT1(19));
   U18 : TINV_X1 port map( I => n1462, EN => n6685, ZN => OUT1(18));
   U19 : TINV_X1 port map( I => n1463, EN => n6687, ZN => OUT1(17));
   U20 : TINV_X1 port map( I => n1464, EN => n6689, ZN => OUT1(16));
   U21 : TINV_X1 port map( I => n1465, EN => n6691, ZN => OUT1(15));
   U22 : TINV_X1 port map( I => n1466, EN => n6693, ZN => OUT1(14));
   U23 : TINV_X1 port map( I => n1467, EN => n6695, ZN => OUT1(13));
   U24 : TINV_X1 port map( I => n1468, EN => n6697, ZN => OUT1(12));
   U25 : TINV_X1 port map( I => n1469, EN => n6699, ZN => OUT1(11));
   U26 : TINV_X1 port map( I => n1470, EN => n6701, ZN => OUT1(10));
   U27 : TINV_X1 port map( I => n1471, EN => n6703, ZN => OUT1(9));
   U28 : TINV_X1 port map( I => n1472, EN => n6705, ZN => OUT1(8));
   U29 : TINV_X1 port map( I => n1473, EN => n6707, ZN => OUT1(7));
   U30 : TINV_X1 port map( I => n1474, EN => n6709, ZN => OUT1(6));
   U31 : TINV_X1 port map( I => n1475, EN => n6711, ZN => OUT1(5));
   U32 : TINV_X1 port map( I => n1476, EN => n6713, ZN => OUT1(4));
   U33 : TINV_X1 port map( I => n1477, EN => n6715, ZN => OUT1(3));
   U34 : TINV_X1 port map( I => n1478, EN => n6717, ZN => OUT1(2));
   U35 : TINV_X1 port map( I => n1479, EN => n6719, ZN => OUT1(1));
   U36 : TINV_X1 port map( I => n1480, EN => n6721, ZN => OUT1(0));
   U37 : TINV_X1 port map( I => n1481, EN => n6723, ZN => OUT2(31));
   U38 : TINV_X1 port map( I => n1482, EN => n6725, ZN => OUT2(30));
   U39 : TINV_X1 port map( I => n1483, EN => n6727, ZN => OUT2(29));
   U40 : TINV_X1 port map( I => n1484, EN => n6729, ZN => OUT2(28));
   U41 : TINV_X1 port map( I => n1485, EN => n6731, ZN => OUT2(27));
   U42 : TINV_X1 port map( I => n1486, EN => n6733, ZN => OUT2(26));
   U43 : TINV_X1 port map( I => n1487, EN => n6735, ZN => OUT2(25));
   U44 : TINV_X1 port map( I => n1488, EN => n6737, ZN => OUT2(24));
   U45 : TINV_X1 port map( I => n1489, EN => n6739, ZN => OUT2(23));
   U46 : TINV_X1 port map( I => n1490, EN => n6741, ZN => OUT2(22));
   U47 : TINV_X1 port map( I => n1491, EN => n6743, ZN => OUT2(21));
   U48 : TINV_X1 port map( I => n1492, EN => n6745, ZN => OUT2(20));
   U49 : TINV_X1 port map( I => n1493, EN => n6747, ZN => OUT2(19));
   U50 : TINV_X1 port map( I => n1494, EN => n6749, ZN => OUT2(18));
   U51 : TINV_X1 port map( I => n1495, EN => n6751, ZN => OUT2(17));
   U52 : TINV_X1 port map( I => n1496, EN => n6753, ZN => OUT2(16));
   U53 : TINV_X1 port map( I => n1497, EN => n6755, ZN => OUT2(15));
   U54 : TINV_X1 port map( I => n1498, EN => n6757, ZN => OUT2(14));
   U55 : TINV_X1 port map( I => n1499, EN => n6759, ZN => OUT2(13));
   U56 : TINV_X1 port map( I => n1500, EN => n6761, ZN => OUT2(12));
   U57 : TINV_X1 port map( I => n1501, EN => n6763, ZN => OUT2(11));
   U58 : TINV_X1 port map( I => n1502, EN => n6765, ZN => OUT2(10));
   U59 : TINV_X1 port map( I => n1503, EN => n6767, ZN => OUT2(9));
   U60 : TINV_X1 port map( I => n1504, EN => n6769, ZN => OUT2(8));
   U61 : TINV_X1 port map( I => n1505, EN => n6771, ZN => OUT2(7));
   U62 : TINV_X1 port map( I => n1506, EN => n6773, ZN => OUT2(6));
   U63 : TINV_X1 port map( I => n1507, EN => n6775, ZN => OUT2(5));
   U64 : TINV_X1 port map( I => n1508, EN => n6777, ZN => OUT2(4));
   U65 : TINV_X1 port map( I => n1509, EN => n6779, ZN => OUT2(3));
   U66 : TINV_X1 port map( I => n1510, EN => n6781, ZN => OUT2(2));
   U67 : TINV_X1 port map( I => n1511, EN => n6783, ZN => OUT2(1));
   U68 : TINV_X1 port map( I => n1512, EN => n6785, ZN => OUT2(0));
   U3817 : NOR4_X2 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), A3 => 
                           ADD_RD1(5), A4 => ADD_RD1(6), ZN => n4282);
   U5158 : NOR4_X2 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), A3 => 
                           ADD_RD2(5), A4 => ADD_RD2(6), ZN => n5679);
   U5252 : NOR3_X2 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), A3 => 
                           ADD_RD2(0), ZN => n5660);
   U7617 : XOR2_X1 port map( A => ADD_WR(6), B => ADD_RD1(6), Z => n4320);
   U7618 : XOR2_X1 port map( A => ADD_WR(5), B => ADD_RD1(5), Z => n4319);
   U7619 : XOR2_X1 port map( A => ADD_WR(4), B => ADD_RD1(4), Z => n4318);
   U7620 : XOR2_X1 port map( A => ADD_WR(3), B => ADD_RD1(3), Z => n4317);
   U7621 : XOR2_X1 port map( A => ADD_WR(0), B => ADD_RD1(0), Z => n4321);
   U7622 : XOR2_X1 port map( A => n16071, B => ADD_RD1(1), Z => n4314);
   U7623 : XOR2_X1 port map( A => n16072, B => ADD_RD1(2), Z => n4313);
   U7624 : XOR2_X1 port map( A => ADD_WR(6), B => ADD_RD2(6), Z => n5752);
   U7625 : XOR2_X1 port map( A => ADD_WR(5), B => ADD_RD2(5), Z => n5750);
   U7626 : XOR2_X1 port map( A => ADD_WR(4), B => ADD_RD2(4), Z => n5748);
   U7627 : XOR2_X1 port map( A => ADD_WR(3), B => ADD_RD2(3), Z => n5746);
   U7628 : XOR2_X1 port map( A => ADD_WR(0), B => ADD_RD2(0), Z => n5754);
   U7629 : XOR2_X1 port map( A => n16071, B => ADD_RD2(1), Z => n5740);
   U7630 : XOR2_X1 port map( A => n16072, B => ADD_RD2(2), Z => n5738);
   REGISTERS_reg_68_31_inst : DFF_X1 port map( D => n7801, CK => CLK, Q => 
                           n15430, QN => n6973);
   REGISTERS_reg_68_30_inst : DFF_X1 port map( D => n7800, CK => CLK, Q => 
                           n15431, QN => n6972);
   REGISTERS_reg_68_29_inst : DFF_X1 port map( D => n7799, CK => CLK, Q => 
                           n15432, QN => n6971);
   REGISTERS_reg_68_28_inst : DFF_X1 port map( D => n7798, CK => CLK, Q => 
                           n15433, QN => n6970);
   REGISTERS_reg_68_27_inst : DFF_X1 port map( D => n7797, CK => CLK, Q => 
                           n15434, QN => n6969);
   REGISTERS_reg_68_26_inst : DFF_X1 port map( D => n7796, CK => CLK, Q => 
                           n15435, QN => n6968);
   REGISTERS_reg_68_25_inst : DFF_X1 port map( D => n7795, CK => CLK, Q => 
                           n15436, QN => n6967);
   REGISTERS_reg_68_24_inst : DFF_X1 port map( D => n7794, CK => CLK, Q => 
                           n15437, QN => n6966);
   REGISTERS_reg_67_31_inst : DFF_X1 port map( D => n7833, CK => CLK, Q => 
                           n15398, QN => n7191);
   REGISTERS_reg_67_30_inst : DFF_X1 port map( D => n7832, CK => CLK, Q => 
                           n15399, QN => n7190);
   REGISTERS_reg_67_29_inst : DFF_X1 port map( D => n7831, CK => CLK, Q => 
                           n15400, QN => n7189);
   REGISTERS_reg_67_28_inst : DFF_X1 port map( D => n7830, CK => CLK, Q => 
                           n15401, QN => n7188);
   REGISTERS_reg_67_27_inst : DFF_X1 port map( D => n7829, CK => CLK, Q => 
                           n15402, QN => n7187);
   REGISTERS_reg_67_26_inst : DFF_X1 port map( D => n7828, CK => CLK, Q => 
                           n15403, QN => n7186);
   REGISTERS_reg_67_25_inst : DFF_X1 port map( D => n7827, CK => CLK, Q => 
                           n15404, QN => n7185);
   REGISTERS_reg_67_24_inst : DFF_X1 port map( D => n7826, CK => CLK, Q => 
                           n15405, QN => n7184);
   REGISTERS_reg_63_31_inst : DFF_X1 port map( D => n7961, CK => CLK, Q => 
                           n15302, QN => n7223);
   REGISTERS_reg_63_30_inst : DFF_X1 port map( D => n7960, CK => CLK, Q => 
                           n15303, QN => n7222);
   REGISTERS_reg_63_29_inst : DFF_X1 port map( D => n7959, CK => CLK, Q => 
                           n15304, QN => n7221);
   REGISTERS_reg_63_28_inst : DFF_X1 port map( D => n7958, CK => CLK, Q => 
                           n15305, QN => n7220);
   REGISTERS_reg_63_27_inst : DFF_X1 port map( D => n7957, CK => CLK, Q => 
                           n15306, QN => n7219);
   REGISTERS_reg_63_26_inst : DFF_X1 port map( D => n7956, CK => CLK, Q => 
                           n15307, QN => n7218);
   REGISTERS_reg_63_25_inst : DFF_X1 port map( D => n7955, CK => CLK, Q => 
                           n15308, QN => n7217);
   REGISTERS_reg_63_24_inst : DFF_X1 port map( D => n7954, CK => CLK, Q => 
                           n15309, QN => n7216);
   REGISTERS_reg_58_31_inst : DFF_X1 port map( D => n8121, CK => CLK, Q => 
                           n15174, QN => n7255);
   REGISTERS_reg_58_30_inst : DFF_X1 port map( D => n8120, CK => CLK, Q => 
                           n15175, QN => n7254);
   REGISTERS_reg_58_29_inst : DFF_X1 port map( D => n8119, CK => CLK, Q => 
                           n15176, QN => n7253);
   REGISTERS_reg_58_28_inst : DFF_X1 port map( D => n8118, CK => CLK, Q => 
                           n15177, QN => n7252);
   REGISTERS_reg_58_27_inst : DFF_X1 port map( D => n8117, CK => CLK, Q => 
                           n15178, QN => n7251);
   REGISTERS_reg_58_26_inst : DFF_X1 port map( D => n8116, CK => CLK, Q => 
                           n15179, QN => n7250);
   REGISTERS_reg_58_25_inst : DFF_X1 port map( D => n8115, CK => CLK, Q => 
                           n15180, QN => n7249);
   REGISTERS_reg_58_24_inst : DFF_X1 port map( D => n8114, CK => CLK, Q => 
                           n15181, QN => n7248);
   REGISTERS_reg_50_31_inst : DFF_X1 port map( D => n8377, CK => CLK, Q => 
                           n14982, QN => n6981);
   REGISTERS_reg_50_30_inst : DFF_X1 port map( D => n8376, CK => CLK, Q => 
                           n14983, QN => n6980);
   REGISTERS_reg_50_29_inst : DFF_X1 port map( D => n8375, CK => CLK, Q => 
                           n14984, QN => n6979);
   REGISTERS_reg_50_28_inst : DFF_X1 port map( D => n8374, CK => CLK, Q => 
                           n14985, QN => n6978);
   REGISTERS_reg_50_27_inst : DFF_X1 port map( D => n8373, CK => CLK, Q => 
                           n14986, QN => n6977);
   REGISTERS_reg_50_26_inst : DFF_X1 port map( D => n8372, CK => CLK, Q => 
                           n14987, QN => n6976);
   REGISTERS_reg_50_25_inst : DFF_X1 port map( D => n8371, CK => CLK, Q => 
                           n14988, QN => n6975);
   REGISTERS_reg_50_24_inst : DFF_X1 port map( D => n8370, CK => CLK, Q => 
                           n14989, QN => n6974);
   REGISTERS_reg_49_31_inst : DFF_X1 port map( D => n8409, CK => CLK, Q => 
                           n15634, QN => n969);
   REGISTERS_reg_49_30_inst : DFF_X1 port map( D => n8408, CK => CLK, Q => 
                           n15635, QN => n970);
   REGISTERS_reg_49_29_inst : DFF_X1 port map( D => n8407, CK => CLK, Q => 
                           n15636, QN => n971);
   REGISTERS_reg_49_28_inst : DFF_X1 port map( D => n8406, CK => CLK, Q => 
                           n15637, QN => n972);
   REGISTERS_reg_49_27_inst : DFF_X1 port map( D => n8405, CK => CLK, Q => 
                           n15638, QN => n973);
   REGISTERS_reg_49_26_inst : DFF_X1 port map( D => n8404, CK => CLK, Q => 
                           n15639, QN => n974);
   REGISTERS_reg_49_25_inst : DFF_X1 port map( D => n8403, CK => CLK, Q => 
                           n15640, QN => n975);
   REGISTERS_reg_49_24_inst : DFF_X1 port map( D => n8402, CK => CLK, Q => 
                           n15641, QN => n976);
   REGISTERS_reg_45_31_inst : DFF_X1 port map( D => n8537, CK => CLK, Q => 
                           n14948, QN => n7257);
   REGISTERS_reg_45_30_inst : DFF_X1 port map( D => n8536, CK => CLK, Q => 
                           n15613, QN => n622);
   REGISTERS_reg_45_29_inst : DFF_X1 port map( D => n8535, CK => CLK, Q => 
                           n15614, QN => n625);
   REGISTERS_reg_45_28_inst : DFF_X1 port map( D => n8534, CK => CLK, Q => 
                           n15615, QN => n628);
   REGISTERS_reg_45_27_inst : DFF_X1 port map( D => n8533, CK => CLK, Q => 
                           n15616, QN => n631);
   REGISTERS_reg_45_26_inst : DFF_X1 port map( D => n8532, CK => CLK, Q => 
                           n15617, QN => n634);
   REGISTERS_reg_45_25_inst : DFF_X1 port map( D => n8531, CK => CLK, Q => 
                           n15618, QN => n637);
   REGISTERS_reg_45_24_inst : DFF_X1 port map( D => n8530, CK => CLK, Q => 
                           n15619, QN => n640);
   REGISTERS_reg_40_31_inst : DFF_X1 port map( D => n8697, CK => CLK, Q => 
                           n15558, QN => n937);
   REGISTERS_reg_40_30_inst : DFF_X1 port map( D => n8696, CK => CLK, Q => 
                           n15559, QN => n938);
   REGISTERS_reg_40_29_inst : DFF_X1 port map( D => n8695, CK => CLK, Q => 
                           n15560, QN => n939);
   REGISTERS_reg_40_28_inst : DFF_X1 port map( D => n8694, CK => CLK, Q => 
                           n15561, QN => n940);
   REGISTERS_reg_40_27_inst : DFF_X1 port map( D => n8693, CK => CLK, Q => 
                           n15562, QN => n941);
   REGISTERS_reg_40_26_inst : DFF_X1 port map( D => n8692, CK => CLK, Q => 
                           n15563, QN => n942);
   REGISTERS_reg_40_25_inst : DFF_X1 port map( D => n8691, CK => CLK, Q => 
                           n15564, QN => n943);
   REGISTERS_reg_40_24_inst : DFF_X1 port map( D => n8690, CK => CLK, Q => 
                           n15565, QN => n944);
   REGISTERS_reg_32_31_inst : DFF_X1 port map( D => n8953, CK => CLK, Q => 
                           n14660, QN => n6989);
   REGISTERS_reg_32_30_inst : DFF_X1 port map( D => n8952, CK => CLK, Q => 
                           n14661, QN => n6988);
   REGISTERS_reg_32_29_inst : DFF_X1 port map( D => n8951, CK => CLK, Q => 
                           n14662, QN => n6987);
   REGISTERS_reg_32_28_inst : DFF_X1 port map( D => n8950, CK => CLK, Q => 
                           n14663, QN => n6986);
   REGISTERS_reg_32_27_inst : DFF_X1 port map( D => n8949, CK => CLK, Q => 
                           n14664, QN => n6985);
   REGISTERS_reg_32_26_inst : DFF_X1 port map( D => n8948, CK => CLK, Q => 
                           n14665, QN => n6984);
   REGISTERS_reg_32_25_inst : DFF_X1 port map( D => n8947, CK => CLK, Q => 
                           n14666, QN => n6983);
   REGISTERS_reg_32_24_inst : DFF_X1 port map( D => n8946, CK => CLK, Q => 
                           n14667, QN => n6982);
   REGISTERS_reg_31_31_inst : DFF_X1 port map( D => n8985, CK => CLK, Q => 
                           n15566, QN => n905);
   REGISTERS_reg_31_30_inst : DFF_X1 port map( D => n8984, CK => CLK, Q => 
                           n15567, QN => n906);
   REGISTERS_reg_31_29_inst : DFF_X1 port map( D => n8983, CK => CLK, Q => 
                           n15568, QN => n907);
   REGISTERS_reg_31_28_inst : DFF_X1 port map( D => n8982, CK => CLK, Q => 
                           n15569, QN => n908);
   REGISTERS_reg_31_27_inst : DFF_X1 port map( D => n8981, CK => CLK, Q => 
                           n15570, QN => n909);
   REGISTERS_reg_31_26_inst : DFF_X1 port map( D => n8980, CK => CLK, Q => 
                           n15571, QN => n910);
   REGISTERS_reg_31_25_inst : DFF_X1 port map( D => n8979, CK => CLK, Q => 
                           n15572, QN => n911);
   REGISTERS_reg_31_24_inst : DFF_X1 port map( D => n8978, CK => CLK, Q => 
                           n15573, QN => n912);
   REGISTERS_reg_30_31_inst : DFF_X1 port map( D => n9017, CK => CLK, Q => 
                           n15574, QN => n5693);
   REGISTERS_reg_30_30_inst : DFF_X1 port map( D => n9016, CK => CLK, Q => 
                           n15575, QN => n5683);
   REGISTERS_reg_30_29_inst : DFF_X1 port map( D => n9015, CK => CLK, Q => 
                           n15576, QN => n5673);
   REGISTERS_reg_30_28_inst : DFF_X1 port map( D => n9014, CK => CLK, Q => 
                           n15577, QN => n5663);
   REGISTERS_reg_30_27_inst : DFF_X1 port map( D => n9013, CK => CLK, Q => 
                           n15578, QN => n5653);
   REGISTERS_reg_30_26_inst : DFF_X1 port map( D => n9012, CK => CLK, Q => 
                           n15579, QN => n5643);
   REGISTERS_reg_30_25_inst : DFF_X1 port map( D => n9011, CK => CLK, Q => 
                           n15580, QN => n5633);
   REGISTERS_reg_30_24_inst : DFF_X1 port map( D => n9010, CK => CLK, Q => 
                           n15581, QN => n5623);
   REGISTERS_reg_29_31_inst : DFF_X1 port map( D => n9049, CK => CLK, Q => 
                           n15790, QN => n5692);
   REGISTERS_reg_29_30_inst : DFF_X1 port map( D => n9048, CK => CLK, Q => 
                           n15791, QN => n5682);
   REGISTERS_reg_29_29_inst : DFF_X1 port map( D => n9047, CK => CLK, Q => 
                           n15792, QN => n5672);
   REGISTERS_reg_29_28_inst : DFF_X1 port map( D => n9046, CK => CLK, Q => 
                           n15793, QN => n5662);
   REGISTERS_reg_29_27_inst : DFF_X1 port map( D => n9045, CK => CLK, Q => 
                           n15794, QN => n5652);
   REGISTERS_reg_29_26_inst : DFF_X1 port map( D => n9044, CK => CLK, Q => 
                           n15795, QN => n5642);
   REGISTERS_reg_29_25_inst : DFF_X1 port map( D => n9043, CK => CLK, Q => 
                           n15796, QN => n5632);
   REGISTERS_reg_29_24_inst : DFF_X1 port map( D => n9042, CK => CLK, Q => 
                           n15797, QN => n5622);
   REGISTERS_reg_23_31_inst : DFF_X1 port map( D => n9241, CK => CLK, Q => 
                           n14461, QN => n6997);
   REGISTERS_reg_23_30_inst : DFF_X1 port map( D => n9240, CK => CLK, Q => 
                           n14462, QN => n6996);
   REGISTERS_reg_23_29_inst : DFF_X1 port map( D => n9239, CK => CLK, Q => 
                           n14463, QN => n6995);
   REGISTERS_reg_23_28_inst : DFF_X1 port map( D => n9238, CK => CLK, Q => 
                           n14464, QN => n6994);
   REGISTERS_reg_23_27_inst : DFF_X1 port map( D => n9237, CK => CLK, Q => 
                           n14465, QN => n6993);
   REGISTERS_reg_23_26_inst : DFF_X1 port map( D => n9236, CK => CLK, Q => 
                           n14466, QN => n6992);
   REGISTERS_reg_23_25_inst : DFF_X1 port map( D => n9235, CK => CLK, Q => 
                           n14467, QN => n6991);
   REGISTERS_reg_23_24_inst : DFF_X1 port map( D => n9234, CK => CLK, Q => 
                           n14468, QN => n6990);
   REGISTERS_reg_22_31_inst : DFF_X1 port map( D => n9273, CK => CLK, Q => 
                           n15582, QN => n873);
   REGISTERS_reg_22_30_inst : DFF_X1 port map( D => n9272, CK => CLK, Q => 
                           n15583, QN => n874);
   REGISTERS_reg_22_29_inst : DFF_X1 port map( D => n9271, CK => CLK, Q => 
                           n15584, QN => n875);
   REGISTERS_reg_22_28_inst : DFF_X1 port map( D => n9270, CK => CLK, Q => 
                           n15585, QN => n876);
   REGISTERS_reg_22_27_inst : DFF_X1 port map( D => n9269, CK => CLK, Q => 
                           n15586, QN => n877);
   REGISTERS_reg_22_26_inst : DFF_X1 port map( D => n9268, CK => CLK, Q => 
                           n15587, QN => n878);
   REGISTERS_reg_22_25_inst : DFF_X1 port map( D => n9267, CK => CLK, Q => 
                           n15588, QN => n879);
   REGISTERS_reg_22_24_inst : DFF_X1 port map( D => n9266, CK => CLK, Q => 
                           n15589, QN => n880);
   REGISTERS_reg_20_31_inst : DFF_X1 port map( D => n9337, CK => CLK, Q => 
                           n15862, QN => n5824);
   REGISTERS_reg_20_30_inst : DFF_X1 port map( D => n9336, CK => CLK, Q => 
                           n15863, QN => n5820);
   REGISTERS_reg_20_29_inst : DFF_X1 port map( D => n9335, CK => CLK, Q => 
                           n15864, QN => n5816);
   REGISTERS_reg_20_28_inst : DFF_X1 port map( D => n9334, CK => CLK, Q => 
                           n15865, QN => n5812);
   REGISTERS_reg_20_27_inst : DFF_X1 port map( D => n9333, CK => CLK, Q => 
                           n15866, QN => n5808);
   REGISTERS_reg_20_26_inst : DFF_X1 port map( D => n9332, CK => CLK, Q => 
                           n15867, QN => n5804);
   REGISTERS_reg_20_25_inst : DFF_X1 port map( D => n9331, CK => CLK, Q => 
                           n15868, QN => n5800);
   REGISTERS_reg_20_24_inst : DFF_X1 port map( D => n9330, CK => CLK, Q => 
                           n15869, QN => n5796);
   REGISTERS_reg_14_31_inst : DFF_X1 port map( D => n9529, CK => CLK, Q => 
                           n14248, QN => n7013);
   REGISTERS_reg_14_30_inst : DFF_X1 port map( D => n9528, CK => CLK, Q => 
                           n14249, QN => n7012);
   REGISTERS_reg_14_29_inst : DFF_X1 port map( D => n9527, CK => CLK, Q => 
                           n14250, QN => n7011);
   REGISTERS_reg_14_28_inst : DFF_X1 port map( D => n9526, CK => CLK, Q => 
                           n14251, QN => n7010);
   REGISTERS_reg_14_27_inst : DFF_X1 port map( D => n9525, CK => CLK, Q => 
                           n14252, QN => n7009);
   REGISTERS_reg_14_26_inst : DFF_X1 port map( D => n9524, CK => CLK, Q => 
                           n14253, QN => n7008);
   REGISTERS_reg_14_25_inst : DFF_X1 port map( D => n9523, CK => CLK, Q => 
                           n14254, QN => n7007);
   REGISTERS_reg_14_24_inst : DFF_X1 port map( D => n9522, CK => CLK, Q => 
                           n14255, QN => n7006);
   REGISTERS_reg_13_31_inst : DFF_X1 port map( D => n9561, CK => CLK, Q => 
                           n15590, QN => n841);
   REGISTERS_reg_13_30_inst : DFF_X1 port map( D => n9560, CK => CLK, Q => 
                           n15591, QN => n842);
   REGISTERS_reg_13_29_inst : DFF_X1 port map( D => n9559, CK => CLK, Q => 
                           n15592, QN => n843);
   REGISTERS_reg_13_28_inst : DFF_X1 port map( D => n9558, CK => CLK, Q => 
                           n15593, QN => n844);
   REGISTERS_reg_13_27_inst : DFF_X1 port map( D => n9557, CK => CLK, Q => 
                           n15594, QN => n845);
   REGISTERS_reg_13_26_inst : DFF_X1 port map( D => n9556, CK => CLK, Q => 
                           n15595, QN => n846);
   REGISTERS_reg_13_25_inst : DFF_X1 port map( D => n9555, CK => CLK, Q => 
                           n15596, QN => n847);
   REGISTERS_reg_13_24_inst : DFF_X1 port map( D => n9554, CK => CLK, Q => 
                           n15597, QN => n848);
   REGISTERS_reg_5_31_inst : DFF_X1 port map( D => n9817, CK => CLK, Q => 
                           n14076, QN => n7021);
   REGISTERS_reg_5_30_inst : DFF_X1 port map( D => n9816, CK => CLK, Q => 
                           n14077, QN => n7020);
   REGISTERS_reg_5_29_inst : DFF_X1 port map( D => n9815, CK => CLK, Q => 
                           n14078, QN => n7019);
   REGISTERS_reg_5_28_inst : DFF_X1 port map( D => n9814, CK => CLK, Q => 
                           n14079, QN => n7018);
   REGISTERS_reg_5_27_inst : DFF_X1 port map( D => n9813, CK => CLK, Q => 
                           n14080, QN => n7017);
   REGISTERS_reg_5_26_inst : DFF_X1 port map( D => n9812, CK => CLK, Q => 
                           n14081, QN => n7016);
   REGISTERS_reg_5_25_inst : DFF_X1 port map( D => n9811, CK => CLK, Q => 
                           n14082, QN => n7015);
   REGISTERS_reg_5_24_inst : DFF_X1 port map( D => n9810, CK => CLK, Q => 
                           n14083, QN => n7014);
   REGISTERS_reg_4_31_inst : DFF_X1 port map( D => n9849, CK => CLK, Q => 
                           n15598, QN => n809);
   REGISTERS_reg_4_30_inst : DFF_X1 port map( D => n9848, CK => CLK, Q => 
                           n15599, QN => n810);
   REGISTERS_reg_4_29_inst : DFF_X1 port map( D => n9847, CK => CLK, Q => 
                           n15600, QN => n811);
   REGISTERS_reg_4_28_inst : DFF_X1 port map( D => n9846, CK => CLK, Q => 
                           n15601, QN => n812);
   REGISTERS_reg_4_27_inst : DFF_X1 port map( D => n9845, CK => CLK, Q => 
                           n15602, QN => n813);
   REGISTERS_reg_4_26_inst : DFF_X1 port map( D => n9844, CK => CLK, Q => 
                           n15603, QN => n814);
   REGISTERS_reg_4_25_inst : DFF_X1 port map( D => n9843, CK => CLK, Q => 
                           n15604, QN => n815);
   REGISTERS_reg_4_24_inst : DFF_X1 port map( D => n9842, CK => CLK, Q => 
                           n15605, QN => n816);
   REGISTERS_reg_39_30_inst : DFF_X1 port map( D => n8728, CK => CLK, Q => 
                           n15620, QN => n5819);
   REGISTERS_reg_39_29_inst : DFF_X1 port map( D => n8727, CK => CLK, Q => 
                           n15621, QN => n5815);
   REGISTERS_reg_39_28_inst : DFF_X1 port map( D => n8726, CK => CLK, Q => 
                           n15622, QN => n5811);
   REGISTERS_reg_39_27_inst : DFF_X1 port map( D => n8725, CK => CLK, Q => 
                           n15623, QN => n5807);
   REGISTERS_reg_39_26_inst : DFF_X1 port map( D => n8724, CK => CLK, Q => 
                           n15624, QN => n5803);
   REGISTERS_reg_39_25_inst : DFF_X1 port map( D => n8723, CK => CLK, Q => 
                           n15625, QN => n5799);
   REGISTERS_reg_39_24_inst : DFF_X1 port map( D => n8722, CK => CLK, Q => 
                           n15626, QN => n5795);
   REGISTERS_reg_21_29_inst : DFF_X1 port map( D => n9303, CK => CLK, Q => 
                           n15627, QN => n5817);
   REGISTERS_reg_21_28_inst : DFF_X1 port map( D => n9302, CK => CLK, Q => 
                           n15628, QN => n5813);
   REGISTERS_reg_21_27_inst : DFF_X1 port map( D => n9301, CK => CLK, Q => 
                           n15629, QN => n5809);
   REGISTERS_reg_21_26_inst : DFF_X1 port map( D => n9300, CK => CLK, Q => 
                           n15630, QN => n5805);
   REGISTERS_reg_21_25_inst : DFF_X1 port map( D => n9299, CK => CLK, Q => 
                           n15631, QN => n5801);
   REGISTERS_reg_21_24_inst : DFF_X1 port map( D => n9298, CK => CLK, Q => 
                           n15632, QN => n5797);
   REGISTERS_reg_68_23_inst : DFF_X1 port map( D => n7793, CK => CLK, Q => 
                           n15438, QN => n6965);
   REGISTERS_reg_68_22_inst : DFF_X1 port map( D => n7792, CK => CLK, Q => 
                           n15439, QN => n6964);
   REGISTERS_reg_68_21_inst : DFF_X1 port map( D => n7791, CK => CLK, Q => 
                           n15440, QN => n6963);
   REGISTERS_reg_68_20_inst : DFF_X1 port map( D => n7790, CK => CLK, Q => 
                           n15441, QN => n6962);
   REGISTERS_reg_68_19_inst : DFF_X1 port map( D => n7789, CK => CLK, Q => 
                           n15442, QN => n6961);
   REGISTERS_reg_68_18_inst : DFF_X1 port map( D => n7788, CK => CLK, Q => 
                           n15443, QN => n6960);
   REGISTERS_reg_68_17_inst : DFF_X1 port map( D => n7787, CK => CLK, Q => 
                           n15444, QN => n6959);
   REGISTERS_reg_68_16_inst : DFF_X1 port map( D => n7786, CK => CLK, Q => 
                           n15445, QN => n6958);
   REGISTERS_reg_68_15_inst : DFF_X1 port map( D => n7785, CK => CLK, Q => 
                           n15446, QN => n6957);
   REGISTERS_reg_68_14_inst : DFF_X1 port map( D => n7784, CK => CLK, Q => 
                           n15447, QN => n6956);
   REGISTERS_reg_68_13_inst : DFF_X1 port map( D => n7783, CK => CLK, Q => 
                           n15448, QN => n6955);
   REGISTERS_reg_68_12_inst : DFF_X1 port map( D => n7782, CK => CLK, Q => 
                           n15449, QN => n6954);
   REGISTERS_reg_68_11_inst : DFF_X1 port map( D => n7781, CK => CLK, Q => 
                           n15450, QN => n6953);
   REGISTERS_reg_68_10_inst : DFF_X1 port map( D => n7780, CK => CLK, Q => 
                           n15451, QN => n6952);
   REGISTERS_reg_68_9_inst : DFF_X1 port map( D => n7779, CK => CLK, Q => 
                           n15452, QN => n6951);
   REGISTERS_reg_68_8_inst : DFF_X1 port map( D => n7778, CK => CLK, Q => 
                           n15453, QN => n6950);
   REGISTERS_reg_68_7_inst : DFF_X1 port map( D => n7777, CK => CLK, Q => 
                           n15454, QN => n6949);
   REGISTERS_reg_68_6_inst : DFF_X1 port map( D => n7776, CK => CLK, Q => 
                           n15455, QN => n6948);
   REGISTERS_reg_68_5_inst : DFF_X1 port map( D => n7775, CK => CLK, Q => 
                           n15456, QN => n6947);
   REGISTERS_reg_68_4_inst : DFF_X1 port map( D => n7774, CK => CLK, Q => 
                           n15457, QN => n6946);
   REGISTERS_reg_68_3_inst : DFF_X1 port map( D => n7773, CK => CLK, Q => 
                           n15458, QN => n6945);
   REGISTERS_reg_68_2_inst : DFF_X1 port map( D => n7772, CK => CLK, Q => 
                           n15459, QN => n6944);
   REGISTERS_reg_68_1_inst : DFF_X1 port map( D => n7771, CK => CLK, Q => 
                           n15460, QN => n6943);
   REGISTERS_reg_68_0_inst : DFF_X1 port map( D => n7770, CK => CLK, Q => 
                           n15461, QN => n6942);
   REGISTERS_reg_67_23_inst : DFF_X1 port map( D => n7825, CK => CLK, Q => 
                           n15406, QN => n7183);
   REGISTERS_reg_67_22_inst : DFF_X1 port map( D => n7824, CK => CLK, Q => 
                           n15407, QN => n7182);
   REGISTERS_reg_67_21_inst : DFF_X1 port map( D => n7823, CK => CLK, Q => 
                           n15408, QN => n7181);
   REGISTERS_reg_67_20_inst : DFF_X1 port map( D => n7822, CK => CLK, Q => 
                           n15409, QN => n7180);
   REGISTERS_reg_67_19_inst : DFF_X1 port map( D => n7821, CK => CLK, Q => 
                           n15410, QN => n7179);
   REGISTERS_reg_67_18_inst : DFF_X1 port map( D => n7820, CK => CLK, Q => 
                           n15411, QN => n7178);
   REGISTERS_reg_67_17_inst : DFF_X1 port map( D => n7819, CK => CLK, Q => 
                           n15412, QN => n7177);
   REGISTERS_reg_67_16_inst : DFF_X1 port map( D => n7818, CK => CLK, Q => 
                           n15413, QN => n7176);
   REGISTERS_reg_67_15_inst : DFF_X1 port map( D => n7817, CK => CLK, Q => 
                           n15414, QN => n7175);
   REGISTERS_reg_67_14_inst : DFF_X1 port map( D => n7816, CK => CLK, Q => 
                           n15415, QN => n7174);
   REGISTERS_reg_67_13_inst : DFF_X1 port map( D => n7815, CK => CLK, Q => 
                           n15416, QN => n7173);
   REGISTERS_reg_67_12_inst : DFF_X1 port map( D => n7814, CK => CLK, Q => 
                           n15417, QN => n7172);
   REGISTERS_reg_67_11_inst : DFF_X1 port map( D => n7813, CK => CLK, Q => 
                           n15418, QN => n7171);
   REGISTERS_reg_67_10_inst : DFF_X1 port map( D => n7812, CK => CLK, Q => 
                           n15419, QN => n7170);
   REGISTERS_reg_67_9_inst : DFF_X1 port map( D => n7811, CK => CLK, Q => 
                           n15420, QN => n7169);
   REGISTERS_reg_67_8_inst : DFF_X1 port map( D => n7810, CK => CLK, Q => 
                           n15421, QN => n7168);
   REGISTERS_reg_67_7_inst : DFF_X1 port map( D => n7809, CK => CLK, Q => 
                           n15422, QN => n7167);
   REGISTERS_reg_67_6_inst : DFF_X1 port map( D => n7808, CK => CLK, Q => 
                           n15423, QN => n7166);
   REGISTERS_reg_67_5_inst : DFF_X1 port map( D => n7807, CK => CLK, Q => 
                           n15424, QN => n7165);
   REGISTERS_reg_67_4_inst : DFF_X1 port map( D => n7806, CK => CLK, Q => 
                           n15425, QN => n7164);
   REGISTERS_reg_67_3_inst : DFF_X1 port map( D => n7805, CK => CLK, Q => 
                           n15426, QN => n7163);
   REGISTERS_reg_67_2_inst : DFF_X1 port map( D => n7804, CK => CLK, Q => 
                           n15427, QN => n7162);
   REGISTERS_reg_67_1_inst : DFF_X1 port map( D => n7803, CK => CLK, Q => 
                           n15428, QN => n7161);
   REGISTERS_reg_67_0_inst : DFF_X1 port map( D => n7802, CK => CLK, Q => 
                           n15429, QN => n7160);
   REGISTERS_reg_63_23_inst : DFF_X1 port map( D => n7953, CK => CLK, Q => 
                           n15310, QN => n7215);
   REGISTERS_reg_63_22_inst : DFF_X1 port map( D => n7952, CK => CLK, Q => 
                           n15311, QN => n7214);
   REGISTERS_reg_63_21_inst : DFF_X1 port map( D => n7951, CK => CLK, Q => 
                           n15312, QN => n7213);
   REGISTERS_reg_63_20_inst : DFF_X1 port map( D => n7950, CK => CLK, Q => 
                           n15313, QN => n7212);
   REGISTERS_reg_63_19_inst : DFF_X1 port map( D => n7949, CK => CLK, Q => 
                           n15314, QN => n7211);
   REGISTERS_reg_63_18_inst : DFF_X1 port map( D => n7948, CK => CLK, Q => 
                           n15315, QN => n7210);
   REGISTERS_reg_63_17_inst : DFF_X1 port map( D => n7947, CK => CLK, Q => 
                           n15316, QN => n7209);
   REGISTERS_reg_63_16_inst : DFF_X1 port map( D => n7946, CK => CLK, Q => 
                           n15317, QN => n7208);
   REGISTERS_reg_63_15_inst : DFF_X1 port map( D => n7945, CK => CLK, Q => 
                           n15318, QN => n7207);
   REGISTERS_reg_63_14_inst : DFF_X1 port map( D => n7944, CK => CLK, Q => 
                           n15319, QN => n7206);
   REGISTERS_reg_63_13_inst : DFF_X1 port map( D => n7943, CK => CLK, Q => 
                           n15320, QN => n7205);
   REGISTERS_reg_63_12_inst : DFF_X1 port map( D => n7942, CK => CLK, Q => 
                           n15321, QN => n7204);
   REGISTERS_reg_63_11_inst : DFF_X1 port map( D => n7941, CK => CLK, Q => 
                           n15322, QN => n7203);
   REGISTERS_reg_63_10_inst : DFF_X1 port map( D => n7940, CK => CLK, Q => 
                           n15323, QN => n7202);
   REGISTERS_reg_63_9_inst : DFF_X1 port map( D => n7939, CK => CLK, Q => 
                           n15324, QN => n7201);
   REGISTERS_reg_63_8_inst : DFF_X1 port map( D => n7938, CK => CLK, Q => 
                           n15325, QN => n7200);
   REGISTERS_reg_63_7_inst : DFF_X1 port map( D => n7937, CK => CLK, Q => 
                           n15326, QN => n7199);
   REGISTERS_reg_63_6_inst : DFF_X1 port map( D => n7936, CK => CLK, Q => 
                           n15327, QN => n7198);
   REGISTERS_reg_63_5_inst : DFF_X1 port map( D => n7935, CK => CLK, Q => 
                           n15328, QN => n7197);
   REGISTERS_reg_63_4_inst : DFF_X1 port map( D => n7934, CK => CLK, Q => 
                           n15329, QN => n7196);
   REGISTERS_reg_63_3_inst : DFF_X1 port map( D => n7933, CK => CLK, Q => 
                           n15330, QN => n7195);
   REGISTERS_reg_63_2_inst : DFF_X1 port map( D => n7932, CK => CLK, Q => 
                           n15331, QN => n7194);
   REGISTERS_reg_63_1_inst : DFF_X1 port map( D => n7931, CK => CLK, Q => 
                           n15332, QN => n7193);
   REGISTERS_reg_63_0_inst : DFF_X1 port map( D => n7930, CK => CLK, Q => 
                           n15333, QN => n7192);
   REGISTERS_reg_58_23_inst : DFF_X1 port map( D => n8113, CK => CLK, Q => 
                           n15182, QN => n7247);
   REGISTERS_reg_58_22_inst : DFF_X1 port map( D => n8112, CK => CLK, Q => 
                           n15183, QN => n7246);
   REGISTERS_reg_58_21_inst : DFF_X1 port map( D => n8111, CK => CLK, Q => 
                           n15184, QN => n7245);
   REGISTERS_reg_58_20_inst : DFF_X1 port map( D => n8110, CK => CLK, Q => 
                           n15185, QN => n7244);
   REGISTERS_reg_58_19_inst : DFF_X1 port map( D => n8109, CK => CLK, Q => 
                           n15186, QN => n7243);
   REGISTERS_reg_58_18_inst : DFF_X1 port map( D => n8108, CK => CLK, Q => 
                           n15187, QN => n7242);
   REGISTERS_reg_58_17_inst : DFF_X1 port map( D => n8107, CK => CLK, Q => 
                           n15188, QN => n7241);
   REGISTERS_reg_58_16_inst : DFF_X1 port map( D => n8106, CK => CLK, Q => 
                           n15189, QN => n7240);
   REGISTERS_reg_58_15_inst : DFF_X1 port map( D => n8105, CK => CLK, Q => 
                           n15190, QN => n7239);
   REGISTERS_reg_58_14_inst : DFF_X1 port map( D => n8104, CK => CLK, Q => 
                           n15191, QN => n7238);
   REGISTERS_reg_58_13_inst : DFF_X1 port map( D => n8103, CK => CLK, Q => 
                           n15192, QN => n7237);
   REGISTERS_reg_58_12_inst : DFF_X1 port map( D => n8102, CK => CLK, Q => 
                           n15193, QN => n7236);
   REGISTERS_reg_58_11_inst : DFF_X1 port map( D => n8101, CK => CLK, Q => 
                           n15194, QN => n7235);
   REGISTERS_reg_58_10_inst : DFF_X1 port map( D => n8100, CK => CLK, Q => 
                           n15195, QN => n7234);
   REGISTERS_reg_58_9_inst : DFF_X1 port map( D => n8099, CK => CLK, Q => 
                           n15196, QN => n7233);
   REGISTERS_reg_58_8_inst : DFF_X1 port map( D => n8098, CK => CLK, Q => 
                           n15197, QN => n7232);
   REGISTERS_reg_58_7_inst : DFF_X1 port map( D => n8097, CK => CLK, Q => 
                           n15198, QN => n7231);
   REGISTERS_reg_58_6_inst : DFF_X1 port map( D => n8096, CK => CLK, Q => 
                           n15199, QN => n7230);
   REGISTERS_reg_58_5_inst : DFF_X1 port map( D => n8095, CK => CLK, Q => 
                           n15200, QN => n7229);
   REGISTERS_reg_58_4_inst : DFF_X1 port map( D => n8094, CK => CLK, Q => 
                           n15201, QN => n7228);
   REGISTERS_reg_58_3_inst : DFF_X1 port map( D => n8093, CK => CLK, Q => 
                           n15202, QN => n7227);
   REGISTERS_reg_58_2_inst : DFF_X1 port map( D => n8092, CK => CLK, Q => 
                           n15203, QN => n7226);
   REGISTERS_reg_58_1_inst : DFF_X1 port map( D => n8091, CK => CLK, Q => 
                           n15204, QN => n7225);
   REGISTERS_reg_58_0_inst : DFF_X1 port map( D => n8090, CK => CLK, Q => 
                           n15205, QN => n7224);
   REGISTERS_reg_50_23_inst : DFF_X1 port map( D => n8369, CK => CLK, Q => 
                           n14990, QN => n7045);
   REGISTERS_reg_50_22_inst : DFF_X1 port map( D => n8368, CK => CLK, Q => 
                           n14991, QN => n7044);
   REGISTERS_reg_50_21_inst : DFF_X1 port map( D => n8367, CK => CLK, Q => 
                           n14992, QN => n7043);
   REGISTERS_reg_50_20_inst : DFF_X1 port map( D => n8366, CK => CLK, Q => 
                           n14993, QN => n7042);
   REGISTERS_reg_50_19_inst : DFF_X1 port map( D => n8365, CK => CLK, Q => 
                           n14994, QN => n7041);
   REGISTERS_reg_50_18_inst : DFF_X1 port map( D => n8364, CK => CLK, Q => 
                           n14995, QN => n7040);
   REGISTERS_reg_50_17_inst : DFF_X1 port map( D => n8363, CK => CLK, Q => 
                           n14996, QN => n7039);
   REGISTERS_reg_50_16_inst : DFF_X1 port map( D => n8362, CK => CLK, Q => 
                           n14997, QN => n7038);
   REGISTERS_reg_50_15_inst : DFF_X1 port map( D => n8361, CK => CLK, Q => 
                           n14998, QN => n7037);
   REGISTERS_reg_50_14_inst : DFF_X1 port map( D => n8360, CK => CLK, Q => 
                           n14999, QN => n7036);
   REGISTERS_reg_50_13_inst : DFF_X1 port map( D => n8359, CK => CLK, Q => 
                           n15000, QN => n7035);
   REGISTERS_reg_50_12_inst : DFF_X1 port map( D => n8358, CK => CLK, Q => 
                           n15001, QN => n7034);
   REGISTERS_reg_50_11_inst : DFF_X1 port map( D => n8357, CK => CLK, Q => 
                           n15002, QN => n7033);
   REGISTERS_reg_50_10_inst : DFF_X1 port map( D => n8356, CK => CLK, Q => 
                           n15003, QN => n7032);
   REGISTERS_reg_50_9_inst : DFF_X1 port map( D => n8355, CK => CLK, Q => 
                           n15004, QN => n7031);
   REGISTERS_reg_50_8_inst : DFF_X1 port map( D => n8354, CK => CLK, Q => 
                           n15005, QN => n7030);
   REGISTERS_reg_50_7_inst : DFF_X1 port map( D => n8353, CK => CLK, Q => 
                           n15006, QN => n7029);
   REGISTERS_reg_50_6_inst : DFF_X1 port map( D => n8352, CK => CLK, Q => 
                           n15007, QN => n7028);
   REGISTERS_reg_50_5_inst : DFF_X1 port map( D => n8351, CK => CLK, Q => 
                           n15008, QN => n7027);
   REGISTERS_reg_50_4_inst : DFF_X1 port map( D => n8350, CK => CLK, Q => 
                           n15009, QN => n7026);
   REGISTERS_reg_50_3_inst : DFF_X1 port map( D => n8349, CK => CLK, Q => 
                           n15010, QN => n7025);
   REGISTERS_reg_50_2_inst : DFF_X1 port map( D => n8348, CK => CLK, Q => 
                           n15011, QN => n7024);
   REGISTERS_reg_50_1_inst : DFF_X1 port map( D => n8347, CK => CLK, Q => 
                           n15012, QN => n7023);
   REGISTERS_reg_50_0_inst : DFF_X1 port map( D => n8346, CK => CLK, Q => 
                           n15013, QN => n7022);
   REGISTERS_reg_49_23_inst : DFF_X1 port map( D => n8401, CK => CLK, Q => 
                           n15642, QN => n977);
   REGISTERS_reg_49_22_inst : DFF_X1 port map( D => n8400, CK => CLK, Q => 
                           n15643, QN => n978);
   REGISTERS_reg_49_21_inst : DFF_X1 port map( D => n8399, CK => CLK, Q => 
                           n15644, QN => n979);
   REGISTERS_reg_49_20_inst : DFF_X1 port map( D => n8398, CK => CLK, Q => 
                           n15645, QN => n980);
   REGISTERS_reg_49_19_inst : DFF_X1 port map( D => n8397, CK => CLK, Q => 
                           n15646, QN => n981);
   REGISTERS_reg_49_18_inst : DFF_X1 port map( D => n8396, CK => CLK, Q => 
                           n15647, QN => n982);
   REGISTERS_reg_49_17_inst : DFF_X1 port map( D => n8395, CK => CLK, Q => 
                           n15648, QN => n983);
   REGISTERS_reg_49_16_inst : DFF_X1 port map( D => n8394, CK => CLK, Q => 
                           n15649, QN => n984);
   REGISTERS_reg_49_15_inst : DFF_X1 port map( D => n8393, CK => CLK, Q => 
                           n15650, QN => n985);
   REGISTERS_reg_49_14_inst : DFF_X1 port map( D => n8392, CK => CLK, Q => 
                           n15651, QN => n986);
   REGISTERS_reg_49_13_inst : DFF_X1 port map( D => n8391, CK => CLK, Q => 
                           n15652, QN => n987);
   REGISTERS_reg_49_12_inst : DFF_X1 port map( D => n8390, CK => CLK, Q => 
                           n15653, QN => n988);
   REGISTERS_reg_49_11_inst : DFF_X1 port map( D => n8389, CK => CLK, Q => 
                           n15654, QN => n989);
   REGISTERS_reg_49_10_inst : DFF_X1 port map( D => n8388, CK => CLK, Q => 
                           n15655, QN => n990);
   REGISTERS_reg_49_9_inst : DFF_X1 port map( D => n8387, CK => CLK, Q => 
                           n15656, QN => n991);
   REGISTERS_reg_49_8_inst : DFF_X1 port map( D => n8386, CK => CLK, Q => 
                           n15657, QN => n992);
   REGISTERS_reg_49_7_inst : DFF_X1 port map( D => n8385, CK => CLK, Q => 
                           n15606, QN => n993);
   REGISTERS_reg_49_6_inst : DFF_X1 port map( D => n8384, CK => CLK, Q => 
                           n15607, QN => n994);
   REGISTERS_reg_49_5_inst : DFF_X1 port map( D => n8383, CK => CLK, Q => 
                           n15608, QN => n995);
   REGISTERS_reg_49_4_inst : DFF_X1 port map( D => n8382, CK => CLK, Q => 
                           n15609, QN => n996);
   REGISTERS_reg_49_3_inst : DFF_X1 port map( D => n8381, CK => CLK, Q => 
                           n15610, QN => n997);
   REGISTERS_reg_49_2_inst : DFF_X1 port map( D => n8380, CK => CLK, Q => 
                           n15611, QN => n998);
   REGISTERS_reg_49_1_inst : DFF_X1 port map( D => n8379, CK => CLK, Q => 
                           n15612, QN => n999);
   REGISTERS_reg_49_0_inst : DFF_X1 port map( D => n8378, CK => CLK, Q => 
                           n14981, QN => n7256);
   REGISTERS_reg_45_23_inst : DFF_X1 port map( D => n8529, CK => CLK, Q => 
                           n15658, QN => n643);
   REGISTERS_reg_45_22_inst : DFF_X1 port map( D => n8528, CK => CLK, Q => 
                           n15659, QN => n646);
   REGISTERS_reg_45_21_inst : DFF_X1 port map( D => n8527, CK => CLK, Q => 
                           n15660, QN => n649);
   REGISTERS_reg_45_20_inst : DFF_X1 port map( D => n8526, CK => CLK, Q => 
                           n15661, QN => n652);
   REGISTERS_reg_45_19_inst : DFF_X1 port map( D => n8525, CK => CLK, Q => 
                           n15662, QN => n655);
   REGISTERS_reg_45_18_inst : DFF_X1 port map( D => n8524, CK => CLK, Q => 
                           n15663, QN => n658);
   REGISTERS_reg_45_17_inst : DFF_X1 port map( D => n8523, CK => CLK, Q => 
                           n15664, QN => n661);
   REGISTERS_reg_45_16_inst : DFF_X1 port map( D => n8522, CK => CLK, Q => 
                           n15665, QN => n664);
   REGISTERS_reg_45_15_inst : DFF_X1 port map( D => n8521, CK => CLK, Q => 
                           n15666, QN => n667);
   REGISTERS_reg_45_14_inst : DFF_X1 port map( D => n8520, CK => CLK, Q => 
                           n15667, QN => n670);
   REGISTERS_reg_45_13_inst : DFF_X1 port map( D => n8519, CK => CLK, Q => 
                           n15668, QN => n673);
   REGISTERS_reg_45_12_inst : DFF_X1 port map( D => n8518, CK => CLK, Q => 
                           n15669, QN => n676);
   REGISTERS_reg_45_11_inst : DFF_X1 port map( D => n8517, CK => CLK, Q => 
                           n15670, QN => n679);
   REGISTERS_reg_45_10_inst : DFF_X1 port map( D => n8516, CK => CLK, Q => 
                           n15671, QN => n682);
   REGISTERS_reg_45_9_inst : DFF_X1 port map( D => n8515, CK => CLK, Q => 
                           n15672, QN => n685);
   REGISTERS_reg_45_8_inst : DFF_X1 port map( D => n8514, CK => CLK, Q => 
                           n15673, QN => n688);
   REGISTERS_reg_45_7_inst : DFF_X1 port map( D => n8513, CK => CLK, Q => 
                           n15674, QN => n691);
   REGISTERS_reg_45_6_inst : DFF_X1 port map( D => n8512, CK => CLK, Q => 
                           n15675, QN => n694);
   REGISTERS_reg_45_5_inst : DFF_X1 port map( D => n8511, CK => CLK, Q => 
                           n15676, QN => n697);
   REGISTERS_reg_45_4_inst : DFF_X1 port map( D => n8510, CK => CLK, Q => 
                           n15677, QN => n700);
   REGISTERS_reg_45_3_inst : DFF_X1 port map( D => n8509, CK => CLK, Q => 
                           n15678, QN => n703);
   REGISTERS_reg_45_2_inst : DFF_X1 port map( D => n8508, CK => CLK, Q => 
                           n15679, QN => n706);
   REGISTERS_reg_45_1_inst : DFF_X1 port map( D => n8507, CK => CLK, Q => 
                           n15680, QN => n709);
   REGISTERS_reg_45_0_inst : DFF_X1 port map( D => n8506, CK => CLK, Q => 
                           n15681, QN => n712);
   REGISTERS_reg_40_23_inst : DFF_X1 port map( D => n8689, CK => CLK, Q => 
                           n15682, QN => n945);
   REGISTERS_reg_40_22_inst : DFF_X1 port map( D => n8688, CK => CLK, Q => 
                           n15683, QN => n946);
   REGISTERS_reg_40_21_inst : DFF_X1 port map( D => n8687, CK => CLK, Q => 
                           n15684, QN => n947);
   REGISTERS_reg_40_20_inst : DFF_X1 port map( D => n8686, CK => CLK, Q => 
                           n15685, QN => n948);
   REGISTERS_reg_40_19_inst : DFF_X1 port map( D => n8685, CK => CLK, Q => 
                           n15686, QN => n949);
   REGISTERS_reg_40_18_inst : DFF_X1 port map( D => n8684, CK => CLK, Q => 
                           n15687, QN => n950);
   REGISTERS_reg_40_17_inst : DFF_X1 port map( D => n8683, CK => CLK, Q => 
                           n15688, QN => n951);
   REGISTERS_reg_40_16_inst : DFF_X1 port map( D => n8682, CK => CLK, Q => 
                           n15689, QN => n952);
   REGISTERS_reg_40_15_inst : DFF_X1 port map( D => n8681, CK => CLK, Q => 
                           n15690, QN => n953);
   REGISTERS_reg_40_14_inst : DFF_X1 port map( D => n8680, CK => CLK, Q => 
                           n15691, QN => n954);
   REGISTERS_reg_40_13_inst : DFF_X1 port map( D => n8679, CK => CLK, Q => 
                           n15692, QN => n955);
   REGISTERS_reg_40_12_inst : DFF_X1 port map( D => n8678, CK => CLK, Q => 
                           n15693, QN => n956);
   REGISTERS_reg_40_11_inst : DFF_X1 port map( D => n8677, CK => CLK, Q => 
                           n15694, QN => n957);
   REGISTERS_reg_40_10_inst : DFF_X1 port map( D => n8676, CK => CLK, Q => 
                           n15695, QN => n958);
   REGISTERS_reg_40_9_inst : DFF_X1 port map( D => n8675, CK => CLK, Q => 
                           n15696, QN => n959);
   REGISTERS_reg_40_8_inst : DFF_X1 port map( D => n8674, CK => CLK, Q => 
                           n15697, QN => n960);
   REGISTERS_reg_40_7_inst : DFF_X1 port map( D => n8673, CK => CLK, Q => 
                           n15698, QN => n961);
   REGISTERS_reg_40_6_inst : DFF_X1 port map( D => n8672, CK => CLK, Q => 
                           n15699, QN => n962);
   REGISTERS_reg_40_5_inst : DFF_X1 port map( D => n8671, CK => CLK, Q => 
                           n15700, QN => n963);
   REGISTERS_reg_40_4_inst : DFF_X1 port map( D => n8670, CK => CLK, Q => 
                           n15701, QN => n964);
   REGISTERS_reg_40_3_inst : DFF_X1 port map( D => n8669, CK => CLK, Q => 
                           n15702, QN => n965);
   REGISTERS_reg_40_2_inst : DFF_X1 port map( D => n8668, CK => CLK, Q => 
                           n15703, QN => n966);
   REGISTERS_reg_40_1_inst : DFF_X1 port map( D => n8667, CK => CLK, Q => 
                           n15704, QN => n967);
   REGISTERS_reg_40_0_inst : DFF_X1 port map( D => n8666, CK => CLK, Q => 
                           n15705, QN => n968);
   REGISTERS_reg_39_23_inst : DFF_X1 port map( D => n8721, CK => CLK, Q => 
                           n15706, QN => n5791);
   REGISTERS_reg_39_22_inst : DFF_X1 port map( D => n8720, CK => CLK, Q => 
                           n15707, QN => n5787);
   REGISTERS_reg_39_21_inst : DFF_X1 port map( D => n8719, CK => CLK, Q => 
                           n15708, QN => n5783);
   REGISTERS_reg_39_20_inst : DFF_X1 port map( D => n8718, CK => CLK, Q => 
                           n15709, QN => n5779);
   REGISTERS_reg_39_19_inst : DFF_X1 port map( D => n8717, CK => CLK, Q => 
                           n15710, QN => n5775);
   REGISTERS_reg_39_18_inst : DFF_X1 port map( D => n8716, CK => CLK, Q => 
                           n15711, QN => n5771);
   REGISTERS_reg_39_17_inst : DFF_X1 port map( D => n8715, CK => CLK, Q => 
                           n15712, QN => n5767);
   REGISTERS_reg_39_16_inst : DFF_X1 port map( D => n8714, CK => CLK, Q => 
                           n15713, QN => n5763);
   REGISTERS_reg_39_15_inst : DFF_X1 port map( D => n8713, CK => CLK, Q => 
                           n15714, QN => n5759);
   REGISTERS_reg_39_14_inst : DFF_X1 port map( D => n8712, CK => CLK, Q => 
                           n15715, QN => n5755);
   REGISTERS_reg_39_13_inst : DFF_X1 port map( D => n8711, CK => CLK, Q => 
                           n15716, QN => n5751);
   REGISTERS_reg_39_12_inst : DFF_X1 port map( D => n8710, CK => CLK, Q => 
                           n15717, QN => n5747);
   REGISTERS_reg_39_11_inst : DFF_X1 port map( D => n8709, CK => CLK, Q => 
                           n15718, QN => n5743);
   REGISTERS_reg_39_10_inst : DFF_X1 port map( D => n8708, CK => CLK, Q => 
                           n15719, QN => n5739);
   REGISTERS_reg_39_9_inst : DFF_X1 port map( D => n8707, CK => CLK, Q => 
                           n15720, QN => n5735);
   REGISTERS_reg_39_8_inst : DFF_X1 port map( D => n8706, CK => CLK, Q => 
                           n15721, QN => n5731);
   REGISTERS_reg_39_7_inst : DFF_X1 port map( D => n8705, CK => CLK, Q => 
                           n15722, QN => n5727);
   REGISTERS_reg_39_6_inst : DFF_X1 port map( D => n8704, CK => CLK, Q => 
                           n15723, QN => n5723);
   REGISTERS_reg_39_5_inst : DFF_X1 port map( D => n8703, CK => CLK, Q => 
                           n15724, QN => n5719);
   REGISTERS_reg_39_4_inst : DFF_X1 port map( D => n8702, CK => CLK, Q => 
                           n15725, QN => n5715);
   REGISTERS_reg_39_3_inst : DFF_X1 port map( D => n8701, CK => CLK, Q => 
                           n15726, QN => n5711);
   REGISTERS_reg_39_2_inst : DFF_X1 port map( D => n8700, CK => CLK, Q => 
                           n15727, QN => n5707);
   REGISTERS_reg_39_1_inst : DFF_X1 port map( D => n8699, CK => CLK, Q => 
                           n15728, QN => n5703);
   REGISTERS_reg_39_0_inst : DFF_X1 port map( D => n8698, CK => CLK, Q => 
                           n15729, QN => n5699);
   REGISTERS_reg_38_31_inst : DFF_X1 port map( D => n8761, CK => CLK, Q => 
                           n15730, QN => n5822);
   REGISTERS_reg_38_30_inst : DFF_X1 port map( D => n8760, CK => CLK, Q => 
                           n15731, QN => n5818);
   REGISTERS_reg_38_29_inst : DFF_X1 port map( D => n8759, CK => CLK, Q => 
                           n15732, QN => n5814);
   REGISTERS_reg_38_28_inst : DFF_X1 port map( D => n8758, CK => CLK, Q => 
                           n15733, QN => n5810);
   REGISTERS_reg_38_27_inst : DFF_X1 port map( D => n8757, CK => CLK, Q => 
                           n15734, QN => n5806);
   REGISTERS_reg_38_26_inst : DFF_X1 port map( D => n8756, CK => CLK, Q => 
                           n15735, QN => n5802);
   REGISTERS_reg_38_25_inst : DFF_X1 port map( D => n8755, CK => CLK, Q => 
                           n15736, QN => n5798);
   REGISTERS_reg_38_24_inst : DFF_X1 port map( D => n8754, CK => CLK, Q => 
                           n15737, QN => n5794);
   REGISTERS_reg_38_23_inst : DFF_X1 port map( D => n8753, CK => CLK, Q => 
                           n15738, QN => n5790);
   REGISTERS_reg_38_22_inst : DFF_X1 port map( D => n8752, CK => CLK, Q => 
                           n15739, QN => n5786);
   REGISTERS_reg_38_21_inst : DFF_X1 port map( D => n8751, CK => CLK, Q => 
                           n15740, QN => n5782);
   REGISTERS_reg_38_20_inst : DFF_X1 port map( D => n8750, CK => CLK, Q => 
                           n15741, QN => n5778);
   REGISTERS_reg_32_23_inst : DFF_X1 port map( D => n8945, CK => CLK, Q => 
                           n14668, QN => n7069);
   REGISTERS_reg_32_22_inst : DFF_X1 port map( D => n8944, CK => CLK, Q => 
                           n14669, QN => n7068);
   REGISTERS_reg_32_21_inst : DFF_X1 port map( D => n8943, CK => CLK, Q => 
                           n14670, QN => n7067);
   REGISTERS_reg_32_20_inst : DFF_X1 port map( D => n8942, CK => CLK, Q => 
                           n14671, QN => n7066);
   REGISTERS_reg_32_19_inst : DFF_X1 port map( D => n8941, CK => CLK, Q => 
                           n14672, QN => n7065);
   REGISTERS_reg_32_18_inst : DFF_X1 port map( D => n8940, CK => CLK, Q => 
                           n14673, QN => n7064);
   REGISTERS_reg_32_17_inst : DFF_X1 port map( D => n8939, CK => CLK, Q => 
                           n14674, QN => n7063);
   REGISTERS_reg_32_16_inst : DFF_X1 port map( D => n8938, CK => CLK, Q => 
                           n14675, QN => n7062);
   REGISTERS_reg_32_15_inst : DFF_X1 port map( D => n8937, CK => CLK, Q => 
                           n14676, QN => n7061);
   REGISTERS_reg_32_14_inst : DFF_X1 port map( D => n8936, CK => CLK, Q => 
                           n14677, QN => n7060);
   REGISTERS_reg_32_13_inst : DFF_X1 port map( D => n8935, CK => CLK, Q => 
                           n14678, QN => n7059);
   REGISTERS_reg_32_12_inst : DFF_X1 port map( D => n8934, CK => CLK, Q => 
                           n14679, QN => n7058);
   REGISTERS_reg_32_11_inst : DFF_X1 port map( D => n8933, CK => CLK, Q => 
                           n14680, QN => n7057);
   REGISTERS_reg_32_10_inst : DFF_X1 port map( D => n8932, CK => CLK, Q => 
                           n14681, QN => n7056);
   REGISTERS_reg_32_9_inst : DFF_X1 port map( D => n8931, CK => CLK, Q => 
                           n14682, QN => n7055);
   REGISTERS_reg_32_8_inst : DFF_X1 port map( D => n8930, CK => CLK, Q => 
                           n14683, QN => n7054);
   REGISTERS_reg_32_7_inst : DFF_X1 port map( D => n8929, CK => CLK, Q => 
                           n14684, QN => n7053);
   REGISTERS_reg_32_6_inst : DFF_X1 port map( D => n8928, CK => CLK, Q => 
                           n14685, QN => n7052);
   REGISTERS_reg_32_5_inst : DFF_X1 port map( D => n8927, CK => CLK, Q => 
                           n14686, QN => n7051);
   REGISTERS_reg_32_4_inst : DFF_X1 port map( D => n8926, CK => CLK, Q => 
                           n14687, QN => n7050);
   REGISTERS_reg_32_3_inst : DFF_X1 port map( D => n8925, CK => CLK, Q => 
                           n14688, QN => n7049);
   REGISTERS_reg_32_2_inst : DFF_X1 port map( D => n8924, CK => CLK, Q => 
                           n14689, QN => n7048);
   REGISTERS_reg_32_1_inst : DFF_X1 port map( D => n8923, CK => CLK, Q => 
                           n14690, QN => n7047);
   REGISTERS_reg_32_0_inst : DFF_X1 port map( D => n8922, CK => CLK, Q => 
                           n14691, QN => n7046);
   REGISTERS_reg_31_23_inst : DFF_X1 port map( D => n8977, CK => CLK, Q => 
                           n15742, QN => n913);
   REGISTERS_reg_31_22_inst : DFF_X1 port map( D => n8976, CK => CLK, Q => 
                           n15743, QN => n914);
   REGISTERS_reg_31_21_inst : DFF_X1 port map( D => n8975, CK => CLK, Q => 
                           n15744, QN => n915);
   REGISTERS_reg_31_20_inst : DFF_X1 port map( D => n8974, CK => CLK, Q => 
                           n15745, QN => n916);
   REGISTERS_reg_31_19_inst : DFF_X1 port map( D => n8973, CK => CLK, Q => 
                           n15746, QN => n917);
   REGISTERS_reg_31_18_inst : DFF_X1 port map( D => n8972, CK => CLK, Q => 
                           n15747, QN => n918);
   REGISTERS_reg_31_17_inst : DFF_X1 port map( D => n8971, CK => CLK, Q => 
                           n15748, QN => n919);
   REGISTERS_reg_31_16_inst : DFF_X1 port map( D => n8970, CK => CLK, Q => 
                           n15749, QN => n920);
   REGISTERS_reg_31_15_inst : DFF_X1 port map( D => n8969, CK => CLK, Q => 
                           n15750, QN => n921);
   REGISTERS_reg_31_14_inst : DFF_X1 port map( D => n8968, CK => CLK, Q => 
                           n15751, QN => n922);
   REGISTERS_reg_31_13_inst : DFF_X1 port map( D => n8967, CK => CLK, Q => 
                           n15752, QN => n923);
   REGISTERS_reg_31_12_inst : DFF_X1 port map( D => n8966, CK => CLK, Q => 
                           n15753, QN => n924);
   REGISTERS_reg_31_11_inst : DFF_X1 port map( D => n8965, CK => CLK, Q => 
                           n15754, QN => n925);
   REGISTERS_reg_31_10_inst : DFF_X1 port map( D => n8964, CK => CLK, Q => 
                           n15755, QN => n926);
   REGISTERS_reg_31_9_inst : DFF_X1 port map( D => n8963, CK => CLK, Q => 
                           n15756, QN => n927);
   REGISTERS_reg_31_8_inst : DFF_X1 port map( D => n8962, CK => CLK, Q => 
                           n15757, QN => n928);
   REGISTERS_reg_31_7_inst : DFF_X1 port map( D => n8961, CK => CLK, Q => 
                           n15758, QN => n929);
   REGISTERS_reg_31_6_inst : DFF_X1 port map( D => n8960, CK => CLK, Q => 
                           n15759, QN => n930);
   REGISTERS_reg_31_5_inst : DFF_X1 port map( D => n8959, CK => CLK, Q => 
                           n15760, QN => n931);
   REGISTERS_reg_31_4_inst : DFF_X1 port map( D => n8958, CK => CLK, Q => 
                           n15761, QN => n932);
   REGISTERS_reg_31_3_inst : DFF_X1 port map( D => n8957, CK => CLK, Q => 
                           n15762, QN => n933);
   REGISTERS_reg_31_2_inst : DFF_X1 port map( D => n8956, CK => CLK, Q => 
                           n15763, QN => n934);
   REGISTERS_reg_31_1_inst : DFF_X1 port map( D => n8955, CK => CLK, Q => 
                           n15764, QN => n935);
   REGISTERS_reg_31_0_inst : DFF_X1 port map( D => n8954, CK => CLK, Q => 
                           n15765, QN => n936);
   REGISTERS_reg_30_23_inst : DFF_X1 port map( D => n9009, CK => CLK, Q => 
                           n15766, QN => n5613);
   REGISTERS_reg_30_22_inst : DFF_X1 port map( D => n9008, CK => CLK, Q => 
                           n15767, QN => n5603);
   REGISTERS_reg_30_21_inst : DFF_X1 port map( D => n9007, CK => CLK, Q => 
                           n15768, QN => n5593);
   REGISTERS_reg_30_20_inst : DFF_X1 port map( D => n9006, CK => CLK, Q => 
                           n15769, QN => n5583);
   REGISTERS_reg_30_19_inst : DFF_X1 port map( D => n9005, CK => CLK, Q => 
                           n15770, QN => n5573);
   REGISTERS_reg_30_18_inst : DFF_X1 port map( D => n9004, CK => CLK, Q => 
                           n15771, QN => n5563);
   REGISTERS_reg_30_17_inst : DFF_X1 port map( D => n9003, CK => CLK, Q => 
                           n15772, QN => n5553);
   REGISTERS_reg_30_16_inst : DFF_X1 port map( D => n9002, CK => CLK, Q => 
                           n15773, QN => n5543);
   REGISTERS_reg_30_15_inst : DFF_X1 port map( D => n9001, CK => CLK, Q => 
                           n15774, QN => n5533);
   REGISTERS_reg_30_14_inst : DFF_X1 port map( D => n9000, CK => CLK, Q => 
                           n15775, QN => n5523);
   REGISTERS_reg_30_13_inst : DFF_X1 port map( D => n8999, CK => CLK, Q => 
                           n15776, QN => n5513);
   REGISTERS_reg_30_12_inst : DFF_X1 port map( D => n8998, CK => CLK, Q => 
                           n15777, QN => n5503);
   REGISTERS_reg_30_11_inst : DFF_X1 port map( D => n8997, CK => CLK, Q => 
                           n15778, QN => n5493);
   REGISTERS_reg_30_10_inst : DFF_X1 port map( D => n8996, CK => CLK, Q => 
                           n15779, QN => n5483);
   REGISTERS_reg_30_9_inst : DFF_X1 port map( D => n8995, CK => CLK, Q => 
                           n15780, QN => n5473);
   REGISTERS_reg_30_8_inst : DFF_X1 port map( D => n8994, CK => CLK, Q => 
                           n15781, QN => n5463);
   REGISTERS_reg_30_7_inst : DFF_X1 port map( D => n8993, CK => CLK, Q => 
                           n15782, QN => n5453);
   REGISTERS_reg_30_6_inst : DFF_X1 port map( D => n8992, CK => CLK, Q => 
                           n15783, QN => n5443);
   REGISTERS_reg_30_5_inst : DFF_X1 port map( D => n8991, CK => CLK, Q => 
                           n15784, QN => n5433);
   REGISTERS_reg_30_4_inst : DFF_X1 port map( D => n8990, CK => CLK, Q => 
                           n15785, QN => n5423);
   REGISTERS_reg_30_3_inst : DFF_X1 port map( D => n8989, CK => CLK, Q => 
                           n15786, QN => n5413);
   REGISTERS_reg_30_2_inst : DFF_X1 port map( D => n8988, CK => CLK, Q => 
                           n15787, QN => n5403);
   REGISTERS_reg_30_1_inst : DFF_X1 port map( D => n8987, CK => CLK, Q => 
                           n15788, QN => n5393);
   REGISTERS_reg_30_0_inst : DFF_X1 port map( D => n8986, CK => CLK, Q => 
                           n15789, QN => n5383);
   REGISTERS_reg_29_23_inst : DFF_X1 port map( D => n9041, CK => CLK, Q => 
                           n15798, QN => n5612);
   REGISTERS_reg_29_22_inst : DFF_X1 port map( D => n9040, CK => CLK, Q => 
                           n15799, QN => n5602);
   REGISTERS_reg_29_21_inst : DFF_X1 port map( D => n9039, CK => CLK, Q => 
                           n15800, QN => n5592);
   REGISTERS_reg_29_20_inst : DFF_X1 port map( D => n9038, CK => CLK, Q => 
                           n15801, QN => n5582);
   REGISTERS_reg_29_19_inst : DFF_X1 port map( D => n9037, CK => CLK, Q => 
                           n15802, QN => n5572);
   REGISTERS_reg_29_18_inst : DFF_X1 port map( D => n9036, CK => CLK, Q => 
                           n15803, QN => n5562);
   REGISTERS_reg_29_17_inst : DFF_X1 port map( D => n9035, CK => CLK, Q => 
                           n15804, QN => n5552);
   REGISTERS_reg_29_16_inst : DFF_X1 port map( D => n9034, CK => CLK, Q => 
                           n15805, QN => n5542);
   REGISTERS_reg_29_15_inst : DFF_X1 port map( D => n9033, CK => CLK, Q => 
                           n15806, QN => n5532);
   REGISTERS_reg_29_14_inst : DFF_X1 port map( D => n9032, CK => CLK, Q => 
                           n15807, QN => n5522);
   REGISTERS_reg_29_13_inst : DFF_X1 port map( D => n9031, CK => CLK, Q => 
                           n15808, QN => n5512);
   REGISTERS_reg_29_12_inst : DFF_X1 port map( D => n9030, CK => CLK, Q => 
                           n15809, QN => n5502);
   REGISTERS_reg_29_11_inst : DFF_X1 port map( D => n9029, CK => CLK, Q => 
                           n15810, QN => n5492);
   REGISTERS_reg_29_10_inst : DFF_X1 port map( D => n9028, CK => CLK, Q => 
                           n15811, QN => n5482);
   REGISTERS_reg_29_9_inst : DFF_X1 port map( D => n9027, CK => CLK, Q => 
                           n15812, QN => n5472);
   REGISTERS_reg_29_8_inst : DFF_X1 port map( D => n9026, CK => CLK, Q => 
                           n15813, QN => n5462);
   REGISTERS_reg_29_7_inst : DFF_X1 port map( D => n9025, CK => CLK, Q => 
                           n15633, QN => n5452);
   REGISTERS_reg_29_6_inst : DFF_X1 port map( D => n9024, CK => CLK, Q => 
                           n14653, QN => n7159);
   REGISTERS_reg_29_5_inst : DFF_X1 port map( D => n9023, CK => CLK, Q => 
                           n14654, QN => n7158);
   REGISTERS_reg_29_4_inst : DFF_X1 port map( D => n9022, CK => CLK, Q => 
                           n14655, QN => n7157);
   REGISTERS_reg_29_3_inst : DFF_X1 port map( D => n9021, CK => CLK, Q => 
                           n14656, QN => n7156);
   REGISTERS_reg_29_2_inst : DFF_X1 port map( D => n9020, CK => CLK, Q => 
                           n14657, QN => n7155);
   REGISTERS_reg_29_1_inst : DFF_X1 port map( D => n9019, CK => CLK, Q => 
                           n14658, QN => n7154);
   REGISTERS_reg_29_0_inst : DFF_X1 port map( D => n9018, CK => CLK, Q => 
                           n14659, QN => n7153);
   REGISTERS_reg_23_23_inst : DFF_X1 port map( D => n9233, CK => CLK, Q => 
                           n14469, QN => n7093);
   REGISTERS_reg_23_22_inst : DFF_X1 port map( D => n9232, CK => CLK, Q => 
                           n14470, QN => n7092);
   REGISTERS_reg_23_21_inst : DFF_X1 port map( D => n9231, CK => CLK, Q => 
                           n14471, QN => n7091);
   REGISTERS_reg_23_20_inst : DFF_X1 port map( D => n9230, CK => CLK, Q => 
                           n14472, QN => n7090);
   REGISTERS_reg_23_19_inst : DFF_X1 port map( D => n9229, CK => CLK, Q => 
                           n14473, QN => n7089);
   REGISTERS_reg_23_18_inst : DFF_X1 port map( D => n9228, CK => CLK, Q => 
                           n14474, QN => n7088);
   REGISTERS_reg_23_17_inst : DFF_X1 port map( D => n9227, CK => CLK, Q => 
                           n14475, QN => n7087);
   REGISTERS_reg_23_16_inst : DFF_X1 port map( D => n9226, CK => CLK, Q => 
                           n14476, QN => n7086);
   REGISTERS_reg_23_15_inst : DFF_X1 port map( D => n9225, CK => CLK, Q => 
                           n14477, QN => n7085);
   REGISTERS_reg_23_14_inst : DFF_X1 port map( D => n9224, CK => CLK, Q => 
                           n14478, QN => n7084);
   REGISTERS_reg_23_13_inst : DFF_X1 port map( D => n9223, CK => CLK, Q => 
                           n14479, QN => n7083);
   REGISTERS_reg_23_12_inst : DFF_X1 port map( D => n9222, CK => CLK, Q => 
                           n14480, QN => n7082);
   REGISTERS_reg_23_11_inst : DFF_X1 port map( D => n9221, CK => CLK, Q => 
                           n14481, QN => n7081);
   REGISTERS_reg_23_10_inst : DFF_X1 port map( D => n9220, CK => CLK, Q => 
                           n14482, QN => n7080);
   REGISTERS_reg_23_9_inst : DFF_X1 port map( D => n9219, CK => CLK, Q => 
                           n14483, QN => n7079);
   REGISTERS_reg_23_8_inst : DFF_X1 port map( D => n9218, CK => CLK, Q => 
                           n14484, QN => n7078);
   REGISTERS_reg_23_7_inst : DFF_X1 port map( D => n9217, CK => CLK, Q => 
                           n14485, QN => n7077);
   REGISTERS_reg_23_6_inst : DFF_X1 port map( D => n9216, CK => CLK, Q => 
                           n14486, QN => n7076);
   REGISTERS_reg_23_5_inst : DFF_X1 port map( D => n9215, CK => CLK, Q => 
                           n14487, QN => n7075);
   REGISTERS_reg_23_4_inst : DFF_X1 port map( D => n9214, CK => CLK, Q => 
                           n14488, QN => n7074);
   REGISTERS_reg_23_3_inst : DFF_X1 port map( D => n9213, CK => CLK, Q => 
                           n14489, QN => n7073);
   REGISTERS_reg_23_2_inst : DFF_X1 port map( D => n9212, CK => CLK, Q => 
                           n14490, QN => n7072);
   REGISTERS_reg_23_1_inst : DFF_X1 port map( D => n9211, CK => CLK, Q => 
                           n14491, QN => n7071);
   REGISTERS_reg_23_0_inst : DFF_X1 port map( D => n9210, CK => CLK, Q => 
                           n14492, QN => n7070);
   REGISTERS_reg_22_23_inst : DFF_X1 port map( D => n9265, CK => CLK, Q => 
                           n15814, QN => n881);
   REGISTERS_reg_22_22_inst : DFF_X1 port map( D => n9264, CK => CLK, Q => 
                           n15815, QN => n882);
   REGISTERS_reg_22_21_inst : DFF_X1 port map( D => n9263, CK => CLK, Q => 
                           n15816, QN => n883);
   REGISTERS_reg_22_20_inst : DFF_X1 port map( D => n9262, CK => CLK, Q => 
                           n15817, QN => n884);
   REGISTERS_reg_22_19_inst : DFF_X1 port map( D => n9261, CK => CLK, Q => 
                           n15818, QN => n885);
   REGISTERS_reg_22_18_inst : DFF_X1 port map( D => n9260, CK => CLK, Q => 
                           n15819, QN => n886);
   REGISTERS_reg_22_17_inst : DFF_X1 port map( D => n9259, CK => CLK, Q => 
                           n15820, QN => n887);
   REGISTERS_reg_22_16_inst : DFF_X1 port map( D => n9258, CK => CLK, Q => 
                           n15821, QN => n888);
   REGISTERS_reg_22_15_inst : DFF_X1 port map( D => n9257, CK => CLK, Q => 
                           n15822, QN => n889);
   REGISTERS_reg_22_14_inst : DFF_X1 port map( D => n9256, CK => CLK, Q => 
                           n15823, QN => n890);
   REGISTERS_reg_22_13_inst : DFF_X1 port map( D => n9255, CK => CLK, Q => 
                           n15824, QN => n891);
   REGISTERS_reg_22_12_inst : DFF_X1 port map( D => n9254, CK => CLK, Q => 
                           n15825, QN => n892);
   REGISTERS_reg_22_11_inst : DFF_X1 port map( D => n9253, CK => CLK, Q => 
                           n15826, QN => n893);
   REGISTERS_reg_22_10_inst : DFF_X1 port map( D => n9252, CK => CLK, Q => 
                           n15827, QN => n894);
   REGISTERS_reg_22_9_inst : DFF_X1 port map( D => n9251, CK => CLK, Q => 
                           n15828, QN => n895);
   REGISTERS_reg_22_8_inst : DFF_X1 port map( D => n9250, CK => CLK, Q => 
                           n15829, QN => n896);
   REGISTERS_reg_22_7_inst : DFF_X1 port map( D => n9249, CK => CLK, Q => 
                           n15830, QN => n897);
   REGISTERS_reg_22_6_inst : DFF_X1 port map( D => n9248, CK => CLK, Q => 
                           n15831, QN => n898);
   REGISTERS_reg_22_5_inst : DFF_X1 port map( D => n9247, CK => CLK, Q => 
                           n15832, QN => n899);
   REGISTERS_reg_22_4_inst : DFF_X1 port map( D => n9246, CK => CLK, Q => 
                           n15833, QN => n900);
   REGISTERS_reg_22_3_inst : DFF_X1 port map( D => n9245, CK => CLK, Q => 
                           n15834, QN => n901);
   REGISTERS_reg_22_2_inst : DFF_X1 port map( D => n9244, CK => CLK, Q => 
                           n15835, QN => n902);
   REGISTERS_reg_22_1_inst : DFF_X1 port map( D => n9243, CK => CLK, Q => 
                           n15836, QN => n903);
   REGISTERS_reg_22_0_inst : DFF_X1 port map( D => n9242, CK => CLK, Q => 
                           n15837, QN => n904);
   REGISTERS_reg_21_23_inst : DFF_X1 port map( D => n9297, CK => CLK, Q => 
                           n15838, QN => n5793);
   REGISTERS_reg_21_22_inst : DFF_X1 port map( D => n9296, CK => CLK, Q => 
                           n15839, QN => n5789);
   REGISTERS_reg_21_21_inst : DFF_X1 port map( D => n9295, CK => CLK, Q => 
                           n15840, QN => n5785);
   REGISTERS_reg_21_20_inst : DFF_X1 port map( D => n9294, CK => CLK, Q => 
                           n15841, QN => n5781);
   REGISTERS_reg_21_19_inst : DFF_X1 port map( D => n9293, CK => CLK, Q => 
                           n15842, QN => n5777);
   REGISTERS_reg_21_18_inst : DFF_X1 port map( D => n9292, CK => CLK, Q => 
                           n15843, QN => n5773);
   REGISTERS_reg_21_17_inst : DFF_X1 port map( D => n9291, CK => CLK, Q => 
                           n15844, QN => n5769);
   REGISTERS_reg_21_16_inst : DFF_X1 port map( D => n9290, CK => CLK, Q => 
                           n15845, QN => n5765);
   REGISTERS_reg_21_15_inst : DFF_X1 port map( D => n9289, CK => CLK, Q => 
                           n15846, QN => n5761);
   REGISTERS_reg_21_14_inst : DFF_X1 port map( D => n9288, CK => CLK, Q => 
                           n15847, QN => n5757);
   REGISTERS_reg_21_13_inst : DFF_X1 port map( D => n9287, CK => CLK, Q => 
                           n15848, QN => n5753);
   REGISTERS_reg_21_12_inst : DFF_X1 port map( D => n9286, CK => CLK, Q => 
                           n15849, QN => n5749);
   REGISTERS_reg_21_11_inst : DFF_X1 port map( D => n9285, CK => CLK, Q => 
                           n15850, QN => n5745);
   REGISTERS_reg_21_10_inst : DFF_X1 port map( D => n9284, CK => CLK, Q => 
                           n15851, QN => n5741);
   REGISTERS_reg_21_9_inst : DFF_X1 port map( D => n9283, CK => CLK, Q => 
                           n15852, QN => n5737);
   REGISTERS_reg_21_8_inst : DFF_X1 port map( D => n9282, CK => CLK, Q => 
                           n15853, QN => n5733);
   REGISTERS_reg_21_7_inst : DFF_X1 port map( D => n9281, CK => CLK, Q => 
                           n15854, QN => n5729);
   REGISTERS_reg_21_6_inst : DFF_X1 port map( D => n9280, CK => CLK, Q => 
                           n15855, QN => n5725);
   REGISTERS_reg_21_5_inst : DFF_X1 port map( D => n9279, CK => CLK, Q => 
                           n15856, QN => n5721);
   REGISTERS_reg_21_4_inst : DFF_X1 port map( D => n9278, CK => CLK, Q => 
                           n15857, QN => n5717);
   REGISTERS_reg_21_3_inst : DFF_X1 port map( D => n9277, CK => CLK, Q => 
                           n15858, QN => n5713);
   REGISTERS_reg_21_2_inst : DFF_X1 port map( D => n9276, CK => CLK, Q => 
                           n15859, QN => n5709);
   REGISTERS_reg_21_1_inst : DFF_X1 port map( D => n9275, CK => CLK, Q => 
                           n15860, QN => n5705);
   REGISTERS_reg_21_0_inst : DFF_X1 port map( D => n9274, CK => CLK, Q => 
                           n15861, QN => n5701);
   REGISTERS_reg_20_23_inst : DFF_X1 port map( D => n9329, CK => CLK, Q => 
                           n15870, QN => n5792);
   REGISTERS_reg_20_22_inst : DFF_X1 port map( D => n9328, CK => CLK, Q => 
                           n15871, QN => n5788);
   REGISTERS_reg_20_21_inst : DFF_X1 port map( D => n9327, CK => CLK, Q => 
                           n15872, QN => n5784);
   REGISTERS_reg_20_20_inst : DFF_X1 port map( D => n9326, CK => CLK, Q => 
                           n15873, QN => n5780);
   REGISTERS_reg_20_19_inst : DFF_X1 port map( D => n9325, CK => CLK, Q => 
                           n15922, QN => n5776);
   REGISTERS_reg_20_18_inst : DFF_X1 port map( D => n9324, CK => CLK, Q => 
                           n14440, QN => n7104);
   REGISTERS_reg_20_17_inst : DFF_X1 port map( D => n9323, CK => CLK, Q => 
                           n14441, QN => n7103);
   REGISTERS_reg_20_16_inst : DFF_X1 port map( D => n9322, CK => CLK, Q => 
                           n14442, QN => n7102);
   REGISTERS_reg_20_15_inst : DFF_X1 port map( D => n9321, CK => CLK, Q => 
                           n14443, QN => n7101);
   REGISTERS_reg_20_14_inst : DFF_X1 port map( D => n9320, CK => CLK, Q => 
                           n14444, QN => n7100);
   REGISTERS_reg_20_13_inst : DFF_X1 port map( D => n9319, CK => CLK, Q => 
                           n14445, QN => n7099);
   REGISTERS_reg_20_12_inst : DFF_X1 port map( D => n9318, CK => CLK, Q => 
                           n14446, QN => n7098);
   REGISTERS_reg_20_11_inst : DFF_X1 port map( D => n9317, CK => CLK, Q => 
                           n14447, QN => n7097);
   REGISTERS_reg_20_10_inst : DFF_X1 port map( D => n9316, CK => CLK, Q => 
                           n14448, QN => n7096);
   REGISTERS_reg_20_9_inst : DFF_X1 port map( D => n9315, CK => CLK, Q => 
                           n14449, QN => n7095);
   REGISTERS_reg_20_8_inst : DFF_X1 port map( D => n9314, CK => CLK, Q => 
                           n14450, QN => n7094);
   REGISTERS_reg_20_7_inst : DFF_X1 port map( D => n9313, CK => CLK, Q => 
                           n14451, QN => n7005);
   REGISTERS_reg_20_6_inst : DFF_X1 port map( D => n9312, CK => CLK, Q => 
                           n14452, QN => n7004);
   REGISTERS_reg_20_5_inst : DFF_X1 port map( D => n9311, CK => CLK, Q => 
                           n14453, QN => n7003);
   REGISTERS_reg_20_4_inst : DFF_X1 port map( D => n9310, CK => CLK, Q => 
                           n14454, QN => n7002);
   REGISTERS_reg_20_3_inst : DFF_X1 port map( D => n9309, CK => CLK, Q => 
                           n14455, QN => n7001);
   REGISTERS_reg_20_2_inst : DFF_X1 port map( D => n9308, CK => CLK, Q => 
                           n14456, QN => n7000);
   REGISTERS_reg_20_1_inst : DFF_X1 port map( D => n9307, CK => CLK, Q => 
                           n14457, QN => n6999);
   REGISTERS_reg_20_0_inst : DFF_X1 port map( D => n9306, CK => CLK, Q => 
                           n14458, QN => n6998);
   REGISTERS_reg_14_23_inst : DFF_X1 port map( D => n9521, CK => CLK, Q => 
                           n14256, QN => n7128);
   REGISTERS_reg_14_22_inst : DFF_X1 port map( D => n9520, CK => CLK, Q => 
                           n14257, QN => n7127);
   REGISTERS_reg_14_21_inst : DFF_X1 port map( D => n9519, CK => CLK, Q => 
                           n14258, QN => n7126);
   REGISTERS_reg_14_20_inst : DFF_X1 port map( D => n9518, CK => CLK, Q => 
                           n14259, QN => n7125);
   REGISTERS_reg_14_19_inst : DFF_X1 port map( D => n9517, CK => CLK, Q => 
                           n14260, QN => n7124);
   REGISTERS_reg_14_18_inst : DFF_X1 port map( D => n9516, CK => CLK, Q => 
                           n14261, QN => n7123);
   REGISTERS_reg_14_17_inst : DFF_X1 port map( D => n9515, CK => CLK, Q => 
                           n14262, QN => n7122);
   REGISTERS_reg_14_16_inst : DFF_X1 port map( D => n9514, CK => CLK, Q => 
                           n14263, QN => n7121);
   REGISTERS_reg_14_15_inst : DFF_X1 port map( D => n9513, CK => CLK, Q => 
                           n14264, QN => n7120);
   REGISTERS_reg_14_14_inst : DFF_X1 port map( D => n9512, CK => CLK, Q => 
                           n14265, QN => n7119);
   REGISTERS_reg_14_13_inst : DFF_X1 port map( D => n9511, CK => CLK, Q => 
                           n14266, QN => n7118);
   REGISTERS_reg_14_12_inst : DFF_X1 port map( D => n9510, CK => CLK, Q => 
                           n14267, QN => n7117);
   REGISTERS_reg_14_11_inst : DFF_X1 port map( D => n9509, CK => CLK, Q => 
                           n14268, QN => n7116);
   REGISTERS_reg_14_10_inst : DFF_X1 port map( D => n9508, CK => CLK, Q => 
                           n14269, QN => n7115);
   REGISTERS_reg_14_9_inst : DFF_X1 port map( D => n9507, CK => CLK, Q => 
                           n14270, QN => n7114);
   REGISTERS_reg_14_8_inst : DFF_X1 port map( D => n9506, CK => CLK, Q => 
                           n14271, QN => n7113);
   REGISTERS_reg_14_7_inst : DFF_X1 port map( D => n9505, CK => CLK, Q => 
                           n14272, QN => n7112);
   REGISTERS_reg_14_6_inst : DFF_X1 port map( D => n9504, CK => CLK, Q => 
                           n14273, QN => n7111);
   REGISTERS_reg_14_5_inst : DFF_X1 port map( D => n9503, CK => CLK, Q => 
                           n14274, QN => n7110);
   REGISTERS_reg_14_4_inst : DFF_X1 port map( D => n9502, CK => CLK, Q => 
                           n14275, QN => n7109);
   REGISTERS_reg_14_3_inst : DFF_X1 port map( D => n9501, CK => CLK, Q => 
                           n14276, QN => n7108);
   REGISTERS_reg_14_2_inst : DFF_X1 port map( D => n9500, CK => CLK, Q => 
                           n14277, QN => n7107);
   REGISTERS_reg_14_1_inst : DFF_X1 port map( D => n9499, CK => CLK, Q => 
                           n14278, QN => n7106);
   REGISTERS_reg_14_0_inst : DFF_X1 port map( D => n9498, CK => CLK, Q => 
                           n14279, QN => n7105);
   REGISTERS_reg_13_23_inst : DFF_X1 port map( D => n9553, CK => CLK, Q => 
                           n15874, QN => n849);
   REGISTERS_reg_13_22_inst : DFF_X1 port map( D => n9552, CK => CLK, Q => 
                           n15875, QN => n850);
   REGISTERS_reg_13_21_inst : DFF_X1 port map( D => n9551, CK => CLK, Q => 
                           n15876, QN => n851);
   REGISTERS_reg_13_20_inst : DFF_X1 port map( D => n9550, CK => CLK, Q => 
                           n15877, QN => n852);
   REGISTERS_reg_13_19_inst : DFF_X1 port map( D => n9549, CK => CLK, Q => 
                           n15878, QN => n853);
   REGISTERS_reg_13_18_inst : DFF_X1 port map( D => n9548, CK => CLK, Q => 
                           n15879, QN => n854);
   REGISTERS_reg_13_17_inst : DFF_X1 port map( D => n9547, CK => CLK, Q => 
                           n15880, QN => n855);
   REGISTERS_reg_13_16_inst : DFF_X1 port map( D => n9546, CK => CLK, Q => 
                           n15881, QN => n856);
   REGISTERS_reg_13_15_inst : DFF_X1 port map( D => n9545, CK => CLK, Q => 
                           n15882, QN => n857);
   REGISTERS_reg_13_14_inst : DFF_X1 port map( D => n9544, CK => CLK, Q => 
                           n15883, QN => n858);
   REGISTERS_reg_13_13_inst : DFF_X1 port map( D => n9543, CK => CLK, Q => 
                           n15884, QN => n859);
   REGISTERS_reg_13_12_inst : DFF_X1 port map( D => n9542, CK => CLK, Q => 
                           n15885, QN => n860);
   REGISTERS_reg_13_11_inst : DFF_X1 port map( D => n9541, CK => CLK, Q => 
                           n15886, QN => n861);
   REGISTERS_reg_13_10_inst : DFF_X1 port map( D => n9540, CK => CLK, Q => 
                           n15887, QN => n862);
   REGISTERS_reg_13_9_inst : DFF_X1 port map( D => n9539, CK => CLK, Q => 
                           n15888, QN => n863);
   REGISTERS_reg_13_8_inst : DFF_X1 port map( D => n9538, CK => CLK, Q => 
                           n15889, QN => n864);
   REGISTERS_reg_13_7_inst : DFF_X1 port map( D => n9537, CK => CLK, Q => 
                           n15890, QN => n865);
   REGISTERS_reg_13_6_inst : DFF_X1 port map( D => n9536, CK => CLK, Q => 
                           n15891, QN => n866);
   REGISTERS_reg_13_5_inst : DFF_X1 port map( D => n9535, CK => CLK, Q => 
                           n15892, QN => n867);
   REGISTERS_reg_13_4_inst : DFF_X1 port map( D => n9534, CK => CLK, Q => 
                           n15893, QN => n868);
   REGISTERS_reg_13_3_inst : DFF_X1 port map( D => n9533, CK => CLK, Q => 
                           n15894, QN => n869);
   REGISTERS_reg_13_2_inst : DFF_X1 port map( D => n9532, CK => CLK, Q => 
                           n15895, QN => n870);
   REGISTERS_reg_13_1_inst : DFF_X1 port map( D => n9531, CK => CLK, Q => 
                           n15896, QN => n871);
   REGISTERS_reg_13_0_inst : DFF_X1 port map( D => n9530, CK => CLK, Q => 
                           n15897, QN => n872);
   REGISTERS_reg_5_23_inst : DFF_X1 port map( D => n9809, CK => CLK, Q => 
                           n14084, QN => n7152);
   REGISTERS_reg_5_22_inst : DFF_X1 port map( D => n9808, CK => CLK, Q => 
                           n14085, QN => n7151);
   REGISTERS_reg_5_21_inst : DFF_X1 port map( D => n9807, CK => CLK, Q => 
                           n14086, QN => n7150);
   REGISTERS_reg_5_20_inst : DFF_X1 port map( D => n9806, CK => CLK, Q => 
                           n14087, QN => n7149);
   REGISTERS_reg_5_19_inst : DFF_X1 port map( D => n9805, CK => CLK, Q => 
                           n14088, QN => n7148);
   REGISTERS_reg_5_18_inst : DFF_X1 port map( D => n9804, CK => CLK, Q => 
                           n14089, QN => n7147);
   REGISTERS_reg_5_17_inst : DFF_X1 port map( D => n9803, CK => CLK, Q => 
                           n14090, QN => n7146);
   REGISTERS_reg_5_16_inst : DFF_X1 port map( D => n9802, CK => CLK, Q => 
                           n14091, QN => n7145);
   REGISTERS_reg_5_15_inst : DFF_X1 port map( D => n9801, CK => CLK, Q => 
                           n14092, QN => n7144);
   REGISTERS_reg_5_14_inst : DFF_X1 port map( D => n9800, CK => CLK, Q => 
                           n14093, QN => n7143);
   REGISTERS_reg_5_13_inst : DFF_X1 port map( D => n9799, CK => CLK, Q => 
                           n14094, QN => n7142);
   REGISTERS_reg_5_12_inst : DFF_X1 port map( D => n9798, CK => CLK, Q => 
                           n14095, QN => n7141);
   REGISTERS_reg_5_11_inst : DFF_X1 port map( D => n9797, CK => CLK, Q => 
                           n14096, QN => n7140);
   REGISTERS_reg_5_10_inst : DFF_X1 port map( D => n9796, CK => CLK, Q => 
                           n14097, QN => n7139);
   REGISTERS_reg_5_9_inst : DFF_X1 port map( D => n9795, CK => CLK, Q => n14098
                           , QN => n7138);
   REGISTERS_reg_5_8_inst : DFF_X1 port map( D => n9794, CK => CLK, Q => n14099
                           , QN => n7137);
   REGISTERS_reg_5_7_inst : DFF_X1 port map( D => n9793, CK => CLK, Q => n14100
                           , QN => n7136);
   REGISTERS_reg_5_6_inst : DFF_X1 port map( D => n9792, CK => CLK, Q => n14101
                           , QN => n7135);
   REGISTERS_reg_5_5_inst : DFF_X1 port map( D => n9791, CK => CLK, Q => n14102
                           , QN => n7134);
   REGISTERS_reg_5_4_inst : DFF_X1 port map( D => n9790, CK => CLK, Q => n14103
                           , QN => n7133);
   REGISTERS_reg_5_3_inst : DFF_X1 port map( D => n9789, CK => CLK, Q => n14104
                           , QN => n7132);
   REGISTERS_reg_5_2_inst : DFF_X1 port map( D => n9788, CK => CLK, Q => n14105
                           , QN => n7131);
   REGISTERS_reg_5_1_inst : DFF_X1 port map( D => n9787, CK => CLK, Q => n14106
                           , QN => n7130);
   REGISTERS_reg_5_0_inst : DFF_X1 port map( D => n9786, CK => CLK, Q => n14107
                           , QN => n7129);
   REGISTERS_reg_4_23_inst : DFF_X1 port map( D => n9841, CK => CLK, Q => 
                           n15898, QN => n817);
   REGISTERS_reg_4_22_inst : DFF_X1 port map( D => n9840, CK => CLK, Q => 
                           n15899, QN => n818);
   REGISTERS_reg_4_21_inst : DFF_X1 port map( D => n9839, CK => CLK, Q => 
                           n15900, QN => n819);
   REGISTERS_reg_4_20_inst : DFF_X1 port map( D => n9838, CK => CLK, Q => 
                           n15901, QN => n820);
   REGISTERS_reg_4_19_inst : DFF_X1 port map( D => n9837, CK => CLK, Q => 
                           n15902, QN => n821);
   REGISTERS_reg_4_18_inst : DFF_X1 port map( D => n9836, CK => CLK, Q => 
                           n15903, QN => n822);
   REGISTERS_reg_4_17_inst : DFF_X1 port map( D => n9835, CK => CLK, Q => 
                           n15904, QN => n823);
   REGISTERS_reg_4_16_inst : DFF_X1 port map( D => n9834, CK => CLK, Q => 
                           n15905, QN => n824);
   REGISTERS_reg_4_15_inst : DFF_X1 port map( D => n9833, CK => CLK, Q => 
                           n15906, QN => n825);
   REGISTERS_reg_4_14_inst : DFF_X1 port map( D => n9832, CK => CLK, Q => 
                           n15907, QN => n826);
   REGISTERS_reg_4_13_inst : DFF_X1 port map( D => n9831, CK => CLK, Q => 
                           n15908, QN => n827);
   REGISTERS_reg_4_12_inst : DFF_X1 port map( D => n9830, CK => CLK, Q => 
                           n15909, QN => n828);
   REGISTERS_reg_4_11_inst : DFF_X1 port map( D => n9829, CK => CLK, Q => 
                           n15910, QN => n829);
   REGISTERS_reg_4_10_inst : DFF_X1 port map( D => n9828, CK => CLK, Q => 
                           n15911, QN => n830);
   REGISTERS_reg_4_9_inst : DFF_X1 port map( D => n9827, CK => CLK, Q => n15912
                           , QN => n831);
   REGISTERS_reg_4_8_inst : DFF_X1 port map( D => n9826, CK => CLK, Q => n15913
                           , QN => n832);
   REGISTERS_reg_4_7_inst : DFF_X1 port map( D => n9825, CK => CLK, Q => n15914
                           , QN => n833);
   REGISTERS_reg_4_6_inst : DFF_X1 port map( D => n9824, CK => CLK, Q => n15915
                           , QN => n834);
   REGISTERS_reg_4_5_inst : DFF_X1 port map( D => n9823, CK => CLK, Q => n15916
                           , QN => n835);
   REGISTERS_reg_4_4_inst : DFF_X1 port map( D => n9822, CK => CLK, Q => n15917
                           , QN => n836);
   REGISTERS_reg_4_3_inst : DFF_X1 port map( D => n9821, CK => CLK, Q => n15918
                           , QN => n837);
   REGISTERS_reg_4_2_inst : DFF_X1 port map( D => n9820, CK => CLK, Q => n15919
                           , QN => n838);
   REGISTERS_reg_4_1_inst : DFF_X1 port map( D => n9819, CK => CLK, Q => n15920
                           , QN => n839);
   REGISTERS_reg_4_0_inst : DFF_X1 port map( D => n9818, CK => CLK, Q => n15921
                           , QN => n840);
   REGISTERS_reg_12_31_inst : DFF_X1 port map( D => n9593, CK => CLK, Q => 
                           n15931, QN => n5695);
   REGISTERS_reg_12_30_inst : DFF_X1 port map( D => n9592, CK => CLK, Q => 
                           n15932, QN => n5685);
   REGISTERS_reg_12_29_inst : DFF_X1 port map( D => n9591, CK => CLK, Q => 
                           n15933, QN => n5675);
   REGISTERS_reg_12_28_inst : DFF_X1 port map( D => n9590, CK => CLK, Q => 
                           n15934, QN => n5665);
   REGISTERS_reg_12_27_inst : DFF_X1 port map( D => n9589, CK => CLK, Q => 
                           n15935, QN => n5655);
   REGISTERS_reg_12_26_inst : DFF_X1 port map( D => n9588, CK => CLK, Q => 
                           n15936, QN => n5645);
   REGISTERS_reg_12_25_inst : DFF_X1 port map( D => n9587, CK => CLK, Q => 
                           n15937, QN => n5635);
   REGISTERS_reg_12_24_inst : DFF_X1 port map( D => n9586, CK => CLK, Q => 
                           n15938, QN => n5625);
   REGISTERS_reg_9_31_inst : DFF_X1 port map( D => n9689, CK => CLK, Q => 
                           n14204, QN => n6921);
   REGISTERS_reg_9_30_inst : DFF_X1 port map( D => n9688, CK => CLK, Q => 
                           n14205, QN => n6920);
   REGISTERS_reg_9_29_inst : DFF_X1 port map( D => n9687, CK => CLK, Q => 
                           n14206, QN => n6919);
   REGISTERS_reg_9_28_inst : DFF_X1 port map( D => n9686, CK => CLK, Q => 
                           n14207, QN => n6918);
   REGISTERS_reg_9_27_inst : DFF_X1 port map( D => n9685, CK => CLK, Q => 
                           n14208, QN => n6917);
   REGISTERS_reg_9_26_inst : DFF_X1 port map( D => n9684, CK => CLK, Q => 
                           n14209, QN => n6916);
   REGISTERS_reg_9_25_inst : DFF_X1 port map( D => n9683, CK => CLK, Q => 
                           n14210, QN => n6915);
   REGISTERS_reg_9_24_inst : DFF_X1 port map( D => n9682, CK => CLK, Q => 
                           n14211, QN => n6914);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n9881, CK => CLK, Q => 
                           n15939, QN => n5697);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n9880, CK => CLK, Q => 
                           n15940, QN => n5687);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n9879, CK => CLK, Q => 
                           n15941, QN => n5677);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n9878, CK => CLK, Q => 
                           n15942, QN => n5667);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n9877, CK => CLK, Q => 
                           n15943, QN => n5657);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n9876, CK => CLK, Q => 
                           n15944, QN => n5647);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n9875, CK => CLK, Q => 
                           n15945, QN => n5637);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n9874, CK => CLK, Q => 
                           n15946, QN => n5627);
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n9977, CK => CLK, Q => 
                           n14028, QN => n6937);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n9976, CK => CLK, Q => 
                           n14029, QN => n6936);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n9975, CK => CLK, Q => 
                           n14030, QN => n6935);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n9974, CK => CLK, Q => 
                           n14031, QN => n6934);
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n9973, CK => CLK, Q => 
                           n14032, QN => n6933);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n9972, CK => CLK, Q => 
                           n14033, QN => n6932);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n9971, CK => CLK, Q => 
                           n14034, QN => n6931);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n9970, CK => CLK, Q => 
                           n14035, QN => n6930);
   REGISTERS_reg_10_31_inst : DFF_X1 port map( D => n9657, CK => CLK, Q => 
                           n14216, QN => n6793);
   REGISTERS_reg_10_30_inst : DFF_X1 port map( D => n9656, CK => CLK, Q => 
                           n14217, QN => n6792);
   REGISTERS_reg_10_29_inst : DFF_X1 port map( D => n9655, CK => CLK, Q => 
                           n14218, QN => n6791);
   REGISTERS_reg_10_28_inst : DFF_X1 port map( D => n9654, CK => CLK, Q => 
                           n14219, QN => n6790);
   REGISTERS_reg_10_27_inst : DFF_X1 port map( D => n9653, CK => CLK, Q => 
                           n14220, QN => n6789);
   REGISTERS_reg_10_26_inst : DFF_X1 port map( D => n9652, CK => CLK, Q => 
                           n14221, QN => n6788);
   REGISTERS_reg_10_25_inst : DFF_X1 port map( D => n9651, CK => CLK, Q => 
                           n14222, QN => n6787);
   REGISTERS_reg_10_24_inst : DFF_X1 port map( D => n9650, CK => CLK, Q => 
                           n14223, QN => n6786);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n9945, CK => CLK, Q => 
                           n14044, QN => n6809);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n9944, CK => CLK, Q => 
                           n14045, QN => n6808);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n9943, CK => CLK, Q => 
                           n14046, QN => n6807);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n9942, CK => CLK, Q => 
                           n14047, QN => n6806);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n9941, CK => CLK, Q => 
                           n14048, QN => n6805);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n9940, CK => CLK, Q => 
                           n14049, QN => n6804);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n9939, CK => CLK, Q => 
                           n14050, QN => n6803);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n9938, CK => CLK, Q => 
                           n14051, QN => n6802);
   REGISTERS_reg_12_23_inst : DFF_X1 port map( D => n9585, CK => CLK, Q => 
                           n15971, QN => n5615);
   REGISTERS_reg_12_22_inst : DFF_X1 port map( D => n9584, CK => CLK, Q => 
                           n15972, QN => n5605);
   REGISTERS_reg_12_21_inst : DFF_X1 port map( D => n9583, CK => CLK, Q => 
                           n15973, QN => n5595);
   REGISTERS_reg_12_20_inst : DFF_X1 port map( D => n9582, CK => CLK, Q => 
                           n15974, QN => n5585);
   REGISTERS_reg_12_19_inst : DFF_X1 port map( D => n9581, CK => CLK, Q => 
                           n15975, QN => n5575);
   REGISTERS_reg_12_18_inst : DFF_X1 port map( D => n9580, CK => CLK, Q => 
                           n15976, QN => n5565);
   REGISTERS_reg_12_17_inst : DFF_X1 port map( D => n9579, CK => CLK, Q => 
                           n15977, QN => n5555);
   REGISTERS_reg_12_16_inst : DFF_X1 port map( D => n9578, CK => CLK, Q => 
                           n15978, QN => n5545);
   REGISTERS_reg_12_15_inst : DFF_X1 port map( D => n9577, CK => CLK, Q => 
                           n15979, QN => n5535);
   REGISTERS_reg_12_14_inst : DFF_X1 port map( D => n9576, CK => CLK, Q => 
                           n15980, QN => n5525);
   REGISTERS_reg_12_13_inst : DFF_X1 port map( D => n9575, CK => CLK, Q => 
                           n15981, QN => n5515);
   REGISTERS_reg_12_12_inst : DFF_X1 port map( D => n9574, CK => CLK, Q => 
                           n15982, QN => n5505);
   REGISTERS_reg_12_11_inst : DFF_X1 port map( D => n9573, CK => CLK, Q => 
                           n15983, QN => n5495);
   REGISTERS_reg_12_10_inst : DFF_X1 port map( D => n9572, CK => CLK, Q => 
                           n15984, QN => n5485);
   REGISTERS_reg_12_9_inst : DFF_X1 port map( D => n9571, CK => CLK, Q => 
                           n15985, QN => n5475);
   REGISTERS_reg_12_8_inst : DFF_X1 port map( D => n9570, CK => CLK, Q => 
                           n15986, QN => n5465);
   REGISTERS_reg_12_7_inst : DFF_X1 port map( D => n9569, CK => CLK, Q => 
                           n15987, QN => n5455);
   REGISTERS_reg_12_6_inst : DFF_X1 port map( D => n9568, CK => CLK, Q => 
                           n15988, QN => n5445);
   REGISTERS_reg_12_5_inst : DFF_X1 port map( D => n9567, CK => CLK, Q => 
                           n15989, QN => n5435);
   REGISTERS_reg_12_4_inst : DFF_X1 port map( D => n9566, CK => CLK, Q => 
                           n15990, QN => n5425);
   REGISTERS_reg_12_3_inst : DFF_X1 port map( D => n9565, CK => CLK, Q => 
                           n15991, QN => n5415);
   REGISTERS_reg_12_2_inst : DFF_X1 port map( D => n9564, CK => CLK, Q => 
                           n15992, QN => n5405);
   REGISTERS_reg_12_1_inst : DFF_X1 port map( D => n9563, CK => CLK, Q => 
                           n15993, QN => n5395);
   REGISTERS_reg_12_0_inst : DFF_X1 port map( D => n9562, CK => CLK, Q => 
                           n15994, QN => n5385);
   REGISTERS_reg_9_23_inst : DFF_X1 port map( D => n9681, CK => CLK, Q => 
                           n14212, QN => n6941);
   REGISTERS_reg_9_22_inst : DFF_X1 port map( D => n9680, CK => CLK, Q => 
                           n14213, QN => n6940);
   REGISTERS_reg_9_21_inst : DFF_X1 port map( D => n9679, CK => CLK, Q => 
                           n14214, QN => n6939);
   REGISTERS_reg_9_20_inst : DFF_X1 port map( D => n9678, CK => CLK, Q => 
                           n14215, QN => n6938);
   REGISTERS_reg_9_19_inst : DFF_X1 port map( D => n9677, CK => CLK, Q => 
                           n16043, QN => n653);
   REGISTERS_reg_9_18_inst : DFF_X1 port map( D => n9676, CK => CLK, Q => 
                           n16044, QN => n656);
   REGISTERS_reg_9_17_inst : DFF_X1 port map( D => n9675, CK => CLK, Q => 
                           n16045, QN => n659);
   REGISTERS_reg_9_16_inst : DFF_X1 port map( D => n9674, CK => CLK, Q => 
                           n16046, QN => n662);
   REGISTERS_reg_9_15_inst : DFF_X1 port map( D => n9673, CK => CLK, Q => 
                           n16047, QN => n665);
   REGISTERS_reg_9_14_inst : DFF_X1 port map( D => n9672, CK => CLK, Q => 
                           n16048, QN => n668);
   REGISTERS_reg_9_13_inst : DFF_X1 port map( D => n9671, CK => CLK, Q => 
                           n16049, QN => n671);
   REGISTERS_reg_9_12_inst : DFF_X1 port map( D => n9670, CK => CLK, Q => 
                           n16050, QN => n674);
   REGISTERS_reg_9_11_inst : DFF_X1 port map( D => n9669, CK => CLK, Q => 
                           n15995, QN => n677);
   REGISTERS_reg_9_10_inst : DFF_X1 port map( D => n9668, CK => CLK, Q => 
                           n15996, QN => n680);
   REGISTERS_reg_9_9_inst : DFF_X1 port map( D => n9667, CK => CLK, Q => n15997
                           , QN => n683);
   REGISTERS_reg_9_8_inst : DFF_X1 port map( D => n9666, CK => CLK, Q => n15998
                           , QN => n686);
   REGISTERS_reg_9_7_inst : DFF_X1 port map( D => n9665, CK => CLK, Q => n15999
                           , QN => n689);
   REGISTERS_reg_9_6_inst : DFF_X1 port map( D => n9664, CK => CLK, Q => n16000
                           , QN => n692);
   REGISTERS_reg_9_5_inst : DFF_X1 port map( D => n9663, CK => CLK, Q => n16001
                           , QN => n695);
   REGISTERS_reg_9_4_inst : DFF_X1 port map( D => n9662, CK => CLK, Q => n16002
                           , QN => n698);
   REGISTERS_reg_9_3_inst : DFF_X1 port map( D => n9661, CK => CLK, Q => n16003
                           , QN => n701);
   REGISTERS_reg_9_2_inst : DFF_X1 port map( D => n9660, CK => CLK, Q => n16004
                           , QN => n704);
   REGISTERS_reg_9_1_inst : DFF_X1 port map( D => n9659, CK => CLK, Q => n16005
                           , QN => n707);
   REGISTERS_reg_9_0_inst : DFF_X1 port map( D => n9658, CK => CLK, Q => n16006
                           , QN => n710);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n9873, CK => CLK, Q => 
                           n16007, QN => n5617);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n9872, CK => CLK, Q => 
                           n16008, QN => n5607);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n9871, CK => CLK, Q => 
                           n16009, QN => n5597);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n9870, CK => CLK, Q => 
                           n16010, QN => n5587);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n9869, CK => CLK, Q => 
                           n16011, QN => n5577);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n9868, CK => CLK, Q => 
                           n16012, QN => n5567);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n9867, CK => CLK, Q => 
                           n16013, QN => n5557);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n9866, CK => CLK, Q => 
                           n16014, QN => n5547);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n9865, CK => CLK, Q => 
                           n16015, QN => n5537);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n9864, CK => CLK, Q => 
                           n16016, QN => n5527);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n9863, CK => CLK, Q => 
                           n16017, QN => n5517);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n9862, CK => CLK, Q => 
                           n16018, QN => n5507);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n9861, CK => CLK, Q => 
                           n16019, QN => n5497);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n9860, CK => CLK, Q => 
                           n16020, QN => n5487);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n9859, CK => CLK, Q => n16021
                           , QN => n5477);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n9858, CK => CLK, Q => n16022
                           , QN => n5467);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n9857, CK => CLK, Q => n16023
                           , QN => n5457);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n9856, CK => CLK, Q => n16024
                           , QN => n5447);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n9855, CK => CLK, Q => n16025
                           , QN => n5437);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n9854, CK => CLK, Q => n16026
                           , QN => n5427);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n9853, CK => CLK, Q => n16027
                           , QN => n5417);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n9852, CK => CLK, Q => n16028
                           , QN => n5407);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n9851, CK => CLK, Q => n16029
                           , QN => n5397);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n9850, CK => CLK, Q => n16030
                           , QN => n5387);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n9969, CK => CLK, Q => 
                           n14036, QN => n6929);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n9968, CK => CLK, Q => 
                           n14037, QN => n6928);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n9967, CK => CLK, Q => 
                           n14038, QN => n6927);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n9966, CK => CLK, Q => 
                           n14039, QN => n6926);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n9965, CK => CLK, Q => 
                           n14040, QN => n6925);
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n9964, CK => CLK, Q => 
                           n14041, QN => n6924);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n9963, CK => CLK, Q => 
                           n14042, QN => n6923);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n9962, CK => CLK, Q => 
                           n14043, QN => n6922);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n9961, CK => CLK, Q => 
                           n16051, QN => n666);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n9960, CK => CLK, Q => 
                           n16052, QN => n669);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n9959, CK => CLK, Q => 
                           n16053, QN => n672);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n9958, CK => CLK, Q => 
                           n16054, QN => n675);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n9957, CK => CLK, Q => 
                           n16031, QN => n678);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n9956, CK => CLK, Q => 
                           n16032, QN => n681);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n9955, CK => CLK, Q => n16033
                           , QN => n684);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n9954, CK => CLK, Q => n16034
                           , QN => n687);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n9953, CK => CLK, Q => n16035
                           , QN => n690);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n9952, CK => CLK, Q => n16036
                           , QN => n693);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n9951, CK => CLK, Q => n16037
                           , QN => n696);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n9950, CK => CLK, Q => n16038
                           , QN => n699);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n9949, CK => CLK, Q => n16039
                           , QN => n702);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n9948, CK => CLK, Q => n16040
                           , QN => n705);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n9947, CK => CLK, Q => n16041
                           , QN => n708);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n9946, CK => CLK, Q => n16042
                           , QN => n711);
   REGISTERS_reg_10_23_inst : DFF_X1 port map( D => n9649, CK => CLK, Q => 
                           n14224, QN => n6813);
   REGISTERS_reg_10_22_inst : DFF_X1 port map( D => n9648, CK => CLK, Q => 
                           n14225, QN => n6812);
   REGISTERS_reg_10_21_inst : DFF_X1 port map( D => n9647, CK => CLK, Q => 
                           n14226, QN => n6811);
   REGISTERS_reg_10_20_inst : DFF_X1 port map( D => n9646, CK => CLK, Q => 
                           n14227, QN => n6810);
   REGISTERS_reg_10_19_inst : DFF_X1 port map( D => n9645, CK => CLK, Q => 
                           n14228, QN => n6893);
   REGISTERS_reg_10_18_inst : DFF_X1 port map( D => n9644, CK => CLK, Q => 
                           n14229, QN => n6892);
   REGISTERS_reg_10_17_inst : DFF_X1 port map( D => n9643, CK => CLK, Q => 
                           n14230, QN => n6891);
   REGISTERS_reg_10_16_inst : DFF_X1 port map( D => n9642, CK => CLK, Q => 
                           n14231, QN => n6890);
   REGISTERS_reg_10_15_inst : DFF_X1 port map( D => n9641, CK => CLK, Q => 
                           n14232, QN => n6888);
   REGISTERS_reg_10_14_inst : DFF_X1 port map( D => n9640, CK => CLK, Q => 
                           n14233, QN => n6886);
   REGISTERS_reg_10_13_inst : DFF_X1 port map( D => n9639, CK => CLK, Q => 
                           n14234, QN => n6884);
   REGISTERS_reg_10_12_inst : DFF_X1 port map( D => n9638, CK => CLK, Q => 
                           n14235, QN => n6882);
   REGISTERS_reg_10_11_inst : DFF_X1 port map( D => n9637, CK => CLK, Q => 
                           n14236, QN => n6881);
   REGISTERS_reg_10_10_inst : DFF_X1 port map( D => n9636, CK => CLK, Q => 
                           n14237, QN => n6880);
   REGISTERS_reg_10_9_inst : DFF_X1 port map( D => n9635, CK => CLK, Q => 
                           n14238, QN => n6879);
   REGISTERS_reg_10_8_inst : DFF_X1 port map( D => n9634, CK => CLK, Q => 
                           n14239, QN => n6878);
   REGISTERS_reg_10_7_inst : DFF_X1 port map( D => n9633, CK => CLK, Q => 
                           n14240, QN => n6877);
   REGISTERS_reg_10_6_inst : DFF_X1 port map( D => n9632, CK => CLK, Q => 
                           n14241, QN => n6876);
   REGISTERS_reg_10_5_inst : DFF_X1 port map( D => n9631, CK => CLK, Q => 
                           n14242, QN => n6875);
   REGISTERS_reg_10_4_inst : DFF_X1 port map( D => n9630, CK => CLK, Q => 
                           n14243, QN => n6874);
   REGISTERS_reg_10_3_inst : DFF_X1 port map( D => n9629, CK => CLK, Q => 
                           n14244, QN => n6873);
   REGISTERS_reg_10_2_inst : DFF_X1 port map( D => n9628, CK => CLK, Q => 
                           n14245, QN => n6872);
   REGISTERS_reg_10_1_inst : DFF_X1 port map( D => n9627, CK => CLK, Q => 
                           n14246, QN => n6871);
   REGISTERS_reg_10_0_inst : DFF_X1 port map( D => n9626, CK => CLK, Q => 
                           n14247, QN => n6870);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n9937, CK => CLK, Q => 
                           n14052, QN => n6801);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n9936, CK => CLK, Q => 
                           n14053, QN => n6800);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n9935, CK => CLK, Q => 
                           n14054, QN => n6799);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n9934, CK => CLK, Q => 
                           n14055, QN => n6798);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n9933, CK => CLK, Q => 
                           n14056, QN => n6797);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n9932, CK => CLK, Q => 
                           n14057, QN => n6796);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n9931, CK => CLK, Q => 
                           n14058, QN => n6795);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n9930, CK => CLK, Q => 
                           n14059, QN => n6794);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n9929, CK => CLK, Q => 
                           n14060, QN => n6889);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n9928, CK => CLK, Q => 
                           n14061, QN => n6887);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n9927, CK => CLK, Q => 
                           n14062, QN => n6885);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n9926, CK => CLK, Q => 
                           n14063, QN => n6883);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n9925, CK => CLK, Q => 
                           n14064, QN => n6841);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n9924, CK => CLK, Q => 
                           n14065, QN => n6840);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n9923, CK => CLK, Q => n14066
                           , QN => n6839);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n9922, CK => CLK, Q => n14067
                           , QN => n6838);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n9921, CK => CLK, Q => n14068
                           , QN => n6837);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n9920, CK => CLK, Q => n14069
                           , QN => n6836);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n9919, CK => CLK, Q => n14070
                           , QN => n6835);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n9918, CK => CLK, Q => n14071
                           , QN => n6834);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n9917, CK => CLK, Q => n14072
                           , QN => n6833);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n9916, CK => CLK, Q => n14073
                           , QN => n6832);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n9915, CK => CLK, Q => n14074
                           , QN => n6831);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n9914, CK => CLK, Q => n14075
                           , QN => n6830);
   OUT2_reg_31_inst : DFF_X1 port map( D => n7609, CK => CLK, Q => n_2202, QN 
                           => n1481);
   OUT2_reg_30_inst : DFF_X1 port map( D => n7607, CK => CLK, Q => n_2203, QN 
                           => n1482);
   OUT2_reg_29_inst : DFF_X1 port map( D => n7605, CK => CLK, Q => n_2204, QN 
                           => n1483);
   OUT2_reg_28_inst : DFF_X1 port map( D => n7603, CK => CLK, Q => n_2205, QN 
                           => n1484);
   OUT2_reg_27_inst : DFF_X1 port map( D => n7601, CK => CLK, Q => n_2206, QN 
                           => n1485);
   OUT2_reg_26_inst : DFF_X1 port map( D => n7599, CK => CLK, Q => n_2207, QN 
                           => n1486);
   OUT2_reg_25_inst : DFF_X1 port map( D => n7597, CK => CLK, Q => n_2208, QN 
                           => n1487);
   OUT1_reg_31_inst : DFF_X1 port map( D => n7673, CK => CLK, Q => n_2209, QN 
                           => n1449);
   OUT1_reg_30_inst : DFF_X1 port map( D => n7671, CK => CLK, Q => n_2210, QN 
                           => n1450);
   OUT1_reg_29_inst : DFF_X1 port map( D => n7669, CK => CLK, Q => n_2211, QN 
                           => n1451);
   OUT1_reg_28_inst : DFF_X1 port map( D => n7667, CK => CLK, Q => n_2212, QN 
                           => n1452);
   OUT1_reg_27_inst : DFF_X1 port map( D => n7665, CK => CLK, Q => n_2213, QN 
                           => n1453);
   OUT1_reg_26_inst : DFF_X1 port map( D => n7663, CK => CLK, Q => n_2214, QN 
                           => n1454);
   OUT1_reg_25_inst : DFF_X1 port map( D => n7661, CK => CLK, Q => n_2215, QN 
                           => n1455);
   OUT2_reg_24_inst : DFF_X1 port map( D => n7595, CK => CLK, Q => n_2216, QN 
                           => n1488);
   OUT1_reg_24_inst : DFF_X1 port map( D => n7659, CK => CLK, Q => n_2217, QN 
                           => n1456);
   U3 : NOR3_X1 port map( A1 => n16058, A2 => ADD_RD2(3), A3 => n16057, ZN => 
                           n5710);
   U4 : NOR3_X1 port map( A1 => n16068, A2 => ADD_RD2(0), A3 => n16069, ZN => 
                           n5669);
   U69 : NOR3_X2 port map( A1 => n16064, A2 => ADD_RD1(2), A3 => n16065, ZN => 
                           n4279);
   U70 : NOR3_X1 port map( A1 => n16056, A2 => ADD_RD1(3), A3 => n16055, ZN => 
                           n4299);
   U71 : NOR3_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), A3 => n16064, ZN
                           => n4274);
   U72 : NOR3_X1 port map( A1 => n16065, A2 => ADD_RD1(0), A3 => n16066, ZN => 
                           n4276);
   U73 : NOR3_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), A3 => ADD_RD1(0)
                           , ZN => n4271);
   U74 : NOR3_X1 port map( A1 => n16067, A2 => ADD_RD2(1), A3 => n16069, ZN => 
                           n5668);
   U75 : NOR3_X1 port map( A1 => n16064, A2 => ADD_RD1(1), A3 => n16066, ZN => 
                           n4275);
   U76 : BUF_X1 port map( A => n2875, Z => n13797);
   U77 : BUF_X1 port map( A => n2902, Z => n13743);
   U78 : BUF_X1 port map( A => n2878, Z => n13791);
   U79 : BUF_X1 port map( A => n2905, Z => n13737);
   U80 : BUF_X1 port map( A => n2911, Z => n13725);
   U81 : BUF_X1 port map( A => n2908, Z => n13731);
   U82 : BUF_X1 port map( A => n2899, Z => n13749);
   U83 : BUF_X1 port map( A => n2896, Z => n13755);
   U84 : BUF_X1 port map( A => n2893, Z => n13761);
   U85 : BUF_X1 port map( A => n2890, Z => n13767);
   U86 : BUF_X1 port map( A => n2887, Z => n13773);
   U87 : BUF_X1 port map( A => n2884, Z => n13779);
   U88 : BUF_X1 port map( A => n2881, Z => n13785);
   U89 : BUF_X1 port map( A => n2872, Z => n13803);
   U90 : BUF_X1 port map( A => n2869, Z => n13809);
   U91 : BUF_X1 port map( A => n2980, Z => n13527);
   U92 : BUF_X1 port map( A => n2927, Z => n13683);
   U93 : BUF_X1 port map( A => n2943, Z => n13635);
   U94 : BUF_X1 port map( A => n2945, Z => n13629);
   U95 : BUF_X1 port map( A => n2964, Z => n13575);
   U96 : BUF_X1 port map( A => n3017, Z => n13437);
   U97 : BUF_X1 port map( A => n3015, Z => n13443);
   U98 : BUF_X1 port map( A => n3013, Z => n13449);
   U99 : BUF_X1 port map( A => n3010, Z => n13455);
   U100 : BUF_X1 port map( A => n3007, Z => n13461);
   U101 : BUF_X1 port map( A => n3004, Z => n13467);
   U102 : BUF_X1 port map( A => n3001, Z => n13473);
   U103 : BUF_X1 port map( A => n2997, Z => n13479);
   U104 : BUF_X1 port map( A => n2995, Z => n13485);
   U105 : BUF_X1 port map( A => n2993, Z => n13491);
   U106 : BUF_X1 port map( A => n2991, Z => n13497);
   U107 : BUF_X1 port map( A => n2989, Z => n13503);
   U108 : BUF_X1 port map( A => n2987, Z => n13509);
   U109 : BUF_X1 port map( A => n2985, Z => n13515);
   U110 : BUF_X1 port map( A => n2983, Z => n13521);
   U111 : BUF_X1 port map( A => n2978, Z => n13533);
   U112 : BUF_X1 port map( A => n2976, Z => n13539);
   U113 : BUF_X1 port map( A => n2974, Z => n13545);
   U114 : BUF_X1 port map( A => n2972, Z => n13551);
   U115 : BUF_X1 port map( A => n2970, Z => n13557);
   U116 : BUF_X1 port map( A => n2968, Z => n13563);
   U117 : BUF_X1 port map( A => n2966, Z => n13569);
   U118 : BUF_X1 port map( A => n2962, Z => n13581);
   U119 : BUF_X1 port map( A => n2960, Z => n13587);
   U120 : BUF_X1 port map( A => n2958, Z => n13593);
   U121 : BUF_X1 port map( A => n2956, Z => n13599);
   U122 : BUF_X1 port map( A => n2954, Z => n13605);
   U123 : BUF_X1 port map( A => n2952, Z => n13611);
   U124 : BUF_X1 port map( A => n2950, Z => n13617);
   U125 : BUF_X1 port map( A => n2947, Z => n13623);
   U126 : BUF_X1 port map( A => n2941, Z => n13641);
   U127 : BUF_X1 port map( A => n2939, Z => n13647);
   U128 : BUF_X1 port map( A => n2937, Z => n13653);
   U129 : BUF_X1 port map( A => n2935, Z => n13659);
   U130 : BUF_X1 port map( A => n2933, Z => n13665);
   U131 : BUF_X1 port map( A => n2931, Z => n13671);
   U132 : BUF_X1 port map( A => n2929, Z => n13677);
   U133 : BUF_X1 port map( A => n2925, Z => n13689);
   U134 : BUF_X1 port map( A => n2923, Z => n13695);
   U135 : BUF_X1 port map( A => n2921, Z => n13701);
   U136 : BUF_X1 port map( A => n2919, Z => n13707);
   U137 : BUF_X1 port map( A => n2917, Z => n13713);
   U138 : BUF_X1 port map( A => n2914, Z => n13719);
   U139 : BUF_X1 port map( A => n3034, Z => n13395);
   U140 : BUF_X1 port map( A => n3032, Z => n13401);
   U141 : BUF_X1 port map( A => n3029, Z => n13407);
   U142 : BUF_X1 port map( A => n3027, Z => n13413);
   U143 : BUF_X1 port map( A => n3025, Z => n13419);
   U144 : BUF_X1 port map( A => n3023, Z => n13425);
   U145 : BUF_X1 port map( A => n3019, Z => n13431);
   U146 : BUF_X1 port map( A => n3037, Z => n13386);
   U147 : BUF_X1 port map( A => n2875, Z => n13796);
   U148 : BUF_X1 port map( A => n2893, Z => n13760);
   U149 : BUF_X1 port map( A => n2902, Z => n13742);
   U150 : BUF_X1 port map( A => n2875, Z => n13795);
   U151 : BUF_X1 port map( A => n2902, Z => n13741);
   U152 : BUF_X1 port map( A => n2878, Z => n13790);
   U153 : BUF_X1 port map( A => n2905, Z => n13736);
   U154 : BUF_X1 port map( A => n2878, Z => n13789);
   U155 : BUF_X1 port map( A => n2905, Z => n13735);
   U156 : BUF_X1 port map( A => n2911, Z => n13724);
   U157 : BUF_X1 port map( A => n2911, Z => n13723);
   U158 : BUF_X1 port map( A => n2908, Z => n13730);
   U159 : BUF_X1 port map( A => n2908, Z => n13729);
   U160 : BUF_X1 port map( A => n2899, Z => n13748);
   U161 : BUF_X1 port map( A => n2899, Z => n13747);
   U162 : BUF_X1 port map( A => n2896, Z => n13754);
   U163 : BUF_X1 port map( A => n2896, Z => n13753);
   U164 : BUF_X1 port map( A => n2893, Z => n13759);
   U165 : BUF_X1 port map( A => n2890, Z => n13766);
   U166 : BUF_X1 port map( A => n2890, Z => n13765);
   U167 : BUF_X1 port map( A => n2887, Z => n13772);
   U168 : BUF_X1 port map( A => n2887, Z => n13771);
   U169 : BUF_X1 port map( A => n2884, Z => n13778);
   U170 : BUF_X1 port map( A => n2884, Z => n13777);
   U171 : BUF_X1 port map( A => n2881, Z => n13784);
   U172 : BUF_X1 port map( A => n2881, Z => n13783);
   U173 : BUF_X1 port map( A => n2872, Z => n13802);
   U174 : BUF_X1 port map( A => n2872, Z => n13801);
   U175 : BUF_X1 port map( A => n2869, Z => n13808);
   U176 : BUF_X1 port map( A => n2869, Z => n13807);
   U177 : BUF_X1 port map( A => n2980, Z => n13526);
   U178 : BUF_X1 port map( A => n2980, Z => n13525);
   U179 : BUF_X1 port map( A => n2923, Z => n13693);
   U180 : BUF_X1 port map( A => n2925, Z => n13688);
   U181 : BUF_X1 port map( A => n2927, Z => n13682);
   U182 : BUF_X1 port map( A => n2941, Z => n13640);
   U183 : BUF_X1 port map( A => n2941, Z => n13639);
   U184 : BUF_X1 port map( A => n2943, Z => n13634);
   U185 : BUF_X1 port map( A => n2945, Z => n13628);
   U186 : BUF_X1 port map( A => n2960, Z => n13585);
   U187 : BUF_X1 port map( A => n2962, Z => n13580);
   U188 : BUF_X1 port map( A => n2964, Z => n13574);
   U189 : BUF_X1 port map( A => n2974, Z => n13544);
   U190 : BUF_X1 port map( A => n2983, Z => n13520);
   U191 : BUF_X1 port map( A => n2983, Z => n13519);
   U192 : BUF_X1 port map( A => n2927, Z => n13681);
   U193 : BUF_X1 port map( A => n2943, Z => n13633);
   U194 : BUF_X1 port map( A => n2945, Z => n13627);
   U195 : BUF_X1 port map( A => n2964, Z => n13573);
   U196 : BUF_X1 port map( A => n3017, Z => n13436);
   U197 : BUF_X1 port map( A => n3017, Z => n13435);
   U198 : BUF_X1 port map( A => n3015, Z => n13442);
   U199 : BUF_X1 port map( A => n3015, Z => n13441);
   U200 : BUF_X1 port map( A => n3013, Z => n13448);
   U201 : BUF_X1 port map( A => n3013, Z => n13447);
   U202 : BUF_X1 port map( A => n3010, Z => n13454);
   U203 : BUF_X1 port map( A => n3010, Z => n13453);
   U204 : BUF_X1 port map( A => n3007, Z => n13460);
   U205 : BUF_X1 port map( A => n3007, Z => n13459);
   U206 : BUF_X1 port map( A => n3004, Z => n13466);
   U207 : BUF_X1 port map( A => n3004, Z => n13465);
   U208 : BUF_X1 port map( A => n3001, Z => n13472);
   U209 : BUF_X1 port map( A => n3001, Z => n13471);
   U210 : BUF_X1 port map( A => n2997, Z => n13478);
   U211 : BUF_X1 port map( A => n2997, Z => n13477);
   U212 : BUF_X1 port map( A => n2995, Z => n13484);
   U213 : BUF_X1 port map( A => n2995, Z => n13483);
   U214 : BUF_X1 port map( A => n2993, Z => n13490);
   U215 : BUF_X1 port map( A => n2993, Z => n13489);
   U216 : BUF_X1 port map( A => n2991, Z => n13496);
   U217 : BUF_X1 port map( A => n2991, Z => n13495);
   U218 : BUF_X1 port map( A => n2989, Z => n13502);
   U219 : BUF_X1 port map( A => n2989, Z => n13501);
   U220 : BUF_X1 port map( A => n2987, Z => n13508);
   U221 : BUF_X1 port map( A => n2987, Z => n13507);
   U222 : BUF_X1 port map( A => n2985, Z => n13514);
   U223 : BUF_X1 port map( A => n2985, Z => n13513);
   U224 : BUF_X1 port map( A => n2978, Z => n13532);
   U225 : BUF_X1 port map( A => n2978, Z => n13531);
   U226 : BUF_X1 port map( A => n2976, Z => n13538);
   U227 : BUF_X1 port map( A => n2976, Z => n13537);
   U228 : BUF_X1 port map( A => n2974, Z => n13543);
   U229 : BUF_X1 port map( A => n2972, Z => n13550);
   U230 : BUF_X1 port map( A => n2972, Z => n13549);
   U231 : BUF_X1 port map( A => n2970, Z => n13556);
   U232 : BUF_X1 port map( A => n2970, Z => n13555);
   U233 : BUF_X1 port map( A => n2968, Z => n13562);
   U234 : BUF_X1 port map( A => n2968, Z => n13561);
   U235 : BUF_X1 port map( A => n2966, Z => n13568);
   U236 : BUF_X1 port map( A => n2966, Z => n13567);
   U237 : BUF_X1 port map( A => n2962, Z => n13579);
   U238 : BUF_X1 port map( A => n2960, Z => n13586);
   U239 : BUF_X1 port map( A => n2958, Z => n13592);
   U240 : BUF_X1 port map( A => n2958, Z => n13591);
   U241 : BUF_X1 port map( A => n2956, Z => n13598);
   U242 : BUF_X1 port map( A => n2956, Z => n13597);
   U243 : BUF_X1 port map( A => n2954, Z => n13604);
   U244 : BUF_X1 port map( A => n2954, Z => n13603);
   U245 : BUF_X1 port map( A => n2952, Z => n13610);
   U246 : BUF_X1 port map( A => n2952, Z => n13609);
   U247 : BUF_X1 port map( A => n2950, Z => n13616);
   U248 : BUF_X1 port map( A => n2950, Z => n13615);
   U249 : BUF_X1 port map( A => n2947, Z => n13622);
   U250 : BUF_X1 port map( A => n2947, Z => n13621);
   U251 : BUF_X1 port map( A => n2939, Z => n13646);
   U252 : BUF_X1 port map( A => n2939, Z => n13645);
   U253 : BUF_X1 port map( A => n2937, Z => n13652);
   U254 : BUF_X1 port map( A => n2937, Z => n13651);
   U255 : BUF_X1 port map( A => n2935, Z => n13658);
   U256 : BUF_X1 port map( A => n2935, Z => n13657);
   U257 : BUF_X1 port map( A => n2933, Z => n13664);
   U258 : BUF_X1 port map( A => n2933, Z => n13663);
   U259 : BUF_X1 port map( A => n2931, Z => n13670);
   U260 : BUF_X1 port map( A => n2931, Z => n13669);
   U261 : BUF_X1 port map( A => n2929, Z => n13676);
   U262 : BUF_X1 port map( A => n2929, Z => n13675);
   U263 : BUF_X1 port map( A => n2925, Z => n13687);
   U264 : BUF_X1 port map( A => n2923, Z => n13694);
   U265 : BUF_X1 port map( A => n2921, Z => n13700);
   U266 : BUF_X1 port map( A => n2921, Z => n13699);
   U267 : BUF_X1 port map( A => n2919, Z => n13706);
   U268 : BUF_X1 port map( A => n2919, Z => n13705);
   U269 : BUF_X1 port map( A => n2917, Z => n13712);
   U270 : BUF_X1 port map( A => n2917, Z => n13711);
   U271 : BUF_X1 port map( A => n2914, Z => n13718);
   U272 : BUF_X1 port map( A => n2914, Z => n13717);
   U273 : BUF_X1 port map( A => n4395, Z => n13012);
   U274 : BUF_X1 port map( A => n4432, Z => n12931);
   U275 : BUF_X1 port map( A => n4395, Z => n13013);
   U276 : BUF_X1 port map( A => n4432, Z => n12932);
   U277 : BUF_X1 port map( A => n3111, Z => n13240);
   U278 : BUF_X1 port map( A => n3111, Z => n13241);
   U279 : BUF_X1 port map( A => n3034, Z => n13394);
   U280 : BUF_X1 port map( A => n3034, Z => n13393);
   U281 : BUF_X1 port map( A => n3032, Z => n13400);
   U282 : BUF_X1 port map( A => n3032, Z => n13399);
   U283 : BUF_X1 port map( A => n3029, Z => n13406);
   U284 : BUF_X1 port map( A => n3029, Z => n13405);
   U285 : BUF_X1 port map( A => n3027, Z => n13412);
   U286 : BUF_X1 port map( A => n3027, Z => n13411);
   U287 : BUF_X1 port map( A => n3025, Z => n13418);
   U288 : BUF_X1 port map( A => n3025, Z => n13417);
   U289 : BUF_X1 port map( A => n3023, Z => n13424);
   U290 : BUF_X1 port map( A => n3023, Z => n13423);
   U291 : BUF_X1 port map( A => n3019, Z => n13430);
   U292 : BUF_X1 port map( A => n3019, Z => n13429);
   U293 : BUF_X1 port map( A => n3037, Z => n13384);
   U294 : BUF_X1 port map( A => n3149, Z => n13156);
   U295 : BUF_X1 port map( A => n3149, Z => n13157);
   U296 : BUF_X1 port map( A => n3037, Z => n13385);
   U297 : BUF_X1 port map( A => n4371, Z => n13060);
   U298 : BUF_X1 port map( A => n4371, Z => n13061);
   U299 : BUF_X1 port map( A => n3087, Z => n13288);
   U300 : BUF_X1 port map( A => n3087, Z => n13289);
   U301 : BUF_X1 port map( A => n2832, Z => n14021);
   U302 : BUF_X1 port map( A => n4361, Z => n13084);
   U303 : BUF_X1 port map( A => n4404, Z => n12988);
   U304 : BUF_X1 port map( A => n4419, Z => n12961);
   U305 : BUF_X1 port map( A => n4361, Z => n13085);
   U306 : BUF_X1 port map( A => n4404, Z => n12989);
   U307 : BUF_X1 port map( A => n4419, Z => n12962);
   U308 : BUF_X1 port map( A => n3077, Z => n13312);
   U309 : BUF_X1 port map( A => n3120, Z => n13216);
   U310 : BUF_X1 port map( A => n3135, Z => n13189);
   U311 : BUF_X1 port map( A => n3077, Z => n13313);
   U312 : BUF_X1 port map( A => n3120, Z => n13217);
   U313 : BUF_X1 port map( A => n3135, Z => n13190);
   U314 : BUF_X1 port map( A => n2832, Z => n14020);
   U315 : BUF_X1 port map( A => n2832, Z => n14019);
   U316 : BUF_X1 port map( A => n4350, Z => n13102);
   U317 : BUF_X1 port map( A => n4350, Z => n13103);
   U318 : BUF_X1 port map( A => n3066, Z => n13330);
   U319 : BUF_X1 port map( A => n3066, Z => n13331);
   U320 : BUF_X1 port map( A => n4395, Z => n13014);
   U321 : BUF_X1 port map( A => n4432, Z => n12933);
   U322 : BUF_X1 port map( A => n3111, Z => n13242);
   U323 : BUF_X1 port map( A => n4324, Z => n13150);
   U324 : BUF_X1 port map( A => n4324, Z => n13151);
   U325 : BUF_X1 port map( A => n3040, Z => n13378);
   U326 : BUF_X1 port map( A => n3040, Z => n13379);
   U327 : BUF_X1 port map( A => n4338, Z => n13132);
   U328 : BUF_X1 port map( A => n4338, Z => n13133);
   U329 : BUF_X1 port map( A => n3054, Z => n13360);
   U330 : BUF_X1 port map( A => n3054, Z => n13361);
   U331 : BUF_X1 port map( A => n3149, Z => n13158);
   U332 : BUF_X1 port map( A => n4371, Z => n13062);
   U333 : BUF_X1 port map( A => n3087, Z => n13290);
   U334 : BUF_X1 port map( A => n4361, Z => n13086);
   U335 : BUF_X1 port map( A => n4404, Z => n12990);
   U336 : BUF_X1 port map( A => n4419, Z => n12963);
   U337 : BUF_X1 port map( A => n3077, Z => n13314);
   U338 : BUF_X1 port map( A => n3120, Z => n13218);
   U339 : BUF_X1 port map( A => n3135, Z => n13191);
   U340 : BUF_X1 port map( A => n4350, Z => n13104);
   U341 : BUF_X1 port map( A => n3066, Z => n13332);
   U342 : BUF_X1 port map( A => n4324, Z => n13152);
   U343 : BUF_X1 port map( A => n3040, Z => n13380);
   U344 : BUF_X1 port map( A => n4338, Z => n13134);
   U345 : BUF_X1 port map( A => n3054, Z => n13362);
   U346 : NOR3_X1 port map( A1 => n16058, A2 => n16062, A3 => n16057, ZN => 
                           n5732);
   U347 : NOR3_X1 port map( A1 => n16056, A2 => n16061, A3 => n16055, ZN => 
                           n4310);
   U348 : INV_X1 port map( A => n13822, ZN => n13813);
   U349 : INV_X1 port map( A => n13822, ZN => n13812);
   U350 : INV_X1 port map( A => n13822, ZN => n13811);
   U351 : NAND2_X1 port map( A1 => n5679, A2 => n5664, ZN => n4350);
   U352 : NAND2_X1 port map( A1 => n4282, A2 => n4273, ZN => n3066);
   U353 : NAND2_X1 port map( A1 => n2982, A2 => n2867, ZN => n2980);
   U354 : NAND2_X1 port map( A1 => n2916, A2 => n2907, ZN => n2941);
   U355 : NAND2_X1 port map( A1 => n2982, A2 => n2871, ZN => n2983);
   U356 : NAND2_X1 port map( A1 => n2916, A2 => n2886, ZN => n2927);
   U357 : NAND2_X1 port map( A1 => n2916, A2 => n2910, ZN => n2943);
   U358 : NAND2_X1 port map( A1 => n2916, A2 => n2913, ZN => n2945);
   U359 : NAND2_X1 port map( A1 => n2949, A2 => n2892, ZN => n2964);
   U360 : NAND2_X1 port map( A1 => n2982, A2 => n2913, ZN => n3017);
   U361 : NAND2_X1 port map( A1 => n2982, A2 => n2910, ZN => n3015);
   U362 : NAND2_X1 port map( A1 => n2982, A2 => n2907, ZN => n3013);
   U363 : NAND2_X1 port map( A1 => n2982, A2 => n2904, ZN => n3010);
   U364 : NAND2_X1 port map( A1 => n2982, A2 => n2901, ZN => n3007);
   U365 : NAND2_X1 port map( A1 => n2982, A2 => n2898, ZN => n3004);
   U366 : NAND2_X1 port map( A1 => n2982, A2 => n2895, ZN => n3001);
   U367 : NAND2_X1 port map( A1 => n2982, A2 => n2892, ZN => n2997);
   U368 : NAND2_X1 port map( A1 => n2982, A2 => n2889, ZN => n2995);
   U369 : NAND2_X1 port map( A1 => n2982, A2 => n2886, ZN => n2993);
   U370 : NAND2_X1 port map( A1 => n2982, A2 => n2883, ZN => n2991);
   U371 : NAND2_X1 port map( A1 => n2982, A2 => n2880, ZN => n2989);
   U372 : NAND2_X1 port map( A1 => n2982, A2 => n2877, ZN => n2987);
   U373 : NAND2_X1 port map( A1 => n2982, A2 => n2874, ZN => n2985);
   U374 : NAND2_X1 port map( A1 => n2949, A2 => n2913, ZN => n2978);
   U375 : NAND2_X1 port map( A1 => n2949, A2 => n2910, ZN => n2976);
   U376 : NAND2_X1 port map( A1 => n2949, A2 => n2907, ZN => n2974);
   U377 : NAND2_X1 port map( A1 => n2949, A2 => n2904, ZN => n2972);
   U378 : NAND2_X1 port map( A1 => n2949, A2 => n2901, ZN => n2970);
   U379 : NAND2_X1 port map( A1 => n2949, A2 => n2898, ZN => n2968);
   U380 : NAND2_X1 port map( A1 => n2949, A2 => n2895, ZN => n2966);
   U381 : NAND2_X1 port map( A1 => n2949, A2 => n2889, ZN => n2962);
   U382 : NAND2_X1 port map( A1 => n2949, A2 => n2886, ZN => n2960);
   U383 : NAND2_X1 port map( A1 => n2949, A2 => n2883, ZN => n2958);
   U384 : NAND2_X1 port map( A1 => n2949, A2 => n2880, ZN => n2956);
   U385 : NAND2_X1 port map( A1 => n2949, A2 => n2877, ZN => n2954);
   U386 : NAND2_X1 port map( A1 => n2949, A2 => n2874, ZN => n2952);
   U387 : NAND2_X1 port map( A1 => n2949, A2 => n2871, ZN => n2950);
   U388 : NAND2_X1 port map( A1 => n2949, A2 => n2867, ZN => n2947);
   U389 : NAND2_X1 port map( A1 => n2916, A2 => n2904, ZN => n2939);
   U390 : NAND2_X1 port map( A1 => n2916, A2 => n2901, ZN => n2937);
   U391 : NAND2_X1 port map( A1 => n2916, A2 => n2898, ZN => n2935);
   U392 : NAND2_X1 port map( A1 => n2916, A2 => n2895, ZN => n2933);
   U393 : NAND2_X1 port map( A1 => n2916, A2 => n2892, ZN => n2931);
   U394 : NAND2_X1 port map( A1 => n2916, A2 => n2889, ZN => n2929);
   U395 : NAND2_X1 port map( A1 => n2916, A2 => n2883, ZN => n2925);
   U396 : NAND2_X1 port map( A1 => n2916, A2 => n2880, ZN => n2923);
   U397 : NAND2_X1 port map( A1 => n2916, A2 => n2877, ZN => n2921);
   U398 : NAND2_X1 port map( A1 => n2916, A2 => n2874, ZN => n2919);
   U399 : NAND2_X1 port map( A1 => n2916, A2 => n2871, ZN => n2917);
   U400 : NAND2_X1 port map( A1 => n2916, A2 => n2867, ZN => n2914);
   U401 : NAND2_X1 port map( A1 => n5710, A2 => n5664, ZN => n4432);
   U402 : NAND2_X1 port map( A1 => n4299, A2 => n4273, ZN => n3149);
   U403 : BUF_X1 port map( A => n2961, Z => n13583);
   U404 : BUF_X1 port map( A => n4354, Z => n13093);
   U405 : BUF_X1 port map( A => n4354, Z => n13094);
   U406 : BUF_X1 port map( A => n3070, Z => n13321);
   U407 : BUF_X1 port map( A => n3070, Z => n13322);
   U408 : BUF_X1 port map( A => n4343, Z => n13120);
   U409 : BUF_X1 port map( A => n4369, Z => n13066);
   U410 : BUF_X1 port map( A => n4380, Z => n13039);
   U411 : BUF_X1 port map( A => n4406, Z => n12985);
   U412 : BUF_X1 port map( A => n4421, Z => n12958);
   U413 : BUF_X1 port map( A => n4343, Z => n13121);
   U414 : BUF_X1 port map( A => n4369, Z => n13067);
   U415 : BUF_X1 port map( A => n4380, Z => n13040);
   U416 : BUF_X1 port map( A => n4406, Z => n12986);
   U417 : BUF_X1 port map( A => n4421, Z => n12959);
   U418 : BUF_X1 port map( A => n3059, Z => n13348);
   U419 : BUF_X1 port map( A => n3085, Z => n13294);
   U420 : BUF_X1 port map( A => n3096, Z => n13267);
   U421 : BUF_X1 port map( A => n3122, Z => n13213);
   U422 : BUF_X1 port map( A => n3137, Z => n13186);
   U423 : BUF_X1 port map( A => n3148, Z => n13159);
   U424 : BUF_X1 port map( A => n3059, Z => n13349);
   U425 : BUF_X1 port map( A => n3085, Z => n13295);
   U426 : BUF_X1 port map( A => n3096, Z => n13268);
   U427 : BUF_X1 port map( A => n3122, Z => n13214);
   U428 : BUF_X1 port map( A => n3137, Z => n13187);
   U429 : BUF_X1 port map( A => n3148, Z => n13160);
   U430 : BUF_X1 port map( A => n2834, Z => n14010);
   U431 : BUF_X1 port map( A => n2876, Z => n13792);
   U432 : BUF_X1 port map( A => n2876, Z => n13793);
   U433 : BUF_X1 port map( A => n2894, Z => n13756);
   U434 : BUF_X1 port map( A => n2903, Z => n13738);
   U435 : BUF_X1 port map( A => n2903, Z => n13739);
   U436 : BUF_X1 port map( A => n2879, Z => n13786);
   U437 : BUF_X1 port map( A => n2879, Z => n13787);
   U438 : BUF_X1 port map( A => n2834, Z => n14011);
   U439 : BUF_X1 port map( A => n2906, Z => n13732);
   U440 : BUF_X1 port map( A => n2906, Z => n13733);
   U441 : BUF_X1 port map( A => n2926, Z => n13684);
   U442 : BUF_X1 port map( A => n2926, Z => n13685);
   U443 : BUF_X1 port map( A => n2928, Z => n13678);
   U444 : BUF_X1 port map( A => n2928, Z => n13679);
   U445 : BUF_X1 port map( A => n2942, Z => n13637);
   U446 : BUF_X1 port map( A => n2944, Z => n13630);
   U447 : BUF_X1 port map( A => n2944, Z => n13631);
   U448 : BUF_X1 port map( A => n2946, Z => n13624);
   U449 : BUF_X1 port map( A => n2946, Z => n13625);
   U450 : BUF_X1 port map( A => n2961, Z => n13582);
   U451 : BUF_X1 port map( A => n2963, Z => n13576);
   U452 : BUF_X1 port map( A => n2963, Z => n13577);
   U453 : BUF_X1 port map( A => n2965, Z => n13570);
   U454 : BUF_X1 port map( A => n2965, Z => n13571);
   U455 : BUF_X1 port map( A => n2975, Z => n13540);
   U456 : BUF_X1 port map( A => n2975, Z => n13541);
   U457 : BUF_X1 port map( A => n2984, Z => n13517);
   U458 : BUF_X1 port map( A => n3030, Z => n13402);
   U459 : BUF_X1 port map( A => n3030, Z => n13403);
   U460 : BUF_X1 port map( A => n3028, Z => n13408);
   U461 : BUF_X1 port map( A => n3028, Z => n13409);
   U462 : BUF_X1 port map( A => n3018, Z => n13432);
   U463 : BUF_X1 port map( A => n3018, Z => n13433);
   U464 : BUF_X1 port map( A => n3005, Z => n13462);
   U465 : BUF_X1 port map( A => n3005, Z => n13463);
   U466 : BUF_X1 port map( A => n2986, Z => n13510);
   U467 : BUF_X1 port map( A => n2986, Z => n13511);
   U468 : BUF_X1 port map( A => n2984, Z => n13516);
   U469 : BUF_X1 port map( A => n2948, Z => n13618);
   U470 : BUF_X1 port map( A => n2948, Z => n13619);
   U471 : BUF_X1 port map( A => n2942, Z => n13636);
   U472 : BUF_X1 port map( A => n2930, Z => n13672);
   U473 : BUF_X1 port map( A => n2930, Z => n13673);
   U474 : BUF_X1 port map( A => n2924, Z => n13690);
   U475 : BUF_X1 port map( A => n2924, Z => n13691);
   U476 : BUF_X1 port map( A => n2909, Z => n13726);
   U477 : BUF_X1 port map( A => n2909, Z => n13727);
   U478 : BUF_X1 port map( A => n2897, Z => n13750);
   U479 : BUF_X1 port map( A => n2897, Z => n13751);
   U480 : BUF_X1 port map( A => n2894, Z => n13757);
   U481 : BUF_X1 port map( A => n2882, Z => n13780);
   U482 : BUF_X1 port map( A => n2882, Z => n13781);
   U483 : BUF_X1 port map( A => n2870, Z => n13804);
   U484 : BUF_X1 port map( A => n2870, Z => n13805);
   U485 : BUF_X1 port map( A => n4355, Z => n13090);
   U486 : BUF_X1 port map( A => n4355, Z => n13091);
   U487 : BUF_X1 port map( A => n3071, Z => n13318);
   U488 : BUF_X1 port map( A => n3071, Z => n13319);
   U489 : BUF_X1 port map( A => n4396, Z => n13009);
   U490 : BUF_X1 port map( A => n4396, Z => n13010);
   U491 : BUF_X1 port map( A => n4344, Z => n13117);
   U492 : BUF_X1 port map( A => n4370, Z => n13063);
   U493 : BUF_X1 port map( A => n4381, Z => n13036);
   U494 : BUF_X1 port map( A => n4407, Z => n12982);
   U495 : BUF_X1 port map( A => n4422, Z => n12955);
   U496 : BUF_X1 port map( A => n4433, Z => n12928);
   U497 : BUF_X1 port map( A => n4344, Z => n13118);
   U498 : BUF_X1 port map( A => n4370, Z => n13064);
   U499 : BUF_X1 port map( A => n4381, Z => n13037);
   U500 : BUF_X1 port map( A => n4407, Z => n12983);
   U501 : BUF_X1 port map( A => n4422, Z => n12956);
   U502 : BUF_X1 port map( A => n4433, Z => n12929);
   U503 : BUF_X1 port map( A => n3060, Z => n13345);
   U504 : BUF_X1 port map( A => n3086, Z => n13291);
   U505 : BUF_X1 port map( A => n3097, Z => n13264);
   U506 : BUF_X1 port map( A => n3112, Z => n13237);
   U507 : BUF_X1 port map( A => n3123, Z => n13210);
   U508 : BUF_X1 port map( A => n3138, Z => n13183);
   U509 : BUF_X1 port map( A => n3060, Z => n13346);
   U510 : BUF_X1 port map( A => n3086, Z => n13292);
   U511 : BUF_X1 port map( A => n3097, Z => n13265);
   U512 : BUF_X1 port map( A => n3112, Z => n13238);
   U513 : BUF_X1 port map( A => n3123, Z => n13211);
   U514 : BUF_X1 port map( A => n3138, Z => n13184);
   U515 : NAND2_X1 port map( A1 => n5661, A2 => n5664, ZN => n4338);
   U516 : NAND2_X1 port map( A1 => n5714, A2 => n5664, ZN => n4395);
   U517 : NAND2_X1 port map( A1 => n4272, A2 => n4273, ZN => n3054);
   U518 : NAND2_X1 port map( A1 => n4301, A2 => n4273, ZN => n3111);
   U519 : BUF_X1 port map( A => n4345, Z => n13114);
   U520 : BUF_X1 port map( A => n4351, Z => n13099);
   U521 : BUF_X1 port map( A => n4345, Z => n13115);
   U522 : BUF_X1 port map( A => n4351, Z => n13100);
   U523 : BUF_X1 port map( A => n3061, Z => n13342);
   U524 : BUF_X1 port map( A => n3067, Z => n13327);
   U525 : BUF_X1 port map( A => n3061, Z => n13343);
   U526 : BUF_X1 port map( A => n3067, Z => n13328);
   U527 : BUF_X1 port map( A => n4334, Z => n13141);
   U528 : BUF_X1 port map( A => n4340, Z => n13126);
   U529 : BUF_X1 port map( A => n4360, Z => n13087);
   U530 : BUF_X1 port map( A => n4366, Z => n13072);
   U531 : BUF_X1 port map( A => n4377, Z => n13045);
   U532 : BUF_X1 port map( A => n4386, Z => n13033);
   U533 : BUF_X1 port map( A => n4397, Z => n13006);
   U534 : BUF_X1 port map( A => n4392, Z => n13018);
   U535 : BUF_X1 port map( A => n4403, Z => n12991);
   U536 : BUF_X1 port map( A => n4412, Z => n12979);
   U537 : BUF_X1 port map( A => n4423, Z => n12952);
   U538 : BUF_X1 port map( A => n4418, Z => n12964);
   U539 : BUF_X1 port map( A => n4429, Z => n12937);
   U540 : BUF_X1 port map( A => n4334, Z => n13142);
   U541 : BUF_X1 port map( A => n4340, Z => n13127);
   U542 : BUF_X1 port map( A => n4360, Z => n13088);
   U543 : BUF_X1 port map( A => n4366, Z => n13073);
   U544 : BUF_X1 port map( A => n4377, Z => n13046);
   U545 : BUF_X1 port map( A => n4386, Z => n13034);
   U546 : BUF_X1 port map( A => n4397, Z => n13007);
   U547 : BUF_X1 port map( A => n4392, Z => n13019);
   U548 : BUF_X1 port map( A => n4403, Z => n12992);
   U549 : BUF_X1 port map( A => n4412, Z => n12980);
   U550 : BUF_X1 port map( A => n4423, Z => n12953);
   U551 : BUF_X1 port map( A => n4418, Z => n12965);
   U552 : BUF_X1 port map( A => n4429, Z => n12938);
   U553 : BUF_X1 port map( A => n3050, Z => n13369);
   U554 : BUF_X1 port map( A => n3056, Z => n13354);
   U555 : BUF_X1 port map( A => n3076, Z => n13315);
   U556 : BUF_X1 port map( A => n3082, Z => n13300);
   U557 : BUF_X1 port map( A => n3093, Z => n13273);
   U558 : BUF_X1 port map( A => n3102, Z => n13261);
   U559 : BUF_X1 port map( A => n3113, Z => n13234);
   U560 : BUF_X1 port map( A => n3108, Z => n13246);
   U561 : BUF_X1 port map( A => n3119, Z => n13219);
   U562 : BUF_X1 port map( A => n3128, Z => n13207);
   U563 : BUF_X1 port map( A => n3139, Z => n13180);
   U564 : BUF_X1 port map( A => n3134, Z => n13192);
   U565 : BUF_X1 port map( A => n3145, Z => n13165);
   U566 : BUF_X1 port map( A => n3050, Z => n13370);
   U567 : BUF_X1 port map( A => n3056, Z => n13355);
   U568 : BUF_X1 port map( A => n3076, Z => n13316);
   U569 : BUF_X1 port map( A => n3082, Z => n13301);
   U570 : BUF_X1 port map( A => n3093, Z => n13274);
   U571 : BUF_X1 port map( A => n3102, Z => n13262);
   U572 : BUF_X1 port map( A => n3113, Z => n13235);
   U573 : BUF_X1 port map( A => n3108, Z => n13247);
   U574 : BUF_X1 port map( A => n3119, Z => n13220);
   U575 : BUF_X1 port map( A => n3128, Z => n13208);
   U576 : BUF_X1 port map( A => n3139, Z => n13181);
   U577 : BUF_X1 port map( A => n3134, Z => n13193);
   U578 : BUF_X1 port map( A => n3145, Z => n13166);
   U579 : BUF_X1 port map( A => n2981, Z => n13522);
   U580 : BUF_X1 port map( A => n2981, Z => n13523);
   U581 : BUF_X1 port map( A => n3035, Z => n13390);
   U582 : BUF_X1 port map( A => n3035, Z => n13391);
   U583 : BUF_X1 port map( A => n3033, Z => n13396);
   U584 : BUF_X1 port map( A => n3033, Z => n13397);
   U585 : BUF_X1 port map( A => n3026, Z => n13414);
   U586 : BUF_X1 port map( A => n3026, Z => n13415);
   U587 : BUF_X1 port map( A => n3024, Z => n13420);
   U588 : BUF_X1 port map( A => n3024, Z => n13421);
   U589 : BUF_X1 port map( A => n3020, Z => n13426);
   U590 : BUF_X1 port map( A => n3020, Z => n13427);
   U591 : BUF_X1 port map( A => n3016, Z => n13438);
   U592 : BUF_X1 port map( A => n3016, Z => n13439);
   U593 : BUF_X1 port map( A => n3014, Z => n13444);
   U594 : BUF_X1 port map( A => n3014, Z => n13445);
   U595 : BUF_X1 port map( A => n3011, Z => n13450);
   U596 : BUF_X1 port map( A => n3011, Z => n13451);
   U597 : BUF_X1 port map( A => n3008, Z => n13456);
   U598 : BUF_X1 port map( A => n3008, Z => n13457);
   U599 : BUF_X1 port map( A => n3002, Z => n13468);
   U600 : BUF_X1 port map( A => n3002, Z => n13469);
   U601 : BUF_X1 port map( A => n2998, Z => n13474);
   U602 : BUF_X1 port map( A => n2998, Z => n13475);
   U603 : BUF_X1 port map( A => n2996, Z => n13480);
   U604 : BUF_X1 port map( A => n2996, Z => n13481);
   U605 : BUF_X1 port map( A => n2994, Z => n13486);
   U606 : BUF_X1 port map( A => n2994, Z => n13487);
   U607 : BUF_X1 port map( A => n2992, Z => n13492);
   U608 : BUF_X1 port map( A => n2992, Z => n13493);
   U609 : BUF_X1 port map( A => n2990, Z => n13498);
   U610 : BUF_X1 port map( A => n2990, Z => n13499);
   U611 : BUF_X1 port map( A => n2988, Z => n13504);
   U612 : BUF_X1 port map( A => n2988, Z => n13505);
   U613 : BUF_X1 port map( A => n2979, Z => n13528);
   U614 : BUF_X1 port map( A => n2979, Z => n13529);
   U615 : BUF_X1 port map( A => n2977, Z => n13534);
   U616 : BUF_X1 port map( A => n2977, Z => n13535);
   U617 : BUF_X1 port map( A => n2973, Z => n13546);
   U618 : BUF_X1 port map( A => n2973, Z => n13547);
   U619 : BUF_X1 port map( A => n2971, Z => n13552);
   U620 : BUF_X1 port map( A => n2971, Z => n13553);
   U621 : BUF_X1 port map( A => n2969, Z => n13558);
   U622 : BUF_X1 port map( A => n2969, Z => n13559);
   U623 : BUF_X1 port map( A => n2967, Z => n13564);
   U624 : BUF_X1 port map( A => n2967, Z => n13565);
   U625 : BUF_X1 port map( A => n2959, Z => n13588);
   U626 : BUF_X1 port map( A => n2959, Z => n13589);
   U627 : BUF_X1 port map( A => n2957, Z => n13594);
   U628 : BUF_X1 port map( A => n2957, Z => n13595);
   U629 : BUF_X1 port map( A => n2955, Z => n13600);
   U630 : BUF_X1 port map( A => n2955, Z => n13601);
   U631 : BUF_X1 port map( A => n2953, Z => n13606);
   U632 : BUF_X1 port map( A => n2953, Z => n13607);
   U633 : BUF_X1 port map( A => n2951, Z => n13612);
   U634 : BUF_X1 port map( A => n2951, Z => n13613);
   U635 : BUF_X1 port map( A => n2940, Z => n13642);
   U636 : BUF_X1 port map( A => n2940, Z => n13643);
   U637 : BUF_X1 port map( A => n2938, Z => n13648);
   U638 : BUF_X1 port map( A => n2938, Z => n13649);
   U639 : BUF_X1 port map( A => n2936, Z => n13654);
   U640 : BUF_X1 port map( A => n2936, Z => n13655);
   U641 : BUF_X1 port map( A => n2934, Z => n13660);
   U642 : BUF_X1 port map( A => n2934, Z => n13661);
   U643 : BUF_X1 port map( A => n2932, Z => n13666);
   U644 : BUF_X1 port map( A => n2932, Z => n13667);
   U645 : BUF_X1 port map( A => n2922, Z => n13696);
   U646 : BUF_X1 port map( A => n2922, Z => n13697);
   U647 : BUF_X1 port map( A => n2920, Z => n13702);
   U648 : BUF_X1 port map( A => n2920, Z => n13703);
   U649 : BUF_X1 port map( A => n2918, Z => n13708);
   U650 : BUF_X1 port map( A => n2918, Z => n13709);
   U651 : BUF_X1 port map( A => n2915, Z => n13714);
   U652 : BUF_X1 port map( A => n2915, Z => n13715);
   U653 : BUF_X1 port map( A => n2912, Z => n13720);
   U654 : BUF_X1 port map( A => n2912, Z => n13721);
   U655 : BUF_X1 port map( A => n2900, Z => n13744);
   U656 : BUF_X1 port map( A => n2900, Z => n13745);
   U657 : BUF_X1 port map( A => n2891, Z => n13762);
   U658 : BUF_X1 port map( A => n2891, Z => n13763);
   U659 : BUF_X1 port map( A => n2888, Z => n13768);
   U660 : BUF_X1 port map( A => n2888, Z => n13769);
   U661 : BUF_X1 port map( A => n2885, Z => n13774);
   U662 : BUF_X1 port map( A => n2885, Z => n13775);
   U663 : BUF_X1 port map( A => n2873, Z => n13798);
   U664 : BUF_X1 port map( A => n2873, Z => n13799);
   U665 : BUF_X1 port map( A => n3036, Z => n13387);
   U666 : BUF_X1 port map( A => n4346, Z => n13111);
   U667 : BUF_X1 port map( A => n4352, Z => n13096);
   U668 : BUF_X1 port map( A => n4346, Z => n13112);
   U669 : BUF_X1 port map( A => n4352, Z => n13097);
   U670 : BUF_X1 port map( A => n3062, Z => n13339);
   U671 : BUF_X1 port map( A => n3068, Z => n13324);
   U672 : BUF_X1 port map( A => n3062, Z => n13340);
   U673 : BUF_X1 port map( A => n3068, Z => n13325);
   U674 : BUF_X1 port map( A => n3036, Z => n13388);
   U675 : BUF_X1 port map( A => n4335, Z => n13138);
   U676 : BUF_X1 port map( A => n4341, Z => n13123);
   U677 : BUF_X1 port map( A => n4372, Z => n13057);
   U678 : BUF_X1 port map( A => n4367, Z => n13069);
   U679 : BUF_X1 port map( A => n4378, Z => n13042);
   U680 : BUF_X1 port map( A => n4387, Z => n13030);
   U681 : BUF_X1 port map( A => n4398, Z => n13003);
   U682 : BUF_X1 port map( A => n4393, Z => n13015);
   U683 : BUF_X1 port map( A => n4413, Z => n12976);
   U684 : BUF_X1 port map( A => n4424, Z => n12949);
   U685 : BUF_X1 port map( A => n4430, Z => n12934);
   U686 : BUF_X1 port map( A => n4335, Z => n13139);
   U687 : BUF_X1 port map( A => n4341, Z => n13124);
   U688 : BUF_X1 port map( A => n4372, Z => n13058);
   U689 : BUF_X1 port map( A => n4367, Z => n13070);
   U690 : BUF_X1 port map( A => n4378, Z => n13043);
   U691 : BUF_X1 port map( A => n4387, Z => n13031);
   U692 : BUF_X1 port map( A => n4398, Z => n13004);
   U693 : BUF_X1 port map( A => n4393, Z => n13016);
   U694 : BUF_X1 port map( A => n4413, Z => n12977);
   U695 : BUF_X1 port map( A => n4424, Z => n12950);
   U696 : BUF_X1 port map( A => n4430, Z => n12935);
   U697 : BUF_X1 port map( A => n3051, Z => n13366);
   U698 : BUF_X1 port map( A => n3057, Z => n13351);
   U699 : BUF_X1 port map( A => n3088, Z => n13285);
   U700 : BUF_X1 port map( A => n3083, Z => n13297);
   U701 : BUF_X1 port map( A => n3094, Z => n13270);
   U702 : BUF_X1 port map( A => n3103, Z => n13258);
   U703 : BUF_X1 port map( A => n3114, Z => n13231);
   U704 : BUF_X1 port map( A => n3109, Z => n13243);
   U705 : BUF_X1 port map( A => n3129, Z => n13204);
   U706 : BUF_X1 port map( A => n3140, Z => n13177);
   U707 : BUF_X1 port map( A => n3146, Z => n13162);
   U708 : BUF_X1 port map( A => n3051, Z => n13367);
   U709 : BUF_X1 port map( A => n3057, Z => n13352);
   U710 : BUF_X1 port map( A => n3088, Z => n13286);
   U711 : BUF_X1 port map( A => n3083, Z => n13298);
   U712 : BUF_X1 port map( A => n3094, Z => n13271);
   U713 : BUF_X1 port map( A => n3103, Z => n13259);
   U714 : BUF_X1 port map( A => n3114, Z => n13232);
   U715 : BUF_X1 port map( A => n3109, Z => n13244);
   U716 : BUF_X1 port map( A => n3129, Z => n13205);
   U717 : BUF_X1 port map( A => n3140, Z => n13178);
   U718 : BUF_X1 port map( A => n3146, Z => n13163);
   U719 : BUF_X1 port map( A => n4339, Z => n13129);
   U720 : BUF_X1 port map( A => n4339, Z => n13130);
   U721 : BUF_X1 port map( A => n4365, Z => n13075);
   U722 : BUF_X1 port map( A => n4376, Z => n13048);
   U723 : BUF_X1 port map( A => n4391, Z => n13021);
   U724 : BUF_X1 port map( A => n4402, Z => n12994);
   U725 : BUF_X1 port map( A => n4417, Z => n12967);
   U726 : BUF_X1 port map( A => n4428, Z => n12940);
   U727 : BUF_X1 port map( A => n4365, Z => n13076);
   U728 : BUF_X1 port map( A => n4376, Z => n13049);
   U729 : BUF_X1 port map( A => n4391, Z => n13022);
   U730 : BUF_X1 port map( A => n4402, Z => n12995);
   U731 : BUF_X1 port map( A => n4417, Z => n12968);
   U732 : BUF_X1 port map( A => n4428, Z => n12941);
   U733 : BUF_X1 port map( A => n3055, Z => n13357);
   U734 : BUF_X1 port map( A => n3081, Z => n13303);
   U735 : BUF_X1 port map( A => n3092, Z => n13276);
   U736 : BUF_X1 port map( A => n3107, Z => n13249);
   U737 : BUF_X1 port map( A => n3118, Z => n13222);
   U738 : BUF_X1 port map( A => n3133, Z => n13195);
   U739 : BUF_X1 port map( A => n3144, Z => n13168);
   U740 : BUF_X1 port map( A => n3055, Z => n13358);
   U741 : BUF_X1 port map( A => n3081, Z => n13304);
   U742 : BUF_X1 port map( A => n3092, Z => n13277);
   U743 : BUF_X1 port map( A => n3107, Z => n13250);
   U744 : BUF_X1 port map( A => n3118, Z => n13223);
   U745 : BUF_X1 port map( A => n3133, Z => n13196);
   U746 : BUF_X1 port map( A => n3144, Z => n13169);
   U747 : BUF_X1 port map( A => n4354, Z => n13095);
   U748 : BUF_X1 port map( A => n3070, Z => n13323);
   U749 : BUF_X1 port map( A => n4343, Z => n13122);
   U750 : BUF_X1 port map( A => n4369, Z => n13068);
   U751 : BUF_X1 port map( A => n4380, Z => n13041);
   U752 : BUF_X1 port map( A => n4406, Z => n12987);
   U753 : BUF_X1 port map( A => n4421, Z => n12960);
   U754 : BUF_X1 port map( A => n3059, Z => n13350);
   U755 : BUF_X1 port map( A => n3085, Z => n13296);
   U756 : BUF_X1 port map( A => n3096, Z => n13269);
   U757 : BUF_X1 port map( A => n3137, Z => n13188);
   U758 : BUF_X1 port map( A => n3148, Z => n13161);
   U759 : BUF_X1 port map( A => n3122, Z => n13215);
   U760 : NAND2_X1 port map( A1 => n2877, A2 => n2868, ZN => n2875);
   U761 : NAND2_X1 port map( A1 => n2904, A2 => n2868, ZN => n2902);
   U762 : NAND2_X1 port map( A1 => n2880, A2 => n2868, ZN => n2878);
   U763 : NAND2_X1 port map( A1 => n2907, A2 => n2868, ZN => n2905);
   U764 : NAND2_X1 port map( A1 => n2913, A2 => n2868, ZN => n2911);
   U765 : NAND2_X1 port map( A1 => n2910, A2 => n2868, ZN => n2908);
   U766 : NAND2_X1 port map( A1 => n2901, A2 => n2868, ZN => n2899);
   U767 : NAND2_X1 port map( A1 => n2898, A2 => n2868, ZN => n2896);
   U768 : NAND2_X1 port map( A1 => n2895, A2 => n2868, ZN => n2893);
   U769 : NAND2_X1 port map( A1 => n2892, A2 => n2868, ZN => n2890);
   U770 : NAND2_X1 port map( A1 => n2889, A2 => n2868, ZN => n2887);
   U771 : NAND2_X1 port map( A1 => n2886, A2 => n2868, ZN => n2884);
   U772 : NAND2_X1 port map( A1 => n2883, A2 => n2868, ZN => n2881);
   U773 : NAND2_X1 port map( A1 => n2874, A2 => n2868, ZN => n2872);
   U774 : NAND2_X1 port map( A1 => n2871, A2 => n2868, ZN => n2869);
   U775 : NAND2_X1 port map( A1 => n2867, A2 => n2868, ZN => n2832);
   U776 : BUF_X1 port map( A => n3030, Z => n13404);
   U777 : BUF_X1 port map( A => n3028, Z => n13410);
   U778 : BUF_X1 port map( A => n2834, Z => n14012);
   U779 : BUF_X1 port map( A => n2876, Z => n13794);
   U780 : BUF_X1 port map( A => n2903, Z => n13740);
   U781 : BUF_X1 port map( A => n2924, Z => n13692);
   U782 : BUF_X1 port map( A => n2942, Z => n13638);
   U783 : BUF_X1 port map( A => n2984, Z => n13518);
   U784 : BUF_X1 port map( A => n2879, Z => n13788);
   U785 : BUF_X1 port map( A => n2906, Z => n13734);
   U786 : BUF_X1 port map( A => n2928, Z => n13680);
   U787 : BUF_X1 port map( A => n2944, Z => n13632);
   U788 : BUF_X1 port map( A => n2946, Z => n13626);
   U789 : BUF_X1 port map( A => n2965, Z => n13572);
   U790 : BUF_X1 port map( A => n3018, Z => n13434);
   U791 : BUF_X1 port map( A => n3005, Z => n13464);
   U792 : BUF_X1 port map( A => n2986, Z => n13512);
   U793 : BUF_X1 port map( A => n2975, Z => n13542);
   U794 : BUF_X1 port map( A => n2948, Z => n13620);
   U795 : BUF_X1 port map( A => n2930, Z => n13674);
   U796 : BUF_X1 port map( A => n2909, Z => n13728);
   U797 : BUF_X1 port map( A => n2897, Z => n13752);
   U798 : BUF_X1 port map( A => n2894, Z => n13758);
   U799 : BUF_X1 port map( A => n2882, Z => n13782);
   U800 : BUF_X1 port map( A => n2870, Z => n13806);
   U801 : BUF_X1 port map( A => n4348, Z => n13108);
   U802 : BUF_X1 port map( A => n4348, Z => n13109);
   U803 : BUF_X1 port map( A => n4337, Z => n13135);
   U804 : BUF_X1 port map( A => n4363, Z => n13081);
   U805 : BUF_X1 port map( A => n4374, Z => n13054);
   U806 : BUF_X1 port map( A => n4389, Z => n13027);
   U807 : BUF_X1 port map( A => n4400, Z => n13000);
   U808 : BUF_X1 port map( A => n4415, Z => n12973);
   U809 : BUF_X1 port map( A => n4426, Z => n12946);
   U810 : BUF_X1 port map( A => n4337, Z => n13136);
   U811 : BUF_X1 port map( A => n4363, Z => n13082);
   U812 : BUF_X1 port map( A => n4374, Z => n13055);
   U813 : BUF_X1 port map( A => n4389, Z => n13028);
   U814 : BUF_X1 port map( A => n4400, Z => n13001);
   U815 : BUF_X1 port map( A => n4415, Z => n12974);
   U816 : BUF_X1 port map( A => n4426, Z => n12947);
   U817 : BUF_X1 port map( A => n3053, Z => n13363);
   U818 : BUF_X1 port map( A => n3064, Z => n13336);
   U819 : BUF_X1 port map( A => n3079, Z => n13309);
   U820 : BUF_X1 port map( A => n3090, Z => n13282);
   U821 : BUF_X1 port map( A => n3105, Z => n13255);
   U822 : BUF_X1 port map( A => n3116, Z => n13228);
   U823 : BUF_X1 port map( A => n3131, Z => n13201);
   U824 : BUF_X1 port map( A => n3142, Z => n13174);
   U825 : BUF_X1 port map( A => n3053, Z => n13364);
   U826 : BUF_X1 port map( A => n3064, Z => n13337);
   U827 : BUF_X1 port map( A => n3079, Z => n13310);
   U828 : BUF_X1 port map( A => n3090, Z => n13283);
   U829 : BUF_X1 port map( A => n3105, Z => n13256);
   U830 : BUF_X1 port map( A => n3116, Z => n13229);
   U831 : BUF_X1 port map( A => n3131, Z => n13202);
   U832 : BUF_X1 port map( A => n3142, Z => n13175);
   U833 : BUF_X1 port map( A => n4349, Z => n13105);
   U834 : BUF_X1 port map( A => n4349, Z => n13106);
   U835 : BUF_X1 port map( A => n3065, Z => n13333);
   U836 : BUF_X1 port map( A => n3065, Z => n13334);
   U837 : BUF_X1 port map( A => n4375, Z => n13051);
   U838 : BUF_X1 port map( A => n4375, Z => n13052);
   U839 : BUF_X1 port map( A => n4364, Z => n13078);
   U840 : BUF_X1 port map( A => n4390, Z => n13024);
   U841 : BUF_X1 port map( A => n4401, Z => n12997);
   U842 : BUF_X1 port map( A => n4416, Z => n12970);
   U843 : BUF_X1 port map( A => n4427, Z => n12943);
   U844 : BUF_X1 port map( A => n4364, Z => n13079);
   U845 : BUF_X1 port map( A => n4390, Z => n13025);
   U846 : BUF_X1 port map( A => n4401, Z => n12998);
   U847 : BUF_X1 port map( A => n4416, Z => n12971);
   U848 : BUF_X1 port map( A => n4427, Z => n12944);
   U849 : BUF_X1 port map( A => n3080, Z => n13306);
   U850 : BUF_X1 port map( A => n3091, Z => n13279);
   U851 : BUF_X1 port map( A => n3106, Z => n13252);
   U852 : BUF_X1 port map( A => n3117, Z => n13225);
   U853 : BUF_X1 port map( A => n3132, Z => n13198);
   U854 : BUF_X1 port map( A => n3143, Z => n13171);
   U855 : BUF_X1 port map( A => n3080, Z => n13307);
   U856 : BUF_X1 port map( A => n3091, Z => n13280);
   U857 : BUF_X1 port map( A => n3106, Z => n13253);
   U858 : BUF_X1 port map( A => n3117, Z => n13226);
   U859 : BUF_X1 port map( A => n3132, Z => n13199);
   U860 : BUF_X1 port map( A => n3143, Z => n13172);
   U861 : BUF_X1 port map( A => n4355, Z => n13092);
   U862 : BUF_X1 port map( A => n3071, Z => n13320);
   U863 : BUF_X1 port map( A => n2963, Z => n13578);
   U864 : BUF_X1 port map( A => n4396, Z => n13011);
   U865 : BUF_X1 port map( A => n4344, Z => n13119);
   U866 : BUF_X1 port map( A => n4370, Z => n13065);
   U867 : BUF_X1 port map( A => n4381, Z => n13038);
   U868 : BUF_X1 port map( A => n4407, Z => n12984);
   U869 : BUF_X1 port map( A => n4422, Z => n12957);
   U870 : BUF_X1 port map( A => n4433, Z => n12930);
   U871 : BUF_X1 port map( A => n3060, Z => n13347);
   U872 : BUF_X1 port map( A => n3086, Z => n13293);
   U873 : BUF_X1 port map( A => n3097, Z => n13266);
   U874 : BUF_X1 port map( A => n3138, Z => n13185);
   U875 : BUF_X1 port map( A => n3112, Z => n13239);
   U876 : BUF_X1 port map( A => n3123, Z => n13212);
   U877 : BUF_X1 port map( A => n2926, Z => n13686);
   U878 : BUF_X1 port map( A => n4345, Z => n13116);
   U879 : BUF_X1 port map( A => n4351, Z => n13101);
   U880 : BUF_X1 port map( A => n3061, Z => n13344);
   U881 : BUF_X1 port map( A => n3067, Z => n13329);
   U882 : BUF_X1 port map( A => n4418, Z => n12966);
   U883 : BUF_X1 port map( A => n4334, Z => n13143);
   U884 : BUF_X1 port map( A => n4340, Z => n13128);
   U885 : BUF_X1 port map( A => n4360, Z => n13089);
   U886 : BUF_X1 port map( A => n4366, Z => n13074);
   U887 : BUF_X1 port map( A => n4377, Z => n13047);
   U888 : BUF_X1 port map( A => n4386, Z => n13035);
   U889 : BUF_X1 port map( A => n4397, Z => n13008);
   U890 : BUF_X1 port map( A => n4392, Z => n13020);
   U891 : BUF_X1 port map( A => n4403, Z => n12993);
   U892 : BUF_X1 port map( A => n4423, Z => n12954);
   U893 : BUF_X1 port map( A => n4429, Z => n12939);
   U894 : BUF_X1 port map( A => n3050, Z => n13371);
   U895 : BUF_X1 port map( A => n3056, Z => n13356);
   U896 : BUF_X1 port map( A => n3076, Z => n13317);
   U897 : BUF_X1 port map( A => n3082, Z => n13302);
   U898 : BUF_X1 port map( A => n3093, Z => n13275);
   U899 : BUF_X1 port map( A => n3102, Z => n13263);
   U900 : BUF_X1 port map( A => n3113, Z => n13236);
   U901 : BUF_X1 port map( A => n3108, Z => n13248);
   U902 : BUF_X1 port map( A => n3119, Z => n13221);
   U903 : BUF_X1 port map( A => n4412, Z => n12981);
   U904 : BUF_X1 port map( A => n3128, Z => n13209);
   U905 : BUF_X1 port map( A => n3139, Z => n13182);
   U906 : BUF_X1 port map( A => n3134, Z => n13194);
   U907 : BUF_X1 port map( A => n3145, Z => n13167);
   U908 : BUF_X1 port map( A => n3035, Z => n13392);
   U909 : BUF_X1 port map( A => n3033, Z => n13398);
   U910 : BUF_X1 port map( A => n3026, Z => n13416);
   U911 : BUF_X1 port map( A => n3024, Z => n13422);
   U912 : BUF_X1 port map( A => n2981, Z => n13524);
   U913 : BUF_X1 port map( A => n3020, Z => n13428);
   U914 : BUF_X1 port map( A => n3016, Z => n13440);
   U915 : BUF_X1 port map( A => n3014, Z => n13446);
   U916 : BUF_X1 port map( A => n3011, Z => n13452);
   U917 : BUF_X1 port map( A => n3008, Z => n13458);
   U918 : BUF_X1 port map( A => n3002, Z => n13470);
   U919 : BUF_X1 port map( A => n2998, Z => n13476);
   U920 : BUF_X1 port map( A => n2996, Z => n13482);
   U921 : BUF_X1 port map( A => n2994, Z => n13488);
   U922 : BUF_X1 port map( A => n2992, Z => n13494);
   U923 : BUF_X1 port map( A => n2990, Z => n13500);
   U924 : BUF_X1 port map( A => n2988, Z => n13506);
   U925 : BUF_X1 port map( A => n2979, Z => n13530);
   U926 : BUF_X1 port map( A => n2977, Z => n13536);
   U927 : BUF_X1 port map( A => n2973, Z => n13548);
   U928 : BUF_X1 port map( A => n2971, Z => n13554);
   U929 : BUF_X1 port map( A => n2969, Z => n13560);
   U930 : BUF_X1 port map( A => n2967, Z => n13566);
   U931 : BUF_X1 port map( A => n2959, Z => n13590);
   U932 : BUF_X1 port map( A => n2957, Z => n13596);
   U933 : BUF_X1 port map( A => n2955, Z => n13602);
   U934 : BUF_X1 port map( A => n2953, Z => n13608);
   U935 : BUF_X1 port map( A => n2951, Z => n13614);
   U936 : BUF_X1 port map( A => n2940, Z => n13644);
   U937 : BUF_X1 port map( A => n2938, Z => n13650);
   U938 : BUF_X1 port map( A => n2936, Z => n13656);
   U939 : BUF_X1 port map( A => n2934, Z => n13662);
   U940 : BUF_X1 port map( A => n2932, Z => n13668);
   U941 : BUF_X1 port map( A => n2922, Z => n13698);
   U942 : BUF_X1 port map( A => n2920, Z => n13704);
   U943 : BUF_X1 port map( A => n2918, Z => n13710);
   U944 : BUF_X1 port map( A => n2915, Z => n13716);
   U945 : BUF_X1 port map( A => n2912, Z => n13722);
   U946 : BUF_X1 port map( A => n2900, Z => n13746);
   U947 : BUF_X1 port map( A => n2891, Z => n13764);
   U948 : BUF_X1 port map( A => n2888, Z => n13770);
   U949 : BUF_X1 port map( A => n2885, Z => n13776);
   U950 : BUF_X1 port map( A => n2873, Z => n13800);
   U951 : BUF_X1 port map( A => n3036, Z => n13389);
   U952 : BUF_X1 port map( A => n4346, Z => n13113);
   U953 : BUF_X1 port map( A => n4352, Z => n13098);
   U954 : BUF_X1 port map( A => n3062, Z => n13341);
   U955 : BUF_X1 port map( A => n3068, Z => n13326);
   U956 : BUF_X1 port map( A => n4335, Z => n13140);
   U957 : BUF_X1 port map( A => n4341, Z => n13125);
   U958 : BUF_X1 port map( A => n4372, Z => n13059);
   U959 : BUF_X1 port map( A => n4367, Z => n13071);
   U960 : BUF_X1 port map( A => n4378, Z => n13044);
   U961 : BUF_X1 port map( A => n4387, Z => n13032);
   U962 : BUF_X1 port map( A => n4398, Z => n13005);
   U963 : BUF_X1 port map( A => n4393, Z => n13017);
   U964 : BUF_X1 port map( A => n4424, Z => n12951);
   U965 : BUF_X1 port map( A => n4430, Z => n12936);
   U966 : BUF_X1 port map( A => n3051, Z => n13368);
   U967 : BUF_X1 port map( A => n3057, Z => n13353);
   U968 : BUF_X1 port map( A => n3088, Z => n13287);
   U969 : BUF_X1 port map( A => n3083, Z => n13299);
   U970 : BUF_X1 port map( A => n3094, Z => n13272);
   U971 : BUF_X1 port map( A => n3103, Z => n13260);
   U972 : BUF_X1 port map( A => n3114, Z => n13233);
   U973 : BUF_X1 port map( A => n3109, Z => n13245);
   U974 : BUF_X1 port map( A => n4413, Z => n12978);
   U975 : BUF_X1 port map( A => n3129, Z => n13206);
   U976 : BUF_X1 port map( A => n3140, Z => n13179);
   U977 : BUF_X1 port map( A => n3146, Z => n13164);
   U978 : AND2_X1 port map( A1 => n3031, A2 => n3009, ZN => n2889);
   U979 : BUF_X1 port map( A => n4339, Z => n13131);
   U980 : BUF_X1 port map( A => n4376, Z => n13050);
   U981 : BUF_X1 port map( A => n3133, Z => n13197);
   U982 : BUF_X1 port map( A => n4365, Z => n13077);
   U983 : BUF_X1 port map( A => n4391, Z => n13023);
   U984 : BUF_X1 port map( A => n4402, Z => n12996);
   U985 : BUF_X1 port map( A => n4417, Z => n12969);
   U986 : BUF_X1 port map( A => n4428, Z => n12942);
   U987 : BUF_X1 port map( A => n3055, Z => n13359);
   U988 : BUF_X1 port map( A => n3092, Z => n13278);
   U989 : BUF_X1 port map( A => n3081, Z => n13305);
   U990 : BUF_X1 port map( A => n3107, Z => n13251);
   U991 : BUF_X1 port map( A => n3118, Z => n13224);
   U992 : BUF_X1 port map( A => n3144, Z => n13170);
   U993 : BUF_X1 port map( A => n4349, Z => n13107);
   U994 : BUF_X1 port map( A => n3065, Z => n13335);
   U995 : BUF_X1 port map( A => n4348, Z => n13110);
   U996 : BUF_X1 port map( A => n4337, Z => n13137);
   U997 : BUF_X1 port map( A => n4374, Z => n13056);
   U998 : BUF_X1 port map( A => n4415, Z => n12975);
   U999 : BUF_X1 port map( A => n4426, Z => n12948);
   U1000 : BUF_X1 port map( A => n3053, Z => n13365);
   U1001 : BUF_X1 port map( A => n3090, Z => n13284);
   U1002 : BUF_X1 port map( A => n3131, Z => n13203);
   U1003 : BUF_X1 port map( A => n3142, Z => n13176);
   U1004 : BUF_X1 port map( A => n4363, Z => n13083);
   U1005 : BUF_X1 port map( A => n4389, Z => n13029);
   U1006 : BUF_X1 port map( A => n4400, Z => n13002);
   U1007 : BUF_X1 port map( A => n3064, Z => n13338);
   U1008 : BUF_X1 port map( A => n3079, Z => n13311);
   U1009 : BUF_X1 port map( A => n3105, Z => n13257);
   U1010 : BUF_X1 port map( A => n3116, Z => n13230);
   U1011 : BUF_X1 port map( A => n4375, Z => n13053);
   U1012 : BUF_X1 port map( A => n4416, Z => n12972);
   U1013 : BUF_X1 port map( A => n3080, Z => n13308);
   U1014 : BUF_X1 port map( A => n3091, Z => n13281);
   U1015 : BUF_X1 port map( A => n3132, Z => n13200);
   U1016 : BUF_X1 port map( A => n4364, Z => n13080);
   U1017 : BUF_X1 port map( A => n4390, Z => n13026);
   U1018 : BUF_X1 port map( A => n4401, Z => n12999);
   U1019 : BUF_X1 port map( A => n4427, Z => n12945);
   U1020 : BUF_X1 port map( A => n3106, Z => n13254);
   U1021 : BUF_X1 port map( A => n3117, Z => n13227);
   U1022 : BUF_X1 port map( A => n3143, Z => n13173);
   U1023 : BUF_X1 port map( A => n2961, Z => n13584);
   U1024 : AND2_X1 port map( A1 => n2999, A2 => n3009, ZN => n2901);
   U1025 : NAND2_X1 port map( A1 => n13149, A2 => n13153, ZN => n4324);
   U1026 : NAND2_X1 port map( A1 => n13377, A2 => n13381, ZN => n3040);
   U1027 : NAND2_X1 port map( A1 => n3021, A2 => n2889, ZN => n3037);
   U1028 : NAND2_X1 port map( A1 => n3021, A2 => n2886, ZN => n3034);
   U1029 : NAND2_X1 port map( A1 => n3021, A2 => n2883, ZN => n3032);
   U1030 : NAND2_X1 port map( A1 => n3021, A2 => n2880, ZN => n3029);
   U1031 : NAND2_X1 port map( A1 => n3021, A2 => n2877, ZN => n3027);
   U1032 : NAND2_X1 port map( A1 => n3021, A2 => n2874, ZN => n3025);
   U1033 : NAND2_X1 port map( A1 => n3021, A2 => n2871, ZN => n3023);
   U1034 : NAND2_X1 port map( A1 => n3021, A2 => n2867, ZN => n3019);
   U1035 : AND2_X1 port map( A1 => n5691, A2 => n5664, ZN => n4361);
   U1036 : AND2_X1 port map( A1 => n5690, A2 => n5664, ZN => n4404);
   U1037 : AND2_X1 port map( A1 => n4290, A2 => n4273, ZN => n3077);
   U1038 : AND2_X1 port map( A1 => n4289, A2 => n4273, ZN => n3120);
   U1039 : AND2_X1 port map( A1 => n5659, A2 => n5664, ZN => n4371);
   U1040 : AND2_X1 port map( A1 => n4270, A2 => n4273, ZN => n3087);
   U1041 : AND2_X1 port map( A1 => n5732, A2 => n5664, ZN => n4419);
   U1042 : AND2_X1 port map( A1 => n4310, A2 => n4273, ZN => n3135);
   U1043 : NOR3_X1 port map( A1 => n16062, A2 => ADD_RD2(5), A3 => n16058, ZN 
                           => n5691);
   U1044 : NOR3_X1 port map( A1 => n16061, A2 => ADD_RD1(5), A3 => n16056, ZN 
                           => n4290);
   U1045 : NOR3_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), A3 => n16057, 
                           ZN => n5690);
   U1046 : NOR3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), A3 => n16055, 
                           ZN => n4289);
   U1047 : NOR3_X1 port map( A1 => ADD_RD2(4), A2 => ADD_RD2(5), A3 => n16062, 
                           ZN => n5661);
   U1048 : NOR3_X1 port map( A1 => ADD_RD1(4), A2 => ADD_RD1(5), A3 => n16061, 
                           ZN => n4272);
   U1049 : NOR3_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(5), A3 => n16058, 
                           ZN => n5659);
   U1050 : NOR3_X1 port map( A1 => n16062, A2 => ADD_RD2(4), A3 => n16057, ZN 
                           => n5714);
   U1051 : NOR3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(5), A3 => n16056, 
                           ZN => n4270);
   U1052 : NOR3_X1 port map( A1 => n16061, A2 => ADD_RD1(4), A3 => n16055, ZN 
                           => n4301);
   U1053 : NOR3_X2 port map( A1 => n16068, A2 => n16067, A3 => n16069, ZN => 
                           n5664);
   U1054 : NOR3_X2 port map( A1 => n16065, A2 => n16064, A3 => n16066, ZN => 
                           n4273);
   U1055 : NOR4_X1 port map( A1 => n5746, A2 => n5748, A3 => n5750, A4 => n5752
                           , ZN => n5744);
   U1056 : NOR4_X1 port map( A1 => n4317, A2 => n4318, A3 => n4319, A4 => n4320
                           , ZN => n4316);
   U1057 : AND3_X1 port map( A1 => n16060, A2 => n16059, A3 => ADD_WR(6), ZN =>
                           n3021);
   U1058 : NAND2_X1 port map( A1 => n5679, A2 => n5669, ZN => n4349);
   U1059 : NAND2_X1 port map( A1 => n5679, A2 => n5666, ZN => n4354);
   U1060 : NAND2_X1 port map( A1 => n5679, A2 => n5660, ZN => n4355);
   U1061 : NAND2_X1 port map( A1 => n4282, A2 => n4276, ZN => n3065);
   U1062 : NAND2_X1 port map( A1 => n4282, A2 => n4280, ZN => n3070);
   U1063 : NAND2_X1 port map( A1 => n4282, A2 => n4279, ZN => n3071);
   U1064 : OAI21_X1 port map( B1 => n14021, B2 => n13810, A => n12927, ZN => 
                           n2834);
   U1065 : OAI21_X1 port map( B1 => n2866, B2 => n13386, A => n12922, ZN => 
                           n3036);
   U1066 : OAI21_X1 port map( B1 => n13810, B2 => n13395, A => n12922, ZN => 
                           n3035);
   U1067 : OAI21_X1 port map( B1 => n2866, B2 => n13401, A => n12922, ZN => 
                           n3033);
   U1068 : OAI21_X1 port map( B1 => n13810, B2 => n13407, A => n12922, ZN => 
                           n3030);
   U1069 : OAI21_X1 port map( B1 => n2866, B2 => n13413, A => n12922, ZN => 
                           n3028);
   U1070 : OAI21_X1 port map( B1 => n13810, B2 => n13419, A => n12922, ZN => 
                           n3026);
   U1071 : OAI21_X1 port map( B1 => n2866, B2 => n13425, A => n12922, ZN => 
                           n3024);
   U1072 : OAI21_X1 port map( B1 => n13810, B2 => n13797, A => n12927, ZN => 
                           n2876);
   U1073 : OAI21_X1 port map( B1 => n2866, B2 => n13743, A => n12926, ZN => 
                           n2903);
   U1074 : OAI21_X1 port map( B1 => n13810, B2 => n13791, A => n12927, ZN => 
                           n2879);
   U1075 : OAI21_X1 port map( B1 => n2866, B2 => n13749, A => n12927, ZN => 
                           n2900);
   U1076 : OAI21_X1 port map( B1 => n13810, B2 => n13755, A => n12927, ZN => 
                           n2897);
   U1077 : OAI21_X1 port map( B1 => n2866, B2 => n13761, A => n12927, ZN => 
                           n2894);
   U1078 : OAI21_X1 port map( B1 => n13810, B2 => n13767, A => n12927, ZN => 
                           n2891);
   U1079 : OAI21_X1 port map( B1 => n2866, B2 => n13773, A => n12927, ZN => 
                           n2888);
   U1080 : OAI21_X1 port map( B1 => n13810, B2 => n13779, A => n12927, ZN => 
                           n2885);
   U1081 : OAI21_X1 port map( B1 => n2866, B2 => n13785, A => n12927, ZN => 
                           n2882);
   U1082 : OAI21_X1 port map( B1 => n13810, B2 => n13803, A => n12927, ZN => 
                           n2873);
   U1083 : OAI21_X1 port map( B1 => n2866, B2 => n13809, A => n12927, ZN => 
                           n2870);
   U1084 : OAI21_X1 port map( B1 => n13812, B2 => n13527, A => n12923, ZN => 
                           n2981);
   U1085 : OAI21_X1 port map( B1 => n2866, B2 => n13737, A => n12926, ZN => 
                           n2906);
   U1086 : OAI21_X1 port map( B1 => n13810, B2 => n13683, A => n12926, ZN => 
                           n2928);
   U1087 : OAI21_X1 port map( B1 => n13811, B2 => n13635, A => n12925, ZN => 
                           n2944);
   U1088 : OAI21_X1 port map( B1 => n13811, B2 => n13629, A => n12925, ZN => 
                           n2946);
   U1089 : OAI21_X1 port map( B1 => n13812, B2 => n13575, A => n12924, ZN => 
                           n2965);
   U1090 : OAI21_X1 port map( B1 => n13813, B2 => n13431, A => n12922, ZN => 
                           n3020);
   U1091 : OAI21_X1 port map( B1 => n13813, B2 => n13437, A => n12922, ZN => 
                           n3018);
   U1092 : OAI21_X1 port map( B1 => n13813, B2 => n13443, A => n12922, ZN => 
                           n3016);
   U1093 : OAI21_X1 port map( B1 => n13813, B2 => n13449, A => n12922, ZN => 
                           n3014);
   U1094 : OAI21_X1 port map( B1 => n13813, B2 => n13455, A => n12922, ZN => 
                           n3011);
   U1095 : OAI21_X1 port map( B1 => n13813, B2 => n13461, A => n12923, ZN => 
                           n3008);
   U1096 : OAI21_X1 port map( B1 => n13813, B2 => n13467, A => n12923, ZN => 
                           n3005);
   U1097 : OAI21_X1 port map( B1 => n13813, B2 => n13473, A => n12923, ZN => 
                           n3002);
   U1098 : OAI21_X1 port map( B1 => n13813, B2 => n13479, A => n12923, ZN => 
                           n2998);
   U1099 : OAI21_X1 port map( B1 => n13813, B2 => n13485, A => n12923, ZN => 
                           n2996);
   U1100 : OAI21_X1 port map( B1 => n13813, B2 => n13491, A => n12923, ZN => 
                           n2994);
   U1101 : OAI21_X1 port map( B1 => n13813, B2 => n13497, A => n12923, ZN => 
                           n2992);
   U1102 : OAI21_X1 port map( B1 => n13813, B2 => n13503, A => n12923, ZN => 
                           n2990);
   U1103 : OAI21_X1 port map( B1 => n13812, B2 => n13509, A => n12923, ZN => 
                           n2988);
   U1104 : OAI21_X1 port map( B1 => n13812, B2 => n13515, A => n12923, ZN => 
                           n2986);
   U1105 : OAI21_X1 port map( B1 => n13812, B2 => n13521, A => n12923, ZN => 
                           n2984);
   U1106 : OAI21_X1 port map( B1 => n13812, B2 => n13533, A => n12924, ZN => 
                           n2979);
   U1107 : OAI21_X1 port map( B1 => n13812, B2 => n13539, A => n12924, ZN => 
                           n2977);
   U1108 : OAI21_X1 port map( B1 => n13812, B2 => n13545, A => n12924, ZN => 
                           n2975);
   U1109 : OAI21_X1 port map( B1 => n13812, B2 => n13551, A => n12924, ZN => 
                           n2973);
   U1110 : OAI21_X1 port map( B1 => n13812, B2 => n13557, A => n12924, ZN => 
                           n2971);
   U1111 : OAI21_X1 port map( B1 => n13812, B2 => n13563, A => n12924, ZN => 
                           n2969);
   U1112 : OAI21_X1 port map( B1 => n13812, B2 => n13569, A => n12924, ZN => 
                           n2967);
   U1113 : OAI21_X1 port map( B1 => n13812, B2 => n13581, A => n12924, ZN => 
                           n2963);
   U1114 : OAI21_X1 port map( B1 => n13811, B2 => n13587, A => n12924, ZN => 
                           n2961);
   U1115 : OAI21_X1 port map( B1 => n13811, B2 => n13593, A => n12924, ZN => 
                           n2959);
   U1116 : OAI21_X1 port map( B1 => n13811, B2 => n13599, A => n12924, ZN => 
                           n2957);
   U1117 : OAI21_X1 port map( B1 => n13811, B2 => n13605, A => n12925, ZN => 
                           n2955);
   U1118 : OAI21_X1 port map( B1 => n13811, B2 => n13611, A => n12925, ZN => 
                           n2953);
   U1119 : OAI21_X1 port map( B1 => n13811, B2 => n13617, A => n12925, ZN => 
                           n2951);
   U1120 : OAI21_X1 port map( B1 => n13811, B2 => n13623, A => n12925, ZN => 
                           n2948);
   U1121 : OAI21_X1 port map( B1 => n13811, B2 => n13641, A => n12925, ZN => 
                           n2942);
   U1122 : OAI21_X1 port map( B1 => n13811, B2 => n13647, A => n12925, ZN => 
                           n2940);
   U1123 : OAI21_X1 port map( B1 => n13811, B2 => n13653, A => n12925, ZN => 
                           n2938);
   U1124 : OAI21_X1 port map( B1 => n13811, B2 => n13659, A => n12925, ZN => 
                           n2936);
   U1125 : OAI21_X1 port map( B1 => n2866, B2 => n13665, A => n12925, ZN => 
                           n2934);
   U1126 : OAI21_X1 port map( B1 => n13810, B2 => n13671, A => n12925, ZN => 
                           n2932);
   U1127 : OAI21_X1 port map( B1 => n2866, B2 => n13677, A => n12926, ZN => 
                           n2930);
   U1128 : OAI21_X1 port map( B1 => n13810, B2 => n13689, A => n12926, ZN => 
                           n2926);
   U1129 : OAI21_X1 port map( B1 => n13813, B2 => n13695, A => n12926, ZN => 
                           n2924);
   U1130 : OAI21_X1 port map( B1 => n13812, B2 => n13701, A => n12926, ZN => 
                           n2922);
   U1131 : OAI21_X1 port map( B1 => n13811, B2 => n13707, A => n12926, ZN => 
                           n2920);
   U1132 : OAI21_X1 port map( B1 => n2866, B2 => n13713, A => n12926, ZN => 
                           n2918);
   U1133 : OAI21_X1 port map( B1 => n13810, B2 => n13719, A => n12926, ZN => 
                           n2915);
   U1134 : OAI21_X1 port map( B1 => n13813, B2 => n13725, A => n12926, ZN => 
                           n2912);
   U1135 : OAI21_X1 port map( B1 => n13812, B2 => n13731, A => n12926, ZN => 
                           n2909);
   U1136 : NAND2_X1 port map( A1 => n5669, A2 => ADD_RD2(6), ZN => n4417);
   U1137 : NAND2_X1 port map( A1 => n4276, A2 => ADD_RD1(6), ZN => n3133);
   U1138 : NAND2_X1 port map( A1 => n4274, A2 => ADD_RD1(6), ZN => n3137);
   U1139 : NAND2_X1 port map( A1 => n5710, A2 => n5674, ZN => n4391);
   U1140 : NAND2_X1 port map( A1 => n5710, A2 => n5668, ZN => n4389);
   U1141 : NAND2_X1 port map( A1 => n5710, A2 => n5676, ZN => n4390);
   U1142 : NAND2_X1 port map( A1 => n5710, A2 => n5660, ZN => n4396);
   U1143 : NAND2_X1 port map( A1 => n5710, A2 => n5669, ZN => n4433);
   U1144 : NAND2_X1 port map( A1 => n4299, A2 => n4278, ZN => n3107);
   U1145 : NAND2_X1 port map( A1 => n4299, A2 => n4275, ZN => n3105);
   U1146 : NAND2_X1 port map( A1 => n4299, A2 => n4279, ZN => n3106);
   U1147 : NAND2_X1 port map( A1 => n4299, A2 => n4271, ZN => n3112);
   U1148 : NAND2_X1 port map( A1 => n4299, A2 => n4276, ZN => n3148);
   U1149 : BUF_X1 port map( A => n4325, Z => n13147);
   U1150 : BUF_X1 port map( A => n4325, Z => n13148);
   U1151 : BUF_X1 port map( A => n3041, Z => n13375);
   U1152 : BUF_X1 port map( A => n3041, Z => n13376);
   U1153 : NAND2_X1 port map( A1 => n5690, A2 => n5671, ZN => n4365);
   U1154 : NAND2_X1 port map( A1 => n5690, A2 => n5676, ZN => n4363);
   U1155 : NAND2_X1 port map( A1 => n5690, A2 => n5666, ZN => n4364);
   U1156 : NAND2_X1 port map( A1 => n5691, A2 => n5666, ZN => n4376);
   U1157 : NAND2_X1 port map( A1 => n5691, A2 => n5671, ZN => n4374);
   U1158 : NAND2_X1 port map( A1 => n5691, A2 => n5660, ZN => n4375);
   U1159 : NAND2_X1 port map( A1 => n5691, A2 => n5674, ZN => n4369);
   U1160 : NAND2_X1 port map( A1 => n5691, A2 => n5676, ZN => n4370);
   U1161 : NAND2_X1 port map( A1 => n5690, A2 => n5668, ZN => n4406);
   U1162 : NAND2_X1 port map( A1 => n5690, A2 => n5674, ZN => n4407);
   U1163 : NAND2_X1 port map( A1 => n4289, A2 => n4280, ZN => n3081);
   U1164 : NAND2_X1 port map( A1 => n4289, A2 => n4279, ZN => n3079);
   U1165 : NAND2_X1 port map( A1 => n4289, A2 => n4274, ZN => n3080);
   U1166 : NAND2_X1 port map( A1 => n4290, A2 => n4274, ZN => n3092);
   U1167 : NAND2_X1 port map( A1 => n4290, A2 => n4280, ZN => n3090);
   U1168 : NAND2_X1 port map( A1 => n4290, A2 => n4271, ZN => n3091);
   U1169 : NAND2_X1 port map( A1 => n4290, A2 => n4279, ZN => n3085);
   U1170 : NAND2_X1 port map( A1 => n4290, A2 => n4278, ZN => n3086);
   U1171 : NAND2_X1 port map( A1 => n4289, A2 => n4275, ZN => n3122);
   U1172 : NAND2_X1 port map( A1 => n4289, A2 => n4278, ZN => n3123);
   U1173 : BUF_X1 port map( A => n4325, Z => n13145);
   U1174 : BUF_X1 port map( A => n4325, Z => n13144);
   U1175 : BUF_X1 port map( A => n3041, Z => n13373);
   U1176 : BUF_X1 port map( A => n3041, Z => n13372);
   U1177 : BUF_X1 port map( A => n4322, Z => n13153);
   U1178 : BUF_X1 port map( A => n3038, Z => n13381);
   U1179 : BUF_X1 port map( A => n4322, Z => n13154);
   U1180 : BUF_X1 port map( A => n3038, Z => n13382);
   U1181 : NAND2_X1 port map( A1 => n5659, A2 => n5660, ZN => n4339);
   U1182 : NAND2_X1 port map( A1 => n5659, A2 => n5666, ZN => n4337);
   U1183 : NAND2_X1 port map( A1 => n5661, A2 => n5660, ZN => n4348);
   U1184 : NAND2_X1 port map( A1 => n5661, A2 => n5671, ZN => n4343);
   U1185 : NAND2_X1 port map( A1 => n5661, A2 => n5666, ZN => n4344);
   U1186 : NAND2_X1 port map( A1 => n5659, A2 => n5676, ZN => n4380);
   U1187 : NAND2_X1 port map( A1 => n5659, A2 => n5671, ZN => n4381);
   U1188 : NAND2_X1 port map( A1 => n5714, A2 => n5676, ZN => n4402);
   U1189 : NAND2_X1 port map( A1 => n5714, A2 => n5674, ZN => n4400);
   U1190 : NAND2_X1 port map( A1 => n5714, A2 => n5671, ZN => n4401);
   U1191 : NAND2_X1 port map( A1 => n4270, A2 => n4271, ZN => n3055);
   U1192 : NAND2_X1 port map( A1 => n4270, A2 => n4274, ZN => n3053);
   U1193 : NAND2_X1 port map( A1 => n4272, A2 => n4271, ZN => n3064);
   U1194 : NAND2_X1 port map( A1 => n4272, A2 => n4279, ZN => n3059);
   U1195 : NAND2_X1 port map( A1 => n4272, A2 => n4278, ZN => n3060);
   U1196 : NAND2_X1 port map( A1 => n4270, A2 => n4279, ZN => n3096);
   U1197 : NAND2_X1 port map( A1 => n4270, A2 => n4280, ZN => n3097);
   U1198 : NAND2_X1 port map( A1 => n4301, A2 => n4279, ZN => n3118);
   U1199 : NAND2_X1 port map( A1 => n4301, A2 => n4278, ZN => n3116);
   U1200 : NAND2_X1 port map( A1 => n4301, A2 => n4280, ZN => n3117);
   U1201 : BUF_X1 port map( A => n4325, Z => n13146);
   U1202 : BUF_X1 port map( A => n3041, Z => n13374);
   U1203 : NAND2_X1 port map( A1 => n5732, A2 => n5668, ZN => n4428);
   U1204 : NAND2_X1 port map( A1 => n5732, A2 => n5669, ZN => n4426);
   U1205 : NAND2_X1 port map( A1 => n5732, A2 => n5674, ZN => n4427);
   U1206 : NAND2_X1 port map( A1 => n4310, A2 => n4275, ZN => n3144);
   U1207 : NAND2_X1 port map( A1 => n4310, A2 => n4276, ZN => n3142);
   U1208 : NAND2_X1 port map( A1 => n4310, A2 => n4278, ZN => n3143);
   U1209 : NOR2_X1 port map( A1 => n16071, A2 => n16070, ZN => n3009);
   U1210 : NOR2_X1 port map( A1 => n16072, A2 => ADD_WR(3), ZN => n3031);
   U1211 : AND2_X1 port map( A1 => n3009, A2 => n3022, ZN => n2877);
   U1212 : AND2_X1 port map( A1 => n3006, A2 => n3022, ZN => n2874);
   U1213 : AND2_X1 port map( A1 => n3003, A2 => n3022, ZN => n2871);
   U1214 : AND2_X1 port map( A1 => n3022, A2 => n3000, ZN => n2867);
   U1215 : AND2_X1 port map( A1 => n3031, A2 => n3000, ZN => n2880);
   U1216 : AND2_X1 port map( A1 => n3031, A2 => n3006, ZN => n2886);
   U1217 : AND2_X1 port map( A1 => n3031, A2 => n3003, ZN => n2883);
   U1218 : NAND2_X1 port map( A1 => n5666, A2 => ADD_RD2(6), ZN => n4421);
   U1219 : NAND2_X1 port map( A1 => n5671, A2 => ADD_RD2(6), ZN => n4422);
   U1220 : NAND2_X1 port map( A1 => n4280, A2 => ADD_RD1(6), ZN => n3138);
   U1221 : NAND2_X1 port map( A1 => n5664, A2 => ADD_RD2(6), ZN => n4415);
   U1222 : NAND2_X1 port map( A1 => n4273, A2 => ADD_RD1(6), ZN => n3131);
   U1223 : NAND2_X1 port map( A1 => n5668, A2 => ADD_RD2(6), ZN => n4416);
   U1224 : NAND2_X1 port map( A1 => n4275, A2 => ADD_RD1(6), ZN => n3132);
   U1225 : BUF_X1 port map( A => n4322, Z => n13155);
   U1226 : BUF_X1 port map( A => n3038, Z => n13383);
   U1227 : AND2_X1 port map( A1 => n3012, A2 => n3000, ZN => n2904);
   U1228 : AND2_X1 port map( A1 => n2999, A2 => n3000, ZN => n2892);
   U1229 : AND2_X1 port map( A1 => n3012, A2 => n3003, ZN => n2907);
   U1230 : AND2_X1 port map( A1 => n3012, A2 => n3009, ZN => n2913);
   U1231 : AND2_X1 port map( A1 => n3012, A2 => n3006, ZN => n2910);
   U1232 : AND2_X1 port map( A1 => n2999, A2 => n3006, ZN => n2898);
   U1233 : AND2_X1 port map( A1 => n2999, A2 => n3003, ZN => n2895);
   U1234 : INV_X1 port map( A => ADD_WR(5), ZN => n16059);
   U1235 : INV_X1 port map( A => ADD_RD2(5), ZN => n16057);
   U1236 : INV_X1 port map( A => ADD_RD1(5), ZN => n16055);
   U1237 : INV_X1 port map( A => ADD_WR(4), ZN => n16060);
   U1238 : INV_X1 port map( A => ADD_RD2(4), ZN => n16058);
   U1239 : INV_X1 port map( A => ADD_RD1(4), ZN => n16056);
   U1240 : INV_X1 port map( A => ADD_RD2(3), ZN => n16062);
   U1241 : INV_X1 port map( A => ADD_RD1(3), ZN => n16061);
   U1242 : BUF_X1 port map( A => n13823, Z => n13822);
   U1243 : AND2_X1 port map( A1 => n5679, A2 => n5668, ZN => n4345);
   U1244 : AND2_X1 port map( A1 => n5679, A2 => n5674, ZN => n4346);
   U1245 : AND2_X1 port map( A1 => n5679, A2 => n5671, ZN => n4351);
   U1246 : AND2_X1 port map( A1 => n5679, A2 => n5676, ZN => n4352);
   U1247 : AND2_X1 port map( A1 => n4282, A2 => n4275, ZN => n3061);
   U1248 : AND2_X1 port map( A1 => n4282, A2 => n4278, ZN => n3062);
   U1249 : AND2_X1 port map( A1 => n4282, A2 => n4274, ZN => n3067);
   U1250 : AND2_X1 port map( A1 => n4282, A2 => n4271, ZN => n3068);
   U1251 : AND2_X1 port map( A1 => n5660, A2 => ADD_RD2(6), ZN => n4418);
   U1252 : AND2_X1 port map( A1 => n5710, A2 => n5671, ZN => n4386);
   U1253 : AND2_X1 port map( A1 => n5710, A2 => n5666, ZN => n4387);
   U1254 : AND2_X1 port map( A1 => n4299, A2 => n4280, ZN => n3102);
   U1255 : AND2_X1 port map( A1 => n4299, A2 => n4274, ZN => n3103);
   U1256 : AND2_X1 port map( A1 => n5690, A2 => n5660, ZN => n4360);
   U1257 : AND2_X1 port map( A1 => n5691, A2 => n5668, ZN => n4366);
   U1258 : AND2_X1 port map( A1 => n5691, A2 => n5669, ZN => n4367);
   U1259 : AND2_X1 port map( A1 => n5690, A2 => n5669, ZN => n4403);
   U1260 : AND2_X1 port map( A1 => n4289, A2 => n4271, ZN => n3076);
   U1261 : AND2_X1 port map( A1 => n4290, A2 => n4276, ZN => n3082);
   U1262 : AND2_X1 port map( A1 => n4290, A2 => n4275, ZN => n3083);
   U1263 : AND2_X1 port map( A1 => n4289, A2 => n4276, ZN => n3119);
   U1264 : AND2_X1 port map( A1 => n5661, A2 => n5669, ZN => n4334);
   U1265 : AND2_X1 port map( A1 => n5661, A2 => n5668, ZN => n4335);
   U1266 : AND2_X1 port map( A1 => n5661, A2 => n5676, ZN => n4340);
   U1267 : AND2_X1 port map( A1 => n5661, A2 => n5674, ZN => n4341);
   U1268 : AND2_X1 port map( A1 => n5659, A2 => n5669, ZN => n4372);
   U1269 : AND2_X1 port map( A1 => n5659, A2 => n5674, ZN => n4377);
   U1270 : AND2_X1 port map( A1 => n5659, A2 => n5668, ZN => n4378);
   U1271 : AND2_X1 port map( A1 => n5714, A2 => n5666, ZN => n4397);
   U1272 : AND2_X1 port map( A1 => n5714, A2 => n5660, ZN => n4398);
   U1273 : AND2_X1 port map( A1 => n5714, A2 => n5669, ZN => n4392);
   U1274 : AND2_X1 port map( A1 => n5714, A2 => n5668, ZN => n4393);
   U1275 : AND2_X1 port map( A1 => n4272, A2 => n4276, ZN => n3050);
   U1276 : AND2_X1 port map( A1 => n4272, A2 => n4275, ZN => n3051);
   U1277 : AND2_X1 port map( A1 => n4272, A2 => n4280, ZN => n3056);
   U1278 : AND2_X1 port map( A1 => n4272, A2 => n4274, ZN => n3057);
   U1279 : AND2_X1 port map( A1 => n4270, A2 => n4276, ZN => n3088);
   U1280 : AND2_X1 port map( A1 => n4270, A2 => n4278, ZN => n3093);
   U1281 : AND2_X1 port map( A1 => n4270, A2 => n4275, ZN => n3094);
   U1282 : AND2_X1 port map( A1 => n4301, A2 => n4274, ZN => n3113);
   U1283 : AND2_X1 port map( A1 => n4301, A2 => n4271, ZN => n3114);
   U1284 : AND2_X1 port map( A1 => n4301, A2 => n4276, ZN => n3108);
   U1285 : AND2_X1 port map( A1 => n4301, A2 => n4275, ZN => n3109);
   U1286 : AND2_X1 port map( A1 => n5732, A2 => n5660, ZN => n4429);
   U1287 : AND2_X1 port map( A1 => n5732, A2 => n5676, ZN => n4423);
   U1288 : AND2_X1 port map( A1 => n5732, A2 => n5671, ZN => n4424);
   U1289 : AND2_X1 port map( A1 => n5732, A2 => n5666, ZN => n4430);
   U1290 : AND2_X1 port map( A1 => n4310, A2 => n4279, ZN => n3139);
   U1291 : AND2_X1 port map( A1 => n4310, A2 => n4280, ZN => n3140);
   U1292 : AND2_X1 port map( A1 => n4310, A2 => n4274, ZN => n3145);
   U1293 : AND2_X1 port map( A1 => n4310, A2 => n4271, ZN => n3146);
   U1294 : AND2_X1 port map( A1 => n4279, A2 => ADD_RD1(6), ZN => n3129);
   U1295 : AND2_X1 port map( A1 => n4278, A2 => ADD_RD1(6), ZN => n3128);
   U1296 : AND2_X1 port map( A1 => n5674, A2 => ADD_RD2(6), ZN => n4412);
   U1297 : AND2_X1 port map( A1 => n5676, A2 => ADD_RD2(6), ZN => n4413);
   U1298 : AND2_X1 port map( A1 => n4271, A2 => ADD_RD1(6), ZN => n3134);
   U1299 : BUF_X1 port map( A => n13823, Z => n13821);
   U1300 : BUF_X1 port map( A => n13823, Z => n13820);
   U1301 : BUF_X1 port map( A => n13816, Z => n13819);
   U1302 : BUF_X1 port map( A => n13814, Z => n13818);
   U1303 : BUF_X1 port map( A => n13821, Z => n13817);
   U1304 : BUF_X1 port map( A => n13823, Z => n13816);
   U1305 : BUF_X1 port map( A => n13823, Z => n13815);
   U1306 : BUF_X1 port map( A => n13823, Z => n13814);
   U1307 : AND2_X1 port map( A1 => ADD_WR(3), A2 => n16072, ZN => n2999);
   U1308 : OAI222_X1 port map( A1 => n14175, A2 => n13338, B1 => n14111, B2 => 
                           n13335, C1 => n14143, C2 => n13332, ZN => n3235);
   U1309 : OAI222_X1 port map( A1 => n14560, A2 => n13284, B1 => n14496, B2 => 
                           n13281, C1 => n14528, C2 => n13278, ZN => n3243);
   U1310 : OAI222_X1 port map( A1 => n14174, A2 => n13338, B1 => n14110, B2 => 
                           n13335, C1 => n14142, C2 => n13332, ZN => n3198);
   U1311 : OAI222_X1 port map( A1 => n14559, A2 => n13284, B1 => n14495, B2 => 
                           n13281, C1 => n14527, C2 => n13278, ZN => n3206);
   U1312 : OAI222_X1 port map( A1 => n14173, A2 => n13338, B1 => n14109, B2 => 
                           n13335, C1 => n14141, C2 => n13332, ZN => n3161);
   U1313 : OAI222_X1 port map( A1 => n14558, A2 => n13284, B1 => n14494, B2 => 
                           n13281, C1 => n14526, C2 => n13278, ZN => n3169);
   U1314 : OAI222_X1 port map( A1 => n14172, A2 => n13338, B1 => n14108, B2 => 
                           n13335, C1 => n14140, C2 => n13332, ZN => n3063);
   U1315 : OAI222_X1 port map( A1 => n14557, A2 => n13284, B1 => n14493, B2 => 
                           n13281, C1 => n14525, C2 => n13278, ZN => n3089);
   U1316 : OAI222_X1 port map( A1 => n14178, A2 => n13110, B1 => n14114, B2 => 
                           n13107, C1 => n14146, C2 => n13104, ZN => n4630);
   U1317 : OAI222_X1 port map( A1 => n14563, A2 => n13056, B1 => n14499, B2 => 
                           n13053, C1 => n14531, C2 => n13050, ZN => n4638);
   U1318 : OAI222_X1 port map( A1 => n14177, A2 => n13110, B1 => n14113, B2 => 
                           n13107, C1 => n14145, C2 => n13104, ZN => n4593);
   U1319 : OAI222_X1 port map( A1 => n14562, A2 => n13056, B1 => n14498, B2 => 
                           n13053, C1 => n14530, C2 => n13050, ZN => n4601);
   U1320 : OAI222_X1 port map( A1 => n14176, A2 => n13110, B1 => n14112, B2 => 
                           n13107, C1 => n14144, C2 => n13104, ZN => n4556);
   U1321 : OAI222_X1 port map( A1 => n14561, A2 => n13056, B1 => n14497, B2 => 
                           n13053, C1 => n14529, C2 => n13050, ZN => n4564);
   U1322 : OAI222_X1 port map( A1 => n14175, A2 => n13110, B1 => n14111, B2 => 
                           n13107, C1 => n14143, C2 => n13104, ZN => n4519);
   U1323 : OAI222_X1 port map( A1 => n14560, A2 => n13056, B1 => n14496, B2 => 
                           n13053, C1 => n14528, C2 => n13050, ZN => n4527);
   U1324 : OAI222_X1 port map( A1 => n14174, A2 => n13110, B1 => n14110, B2 => 
                           n13107, C1 => n14142, C2 => n13104, ZN => n4482);
   U1325 : OAI222_X1 port map( A1 => n14559, A2 => n13056, B1 => n14495, B2 => 
                           n13053, C1 => n14527, C2 => n13050, ZN => n4490);
   U1326 : OAI222_X1 port map( A1 => n14173, A2 => n13110, B1 => n14109, B2 => 
                           n13107, C1 => n14141, C2 => n13104, ZN => n4445);
   U1327 : OAI222_X1 port map( A1 => n14558, A2 => n13056, B1 => n14494, B2 => 
                           n13053, C1 => n14526, C2 => n13050, ZN => n4453);
   U1328 : OAI222_X1 port map( A1 => n14172, A2 => n13110, B1 => n14108, B2 => 
                           n13107, C1 => n14140, C2 => n13104, ZN => n4347);
   U1329 : OAI222_X1 port map( A1 => n14557, A2 => n13056, B1 => n14493, B2 => 
                           n13053, C1 => n14525, C2 => n13050, ZN => n4373);
   U1330 : OAI222_X1 port map( A1 => n14179, A2 => n13110, B1 => n14115, B2 => 
                           n13107, C1 => n14147, C2 => n13104, ZN => n4667);
   U1331 : OAI222_X1 port map( A1 => n14564, A2 => n13056, B1 => n14500, B2 => 
                           n13053, C1 => n14532, C2 => n13050, ZN => n4675);
   U1332 : OAI222_X1 port map( A1 => n14179, A2 => n13338, B1 => n14115, B2 => 
                           n13335, C1 => n14147, C2 => n13332, ZN => n3383);
   U1333 : OAI222_X1 port map( A1 => n14564, A2 => n13284, B1 => n14500, B2 => 
                           n13281, C1 => n14532, C2 => n13278, ZN => n3391);
   U1334 : OAI222_X1 port map( A1 => n14178, A2 => n13338, B1 => n14114, B2 => 
                           n13335, C1 => n14146, C2 => n13332, ZN => n3346);
   U1335 : OAI222_X1 port map( A1 => n14563, A2 => n13284, B1 => n14499, B2 => 
                           n13281, C1 => n14531, C2 => n13278, ZN => n3354);
   U1336 : OAI222_X1 port map( A1 => n14177, A2 => n13338, B1 => n14113, B2 => 
                           n13335, C1 => n14145, C2 => n13332, ZN => n3309);
   U1337 : OAI222_X1 port map( A1 => n14562, A2 => n13284, B1 => n14498, B2 => 
                           n13281, C1 => n14530, C2 => n13278, ZN => n3317);
   U1338 : OAI222_X1 port map( A1 => n14176, A2 => n13338, B1 => n14112, B2 => 
                           n13335, C1 => n14144, C2 => n13332, ZN => n3272);
   U1339 : OAI222_X1 port map( A1 => n14561, A2 => n13284, B1 => n14497, B2 => 
                           n13281, C1 => n14529, C2 => n13278, ZN => n3280);
   U1340 : OAI222_X1 port map( A1 => n14203, A2 => n13108, B1 => n14139, B2 => 
                           n13105, C1 => n14171, C2 => n13102, ZN => n5678);
   U1341 : OAI222_X1 port map( A1 => n14588, A2 => n13054, B1 => n14524, B2 => 
                           n13051, C1 => n14556, C2 => n13048, ZN => n5696);
   U1342 : OAI222_X1 port map( A1 => n14202, A2 => n13108, B1 => n14138, B2 => 
                           n13105, C1 => n14170, C2 => n13102, ZN => n5599);
   U1343 : OAI222_X1 port map( A1 => n14587, A2 => n13054, B1 => n14523, B2 => 
                           n13051, C1 => n14555, C2 => n13048, ZN => n5611);
   U1344 : OAI222_X1 port map( A1 => n14201, A2 => n13108, B1 => n14137, B2 => 
                           n13105, C1 => n14169, C2 => n13102, ZN => n5538);
   U1345 : OAI222_X1 port map( A1 => n14586, A2 => n13054, B1 => n14522, B2 => 
                           n13051, C1 => n14554, C2 => n13048, ZN => n5550);
   U1346 : OAI222_X1 port map( A1 => n14200, A2 => n13108, B1 => n14136, B2 => 
                           n13105, C1 => n14168, C2 => n13102, ZN => n5476);
   U1347 : OAI222_X1 port map( A1 => n14585, A2 => n13054, B1 => n14521, B2 => 
                           n13051, C1 => n14553, C2 => n13048, ZN => n5489);
   U1348 : OAI222_X1 port map( A1 => n14199, A2 => n13108, B1 => n14135, B2 => 
                           n13105, C1 => n14167, C2 => n13102, ZN => n5419);
   U1349 : OAI222_X1 port map( A1 => n14584, A2 => n13054, B1 => n14520, B2 => 
                           n13051, C1 => n14552, C2 => n13048, ZN => n5430);
   U1350 : OAI222_X1 port map( A1 => n14198, A2 => n13108, B1 => n14134, B2 => 
                           n13105, C1 => n14166, C2 => n13102, ZN => n5370);
   U1351 : OAI222_X1 port map( A1 => n14583, A2 => n13054, B1 => n14519, B2 => 
                           n13051, C1 => n14551, C2 => n13048, ZN => n5378);
   U1352 : OAI222_X1 port map( A1 => n14197, A2 => n13108, B1 => n14133, B2 => 
                           n13105, C1 => n14165, C2 => n13102, ZN => n5333);
   U1353 : OAI222_X1 port map( A1 => n14582, A2 => n13054, B1 => n14518, B2 => 
                           n13051, C1 => n14550, C2 => n13048, ZN => n5341);
   U1354 : OAI222_X1 port map( A1 => n14196, A2 => n13108, B1 => n14132, B2 => 
                           n13105, C1 => n14164, C2 => n13102, ZN => n5296);
   U1355 : OAI222_X1 port map( A1 => n14581, A2 => n13054, B1 => n14517, B2 => 
                           n13051, C1 => n14549, C2 => n13048, ZN => n5304);
   U1356 : OAI222_X1 port map( A1 => n14195, A2 => n13108, B1 => n14131, B2 => 
                           n13105, C1 => n14163, C2 => n13102, ZN => n5259);
   U1357 : OAI222_X1 port map( A1 => n14580, A2 => n13054, B1 => n14516, B2 => 
                           n13051, C1 => n14548, C2 => n13048, ZN => n5267);
   U1358 : OAI222_X1 port map( A1 => n14194, A2 => n13108, B1 => n14130, B2 => 
                           n13105, C1 => n14162, C2 => n13102, ZN => n5222);
   U1359 : OAI222_X1 port map( A1 => n14579, A2 => n13054, B1 => n14515, B2 => 
                           n13051, C1 => n14547, C2 => n13048, ZN => n5230);
   U1360 : OAI222_X1 port map( A1 => n14193, A2 => n13108, B1 => n14129, B2 => 
                           n13105, C1 => n14161, C2 => n13102, ZN => n5185);
   U1361 : OAI222_X1 port map( A1 => n14578, A2 => n13054, B1 => n14514, B2 => 
                           n13051, C1 => n14546, C2 => n13048, ZN => n5193);
   U1362 : OAI222_X1 port map( A1 => n14192, A2 => n13108, B1 => n14128, B2 => 
                           n13105, C1 => n14160, C2 => n13102, ZN => n5148);
   U1363 : OAI222_X1 port map( A1 => n14577, A2 => n13054, B1 => n14513, B2 => 
                           n13051, C1 => n14545, C2 => n13048, ZN => n5156);
   U1364 : OAI222_X1 port map( A1 => n14191, A2 => n13109, B1 => n14127, B2 => 
                           n13106, C1 => n14159, C2 => n13103, ZN => n5111);
   U1365 : OAI222_X1 port map( A1 => n14576, A2 => n13055, B1 => n14512, B2 => 
                           n13052, C1 => n14544, C2 => n13049, ZN => n5119);
   U1366 : OAI222_X1 port map( A1 => n14190, A2 => n13109, B1 => n14126, B2 => 
                           n13106, C1 => n14158, C2 => n13103, ZN => n5074);
   U1367 : OAI222_X1 port map( A1 => n14575, A2 => n13055, B1 => n14511, B2 => 
                           n13052, C1 => n14543, C2 => n13049, ZN => n5082);
   U1368 : OAI222_X1 port map( A1 => n14189, A2 => n13109, B1 => n14125, B2 => 
                           n13106, C1 => n14157, C2 => n13103, ZN => n5037);
   U1369 : OAI222_X1 port map( A1 => n14574, A2 => n13055, B1 => n14510, B2 => 
                           n13052, C1 => n14542, C2 => n13049, ZN => n5045);
   U1370 : OAI222_X1 port map( A1 => n14188, A2 => n13109, B1 => n14124, B2 => 
                           n13106, C1 => n14156, C2 => n13103, ZN => n5000);
   U1371 : OAI222_X1 port map( A1 => n14573, A2 => n13055, B1 => n14509, B2 => 
                           n13052, C1 => n14541, C2 => n13049, ZN => n5008);
   U1372 : OAI222_X1 port map( A1 => n14187, A2 => n13109, B1 => n14123, B2 => 
                           n13106, C1 => n14155, C2 => n13103, ZN => n4963);
   U1373 : OAI222_X1 port map( A1 => n14572, A2 => n13055, B1 => n14508, B2 => 
                           n13052, C1 => n14540, C2 => n13049, ZN => n4971);
   U1374 : OAI222_X1 port map( A1 => n14186, A2 => n13109, B1 => n14122, B2 => 
                           n13106, C1 => n14154, C2 => n13103, ZN => n4926);
   U1375 : OAI222_X1 port map( A1 => n14571, A2 => n13055, B1 => n14507, B2 => 
                           n13052, C1 => n14539, C2 => n13049, ZN => n4934);
   U1376 : OAI222_X1 port map( A1 => n14185, A2 => n13109, B1 => n14121, B2 => 
                           n13106, C1 => n14153, C2 => n13103, ZN => n4889);
   U1377 : OAI222_X1 port map( A1 => n14570, A2 => n13055, B1 => n14506, B2 => 
                           n13052, C1 => n14538, C2 => n13049, ZN => n4897);
   U1378 : OAI222_X1 port map( A1 => n14184, A2 => n13109, B1 => n14120, B2 => 
                           n13106, C1 => n14152, C2 => n13103, ZN => n4852);
   U1379 : OAI222_X1 port map( A1 => n14569, A2 => n13055, B1 => n14505, B2 => 
                           n13052, C1 => n14537, C2 => n13049, ZN => n4860);
   U1380 : OAI222_X1 port map( A1 => n14183, A2 => n13109, B1 => n14119, B2 => 
                           n13106, C1 => n14151, C2 => n13103, ZN => n4815);
   U1381 : OAI222_X1 port map( A1 => n14568, A2 => n13055, B1 => n14504, B2 => 
                           n13052, C1 => n14536, C2 => n13049, ZN => n4823);
   U1382 : OAI222_X1 port map( A1 => n14182, A2 => n13109, B1 => n14118, B2 => 
                           n13106, C1 => n14150, C2 => n13103, ZN => n4778);
   U1383 : OAI222_X1 port map( A1 => n14567, A2 => n13055, B1 => n14503, B2 => 
                           n13052, C1 => n14535, C2 => n13049, ZN => n4786);
   U1384 : OAI222_X1 port map( A1 => n14181, A2 => n13109, B1 => n14117, B2 => 
                           n13106, C1 => n14149, C2 => n13103, ZN => n4741);
   U1385 : OAI222_X1 port map( A1 => n14566, A2 => n13055, B1 => n14502, B2 => 
                           n13052, C1 => n14534, C2 => n13049, ZN => n4749);
   U1386 : OAI222_X1 port map( A1 => n14180, A2 => n13109, B1 => n14116, B2 => 
                           n13106, C1 => n14148, C2 => n13103, ZN => n4704);
   U1387 : OAI222_X1 port map( A1 => n14565, A2 => n13055, B1 => n14501, B2 => 
                           n13052, C1 => n14533, C2 => n13049, ZN => n4712);
   U1388 : OAI222_X1 port map( A1 => n14203, A2 => n13336, B1 => n14139, B2 => 
                           n13333, C1 => n14171, C2 => n13330, ZN => n4281);
   U1389 : OAI222_X1 port map( A1 => n14588, A2 => n13282, B1 => n14524, B2 => 
                           n13279, C1 => n14556, C2 => n13276, ZN => n4292);
   U1390 : OAI222_X1 port map( A1 => n14202, A2 => n13336, B1 => n14138, B2 => 
                           n13333, C1 => n14170, C2 => n13330, ZN => n4234);
   U1391 : OAI222_X1 port map( A1 => n14587, A2 => n13282, B1 => n14523, B2 => 
                           n13279, C1 => n14555, C2 => n13276, ZN => n4242);
   U1392 : OAI222_X1 port map( A1 => n14201, A2 => n13336, B1 => n14137, B2 => 
                           n13333, C1 => n14169, C2 => n13330, ZN => n4197);
   U1393 : OAI222_X1 port map( A1 => n14586, A2 => n13282, B1 => n14522, B2 => 
                           n13279, C1 => n14554, C2 => n13276, ZN => n4205);
   U1394 : OAI222_X1 port map( A1 => n14200, A2 => n13336, B1 => n14136, B2 => 
                           n13333, C1 => n14168, C2 => n13330, ZN => n4160);
   U1395 : OAI222_X1 port map( A1 => n14585, A2 => n13282, B1 => n14521, B2 => 
                           n13279, C1 => n14553, C2 => n13276, ZN => n4168);
   U1396 : OAI222_X1 port map( A1 => n14199, A2 => n13336, B1 => n14135, B2 => 
                           n13333, C1 => n14167, C2 => n13330, ZN => n4123);
   U1397 : OAI222_X1 port map( A1 => n14584, A2 => n13282, B1 => n14520, B2 => 
                           n13279, C1 => n14552, C2 => n13276, ZN => n4131);
   U1398 : OAI222_X1 port map( A1 => n14198, A2 => n13336, B1 => n14134, B2 => 
                           n13333, C1 => n14166, C2 => n13330, ZN => n4086);
   U1399 : OAI222_X1 port map( A1 => n14583, A2 => n13282, B1 => n14519, B2 => 
                           n13279, C1 => n14551, C2 => n13276, ZN => n4094);
   U1400 : OAI222_X1 port map( A1 => n14197, A2 => n13336, B1 => n14133, B2 => 
                           n13333, C1 => n14165, C2 => n13330, ZN => n4049);
   U1401 : OAI222_X1 port map( A1 => n14582, A2 => n13282, B1 => n14518, B2 => 
                           n13279, C1 => n14550, C2 => n13276, ZN => n4057);
   U1402 : OAI222_X1 port map( A1 => n14196, A2 => n13336, B1 => n14132, B2 => 
                           n13333, C1 => n14164, C2 => n13330, ZN => n4012);
   U1403 : OAI222_X1 port map( A1 => n14581, A2 => n13282, B1 => n14517, B2 => 
                           n13279, C1 => n14549, C2 => n13276, ZN => n4020);
   U1404 : OAI222_X1 port map( A1 => n14195, A2 => n13336, B1 => n14131, B2 => 
                           n13333, C1 => n14163, C2 => n13330, ZN => n3975);
   U1405 : OAI222_X1 port map( A1 => n14580, A2 => n13282, B1 => n14516, B2 => 
                           n13279, C1 => n14548, C2 => n13276, ZN => n3983);
   U1406 : OAI222_X1 port map( A1 => n14194, A2 => n13336, B1 => n14130, B2 => 
                           n13333, C1 => n14162, C2 => n13330, ZN => n3938);
   U1407 : OAI222_X1 port map( A1 => n14579, A2 => n13282, B1 => n14515, B2 => 
                           n13279, C1 => n14547, C2 => n13276, ZN => n3946);
   U1408 : OAI222_X1 port map( A1 => n14193, A2 => n13336, B1 => n14129, B2 => 
                           n13333, C1 => n14161, C2 => n13330, ZN => n3901);
   U1409 : OAI222_X1 port map( A1 => n14578, A2 => n13282, B1 => n14514, B2 => 
                           n13279, C1 => n14546, C2 => n13276, ZN => n3909);
   U1410 : OAI222_X1 port map( A1 => n14192, A2 => n13336, B1 => n14128, B2 => 
                           n13333, C1 => n14160, C2 => n13330, ZN => n3864);
   U1411 : OAI222_X1 port map( A1 => n14577, A2 => n13282, B1 => n14513, B2 => 
                           n13279, C1 => n14545, C2 => n13276, ZN => n3872);
   U1412 : OAI222_X1 port map( A1 => n14191, A2 => n13337, B1 => n14127, B2 => 
                           n13334, C1 => n14159, C2 => n13331, ZN => n3827);
   U1413 : OAI222_X1 port map( A1 => n14576, A2 => n13283, B1 => n14512, B2 => 
                           n13280, C1 => n14544, C2 => n13277, ZN => n3835);
   U1414 : OAI222_X1 port map( A1 => n14190, A2 => n13337, B1 => n14126, B2 => 
                           n13334, C1 => n14158, C2 => n13331, ZN => n3790);
   U1415 : OAI222_X1 port map( A1 => n14575, A2 => n13283, B1 => n14511, B2 => 
                           n13280, C1 => n14543, C2 => n13277, ZN => n3798);
   U1416 : OAI222_X1 port map( A1 => n14189, A2 => n13337, B1 => n14125, B2 => 
                           n13334, C1 => n14157, C2 => n13331, ZN => n3753);
   U1417 : OAI222_X1 port map( A1 => n14574, A2 => n13283, B1 => n14510, B2 => 
                           n13280, C1 => n14542, C2 => n13277, ZN => n3761);
   U1418 : OAI222_X1 port map( A1 => n14188, A2 => n13337, B1 => n14124, B2 => 
                           n13334, C1 => n14156, C2 => n13331, ZN => n3716);
   U1419 : OAI222_X1 port map( A1 => n14573, A2 => n13283, B1 => n14509, B2 => 
                           n13280, C1 => n14541, C2 => n13277, ZN => n3724);
   U1420 : OAI222_X1 port map( A1 => n14187, A2 => n13337, B1 => n14123, B2 => 
                           n13334, C1 => n14155, C2 => n13331, ZN => n3679);
   U1421 : OAI222_X1 port map( A1 => n14572, A2 => n13283, B1 => n14508, B2 => 
                           n13280, C1 => n14540, C2 => n13277, ZN => n3687);
   U1422 : OAI222_X1 port map( A1 => n14186, A2 => n13337, B1 => n14122, B2 => 
                           n13334, C1 => n14154, C2 => n13331, ZN => n3642);
   U1423 : OAI222_X1 port map( A1 => n14571, A2 => n13283, B1 => n14507, B2 => 
                           n13280, C1 => n14539, C2 => n13277, ZN => n3650);
   U1424 : OAI222_X1 port map( A1 => n14185, A2 => n13337, B1 => n14121, B2 => 
                           n13334, C1 => n14153, C2 => n13331, ZN => n3605);
   U1425 : OAI222_X1 port map( A1 => n14570, A2 => n13283, B1 => n14506, B2 => 
                           n13280, C1 => n14538, C2 => n13277, ZN => n3613);
   U1426 : OAI222_X1 port map( A1 => n14184, A2 => n13337, B1 => n14120, B2 => 
                           n13334, C1 => n14152, C2 => n13331, ZN => n3568);
   U1427 : OAI222_X1 port map( A1 => n14569, A2 => n13283, B1 => n14505, B2 => 
                           n13280, C1 => n14537, C2 => n13277, ZN => n3576);
   U1428 : OAI222_X1 port map( A1 => n14183, A2 => n13337, B1 => n14119, B2 => 
                           n13334, C1 => n14151, C2 => n13331, ZN => n3531);
   U1429 : OAI222_X1 port map( A1 => n14568, A2 => n13283, B1 => n14504, B2 => 
                           n13280, C1 => n14536, C2 => n13277, ZN => n3539);
   U1430 : OAI222_X1 port map( A1 => n14182, A2 => n13337, B1 => n14118, B2 => 
                           n13334, C1 => n14150, C2 => n13331, ZN => n3494);
   U1431 : OAI222_X1 port map( A1 => n14567, A2 => n13283, B1 => n14503, B2 => 
                           n13280, C1 => n14535, C2 => n13277, ZN => n3502);
   U1432 : OAI222_X1 port map( A1 => n14181, A2 => n13337, B1 => n14117, B2 => 
                           n13334, C1 => n14149, C2 => n13331, ZN => n3457);
   U1433 : OAI222_X1 port map( A1 => n14566, A2 => n13283, B1 => n14502, B2 => 
                           n13280, C1 => n14534, C2 => n13277, ZN => n3465);
   U1434 : OAI222_X1 port map( A1 => n14180, A2 => n13337, B1 => n14116, B2 => 
                           n13334, C1 => n14148, C2 => n13331, ZN => n3420);
   U1435 : OAI222_X1 port map( A1 => n14565, A2 => n13283, B1 => n14501, B2 => 
                           n13280, C1 => n14533, C2 => n13277, ZN => n3428);
   U1436 : AOI221_X1 port map( B1 => n13141, B2 => n14279, C1 => n13138, C2 => 
                           n15897, A => n5658, ZN => n5656);
   U1437 : OAI222_X1 port map( A1 => n14375, A2 => n13135, B1 => n14311, B2 => 
                           n13132, C1 => n14343, C2 => n13129, ZN => n5658);
   U1438 : AOI221_X1 port map( B1 => n13033, B2 => n15013, C1 => n13030, C2 => 
                           n14981, A => n5708, ZN => n5706);
   U1439 : OAI222_X1 port map( A1 => n15109, A2 => n13027, B1 => n15045, B2 => 
                           n13024, C1 => n15077, C2 => n13021, ZN => n5708);
   U1440 : AOI221_X1 port map( B1 => n13141, B2 => n14278, C1 => n13138, C2 => 
                           n15896, A => n5596, ZN => n5594);
   U1441 : OAI222_X1 port map( A1 => n14374, A2 => n13135, B1 => n14310, B2 => 
                           n13132, C1 => n14342, C2 => n13129, ZN => n5596);
   U1442 : AOI221_X1 port map( B1 => n13033, B2 => n15012, C1 => n13030, C2 => 
                           n15612, A => n5621, ZN => n5620);
   U1443 : OAI222_X1 port map( A1 => n15108, A2 => n13027, B1 => n15044, B2 => 
                           n13024, C1 => n15076, C2 => n13021, ZN => n5621);
   U1444 : AOI221_X1 port map( B1 => n13141, B2 => n14277, C1 => n13138, C2 => 
                           n15895, A => n5534, ZN => n5531);
   U1445 : OAI222_X1 port map( A1 => n14373, A2 => n13135, B1 => n14309, B2 => 
                           n13132, C1 => n14341, C2 => n13129, ZN => n5534);
   U1446 : AOI221_X1 port map( B1 => n13033, B2 => n15011, C1 => n13030, C2 => 
                           n15611, A => n5560, ZN => n5559);
   U1447 : OAI222_X1 port map( A1 => n15107, A2 => n13027, B1 => n15043, B2 => 
                           n13024, C1 => n15075, C2 => n13021, ZN => n5560);
   U1448 : AOI221_X1 port map( B1 => n13141, B2 => n14276, C1 => n13138, C2 => 
                           n15894, A => n5471, ZN => n5470);
   U1449 : OAI222_X1 port map( A1 => n14372, A2 => n13135, B1 => n14308, B2 => 
                           n13132, C1 => n14340, C2 => n13129, ZN => n5471);
   U1450 : AOI221_X1 port map( B1 => n13033, B2 => n15010, C1 => n13030, C2 => 
                           n15610, A => n5499, ZN => n5498);
   U1451 : OAI222_X1 port map( A1 => n15106, A2 => n13027, B1 => n15042, B2 => 
                           n13024, C1 => n15074, C2 => n13021, ZN => n5499);
   U1452 : AOI221_X1 port map( B1 => n13141, B2 => n14275, C1 => n13138, C2 => 
                           n15893, A => n5416, ZN => n5414);
   U1453 : OAI222_X1 port map( A1 => n14371, A2 => n13135, B1 => n14307, B2 => 
                           n13132, C1 => n14339, C2 => n13129, ZN => n5416);
   U1454 : AOI221_X1 port map( B1 => n13033, B2 => n15009, C1 => n13030, C2 => 
                           n15609, A => n5439, ZN => n5438);
   U1455 : OAI222_X1 port map( A1 => n15105, A2 => n13027, B1 => n15041, B2 => 
                           n13024, C1 => n15073, C2 => n13021, ZN => n5439);
   U1456 : AOI221_X1 port map( B1 => n13141, B2 => n14274, C1 => n13138, C2 => 
                           n15892, A => n5368, ZN => n5367);
   U1457 : OAI222_X1 port map( A1 => n14370, A2 => n13135, B1 => n14306, B2 => 
                           n13132, C1 => n14338, C2 => n13129, ZN => n5368);
   U1458 : AOI221_X1 port map( B1 => n13033, B2 => n15008, C1 => n13030, C2 => 
                           n15608, A => n5386, ZN => n5384);
   U1459 : OAI222_X1 port map( A1 => n15104, A2 => n13027, B1 => n15040, B2 => 
                           n13024, C1 => n15072, C2 => n13021, ZN => n5386);
   U1460 : AOI221_X1 port map( B1 => n13141, B2 => n14273, C1 => n13138, C2 => 
                           n15891, A => n5331, ZN => n5330);
   U1461 : OAI222_X1 port map( A1 => n14369, A2 => n13135, B1 => n14305, B2 => 
                           n13132, C1 => n14337, C2 => n13129, ZN => n5331);
   U1462 : AOI221_X1 port map( B1 => n13033, B2 => n15007, C1 => n13030, C2 => 
                           n15607, A => n5347, ZN => n5346);
   U1463 : OAI222_X1 port map( A1 => n15103, A2 => n13027, B1 => n15039, B2 => 
                           n13024, C1 => n15071, C2 => n13021, ZN => n5347);
   U1464 : AOI221_X1 port map( B1 => n13141, B2 => n14272, C1 => n13138, C2 => 
                           n15890, A => n5294, ZN => n5293);
   U1465 : OAI222_X1 port map( A1 => n14368, A2 => n13135, B1 => n14304, B2 => 
                           n13132, C1 => n14336, C2 => n13129, ZN => n5294);
   U1466 : AOI221_X1 port map( B1 => n13033, B2 => n15006, C1 => n13030, C2 => 
                           n15606, A => n5310, ZN => n5309);
   U1467 : OAI222_X1 port map( A1 => n15102, A2 => n13027, B1 => n15038, B2 => 
                           n13024, C1 => n15070, C2 => n13021, ZN => n5310);
   U1468 : AOI221_X1 port map( B1 => n13141, B2 => n14271, C1 => n13138, C2 => 
                           n15889, A => n5257, ZN => n5256);
   U1469 : OAI222_X1 port map( A1 => n14367, A2 => n13135, B1 => n14303, B2 => 
                           n13132, C1 => n14335, C2 => n13129, ZN => n5257);
   U1470 : AOI221_X1 port map( B1 => n13033, B2 => n15005, C1 => n13030, C2 => 
                           n15657, A => n5273, ZN => n5272);
   U1471 : OAI222_X1 port map( A1 => n15101, A2 => n13027, B1 => n15037, B2 => 
                           n13024, C1 => n15069, C2 => n13021, ZN => n5273);
   U1472 : AOI221_X1 port map( B1 => n13141, B2 => n14270, C1 => n13138, C2 => 
                           n15888, A => n5220, ZN => n5219);
   U1473 : OAI222_X1 port map( A1 => n14366, A2 => n13135, B1 => n14302, B2 => 
                           n13132, C1 => n14334, C2 => n13129, ZN => n5220);
   U1474 : AOI221_X1 port map( B1 => n13033, B2 => n15004, C1 => n13030, C2 => 
                           n15656, A => n5236, ZN => n5235);
   U1475 : OAI222_X1 port map( A1 => n15100, A2 => n13027, B1 => n15036, B2 => 
                           n13024, C1 => n15068, C2 => n13021, ZN => n5236);
   U1476 : AOI221_X1 port map( B1 => n13141, B2 => n14269, C1 => n13138, C2 => 
                           n15887, A => n5183, ZN => n5182);
   U1477 : OAI222_X1 port map( A1 => n14365, A2 => n13135, B1 => n14301, B2 => 
                           n13132, C1 => n14333, C2 => n13129, ZN => n5183);
   U1478 : AOI221_X1 port map( B1 => n13033, B2 => n15003, C1 => n13030, C2 => 
                           n15655, A => n5199, ZN => n5198);
   U1479 : OAI222_X1 port map( A1 => n15099, A2 => n13027, B1 => n15035, B2 => 
                           n13024, C1 => n15067, C2 => n13021, ZN => n5199);
   U1480 : AOI221_X1 port map( B1 => n13141, B2 => n14268, C1 => n13138, C2 => 
                           n15886, A => n5146, ZN => n5145);
   U1481 : OAI222_X1 port map( A1 => n14364, A2 => n13135, B1 => n14300, B2 => 
                           n13132, C1 => n14332, C2 => n13129, ZN => n5146);
   U1482 : AOI221_X1 port map( B1 => n13033, B2 => n15002, C1 => n13030, C2 => 
                           n15654, A => n5162, ZN => n5161);
   U1483 : OAI222_X1 port map( A1 => n15098, A2 => n13027, B1 => n15034, B2 => 
                           n13024, C1 => n15066, C2 => n13021, ZN => n5162);
   U1484 : AOI221_X1 port map( B1 => n12980, B2 => n15449, C1 => n12977, C2 => 
                           n15417, A => n5133, ZN => n5132);
   U1485 : OAI222_X1 port map( A1 => n15545, A2 => n12974, B1 => n15481, B2 => 
                           n12971, C1 => n15513, C2 => n12968, ZN => n5133);
   U1486 : AOI221_X1 port map( B1 => n12980, B2 => n15448, C1 => n12977, C2 => 
                           n15416, A => n5096, ZN => n5095);
   U1487 : OAI222_X1 port map( A1 => n15544, A2 => n12974, B1 => n15480, B2 => 
                           n12971, C1 => n15512, C2 => n12968, ZN => n5096);
   U1488 : AOI221_X1 port map( B1 => n12980, B2 => n15447, C1 => n12977, C2 => 
                           n15415, A => n5059, ZN => n5058);
   U1489 : OAI222_X1 port map( A1 => n15543, A2 => n12974, B1 => n15479, B2 => 
                           n12971, C1 => n15511, C2 => n12968, ZN => n5059);
   U1490 : AOI221_X1 port map( B1 => n12980, B2 => n15446, C1 => n12977, C2 => 
                           n15414, A => n5022, ZN => n5021);
   U1491 : OAI222_X1 port map( A1 => n15542, A2 => n12974, B1 => n15478, B2 => 
                           n12971, C1 => n15510, C2 => n12968, ZN => n5022);
   U1492 : AOI221_X1 port map( B1 => n12980, B2 => n15445, C1 => n12977, C2 => 
                           n15413, A => n4985, ZN => n4984);
   U1493 : OAI222_X1 port map( A1 => n15541, A2 => n12974, B1 => n15477, B2 => 
                           n12971, C1 => n15509, C2 => n12968, ZN => n4985);
   U1494 : AOI221_X1 port map( B1 => n12980, B2 => n15444, C1 => n12977, C2 => 
                           n15412, A => n4948, ZN => n4947);
   U1495 : OAI222_X1 port map( A1 => n15540, A2 => n12974, B1 => n15476, B2 => 
                           n12971, C1 => n15508, C2 => n12968, ZN => n4948);
   U1496 : AOI221_X1 port map( B1 => n12980, B2 => n15443, C1 => n12977, C2 => 
                           n15411, A => n4911, ZN => n4910);
   U1497 : OAI222_X1 port map( A1 => n15539, A2 => n12974, B1 => n15475, B2 => 
                           n12971, C1 => n15507, C2 => n12968, ZN => n4911);
   U1498 : AOI221_X1 port map( B1 => n12980, B2 => n15442, C1 => n12977, C2 => 
                           n15410, A => n4874, ZN => n4873);
   U1499 : OAI222_X1 port map( A1 => n15538, A2 => n12974, B1 => n15474, B2 => 
                           n12971, C1 => n15506, C2 => n12968, ZN => n4874);
   U1500 : AOI221_X1 port map( B1 => n13034, B2 => n14993, C1 => n13031, C2 => 
                           n15645, A => n4829, ZN => n4828);
   U1501 : OAI222_X1 port map( A1 => n15089, A2 => n13028, B1 => n15025, B2 => 
                           n13025, C1 => n15057, C2 => n13022, ZN => n4829);
   U1502 : AOI221_X1 port map( B1 => n12980, B2 => n15441, C1 => n12977, C2 => 
                           n15409, A => n4837, ZN => n4836);
   U1503 : OAI222_X1 port map( A1 => n15537, A2 => n12974, B1 => n15473, B2 => 
                           n12971, C1 => n15505, C2 => n12968, ZN => n4837);
   U1504 : AOI221_X1 port map( B1 => n13034, B2 => n14992, C1 => n13031, C2 => 
                           n15644, A => n4792, ZN => n4791);
   U1505 : OAI222_X1 port map( A1 => n15088, A2 => n13028, B1 => n15024, B2 => 
                           n13025, C1 => n15056, C2 => n13022, ZN => n4792);
   U1506 : AOI221_X1 port map( B1 => n12980, B2 => n15440, C1 => n12977, C2 => 
                           n15408, A => n4800, ZN => n4799);
   U1507 : OAI222_X1 port map( A1 => n15536, A2 => n12974, B1 => n15472, B2 => 
                           n12971, C1 => n15504, C2 => n12968, ZN => n4800);
   U1508 : AOI221_X1 port map( B1 => n13034, B2 => n14991, C1 => n13031, C2 => 
                           n15643, A => n4755, ZN => n4754);
   U1509 : OAI222_X1 port map( A1 => n15087, A2 => n13028, B1 => n15023, B2 => 
                           n13025, C1 => n15055, C2 => n13022, ZN => n4755);
   U1510 : AOI221_X1 port map( B1 => n12980, B2 => n15439, C1 => n12977, C2 => 
                           n15407, A => n4763, ZN => n4762);
   U1511 : OAI222_X1 port map( A1 => n15535, A2 => n12974, B1 => n15471, B2 => 
                           n12971, C1 => n15503, C2 => n12968, ZN => n4763);
   U1512 : AOI221_X1 port map( B1 => n13034, B2 => n14990, C1 => n13031, C2 => 
                           n15642, A => n4718, ZN => n4717);
   U1513 : OAI222_X1 port map( A1 => n15086, A2 => n13028, B1 => n15022, B2 => 
                           n13025, C1 => n15054, C2 => n13022, ZN => n4718);
   U1514 : AOI221_X1 port map( B1 => n12980, B2 => n15438, C1 => n12977, C2 => 
                           n15406, A => n4726, ZN => n4725);
   U1515 : OAI222_X1 port map( A1 => n15534, A2 => n12974, B1 => n15470, B2 => 
                           n12971, C1 => n15502, C2 => n12968, ZN => n4726);
   U1516 : AOI221_X1 port map( B1 => n13369, B2 => n14279, C1 => n13366, C2 => 
                           n15897, A => n4269, ZN => n4268);
   U1517 : OAI222_X1 port map( A1 => n14375, A2 => n13363, B1 => n14311, B2 => 
                           n13360, C1 => n14343, C2 => n13357, ZN => n4269);
   U1518 : AOI221_X1 port map( B1 => n13261, B2 => n15013, C1 => n13258, C2 => 
                           n14981, A => n4298, ZN => n4297);
   U1519 : OAI222_X1 port map( A1 => n15109, A2 => n13255, B1 => n15045, B2 => 
                           n13252, C1 => n15077, C2 => n13249, ZN => n4298);
   U1520 : AOI221_X1 port map( B1 => n13369, B2 => n14278, C1 => n13366, C2 => 
                           n15896, A => n4232, ZN => n4231);
   U1521 : OAI222_X1 port map( A1 => n14374, A2 => n13363, B1 => n14310, B2 => 
                           n13360, C1 => n14342, C2 => n13357, ZN => n4232);
   U1522 : AOI221_X1 port map( B1 => n13261, B2 => n15012, C1 => n13258, C2 => 
                           n15612, A => n4248, ZN => n4247);
   U1523 : OAI222_X1 port map( A1 => n15108, A2 => n13255, B1 => n15044, B2 => 
                           n13252, C1 => n15076, C2 => n13249, ZN => n4248);
   U1524 : AOI221_X1 port map( B1 => n13369, B2 => n14277, C1 => n13366, C2 => 
                           n15895, A => n4195, ZN => n4194);
   U1525 : OAI222_X1 port map( A1 => n14373, A2 => n13363, B1 => n14309, B2 => 
                           n13360, C1 => n14341, C2 => n13357, ZN => n4195);
   U1526 : AOI221_X1 port map( B1 => n13261, B2 => n15011, C1 => n13258, C2 => 
                           n15611, A => n4211, ZN => n4210);
   U1527 : OAI222_X1 port map( A1 => n15107, A2 => n13255, B1 => n15043, B2 => 
                           n13252, C1 => n15075, C2 => n13249, ZN => n4211);
   U1528 : AOI221_X1 port map( B1 => n13369, B2 => n14276, C1 => n13366, C2 => 
                           n15894, A => n4158, ZN => n4157);
   U1529 : OAI222_X1 port map( A1 => n14372, A2 => n13363, B1 => n14308, B2 => 
                           n13360, C1 => n14340, C2 => n13357, ZN => n4158);
   U1530 : AOI221_X1 port map( B1 => n13261, B2 => n15010, C1 => n13258, C2 => 
                           n15610, A => n4174, ZN => n4173);
   U1531 : OAI222_X1 port map( A1 => n15106, A2 => n13255, B1 => n15042, B2 => 
                           n13252, C1 => n15074, C2 => n13249, ZN => n4174);
   U1532 : AOI221_X1 port map( B1 => n13369, B2 => n14275, C1 => n13366, C2 => 
                           n15893, A => n4121, ZN => n4120);
   U1533 : OAI222_X1 port map( A1 => n14371, A2 => n13363, B1 => n14307, B2 => 
                           n13360, C1 => n14339, C2 => n13357, ZN => n4121);
   U1534 : AOI221_X1 port map( B1 => n13261, B2 => n15009, C1 => n13258, C2 => 
                           n15609, A => n4137, ZN => n4136);
   U1535 : OAI222_X1 port map( A1 => n15105, A2 => n13255, B1 => n15041, B2 => 
                           n13252, C1 => n15073, C2 => n13249, ZN => n4137);
   U1536 : AOI221_X1 port map( B1 => n13369, B2 => n14274, C1 => n13366, C2 => 
                           n15892, A => n4084, ZN => n4083);
   U1537 : OAI222_X1 port map( A1 => n14370, A2 => n13363, B1 => n14306, B2 => 
                           n13360, C1 => n14338, C2 => n13357, ZN => n4084);
   U1538 : AOI221_X1 port map( B1 => n13261, B2 => n15008, C1 => n13258, C2 => 
                           n15608, A => n4100, ZN => n4099);
   U1539 : OAI222_X1 port map( A1 => n15104, A2 => n13255, B1 => n15040, B2 => 
                           n13252, C1 => n15072, C2 => n13249, ZN => n4100);
   U1540 : AOI221_X1 port map( B1 => n13369, B2 => n14273, C1 => n13366, C2 => 
                           n15891, A => n4047, ZN => n4046);
   U1541 : OAI222_X1 port map( A1 => n14369, A2 => n13363, B1 => n14305, B2 => 
                           n13360, C1 => n14337, C2 => n13357, ZN => n4047);
   U1542 : AOI221_X1 port map( B1 => n13261, B2 => n15007, C1 => n13258, C2 => 
                           n15607, A => n4063, ZN => n4062);
   U1543 : OAI222_X1 port map( A1 => n15103, A2 => n13255, B1 => n15039, B2 => 
                           n13252, C1 => n15071, C2 => n13249, ZN => n4063);
   U1544 : AOI221_X1 port map( B1 => n13369, B2 => n14272, C1 => n13366, C2 => 
                           n15890, A => n4010, ZN => n4009);
   U1545 : OAI222_X1 port map( A1 => n14368, A2 => n13363, B1 => n14304, B2 => 
                           n13360, C1 => n14336, C2 => n13357, ZN => n4010);
   U1546 : AOI221_X1 port map( B1 => n13261, B2 => n15006, C1 => n13258, C2 => 
                           n15606, A => n4026, ZN => n4025);
   U1547 : OAI222_X1 port map( A1 => n15102, A2 => n13255, B1 => n15038, B2 => 
                           n13252, C1 => n15070, C2 => n13249, ZN => n4026);
   U1548 : AOI221_X1 port map( B1 => n13369, B2 => n14271, C1 => n13366, C2 => 
                           n15889, A => n3973, ZN => n3972);
   U1549 : OAI222_X1 port map( A1 => n14367, A2 => n13363, B1 => n14303, B2 => 
                           n13360, C1 => n14335, C2 => n13357, ZN => n3973);
   U1550 : AOI221_X1 port map( B1 => n13261, B2 => n15005, C1 => n13258, C2 => 
                           n15657, A => n3989, ZN => n3988);
   U1551 : OAI222_X1 port map( A1 => n15101, A2 => n13255, B1 => n15037, B2 => 
                           n13252, C1 => n15069, C2 => n13249, ZN => n3989);
   U1552 : AOI221_X1 port map( B1 => n13369, B2 => n14270, C1 => n13366, C2 => 
                           n15888, A => n3936, ZN => n3935);
   U1553 : OAI222_X1 port map( A1 => n14366, A2 => n13363, B1 => n14302, B2 => 
                           n13360, C1 => n14334, C2 => n13357, ZN => n3936);
   U1554 : AOI221_X1 port map( B1 => n13261, B2 => n15004, C1 => n13258, C2 => 
                           n15656, A => n3952, ZN => n3951);
   U1555 : OAI222_X1 port map( A1 => n15100, A2 => n13255, B1 => n15036, B2 => 
                           n13252, C1 => n15068, C2 => n13249, ZN => n3952);
   U1556 : AOI221_X1 port map( B1 => n13369, B2 => n14269, C1 => n13366, C2 => 
                           n15887, A => n3899, ZN => n3898);
   U1557 : OAI222_X1 port map( A1 => n14365, A2 => n13363, B1 => n14301, B2 => 
                           n13360, C1 => n14333, C2 => n13357, ZN => n3899);
   U1558 : AOI221_X1 port map( B1 => n13261, B2 => n15003, C1 => n13258, C2 => 
                           n15655, A => n3915, ZN => n3914);
   U1559 : OAI222_X1 port map( A1 => n15099, A2 => n13255, B1 => n15035, B2 => 
                           n13252, C1 => n15067, C2 => n13249, ZN => n3915);
   U1560 : AOI221_X1 port map( B1 => n13369, B2 => n14268, C1 => n13366, C2 => 
                           n15886, A => n3862, ZN => n3861);
   U1561 : OAI222_X1 port map( A1 => n14364, A2 => n13363, B1 => n14300, B2 => 
                           n13360, C1 => n14332, C2 => n13357, ZN => n3862);
   U1562 : AOI221_X1 port map( B1 => n13261, B2 => n15002, C1 => n13258, C2 => 
                           n15654, A => n3878, ZN => n3877);
   U1563 : OAI222_X1 port map( A1 => n15098, A2 => n13255, B1 => n15034, B2 => 
                           n13252, C1 => n15066, C2 => n13249, ZN => n3878);
   U1564 : AOI221_X1 port map( B1 => n13208, B2 => n15449, C1 => n13205, C2 => 
                           n15417, A => n3849, ZN => n3848);
   U1565 : OAI222_X1 port map( A1 => n15545, A2 => n13202, B1 => n15481, B2 => 
                           n13199, C1 => n15513, C2 => n13196, ZN => n3849);
   U1566 : AOI221_X1 port map( B1 => n13208, B2 => n15448, C1 => n13205, C2 => 
                           n15416, A => n3812, ZN => n3811);
   U1567 : OAI222_X1 port map( A1 => n15544, A2 => n13202, B1 => n15480, B2 => 
                           n13199, C1 => n15512, C2 => n13196, ZN => n3812);
   U1568 : AOI221_X1 port map( B1 => n13208, B2 => n15447, C1 => n13205, C2 => 
                           n15415, A => n3775, ZN => n3774);
   U1569 : OAI222_X1 port map( A1 => n15543, A2 => n13202, B1 => n15479, B2 => 
                           n13199, C1 => n15511, C2 => n13196, ZN => n3775);
   U1570 : AOI221_X1 port map( B1 => n13208, B2 => n15446, C1 => n13205, C2 => 
                           n15414, A => n3738, ZN => n3737);
   U1571 : OAI222_X1 port map( A1 => n15542, A2 => n13202, B1 => n15478, B2 => 
                           n13199, C1 => n15510, C2 => n13196, ZN => n3738);
   U1572 : AOI221_X1 port map( B1 => n13208, B2 => n15445, C1 => n13205, C2 => 
                           n15413, A => n3701, ZN => n3700);
   U1573 : OAI222_X1 port map( A1 => n15541, A2 => n13202, B1 => n15477, B2 => 
                           n13199, C1 => n15509, C2 => n13196, ZN => n3701);
   U1574 : AOI221_X1 port map( B1 => n13208, B2 => n15444, C1 => n13205, C2 => 
                           n15412, A => n3664, ZN => n3663);
   U1575 : OAI222_X1 port map( A1 => n15540, A2 => n13202, B1 => n15476, B2 => 
                           n13199, C1 => n15508, C2 => n13196, ZN => n3664);
   U1576 : AOI221_X1 port map( B1 => n13208, B2 => n15443, C1 => n13205, C2 => 
                           n15411, A => n3627, ZN => n3626);
   U1577 : OAI222_X1 port map( A1 => n15539, A2 => n13202, B1 => n15475, B2 => 
                           n13199, C1 => n15507, C2 => n13196, ZN => n3627);
   U1578 : AOI221_X1 port map( B1 => n13208, B2 => n15442, C1 => n13205, C2 => 
                           n15410, A => n3590, ZN => n3589);
   U1579 : OAI222_X1 port map( A1 => n15538, A2 => n13202, B1 => n15474, B2 => 
                           n13199, C1 => n15506, C2 => n13196, ZN => n3590);
   U1580 : AOI221_X1 port map( B1 => n13262, B2 => n14993, C1 => n13259, C2 => 
                           n15645, A => n3545, ZN => n3544);
   U1581 : OAI222_X1 port map( A1 => n15089, A2 => n13256, B1 => n15025, B2 => 
                           n13253, C1 => n15057, C2 => n13250, ZN => n3545);
   U1582 : AOI221_X1 port map( B1 => n13208, B2 => n15441, C1 => n13205, C2 => 
                           n15409, A => n3553, ZN => n3552);
   U1583 : OAI222_X1 port map( A1 => n15537, A2 => n13202, B1 => n15473, B2 => 
                           n13199, C1 => n15505, C2 => n13196, ZN => n3553);
   U1584 : AOI221_X1 port map( B1 => n13262, B2 => n14992, C1 => n13259, C2 => 
                           n15644, A => n3508, ZN => n3507);
   U1585 : OAI222_X1 port map( A1 => n15088, A2 => n13256, B1 => n15024, B2 => 
                           n13253, C1 => n15056, C2 => n13250, ZN => n3508);
   U1586 : AOI221_X1 port map( B1 => n13208, B2 => n15440, C1 => n13205, C2 => 
                           n15408, A => n3516, ZN => n3515);
   U1587 : OAI222_X1 port map( A1 => n15536, A2 => n13202, B1 => n15472, B2 => 
                           n13199, C1 => n15504, C2 => n13196, ZN => n3516);
   U1588 : AOI221_X1 port map( B1 => n13262, B2 => n14991, C1 => n13259, C2 => 
                           n15643, A => n3471, ZN => n3470);
   U1589 : OAI222_X1 port map( A1 => n15087, A2 => n13256, B1 => n15023, B2 => 
                           n13253, C1 => n15055, C2 => n13250, ZN => n3471);
   U1590 : AOI221_X1 port map( B1 => n13208, B2 => n15439, C1 => n13205, C2 => 
                           n15407, A => n3479, ZN => n3478);
   U1591 : OAI222_X1 port map( A1 => n15535, A2 => n13202, B1 => n15471, B2 => 
                           n13199, C1 => n15503, C2 => n13196, ZN => n3479);
   U1592 : AOI221_X1 port map( B1 => n13262, B2 => n14990, C1 => n13259, C2 => 
                           n15642, A => n3434, ZN => n3433);
   U1593 : OAI222_X1 port map( A1 => n15086, A2 => n13256, B1 => n15022, B2 => 
                           n13253, C1 => n15054, C2 => n13250, ZN => n3434);
   U1594 : AOI221_X1 port map( B1 => n13208, B2 => n15438, C1 => n13205, C2 => 
                           n15406, A => n3442, ZN => n3441);
   U1595 : OAI222_X1 port map( A1 => n15534, A2 => n13202, B1 => n15470, B2 => 
                           n13199, C1 => n15502, C2 => n13196, ZN => n3442);
   U1596 : AOI221_X1 port map( B1 => n13371, B2 => n14251, C1 => n13368, C2 => 
                           n15593, A => n3233, ZN => n3232);
   U1597 : OAI222_X1 port map( A1 => n14347, A2 => n13365, B1 => n14283, B2 => 
                           n13362, C1 => n14315, C2 => n13359, ZN => n3233);
   U1598 : AOI221_X1 port map( B1 => n13317, B2 => n14663, C1 => n13314, C2 => 
                           n15569, A => n3241, ZN => n3240);
   U1599 : OAI222_X1 port map( A1 => n14759, A2 => n13311, B1 => n14695, B2 => 
                           n13308, C1 => n14727, C2 => n13305, ZN => n3241);
   U1600 : AOI221_X1 port map( B1 => n13263, B2 => n14985, C1 => n13260, C2 => 
                           n15637, A => n3249, ZN => n3248);
   U1601 : OAI222_X1 port map( A1 => n15081, A2 => n13257, B1 => n15017, B2 => 
                           n13254, C1 => n15049, C2 => n13251, ZN => n3249);
   U1602 : AOI221_X1 port map( B1 => n13209, B2 => n15433, C1 => n13206, C2 => 
                           n15401, A => n3257, ZN => n3256);
   U1603 : OAI222_X1 port map( A1 => n15529, A2 => n13203, B1 => n15465, B2 => 
                           n13200, C1 => n15497, C2 => n13197, ZN => n3257);
   U1604 : AOI221_X1 port map( B1 => n13371, B2 => n14250, C1 => n13368, C2 => 
                           n15592, A => n3196, ZN => n3195);
   U1605 : OAI222_X1 port map( A1 => n14346, A2 => n13365, B1 => n14282, B2 => 
                           n13362, C1 => n14314, C2 => n13359, ZN => n3196);
   U1606 : AOI221_X1 port map( B1 => n13317, B2 => n14662, C1 => n13314, C2 => 
                           n15568, A => n3204, ZN => n3203);
   U1607 : OAI222_X1 port map( A1 => n14758, A2 => n13311, B1 => n14694, B2 => 
                           n13308, C1 => n14726, C2 => n13305, ZN => n3204);
   U1608 : AOI221_X1 port map( B1 => n13263, B2 => n14984, C1 => n13260, C2 => 
                           n15636, A => n3212, ZN => n3211);
   U1609 : OAI222_X1 port map( A1 => n15080, A2 => n13257, B1 => n15016, B2 => 
                           n13254, C1 => n15048, C2 => n13251, ZN => n3212);
   U1610 : AOI221_X1 port map( B1 => n13209, B2 => n15432, C1 => n13206, C2 => 
                           n15400, A => n3220, ZN => n3219);
   U1611 : OAI222_X1 port map( A1 => n15528, A2 => n13203, B1 => n15464, B2 => 
                           n13200, C1 => n15496, C2 => n13197, ZN => n3220);
   U1612 : AOI221_X1 port map( B1 => n13371, B2 => n14249, C1 => n13368, C2 => 
                           n15591, A => n3159, ZN => n3158);
   U1613 : OAI222_X1 port map( A1 => n14345, A2 => n13365, B1 => n14281, B2 => 
                           n13362, C1 => n14313, C2 => n13359, ZN => n3159);
   U1614 : AOI221_X1 port map( B1 => n13317, B2 => n14661, C1 => n13314, C2 => 
                           n15567, A => n3167, ZN => n3166);
   U1615 : OAI222_X1 port map( A1 => n14757, A2 => n13311, B1 => n14693, B2 => 
                           n13308, C1 => n14725, C2 => n13305, ZN => n3167);
   U1616 : AOI221_X1 port map( B1 => n13263, B2 => n14983, C1 => n13260, C2 => 
                           n15635, A => n3175, ZN => n3174);
   U1617 : OAI222_X1 port map( A1 => n15079, A2 => n13257, B1 => n15015, B2 => 
                           n13254, C1 => n15047, C2 => n13251, ZN => n3175);
   U1618 : AOI221_X1 port map( B1 => n13209, B2 => n15431, C1 => n13206, C2 => 
                           n15399, A => n3183, ZN => n3182);
   U1619 : OAI222_X1 port map( A1 => n15527, A2 => n13203, B1 => n15463, B2 => 
                           n13200, C1 => n15495, C2 => n13197, ZN => n3183);
   U1620 : AOI221_X1 port map( B1 => n13371, B2 => n14248, C1 => n13368, C2 => 
                           n15590, A => n3052, ZN => n3049);
   U1621 : OAI222_X1 port map( A1 => n14344, A2 => n13365, B1 => n14280, B2 => 
                           n13362, C1 => n14312, C2 => n13359, ZN => n3052);
   U1622 : AOI221_X1 port map( B1 => n13317, B2 => n14660, C1 => n13314, C2 => 
                           n15566, A => n3078, ZN => n3075);
   U1623 : OAI222_X1 port map( A1 => n14756, A2 => n13311, B1 => n14692, B2 => 
                           n13308, C1 => n14724, C2 => n13305, ZN => n3078);
   U1624 : AOI221_X1 port map( B1 => n13263, B2 => n14982, C1 => n13260, C2 => 
                           n15634, A => n3104, ZN => n3101);
   U1625 : OAI222_X1 port map( A1 => n15078, A2 => n13257, B1 => n15014, B2 => 
                           n13254, C1 => n15046, C2 => n13251, ZN => n3104);
   U1626 : AOI221_X1 port map( B1 => n13209, B2 => n15430, C1 => n13206, C2 => 
                           n15398, A => n3130, ZN => n3127);
   U1627 : OAI222_X1 port map( A1 => n15526, A2 => n13203, B1 => n15462, B2 => 
                           n13200, C1 => n15494, C2 => n13197, ZN => n3130);
   U1628 : AOI221_X1 port map( B1 => n13143, B2 => n14254, C1 => n13140, C2 => 
                           n15596, A => n4628, ZN => n4627);
   U1629 : OAI222_X1 port map( A1 => n14350, A2 => n13137, B1 => n14286, B2 => 
                           n13134, C1 => n14318, C2 => n13131, ZN => n4628);
   U1630 : AOI221_X1 port map( B1 => n13089, B2 => n14666, C1 => n13086, C2 => 
                           n15572, A => n4636, ZN => n4635);
   U1631 : OAI222_X1 port map( A1 => n14762, A2 => n13083, B1 => n14698, B2 => 
                           n13080, C1 => n14730, C2 => n13077, ZN => n4636);
   U1632 : AOI221_X1 port map( B1 => n13035, B2 => n14988, C1 => n13032, C2 => 
                           n15640, A => n4644, ZN => n4643);
   U1633 : OAI222_X1 port map( A1 => n15084, A2 => n13029, B1 => n15020, B2 => 
                           n13026, C1 => n15052, C2 => n13023, ZN => n4644);
   U1634 : AOI221_X1 port map( B1 => n12981, B2 => n15436, C1 => n12978, C2 => 
                           n15404, A => n4652, ZN => n4651);
   U1635 : OAI222_X1 port map( A1 => n15532, A2 => n12975, B1 => n15468, B2 => 
                           n12972, C1 => n15500, C2 => n12969, ZN => n4652);
   U1636 : AOI221_X1 port map( B1 => n13143, B2 => n14253, C1 => n13140, C2 => 
                           n15595, A => n4591, ZN => n4590);
   U1637 : OAI222_X1 port map( A1 => n14349, A2 => n13137, B1 => n14285, B2 => 
                           n13134, C1 => n14317, C2 => n13131, ZN => n4591);
   U1638 : AOI221_X1 port map( B1 => n13089, B2 => n14665, C1 => n13086, C2 => 
                           n15571, A => n4599, ZN => n4598);
   U1639 : OAI222_X1 port map( A1 => n14761, A2 => n13083, B1 => n14697, B2 => 
                           n13080, C1 => n14729, C2 => n13077, ZN => n4599);
   U1640 : AOI221_X1 port map( B1 => n13035, B2 => n14987, C1 => n13032, C2 => 
                           n15639, A => n4607, ZN => n4606);
   U1641 : OAI222_X1 port map( A1 => n15083, A2 => n13029, B1 => n15019, B2 => 
                           n13026, C1 => n15051, C2 => n13023, ZN => n4607);
   U1642 : AOI221_X1 port map( B1 => n12981, B2 => n15435, C1 => n12978, C2 => 
                           n15403, A => n4615, ZN => n4614);
   U1643 : OAI222_X1 port map( A1 => n15531, A2 => n12975, B1 => n15467, B2 => 
                           n12972, C1 => n15499, C2 => n12969, ZN => n4615);
   U1644 : AOI221_X1 port map( B1 => n13143, B2 => n14252, C1 => n13140, C2 => 
                           n15594, A => n4554, ZN => n4553);
   U1645 : OAI222_X1 port map( A1 => n14348, A2 => n13137, B1 => n14284, B2 => 
                           n13134, C1 => n14316, C2 => n13131, ZN => n4554);
   U1646 : AOI221_X1 port map( B1 => n13089, B2 => n14664, C1 => n13086, C2 => 
                           n15570, A => n4562, ZN => n4561);
   U1647 : OAI222_X1 port map( A1 => n14760, A2 => n13083, B1 => n14696, B2 => 
                           n13080, C1 => n14728, C2 => n13077, ZN => n4562);
   U1648 : AOI221_X1 port map( B1 => n13035, B2 => n14986, C1 => n13032, C2 => 
                           n15638, A => n4570, ZN => n4569);
   U1649 : OAI222_X1 port map( A1 => n15082, A2 => n13029, B1 => n15018, B2 => 
                           n13026, C1 => n15050, C2 => n13023, ZN => n4570);
   U1650 : AOI221_X1 port map( B1 => n12981, B2 => n15434, C1 => n12978, C2 => 
                           n15402, A => n4578, ZN => n4577);
   U1651 : OAI222_X1 port map( A1 => n15530, A2 => n12975, B1 => n15466, B2 => 
                           n12972, C1 => n15498, C2 => n12969, ZN => n4578);
   U1652 : AOI221_X1 port map( B1 => n13143, B2 => n14251, C1 => n13140, C2 => 
                           n15593, A => n4517, ZN => n4516);
   U1653 : OAI222_X1 port map( A1 => n14347, A2 => n13137, B1 => n14283, B2 => 
                           n13134, C1 => n14315, C2 => n13131, ZN => n4517);
   U1654 : AOI221_X1 port map( B1 => n13089, B2 => n14663, C1 => n13086, C2 => 
                           n15569, A => n4525, ZN => n4524);
   U1655 : OAI222_X1 port map( A1 => n14759, A2 => n13083, B1 => n14695, B2 => 
                           n13080, C1 => n14727, C2 => n13077, ZN => n4525);
   U1656 : AOI221_X1 port map( B1 => n13035, B2 => n14985, C1 => n13032, C2 => 
                           n15637, A => n4533, ZN => n4532);
   U1657 : OAI222_X1 port map( A1 => n15081, A2 => n13029, B1 => n15017, B2 => 
                           n13026, C1 => n15049, C2 => n13023, ZN => n4533);
   U1658 : AOI221_X1 port map( B1 => n12981, B2 => n15433, C1 => n12978, C2 => 
                           n15401, A => n4541, ZN => n4540);
   U1659 : OAI222_X1 port map( A1 => n15529, A2 => n12975, B1 => n15465, B2 => 
                           n12972, C1 => n15497, C2 => n12969, ZN => n4541);
   U1660 : AOI221_X1 port map( B1 => n13143, B2 => n14250, C1 => n13140, C2 => 
                           n15592, A => n4480, ZN => n4479);
   U1661 : OAI222_X1 port map( A1 => n14346, A2 => n13137, B1 => n14282, B2 => 
                           n13134, C1 => n14314, C2 => n13131, ZN => n4480);
   U1662 : AOI221_X1 port map( B1 => n13089, B2 => n14662, C1 => n13086, C2 => 
                           n15568, A => n4488, ZN => n4487);
   U1663 : OAI222_X1 port map( A1 => n14758, A2 => n13083, B1 => n14694, B2 => 
                           n13080, C1 => n14726, C2 => n13077, ZN => n4488);
   U1664 : AOI221_X1 port map( B1 => n13035, B2 => n14984, C1 => n13032, C2 => 
                           n15636, A => n4496, ZN => n4495);
   U1665 : OAI222_X1 port map( A1 => n15080, A2 => n13029, B1 => n15016, B2 => 
                           n13026, C1 => n15048, C2 => n13023, ZN => n4496);
   U1666 : AOI221_X1 port map( B1 => n12981, B2 => n15432, C1 => n12978, C2 => 
                           n15400, A => n4504, ZN => n4503);
   U1667 : OAI222_X1 port map( A1 => n15528, A2 => n12975, B1 => n15464, B2 => 
                           n12972, C1 => n15496, C2 => n12969, ZN => n4504);
   U1668 : AOI221_X1 port map( B1 => n13143, B2 => n14249, C1 => n13140, C2 => 
                           n15591, A => n4443, ZN => n4442);
   U1669 : OAI222_X1 port map( A1 => n14345, A2 => n13137, B1 => n14281, B2 => 
                           n13134, C1 => n14313, C2 => n13131, ZN => n4443);
   U1670 : AOI221_X1 port map( B1 => n13089, B2 => n14661, C1 => n13086, C2 => 
                           n15567, A => n4451, ZN => n4450);
   U1671 : OAI222_X1 port map( A1 => n14757, A2 => n13083, B1 => n14693, B2 => 
                           n13080, C1 => n14725, C2 => n13077, ZN => n4451);
   U1672 : AOI221_X1 port map( B1 => n13035, B2 => n14983, C1 => n13032, C2 => 
                           n15635, A => n4459, ZN => n4458);
   U1673 : OAI222_X1 port map( A1 => n15079, A2 => n13029, B1 => n15015, B2 => 
                           n13026, C1 => n15047, C2 => n13023, ZN => n4459);
   U1674 : AOI221_X1 port map( B1 => n12981, B2 => n15431, C1 => n12978, C2 => 
                           n15399, A => n4467, ZN => n4466);
   U1675 : OAI222_X1 port map( A1 => n15527, A2 => n12975, B1 => n15463, B2 => 
                           n12972, C1 => n15495, C2 => n12969, ZN => n4467);
   U1676 : AOI221_X1 port map( B1 => n13143, B2 => n14248, C1 => n13140, C2 => 
                           n15590, A => n4336, ZN => n4333);
   U1677 : OAI222_X1 port map( A1 => n14344, A2 => n13137, B1 => n14280, B2 => 
                           n13134, C1 => n14312, C2 => n13131, ZN => n4336);
   U1678 : AOI221_X1 port map( B1 => n13089, B2 => n14660, C1 => n13086, C2 => 
                           n15566, A => n4362, ZN => n4359);
   U1679 : OAI222_X1 port map( A1 => n14756, A2 => n13083, B1 => n14692, B2 => 
                           n13080, C1 => n14724, C2 => n13077, ZN => n4362);
   U1680 : AOI221_X1 port map( B1 => n13035, B2 => n14982, C1 => n13032, C2 => 
                           n15634, A => n4388, ZN => n4385);
   U1681 : OAI222_X1 port map( A1 => n15078, A2 => n13029, B1 => n15014, B2 => 
                           n13026, C1 => n15046, C2 => n13023, ZN => n4388);
   U1682 : AOI221_X1 port map( B1 => n12981, B2 => n15430, C1 => n12978, C2 => 
                           n15398, A => n4414, ZN => n4411);
   U1683 : OAI222_X1 port map( A1 => n15526, A2 => n12975, B1 => n15462, B2 => 
                           n12972, C1 => n15494, C2 => n12969, ZN => n4414);
   U1684 : AOI221_X1 port map( B1 => n13087, B2 => n14691, C1 => n13084, C2 => 
                           n15765, A => n5689, ZN => n5688);
   U1685 : OAI222_X1 port map( A1 => n14787, A2 => n13081, B1 => n14723, B2 => 
                           n13078, C1 => n14755, C2 => n13075, ZN => n5689);
   U1686 : AOI221_X1 port map( B1 => n12979, B2 => n15461, C1 => n12976, C2 => 
                           n15429, A => n5728, ZN => n5726);
   U1687 : OAI222_X1 port map( A1 => n15557, A2 => n12973, B1 => n15493, B2 => 
                           n12970, C1 => n15525, C2 => n12967, ZN => n5728);
   U1688 : AOI221_X1 port map( B1 => n13087, B2 => n14690, C1 => n13084, C2 => 
                           n15764, A => n5609, ZN => n5608);
   U1689 : OAI222_X1 port map( A1 => n14786, A2 => n13081, B1 => n14722, B2 => 
                           n13078, C1 => n14754, C2 => n13075, ZN => n5609);
   U1690 : AOI221_X1 port map( B1 => n12979, B2 => n15460, C1 => n12976, C2 => 
                           n15428, A => n5636, ZN => n5634);
   U1691 : OAI222_X1 port map( A1 => n15556, A2 => n12973, B1 => n15492, B2 => 
                           n12970, C1 => n15524, C2 => n12967, ZN => n5636);
   U1692 : AOI221_X1 port map( B1 => n13087, B2 => n14689, C1 => n13084, C2 => 
                           n15763, A => n5548, ZN => n5546);
   U1693 : OAI222_X1 port map( A1 => n14785, A2 => n13081, B1 => n14721, B2 => 
                           n13078, C1 => n14753, C2 => n13075, ZN => n5548);
   U1694 : AOI221_X1 port map( B1 => n12979, B2 => n15459, C1 => n12976, C2 => 
                           n15427, A => n5574, ZN => n5571);
   U1695 : OAI222_X1 port map( A1 => n15555, A2 => n12973, B1 => n15491, B2 => 
                           n12970, C1 => n15523, C2 => n12967, ZN => n5574);
   U1696 : AOI221_X1 port map( B1 => n13087, B2 => n14688, C1 => n13084, C2 => 
                           n15762, A => n5486, ZN => n5484);
   U1697 : OAI222_X1 port map( A1 => n14784, A2 => n13081, B1 => n14720, B2 => 
                           n13078, C1 => n14752, C2 => n13075, ZN => n5486);
   U1698 : AOI221_X1 port map( B1 => n12979, B2 => n15458, C1 => n12976, C2 => 
                           n15426, A => n5511, ZN => n5510);
   U1699 : OAI222_X1 port map( A1 => n15554, A2 => n12973, B1 => n15490, B2 => 
                           n12970, C1 => n15522, C2 => n12967, ZN => n5511);
   U1700 : AOI221_X1 port map( B1 => n13087, B2 => n14687, C1 => n13084, C2 => 
                           n15761, A => n5428, ZN => n5426);
   U1701 : OAI222_X1 port map( A1 => n14783, A2 => n13081, B1 => n14719, B2 => 
                           n13078, C1 => n14751, C2 => n13075, ZN => n5428);
   U1702 : AOI221_X1 port map( B1 => n12979, B2 => n15457, C1 => n12976, C2 => 
                           n15425, A => n5450, ZN => n5449);
   U1703 : OAI222_X1 port map( A1 => n15553, A2 => n12973, B1 => n15489, B2 => 
                           n12970, C1 => n15521, C2 => n12967, ZN => n5450);
   U1704 : AOI221_X1 port map( B1 => n13087, B2 => n14686, C1 => n13084, C2 => 
                           n15760, A => n5376, ZN => n5375);
   U1705 : OAI222_X1 port map( A1 => n14782, A2 => n13081, B1 => n14718, B2 => 
                           n13078, C1 => n14750, C2 => n13075, ZN => n5376);
   U1706 : AOI221_X1 port map( B1 => n12979, B2 => n15456, C1 => n12976, C2 => 
                           n15424, A => n5398, ZN => n5396);
   U1707 : OAI222_X1 port map( A1 => n15552, A2 => n12973, B1 => n15488, B2 => 
                           n12970, C1 => n15520, C2 => n12967, ZN => n5398);
   U1708 : AOI221_X1 port map( B1 => n13087, B2 => n14685, C1 => n13084, C2 => 
                           n15759, A => n5339, ZN => n5338);
   U1709 : OAI222_X1 port map( A1 => n14781, A2 => n13081, B1 => n14717, B2 => 
                           n13078, C1 => n14749, C2 => n13075, ZN => n5339);
   U1710 : AOI221_X1 port map( B1 => n12979, B2 => n15455, C1 => n12976, C2 => 
                           n15423, A => n5355, ZN => n5354);
   U1711 : OAI222_X1 port map( A1 => n15551, A2 => n12973, B1 => n15487, B2 => 
                           n12970, C1 => n15519, C2 => n12967, ZN => n5355);
   U1712 : AOI221_X1 port map( B1 => n13087, B2 => n14684, C1 => n13084, C2 => 
                           n15758, A => n5302, ZN => n5301);
   U1713 : OAI222_X1 port map( A1 => n14780, A2 => n13081, B1 => n14716, B2 => 
                           n13078, C1 => n14748, C2 => n13075, ZN => n5302);
   U1714 : AOI221_X1 port map( B1 => n12979, B2 => n15454, C1 => n12976, C2 => 
                           n15422, A => n5318, ZN => n5317);
   U1715 : OAI222_X1 port map( A1 => n15550, A2 => n12973, B1 => n15486, B2 => 
                           n12970, C1 => n15518, C2 => n12967, ZN => n5318);
   U1716 : AOI221_X1 port map( B1 => n13087, B2 => n14683, C1 => n13084, C2 => 
                           n15757, A => n5265, ZN => n5264);
   U1717 : OAI222_X1 port map( A1 => n14779, A2 => n13081, B1 => n14715, B2 => 
                           n13078, C1 => n14747, C2 => n13075, ZN => n5265);
   U1718 : AOI221_X1 port map( B1 => n12979, B2 => n15453, C1 => n12976, C2 => 
                           n15421, A => n5281, ZN => n5280);
   U1719 : OAI222_X1 port map( A1 => n15549, A2 => n12973, B1 => n15485, B2 => 
                           n12970, C1 => n15517, C2 => n12967, ZN => n5281);
   U1720 : AOI221_X1 port map( B1 => n13087, B2 => n14682, C1 => n13084, C2 => 
                           n15756, A => n5228, ZN => n5227);
   U1721 : OAI222_X1 port map( A1 => n14778, A2 => n13081, B1 => n14714, B2 => 
                           n13078, C1 => n14746, C2 => n13075, ZN => n5228);
   U1722 : AOI221_X1 port map( B1 => n12979, B2 => n15452, C1 => n12976, C2 => 
                           n15420, A => n5244, ZN => n5243);
   U1723 : OAI222_X1 port map( A1 => n15548, A2 => n12973, B1 => n15484, B2 => 
                           n12970, C1 => n15516, C2 => n12967, ZN => n5244);
   U1724 : AOI221_X1 port map( B1 => n13087, B2 => n14681, C1 => n13084, C2 => 
                           n15755, A => n5191, ZN => n5190);
   U1725 : OAI222_X1 port map( A1 => n14777, A2 => n13081, B1 => n14713, B2 => 
                           n13078, C1 => n14745, C2 => n13075, ZN => n5191);
   U1726 : AOI221_X1 port map( B1 => n12979, B2 => n15451, C1 => n12976, C2 => 
                           n15419, A => n5207, ZN => n5206);
   U1727 : OAI222_X1 port map( A1 => n15547, A2 => n12973, B1 => n15483, B2 => 
                           n12970, C1 => n15515, C2 => n12967, ZN => n5207);
   U1728 : AOI221_X1 port map( B1 => n13087, B2 => n14680, C1 => n13084, C2 => 
                           n15754, A => n5154, ZN => n5153);
   U1729 : OAI222_X1 port map( A1 => n14776, A2 => n13081, B1 => n14712, B2 => 
                           n13078, C1 => n14744, C2 => n13075, ZN => n5154);
   U1730 : AOI221_X1 port map( B1 => n12979, B2 => n15450, C1 => n12976, C2 => 
                           n15418, A => n5170, ZN => n5169);
   U1731 : OAI222_X1 port map( A1 => n15546, A2 => n12973, B1 => n15482, B2 => 
                           n12970, C1 => n15514, C2 => n12967, ZN => n5170);
   U1732 : AOI221_X1 port map( B1 => n13142, B2 => n14267, C1 => n13139, C2 => 
                           n15885, A => n5109, ZN => n5108);
   U1733 : OAI222_X1 port map( A1 => n14363, A2 => n13136, B1 => n14299, B2 => 
                           n13133, C1 => n14331, C2 => n13130, ZN => n5109);
   U1734 : AOI221_X1 port map( B1 => n13088, B2 => n14679, C1 => n13085, C2 => 
                           n15753, A => n5117, ZN => n5116);
   U1735 : OAI222_X1 port map( A1 => n14775, A2 => n13082, B1 => n14711, B2 => 
                           n13079, C1 => n14743, C2 => n13076, ZN => n5117);
   U1736 : AOI221_X1 port map( B1 => n13034, B2 => n15001, C1 => n13031, C2 => 
                           n15653, A => n5125, ZN => n5124);
   U1737 : OAI222_X1 port map( A1 => n15097, A2 => n13028, B1 => n15033, B2 => 
                           n13025, C1 => n15065, C2 => n13022, ZN => n5125);
   U1738 : AOI221_X1 port map( B1 => n13142, B2 => n14266, C1 => n13139, C2 => 
                           n15884, A => n5072, ZN => n5071);
   U1739 : OAI222_X1 port map( A1 => n14362, A2 => n13136, B1 => n14298, B2 => 
                           n13133, C1 => n14330, C2 => n13130, ZN => n5072);
   U1740 : AOI221_X1 port map( B1 => n13088, B2 => n14678, C1 => n13085, C2 => 
                           n15752, A => n5080, ZN => n5079);
   U1741 : OAI222_X1 port map( A1 => n14774, A2 => n13082, B1 => n14710, B2 => 
                           n13079, C1 => n14742, C2 => n13076, ZN => n5080);
   U1742 : AOI221_X1 port map( B1 => n13034, B2 => n15000, C1 => n13031, C2 => 
                           n15652, A => n5088, ZN => n5087);
   U1743 : OAI222_X1 port map( A1 => n15096, A2 => n13028, B1 => n15032, B2 => 
                           n13025, C1 => n15064, C2 => n13022, ZN => n5088);
   U1744 : AOI221_X1 port map( B1 => n13142, B2 => n14265, C1 => n13139, C2 => 
                           n15883, A => n5035, ZN => n5034);
   U1745 : OAI222_X1 port map( A1 => n14361, A2 => n13136, B1 => n14297, B2 => 
                           n13133, C1 => n14329, C2 => n13130, ZN => n5035);
   U1746 : AOI221_X1 port map( B1 => n13088, B2 => n14677, C1 => n13085, C2 => 
                           n15751, A => n5043, ZN => n5042);
   U1747 : OAI222_X1 port map( A1 => n14773, A2 => n13082, B1 => n14709, B2 => 
                           n13079, C1 => n14741, C2 => n13076, ZN => n5043);
   U1748 : AOI221_X1 port map( B1 => n13034, B2 => n14999, C1 => n13031, C2 => 
                           n15651, A => n5051, ZN => n5050);
   U1749 : OAI222_X1 port map( A1 => n15095, A2 => n13028, B1 => n15031, B2 => 
                           n13025, C1 => n15063, C2 => n13022, ZN => n5051);
   U1750 : AOI221_X1 port map( B1 => n13142, B2 => n14264, C1 => n13139, C2 => 
                           n15882, A => n4998, ZN => n4997);
   U1751 : OAI222_X1 port map( A1 => n14360, A2 => n13136, B1 => n14296, B2 => 
                           n13133, C1 => n14328, C2 => n13130, ZN => n4998);
   U1752 : AOI221_X1 port map( B1 => n13088, B2 => n14676, C1 => n13085, C2 => 
                           n15750, A => n5006, ZN => n5005);
   U1753 : OAI222_X1 port map( A1 => n14772, A2 => n13082, B1 => n14708, B2 => 
                           n13079, C1 => n14740, C2 => n13076, ZN => n5006);
   U1754 : AOI221_X1 port map( B1 => n13034, B2 => n14998, C1 => n13031, C2 => 
                           n15650, A => n5014, ZN => n5013);
   U1755 : OAI222_X1 port map( A1 => n15094, A2 => n13028, B1 => n15030, B2 => 
                           n13025, C1 => n15062, C2 => n13022, ZN => n5014);
   U1756 : AOI221_X1 port map( B1 => n13142, B2 => n14263, C1 => n13139, C2 => 
                           n15881, A => n4961, ZN => n4960);
   U1757 : OAI222_X1 port map( A1 => n14359, A2 => n13136, B1 => n14295, B2 => 
                           n13133, C1 => n14327, C2 => n13130, ZN => n4961);
   U1758 : AOI221_X1 port map( B1 => n13088, B2 => n14675, C1 => n13085, C2 => 
                           n15749, A => n4969, ZN => n4968);
   U1759 : OAI222_X1 port map( A1 => n14771, A2 => n13082, B1 => n14707, B2 => 
                           n13079, C1 => n14739, C2 => n13076, ZN => n4969);
   U1760 : AOI221_X1 port map( B1 => n13034, B2 => n14997, C1 => n13031, C2 => 
                           n15649, A => n4977, ZN => n4976);
   U1761 : OAI222_X1 port map( A1 => n15093, A2 => n13028, B1 => n15029, B2 => 
                           n13025, C1 => n15061, C2 => n13022, ZN => n4977);
   U1762 : AOI221_X1 port map( B1 => n13142, B2 => n14262, C1 => n13139, C2 => 
                           n15880, A => n4924, ZN => n4923);
   U1763 : OAI222_X1 port map( A1 => n14358, A2 => n13136, B1 => n14294, B2 => 
                           n13133, C1 => n14326, C2 => n13130, ZN => n4924);
   U1764 : AOI221_X1 port map( B1 => n13088, B2 => n14674, C1 => n13085, C2 => 
                           n15748, A => n4932, ZN => n4931);
   U1765 : OAI222_X1 port map( A1 => n14770, A2 => n13082, B1 => n14706, B2 => 
                           n13079, C1 => n14738, C2 => n13076, ZN => n4932);
   U1766 : AOI221_X1 port map( B1 => n13034, B2 => n14996, C1 => n13031, C2 => 
                           n15648, A => n4940, ZN => n4939);
   U1767 : OAI222_X1 port map( A1 => n15092, A2 => n13028, B1 => n15028, B2 => 
                           n13025, C1 => n15060, C2 => n13022, ZN => n4940);
   U1768 : AOI221_X1 port map( B1 => n13142, B2 => n14261, C1 => n13139, C2 => 
                           n15879, A => n4887, ZN => n4886);
   U1769 : OAI222_X1 port map( A1 => n14357, A2 => n13136, B1 => n14293, B2 => 
                           n13133, C1 => n14325, C2 => n13130, ZN => n4887);
   U1770 : AOI221_X1 port map( B1 => n13088, B2 => n14673, C1 => n13085, C2 => 
                           n15747, A => n4895, ZN => n4894);
   U1771 : OAI222_X1 port map( A1 => n14769, A2 => n13082, B1 => n14705, B2 => 
                           n13079, C1 => n14737, C2 => n13076, ZN => n4895);
   U1772 : AOI221_X1 port map( B1 => n13034, B2 => n14995, C1 => n13031, C2 => 
                           n15647, A => n4903, ZN => n4902);
   U1773 : OAI222_X1 port map( A1 => n15091, A2 => n13028, B1 => n15027, B2 => 
                           n13025, C1 => n15059, C2 => n13022, ZN => n4903);
   U1774 : AOI221_X1 port map( B1 => n13142, B2 => n14260, C1 => n13139, C2 => 
                           n15878, A => n4850, ZN => n4849);
   U1775 : OAI222_X1 port map( A1 => n14356, A2 => n13136, B1 => n14292, B2 => 
                           n13133, C1 => n14324, C2 => n13130, ZN => n4850);
   U1776 : AOI221_X1 port map( B1 => n13088, B2 => n14672, C1 => n13085, C2 => 
                           n15746, A => n4858, ZN => n4857);
   U1777 : OAI222_X1 port map( A1 => n14768, A2 => n13082, B1 => n14704, B2 => 
                           n13079, C1 => n14736, C2 => n13076, ZN => n4858);
   U1778 : AOI221_X1 port map( B1 => n13034, B2 => n14994, C1 => n13031, C2 => 
                           n15646, A => n4866, ZN => n4865);
   U1779 : OAI222_X1 port map( A1 => n15090, A2 => n13028, B1 => n15026, B2 => 
                           n13025, C1 => n15058, C2 => n13022, ZN => n4866);
   U1780 : AOI221_X1 port map( B1 => n13142, B2 => n14259, C1 => n13139, C2 => 
                           n15877, A => n4813, ZN => n4812);
   U1781 : OAI222_X1 port map( A1 => n14355, A2 => n13136, B1 => n14291, B2 => 
                           n13133, C1 => n14323, C2 => n13130, ZN => n4813);
   U1782 : AOI221_X1 port map( B1 => n13088, B2 => n14671, C1 => n13085, C2 => 
                           n15745, A => n4821, ZN => n4820);
   U1783 : OAI222_X1 port map( A1 => n14767, A2 => n13082, B1 => n14703, B2 => 
                           n13079, C1 => n14735, C2 => n13076, ZN => n4821);
   U1784 : AOI221_X1 port map( B1 => n13142, B2 => n14258, C1 => n13139, C2 => 
                           n15876, A => n4776, ZN => n4775);
   U1785 : OAI222_X1 port map( A1 => n14354, A2 => n13136, B1 => n14290, B2 => 
                           n13133, C1 => n14322, C2 => n13130, ZN => n4776);
   U1786 : AOI221_X1 port map( B1 => n13088, B2 => n14670, C1 => n13085, C2 => 
                           n15744, A => n4784, ZN => n4783);
   U1787 : OAI222_X1 port map( A1 => n14766, A2 => n13082, B1 => n14702, B2 => 
                           n13079, C1 => n14734, C2 => n13076, ZN => n4784);
   U1788 : AOI221_X1 port map( B1 => n13142, B2 => n14257, C1 => n13139, C2 => 
                           n15875, A => n4739, ZN => n4738);
   U1789 : OAI222_X1 port map( A1 => n14353, A2 => n13136, B1 => n14289, B2 => 
                           n13133, C1 => n14321, C2 => n13130, ZN => n4739);
   U1790 : AOI221_X1 port map( B1 => n13088, B2 => n14669, C1 => n13085, C2 => 
                           n15743, A => n4747, ZN => n4746);
   U1791 : OAI222_X1 port map( A1 => n14765, A2 => n13082, B1 => n14701, B2 => 
                           n13079, C1 => n14733, C2 => n13076, ZN => n4747);
   U1792 : AOI221_X1 port map( B1 => n13142, B2 => n14256, C1 => n13139, C2 => 
                           n15874, A => n4702, ZN => n4701);
   U1793 : OAI222_X1 port map( A1 => n14352, A2 => n13136, B1 => n14288, B2 => 
                           n13133, C1 => n14320, C2 => n13130, ZN => n4702);
   U1794 : AOI221_X1 port map( B1 => n13088, B2 => n14668, C1 => n13085, C2 => 
                           n15742, A => n4710, ZN => n4709);
   U1795 : OAI222_X1 port map( A1 => n14764, A2 => n13082, B1 => n14700, B2 => 
                           n13079, C1 => n14732, C2 => n13076, ZN => n4710);
   U1796 : AOI221_X1 port map( B1 => n13143, B2 => n14255, C1 => n13140, C2 => 
                           n15597, A => n4665, ZN => n4664);
   U1797 : OAI222_X1 port map( A1 => n14351, A2 => n13137, B1 => n14287, B2 => 
                           n13134, C1 => n14319, C2 => n13131, ZN => n4665);
   U1798 : AOI221_X1 port map( B1 => n13089, B2 => n14667, C1 => n13086, C2 => 
                           n15573, A => n4673, ZN => n4672);
   U1799 : OAI222_X1 port map( A1 => n14763, A2 => n13083, B1 => n14699, B2 => 
                           n13080, C1 => n14731, C2 => n13077, ZN => n4673);
   U1800 : AOI221_X1 port map( B1 => n13035, B2 => n14989, C1 => n13032, C2 => 
                           n15641, A => n4681, ZN => n4680);
   U1801 : OAI222_X1 port map( A1 => n15085, A2 => n13029, B1 => n15021, B2 => 
                           n13026, C1 => n15053, C2 => n13023, ZN => n4681);
   U1802 : AOI221_X1 port map( B1 => n12981, B2 => n15437, C1 => n12978, C2 => 
                           n15405, A => n4689, ZN => n4688);
   U1803 : OAI222_X1 port map( A1 => n15533, A2 => n12975, B1 => n15469, B2 => 
                           n12972, C1 => n15501, C2 => n12969, ZN => n4689);
   U1804 : AOI221_X1 port map( B1 => n13315, B2 => n14691, C1 => n13312, C2 => 
                           n15765, A => n4288, ZN => n4287);
   U1805 : OAI222_X1 port map( A1 => n14787, A2 => n13309, B1 => n14723, B2 => 
                           n13306, C1 => n14755, C2 => n13303, ZN => n4288);
   U1806 : AOI221_X1 port map( B1 => n13207, B2 => n15461, C1 => n13204, C2 => 
                           n15429, A => n4308, ZN => n4307);
   U1807 : OAI222_X1 port map( A1 => n15557, A2 => n13201, B1 => n15493, B2 => 
                           n13198, C1 => n15525, C2 => n13195, ZN => n4308);
   U1808 : AOI221_X1 port map( B1 => n13315, B2 => n14690, C1 => n13312, C2 => 
                           n15764, A => n4240, ZN => n4239);
   U1809 : OAI222_X1 port map( A1 => n14786, A2 => n13309, B1 => n14722, B2 => 
                           n13306, C1 => n14754, C2 => n13303, ZN => n4240);
   U1810 : AOI221_X1 port map( B1 => n13207, B2 => n15460, C1 => n13204, C2 => 
                           n15428, A => n4256, ZN => n4255);
   U1811 : OAI222_X1 port map( A1 => n15556, A2 => n13201, B1 => n15492, B2 => 
                           n13198, C1 => n15524, C2 => n13195, ZN => n4256);
   U1812 : AOI221_X1 port map( B1 => n13315, B2 => n14689, C1 => n13312, C2 => 
                           n15763, A => n4203, ZN => n4202);
   U1813 : OAI222_X1 port map( A1 => n14785, A2 => n13309, B1 => n14721, B2 => 
                           n13306, C1 => n14753, C2 => n13303, ZN => n4203);
   U1814 : AOI221_X1 port map( B1 => n13207, B2 => n15459, C1 => n13204, C2 => 
                           n15427, A => n4219, ZN => n4218);
   U1815 : OAI222_X1 port map( A1 => n15555, A2 => n13201, B1 => n15491, B2 => 
                           n13198, C1 => n15523, C2 => n13195, ZN => n4219);
   U1816 : AOI221_X1 port map( B1 => n13315, B2 => n14688, C1 => n13312, C2 => 
                           n15762, A => n4166, ZN => n4165);
   U1817 : OAI222_X1 port map( A1 => n14784, A2 => n13309, B1 => n14720, B2 => 
                           n13306, C1 => n14752, C2 => n13303, ZN => n4166);
   U1818 : AOI221_X1 port map( B1 => n13207, B2 => n15458, C1 => n13204, C2 => 
                           n15426, A => n4182, ZN => n4181);
   U1819 : OAI222_X1 port map( A1 => n15554, A2 => n13201, B1 => n15490, B2 => 
                           n13198, C1 => n15522, C2 => n13195, ZN => n4182);
   U1820 : AOI221_X1 port map( B1 => n13315, B2 => n14687, C1 => n13312, C2 => 
                           n15761, A => n4129, ZN => n4128);
   U1821 : OAI222_X1 port map( A1 => n14783, A2 => n13309, B1 => n14719, B2 => 
                           n13306, C1 => n14751, C2 => n13303, ZN => n4129);
   U1822 : AOI221_X1 port map( B1 => n13207, B2 => n15457, C1 => n13204, C2 => 
                           n15425, A => n4145, ZN => n4144);
   U1823 : OAI222_X1 port map( A1 => n15553, A2 => n13201, B1 => n15489, B2 => 
                           n13198, C1 => n15521, C2 => n13195, ZN => n4145);
   U1824 : AOI221_X1 port map( B1 => n13315, B2 => n14686, C1 => n13312, C2 => 
                           n15760, A => n4092, ZN => n4091);
   U1825 : OAI222_X1 port map( A1 => n14782, A2 => n13309, B1 => n14718, B2 => 
                           n13306, C1 => n14750, C2 => n13303, ZN => n4092);
   U1826 : AOI221_X1 port map( B1 => n13207, B2 => n15456, C1 => n13204, C2 => 
                           n15424, A => n4108, ZN => n4107);
   U1827 : OAI222_X1 port map( A1 => n15552, A2 => n13201, B1 => n15488, B2 => 
                           n13198, C1 => n15520, C2 => n13195, ZN => n4108);
   U1828 : AOI221_X1 port map( B1 => n13315, B2 => n14685, C1 => n13312, C2 => 
                           n15759, A => n4055, ZN => n4054);
   U1829 : OAI222_X1 port map( A1 => n14781, A2 => n13309, B1 => n14717, B2 => 
                           n13306, C1 => n14749, C2 => n13303, ZN => n4055);
   U1830 : AOI221_X1 port map( B1 => n13207, B2 => n15455, C1 => n13204, C2 => 
                           n15423, A => n4071, ZN => n4070);
   U1831 : OAI222_X1 port map( A1 => n15551, A2 => n13201, B1 => n15487, B2 => 
                           n13198, C1 => n15519, C2 => n13195, ZN => n4071);
   U1832 : AOI221_X1 port map( B1 => n13315, B2 => n14684, C1 => n13312, C2 => 
                           n15758, A => n4018, ZN => n4017);
   U1833 : OAI222_X1 port map( A1 => n14780, A2 => n13309, B1 => n14716, B2 => 
                           n13306, C1 => n14748, C2 => n13303, ZN => n4018);
   U1834 : AOI221_X1 port map( B1 => n13207, B2 => n15454, C1 => n13204, C2 => 
                           n15422, A => n4034, ZN => n4033);
   U1835 : OAI222_X1 port map( A1 => n15550, A2 => n13201, B1 => n15486, B2 => 
                           n13198, C1 => n15518, C2 => n13195, ZN => n4034);
   U1836 : AOI221_X1 port map( B1 => n13315, B2 => n14683, C1 => n13312, C2 => 
                           n15757, A => n3981, ZN => n3980);
   U1837 : OAI222_X1 port map( A1 => n14779, A2 => n13309, B1 => n14715, B2 => 
                           n13306, C1 => n14747, C2 => n13303, ZN => n3981);
   U1838 : AOI221_X1 port map( B1 => n13207, B2 => n15453, C1 => n13204, C2 => 
                           n15421, A => n3997, ZN => n3996);
   U1839 : OAI222_X1 port map( A1 => n15549, A2 => n13201, B1 => n15485, B2 => 
                           n13198, C1 => n15517, C2 => n13195, ZN => n3997);
   U1840 : AOI221_X1 port map( B1 => n13315, B2 => n14682, C1 => n13312, C2 => 
                           n15756, A => n3944, ZN => n3943);
   U1841 : OAI222_X1 port map( A1 => n14778, A2 => n13309, B1 => n14714, B2 => 
                           n13306, C1 => n14746, C2 => n13303, ZN => n3944);
   U1842 : AOI221_X1 port map( B1 => n13207, B2 => n15452, C1 => n13204, C2 => 
                           n15420, A => n3960, ZN => n3959);
   U1843 : OAI222_X1 port map( A1 => n15548, A2 => n13201, B1 => n15484, B2 => 
                           n13198, C1 => n15516, C2 => n13195, ZN => n3960);
   U1844 : AOI221_X1 port map( B1 => n13315, B2 => n14681, C1 => n13312, C2 => 
                           n15755, A => n3907, ZN => n3906);
   U1845 : OAI222_X1 port map( A1 => n14777, A2 => n13309, B1 => n14713, B2 => 
                           n13306, C1 => n14745, C2 => n13303, ZN => n3907);
   U1846 : AOI221_X1 port map( B1 => n13207, B2 => n15451, C1 => n13204, C2 => 
                           n15419, A => n3923, ZN => n3922);
   U1847 : OAI222_X1 port map( A1 => n15547, A2 => n13201, B1 => n15483, B2 => 
                           n13198, C1 => n15515, C2 => n13195, ZN => n3923);
   U1848 : AOI221_X1 port map( B1 => n13315, B2 => n14680, C1 => n13312, C2 => 
                           n15754, A => n3870, ZN => n3869);
   U1849 : OAI222_X1 port map( A1 => n14776, A2 => n13309, B1 => n14712, B2 => 
                           n13306, C1 => n14744, C2 => n13303, ZN => n3870);
   U1850 : AOI221_X1 port map( B1 => n13207, B2 => n15450, C1 => n13204, C2 => 
                           n15418, A => n3886, ZN => n3885);
   U1851 : OAI222_X1 port map( A1 => n15546, A2 => n13201, B1 => n15482, B2 => 
                           n13198, C1 => n15514, C2 => n13195, ZN => n3886);
   U1852 : AOI221_X1 port map( B1 => n13370, B2 => n14267, C1 => n13367, C2 => 
                           n15885, A => n3825, ZN => n3824);
   U1853 : OAI222_X1 port map( A1 => n14363, A2 => n13364, B1 => n14299, B2 => 
                           n13361, C1 => n14331, C2 => n13358, ZN => n3825);
   U1854 : AOI221_X1 port map( B1 => n13316, B2 => n14679, C1 => n13313, C2 => 
                           n15753, A => n3833, ZN => n3832);
   U1855 : OAI222_X1 port map( A1 => n14775, A2 => n13310, B1 => n14711, B2 => 
                           n13307, C1 => n14743, C2 => n13304, ZN => n3833);
   U1856 : AOI221_X1 port map( B1 => n13262, B2 => n15001, C1 => n13259, C2 => 
                           n15653, A => n3841, ZN => n3840);
   U1857 : OAI222_X1 port map( A1 => n15097, A2 => n13256, B1 => n15033, B2 => 
                           n13253, C1 => n15065, C2 => n13250, ZN => n3841);
   U1858 : AOI221_X1 port map( B1 => n13370, B2 => n14266, C1 => n13367, C2 => 
                           n15884, A => n3788, ZN => n3787);
   U1859 : OAI222_X1 port map( A1 => n14362, A2 => n13364, B1 => n14298, B2 => 
                           n13361, C1 => n14330, C2 => n13358, ZN => n3788);
   U1860 : AOI221_X1 port map( B1 => n13316, B2 => n14678, C1 => n13313, C2 => 
                           n15752, A => n3796, ZN => n3795);
   U1861 : OAI222_X1 port map( A1 => n14774, A2 => n13310, B1 => n14710, B2 => 
                           n13307, C1 => n14742, C2 => n13304, ZN => n3796);
   U1862 : AOI221_X1 port map( B1 => n13262, B2 => n15000, C1 => n13259, C2 => 
                           n15652, A => n3804, ZN => n3803);
   U1863 : OAI222_X1 port map( A1 => n15096, A2 => n13256, B1 => n15032, B2 => 
                           n13253, C1 => n15064, C2 => n13250, ZN => n3804);
   U1864 : AOI221_X1 port map( B1 => n13370, B2 => n14265, C1 => n13367, C2 => 
                           n15883, A => n3751, ZN => n3750);
   U1865 : OAI222_X1 port map( A1 => n14361, A2 => n13364, B1 => n14297, B2 => 
                           n13361, C1 => n14329, C2 => n13358, ZN => n3751);
   U1866 : AOI221_X1 port map( B1 => n13316, B2 => n14677, C1 => n13313, C2 => 
                           n15751, A => n3759, ZN => n3758);
   U1867 : OAI222_X1 port map( A1 => n14773, A2 => n13310, B1 => n14709, B2 => 
                           n13307, C1 => n14741, C2 => n13304, ZN => n3759);
   U1868 : AOI221_X1 port map( B1 => n13262, B2 => n14999, C1 => n13259, C2 => 
                           n15651, A => n3767, ZN => n3766);
   U1869 : OAI222_X1 port map( A1 => n15095, A2 => n13256, B1 => n15031, B2 => 
                           n13253, C1 => n15063, C2 => n13250, ZN => n3767);
   U1870 : AOI221_X1 port map( B1 => n13370, B2 => n14264, C1 => n13367, C2 => 
                           n15882, A => n3714, ZN => n3713);
   U1871 : OAI222_X1 port map( A1 => n14360, A2 => n13364, B1 => n14296, B2 => 
                           n13361, C1 => n14328, C2 => n13358, ZN => n3714);
   U1872 : AOI221_X1 port map( B1 => n13316, B2 => n14676, C1 => n13313, C2 => 
                           n15750, A => n3722, ZN => n3721);
   U1873 : OAI222_X1 port map( A1 => n14772, A2 => n13310, B1 => n14708, B2 => 
                           n13307, C1 => n14740, C2 => n13304, ZN => n3722);
   U1874 : AOI221_X1 port map( B1 => n13262, B2 => n14998, C1 => n13259, C2 => 
                           n15650, A => n3730, ZN => n3729);
   U1875 : OAI222_X1 port map( A1 => n15094, A2 => n13256, B1 => n15030, B2 => 
                           n13253, C1 => n15062, C2 => n13250, ZN => n3730);
   U1876 : AOI221_X1 port map( B1 => n13370, B2 => n14263, C1 => n13367, C2 => 
                           n15881, A => n3677, ZN => n3676);
   U1877 : OAI222_X1 port map( A1 => n14359, A2 => n13364, B1 => n14295, B2 => 
                           n13361, C1 => n14327, C2 => n13358, ZN => n3677);
   U1878 : AOI221_X1 port map( B1 => n13316, B2 => n14675, C1 => n13313, C2 => 
                           n15749, A => n3685, ZN => n3684);
   U1879 : OAI222_X1 port map( A1 => n14771, A2 => n13310, B1 => n14707, B2 => 
                           n13307, C1 => n14739, C2 => n13304, ZN => n3685);
   U1880 : AOI221_X1 port map( B1 => n13262, B2 => n14997, C1 => n13259, C2 => 
                           n15649, A => n3693, ZN => n3692);
   U1881 : OAI222_X1 port map( A1 => n15093, A2 => n13256, B1 => n15029, B2 => 
                           n13253, C1 => n15061, C2 => n13250, ZN => n3693);
   U1882 : AOI221_X1 port map( B1 => n13370, B2 => n14262, C1 => n13367, C2 => 
                           n15880, A => n3640, ZN => n3639);
   U1883 : OAI222_X1 port map( A1 => n14358, A2 => n13364, B1 => n14294, B2 => 
                           n13361, C1 => n14326, C2 => n13358, ZN => n3640);
   U1884 : AOI221_X1 port map( B1 => n13316, B2 => n14674, C1 => n13313, C2 => 
                           n15748, A => n3648, ZN => n3647);
   U1885 : OAI222_X1 port map( A1 => n14770, A2 => n13310, B1 => n14706, B2 => 
                           n13307, C1 => n14738, C2 => n13304, ZN => n3648);
   U1886 : AOI221_X1 port map( B1 => n13262, B2 => n14996, C1 => n13259, C2 => 
                           n15648, A => n3656, ZN => n3655);
   U1887 : OAI222_X1 port map( A1 => n15092, A2 => n13256, B1 => n15028, B2 => 
                           n13253, C1 => n15060, C2 => n13250, ZN => n3656);
   U1888 : AOI221_X1 port map( B1 => n13370, B2 => n14261, C1 => n13367, C2 => 
                           n15879, A => n3603, ZN => n3602);
   U1889 : OAI222_X1 port map( A1 => n14357, A2 => n13364, B1 => n14293, B2 => 
                           n13361, C1 => n14325, C2 => n13358, ZN => n3603);
   U1890 : AOI221_X1 port map( B1 => n13316, B2 => n14673, C1 => n13313, C2 => 
                           n15747, A => n3611, ZN => n3610);
   U1891 : OAI222_X1 port map( A1 => n14769, A2 => n13310, B1 => n14705, B2 => 
                           n13307, C1 => n14737, C2 => n13304, ZN => n3611);
   U1892 : AOI221_X1 port map( B1 => n13262, B2 => n14995, C1 => n13259, C2 => 
                           n15647, A => n3619, ZN => n3618);
   U1893 : OAI222_X1 port map( A1 => n15091, A2 => n13256, B1 => n15027, B2 => 
                           n13253, C1 => n15059, C2 => n13250, ZN => n3619);
   U1894 : AOI221_X1 port map( B1 => n13370, B2 => n14260, C1 => n13367, C2 => 
                           n15878, A => n3566, ZN => n3565);
   U1895 : OAI222_X1 port map( A1 => n14356, A2 => n13364, B1 => n14292, B2 => 
                           n13361, C1 => n14324, C2 => n13358, ZN => n3566);
   U1896 : AOI221_X1 port map( B1 => n13316, B2 => n14672, C1 => n13313, C2 => 
                           n15746, A => n3574, ZN => n3573);
   U1897 : OAI222_X1 port map( A1 => n14768, A2 => n13310, B1 => n14704, B2 => 
                           n13307, C1 => n14736, C2 => n13304, ZN => n3574);
   U1898 : AOI221_X1 port map( B1 => n13262, B2 => n14994, C1 => n13259, C2 => 
                           n15646, A => n3582, ZN => n3581);
   U1899 : OAI222_X1 port map( A1 => n15090, A2 => n13256, B1 => n15026, B2 => 
                           n13253, C1 => n15058, C2 => n13250, ZN => n3582);
   U1900 : AOI221_X1 port map( B1 => n13370, B2 => n14259, C1 => n13367, C2 => 
                           n15877, A => n3529, ZN => n3528);
   U1901 : OAI222_X1 port map( A1 => n14355, A2 => n13364, B1 => n14291, B2 => 
                           n13361, C1 => n14323, C2 => n13358, ZN => n3529);
   U1902 : AOI221_X1 port map( B1 => n13316, B2 => n14671, C1 => n13313, C2 => 
                           n15745, A => n3537, ZN => n3536);
   U1903 : OAI222_X1 port map( A1 => n14767, A2 => n13310, B1 => n14703, B2 => 
                           n13307, C1 => n14735, C2 => n13304, ZN => n3537);
   U1904 : AOI221_X1 port map( B1 => n13370, B2 => n14258, C1 => n13367, C2 => 
                           n15876, A => n3492, ZN => n3491);
   U1905 : OAI222_X1 port map( A1 => n14354, A2 => n13364, B1 => n14290, B2 => 
                           n13361, C1 => n14322, C2 => n13358, ZN => n3492);
   U1906 : AOI221_X1 port map( B1 => n13316, B2 => n14670, C1 => n13313, C2 => 
                           n15744, A => n3500, ZN => n3499);
   U1907 : OAI222_X1 port map( A1 => n14766, A2 => n13310, B1 => n14702, B2 => 
                           n13307, C1 => n14734, C2 => n13304, ZN => n3500);
   U1908 : AOI221_X1 port map( B1 => n13370, B2 => n14257, C1 => n13367, C2 => 
                           n15875, A => n3455, ZN => n3454);
   U1909 : OAI222_X1 port map( A1 => n14353, A2 => n13364, B1 => n14289, B2 => 
                           n13361, C1 => n14321, C2 => n13358, ZN => n3455);
   U1910 : AOI221_X1 port map( B1 => n13316, B2 => n14669, C1 => n13313, C2 => 
                           n15743, A => n3463, ZN => n3462);
   U1911 : OAI222_X1 port map( A1 => n14765, A2 => n13310, B1 => n14701, B2 => 
                           n13307, C1 => n14733, C2 => n13304, ZN => n3463);
   U1912 : AOI221_X1 port map( B1 => n13370, B2 => n14256, C1 => n13367, C2 => 
                           n15874, A => n3418, ZN => n3417);
   U1913 : OAI222_X1 port map( A1 => n14352, A2 => n13364, B1 => n14288, B2 => 
                           n13361, C1 => n14320, C2 => n13358, ZN => n3418);
   U1914 : AOI221_X1 port map( B1 => n13316, B2 => n14668, C1 => n13313, C2 => 
                           n15742, A => n3426, ZN => n3425);
   U1915 : OAI222_X1 port map( A1 => n14764, A2 => n13310, B1 => n14700, B2 => 
                           n13307, C1 => n14732, C2 => n13304, ZN => n3426);
   U1916 : AOI221_X1 port map( B1 => n13371, B2 => n14255, C1 => n13368, C2 => 
                           n15597, A => n3381, ZN => n3380);
   U1917 : OAI222_X1 port map( A1 => n14351, A2 => n13365, B1 => n14287, B2 => 
                           n13362, C1 => n14319, C2 => n13359, ZN => n3381);
   U1918 : AOI221_X1 port map( B1 => n13317, B2 => n14667, C1 => n13314, C2 => 
                           n15573, A => n3389, ZN => n3388);
   U1919 : OAI222_X1 port map( A1 => n14763, A2 => n13311, B1 => n14699, B2 => 
                           n13308, C1 => n14731, C2 => n13305, ZN => n3389);
   U1920 : AOI221_X1 port map( B1 => n13263, B2 => n14989, C1 => n13260, C2 => 
                           n15641, A => n3397, ZN => n3396);
   U1921 : OAI222_X1 port map( A1 => n15085, A2 => n13257, B1 => n15021, B2 => 
                           n13254, C1 => n15053, C2 => n13251, ZN => n3397);
   U1922 : AOI221_X1 port map( B1 => n13209, B2 => n15437, C1 => n13206, C2 => 
                           n15405, A => n3405, ZN => n3404);
   U1923 : OAI222_X1 port map( A1 => n15533, A2 => n13203, B1 => n15469, B2 => 
                           n13200, C1 => n15501, C2 => n13197, ZN => n3405);
   U1924 : AOI221_X1 port map( B1 => n13371, B2 => n14254, C1 => n13368, C2 => 
                           n15596, A => n3344, ZN => n3343);
   U1925 : OAI222_X1 port map( A1 => n14350, A2 => n13365, B1 => n14286, B2 => 
                           n13362, C1 => n14318, C2 => n13359, ZN => n3344);
   U1926 : AOI221_X1 port map( B1 => n13317, B2 => n14666, C1 => n13314, C2 => 
                           n15572, A => n3352, ZN => n3351);
   U1927 : OAI222_X1 port map( A1 => n14762, A2 => n13311, B1 => n14698, B2 => 
                           n13308, C1 => n14730, C2 => n13305, ZN => n3352);
   U1928 : AOI221_X1 port map( B1 => n13263, B2 => n14988, C1 => n13260, C2 => 
                           n15640, A => n3360, ZN => n3359);
   U1929 : OAI222_X1 port map( A1 => n15084, A2 => n13257, B1 => n15020, B2 => 
                           n13254, C1 => n15052, C2 => n13251, ZN => n3360);
   U1930 : AOI221_X1 port map( B1 => n13209, B2 => n15436, C1 => n13206, C2 => 
                           n15404, A => n3368, ZN => n3367);
   U1931 : OAI222_X1 port map( A1 => n15532, A2 => n13203, B1 => n15468, B2 => 
                           n13200, C1 => n15500, C2 => n13197, ZN => n3368);
   U1932 : AOI221_X1 port map( B1 => n13371, B2 => n14253, C1 => n13368, C2 => 
                           n15595, A => n3307, ZN => n3306);
   U1933 : OAI222_X1 port map( A1 => n14349, A2 => n13365, B1 => n14285, B2 => 
                           n13362, C1 => n14317, C2 => n13359, ZN => n3307);
   U1934 : AOI221_X1 port map( B1 => n13317, B2 => n14665, C1 => n13314, C2 => 
                           n15571, A => n3315, ZN => n3314);
   U1935 : OAI222_X1 port map( A1 => n14761, A2 => n13311, B1 => n14697, B2 => 
                           n13308, C1 => n14729, C2 => n13305, ZN => n3315);
   U1936 : AOI221_X1 port map( B1 => n13263, B2 => n14987, C1 => n13260, C2 => 
                           n15639, A => n3323, ZN => n3322);
   U1937 : OAI222_X1 port map( A1 => n15083, A2 => n13257, B1 => n15019, B2 => 
                           n13254, C1 => n15051, C2 => n13251, ZN => n3323);
   U1938 : AOI221_X1 port map( B1 => n13209, B2 => n15435, C1 => n13206, C2 => 
                           n15403, A => n3331, ZN => n3330);
   U1939 : OAI222_X1 port map( A1 => n15531, A2 => n13203, B1 => n15467, B2 => 
                           n13200, C1 => n15499, C2 => n13197, ZN => n3331);
   U1940 : AOI221_X1 port map( B1 => n13371, B2 => n14252, C1 => n13368, C2 => 
                           n15594, A => n3270, ZN => n3269);
   U1941 : OAI222_X1 port map( A1 => n14348, A2 => n13365, B1 => n14284, B2 => 
                           n13362, C1 => n14316, C2 => n13359, ZN => n3270);
   U1942 : AOI221_X1 port map( B1 => n13317, B2 => n14664, C1 => n13314, C2 => 
                           n15570, A => n3278, ZN => n3277);
   U1943 : OAI222_X1 port map( A1 => n14760, A2 => n13311, B1 => n14696, B2 => 
                           n13308, C1 => n14728, C2 => n13305, ZN => n3278);
   U1944 : AOI221_X1 port map( B1 => n13263, B2 => n14986, C1 => n13260, C2 => 
                           n15638, A => n3286, ZN => n3285);
   U1945 : OAI222_X1 port map( A1 => n15082, A2 => n13257, B1 => n15018, B2 => 
                           n13254, C1 => n15050, C2 => n13251, ZN => n3286);
   U1946 : AOI221_X1 port map( B1 => n13209, B2 => n15434, C1 => n13206, C2 => 
                           n15402, A => n3294, ZN => n3293);
   U1947 : OAI222_X1 port map( A1 => n15530, A2 => n13203, B1 => n15466, B2 => 
                           n13200, C1 => n15498, C2 => n13197, ZN => n3294);
   U1948 : AOI221_X1 port map( B1 => n13221, B2 => n15733, C1 => n13218, C2 => 
                           n15622, A => n3252, ZN => n3245);
   U1949 : OAI22_X1 port map( A1 => n14823, A2 => n13215, B1 => n14791, B2 => 
                           n13212, ZN => n3252);
   U1950 : AOI221_X1 port map( B1 => n13221, B2 => n15732, C1 => n13218, C2 => 
                           n15621, A => n3215, ZN => n3208);
   U1951 : OAI22_X1 port map( A1 => n14822, A2 => n13215, B1 => n14790, B2 => 
                           n13212, ZN => n3215);
   U1952 : AOI221_X1 port map( B1 => n13221, B2 => n15731, C1 => n13218, C2 => 
                           n15620, A => n3178, ZN => n3171);
   U1953 : OAI22_X1 port map( A1 => n14821, A2 => n13215, B1 => n14789, B2 => 
                           n13212, ZN => n3178);
   U1954 : AOI221_X1 port map( B1 => n12993, B2 => n15736, C1 => n12990, C2 => 
                           n15625, A => n4647, ZN => n4640);
   U1955 : OAI22_X1 port map( A1 => n14826, A2 => n12987, B1 => n14794, B2 => 
                           n12984, ZN => n4647);
   U1956 : AOI221_X1 port map( B1 => n12993, B2 => n15735, C1 => n12990, C2 => 
                           n15624, A => n4610, ZN => n4603);
   U1957 : OAI22_X1 port map( A1 => n14825, A2 => n12987, B1 => n14793, B2 => 
                           n12984, ZN => n4610);
   U1958 : AOI221_X1 port map( B1 => n12993, B2 => n15734, C1 => n12990, C2 => 
                           n15623, A => n4573, ZN => n4566);
   U1959 : OAI22_X1 port map( A1 => n14824, A2 => n12987, B1 => n14792, B2 => 
                           n12984, ZN => n4573);
   U1960 : AOI221_X1 port map( B1 => n12993, B2 => n15733, C1 => n12990, C2 => 
                           n15622, A => n4536, ZN => n4529);
   U1961 : OAI22_X1 port map( A1 => n14823, A2 => n12987, B1 => n14791, B2 => 
                           n12984, ZN => n4536);
   U1962 : AOI221_X1 port map( B1 => n12993, B2 => n15732, C1 => n12990, C2 => 
                           n15621, A => n4499, ZN => n4492);
   U1963 : OAI22_X1 port map( A1 => n14822, A2 => n12987, B1 => n14790, B2 => 
                           n12984, ZN => n4499);
   U1964 : AOI221_X1 port map( B1 => n12993, B2 => n15731, C1 => n12990, C2 => 
                           n15620, A => n4462, ZN => n4455);
   U1965 : OAI22_X1 port map( A1 => n14821, A2 => n12987, B1 => n14789, B2 => 
                           n12984, ZN => n4462);
   U1966 : AOI221_X1 port map( B1 => n12993, B2 => n15737, C1 => n12990, C2 => 
                           n15626, A => n4684, ZN => n4677);
   U1967 : OAI22_X1 port map( A1 => n14827, A2 => n12987, B1 => n14795, B2 => 
                           n12984, ZN => n4684);
   U1968 : AOI221_X1 port map( B1 => n13221, B2 => n15737, C1 => n13218, C2 => 
                           n15626, A => n3400, ZN => n3393);
   U1969 : OAI22_X1 port map( A1 => n14827, A2 => n13215, B1 => n14795, B2 => 
                           n13212, ZN => n3400);
   U1970 : AOI221_X1 port map( B1 => n13221, B2 => n15736, C1 => n13218, C2 => 
                           n15625, A => n3363, ZN => n3356);
   U1971 : OAI22_X1 port map( A1 => n14826, A2 => n13215, B1 => n14794, B2 => 
                           n13212, ZN => n3363);
   U1972 : AOI221_X1 port map( B1 => n13221, B2 => n15735, C1 => n13218, C2 => 
                           n15624, A => n3326, ZN => n3319);
   U1973 : OAI22_X1 port map( A1 => n14825, A2 => n13215, B1 => n14793, B2 => 
                           n13212, ZN => n3326);
   U1974 : AOI221_X1 port map( B1 => n13221, B2 => n15734, C1 => n13218, C2 => 
                           n15623, A => n3289, ZN => n3282);
   U1975 : OAI22_X1 port map( A1 => n14824, A2 => n13215, B1 => n14792, B2 => 
                           n13212, ZN => n3289);
   U1976 : OAI22_X1 port map( A1 => n14592, A2 => n13296, B1 => n14624, B2 => 
                           n13293, ZN => n3242);
   U1977 : OAI22_X1 port map( A1 => n14411, A2 => n13269, B1 => n14379, B2 => 
                           n13266, ZN => n3244);
   U1978 : OAI22_X1 port map( A1 => n14591, A2 => n13296, B1 => n14623, B2 => 
                           n13293, ZN => n3205);
   U1979 : OAI22_X1 port map( A1 => n14410, A2 => n13269, B1 => n14378, B2 => 
                           n13266, ZN => n3207);
   U1980 : OAI22_X1 port map( A1 => n14590, A2 => n13296, B1 => n14622, B2 => 
                           n13293, ZN => n3168);
   U1981 : OAI22_X1 port map( A1 => n14409, A2 => n13269, B1 => n14377, B2 => 
                           n13266, ZN => n3170);
   U1982 : OAI22_X1 port map( A1 => n14589, A2 => n13296, B1 => n14621, B2 => 
                           n13293, ZN => n3084);
   U1983 : OAI22_X1 port map( A1 => n14408, A2 => n13269, B1 => n14376, B2 => 
                           n13266, ZN => n3095);
   U1984 : OAI22_X1 port map( A1 => n14627, A2 => n13068, B1 => n14595, B2 => 
                           n13065, ZN => n4637);
   U1985 : OAI22_X1 port map( A1 => n14414, A2 => n13041, B1 => n14382, B2 => 
                           n13038, ZN => n4639);
   U1986 : OAI22_X1 port map( A1 => n14626, A2 => n13068, B1 => n14594, B2 => 
                           n13065, ZN => n4600);
   U1987 : OAI22_X1 port map( A1 => n14413, A2 => n13041, B1 => n14381, B2 => 
                           n13038, ZN => n4602);
   U1988 : OAI22_X1 port map( A1 => n14625, A2 => n13068, B1 => n14593, B2 => 
                           n13065, ZN => n4563);
   U1989 : OAI22_X1 port map( A1 => n14412, A2 => n13041, B1 => n14380, B2 => 
                           n13038, ZN => n4565);
   U1990 : OAI22_X1 port map( A1 => n14624, A2 => n13068, B1 => n14592, B2 => 
                           n13065, ZN => n4526);
   U1991 : OAI22_X1 port map( A1 => n14411, A2 => n13041, B1 => n14379, B2 => 
                           n13038, ZN => n4528);
   U1992 : OAI22_X1 port map( A1 => n14623, A2 => n13068, B1 => n14591, B2 => 
                           n13065, ZN => n4489);
   U1993 : OAI22_X1 port map( A1 => n14410, A2 => n13041, B1 => n14378, B2 => 
                           n13038, ZN => n4491);
   U1994 : OAI22_X1 port map( A1 => n14622, A2 => n13068, B1 => n14590, B2 => 
                           n13065, ZN => n4452);
   U1995 : OAI22_X1 port map( A1 => n14409, A2 => n13041, B1 => n14377, B2 => 
                           n13038, ZN => n4454);
   U1996 : OAI22_X1 port map( A1 => n14621, A2 => n13068, B1 => n14589, B2 => 
                           n13065, ZN => n4368);
   U1997 : OAI22_X1 port map( A1 => n14408, A2 => n13041, B1 => n14376, B2 => 
                           n13038, ZN => n4379);
   U1998 : OAI22_X1 port map( A1 => n14628, A2 => n13068, B1 => n14596, B2 => 
                           n13065, ZN => n4674);
   U1999 : OAI22_X1 port map( A1 => n14415, A2 => n13041, B1 => n14383, B2 => 
                           n13038, ZN => n4676);
   U2000 : OAI22_X1 port map( A1 => n14596, A2 => n13296, B1 => n14628, B2 => 
                           n13293, ZN => n3390);
   U2001 : OAI22_X1 port map( A1 => n14415, A2 => n13269, B1 => n14383, B2 => 
                           n13266, ZN => n3392);
   U2002 : OAI22_X1 port map( A1 => n14595, A2 => n13296, B1 => n14627, B2 => 
                           n13293, ZN => n3353);
   U2003 : OAI22_X1 port map( A1 => n14414, A2 => n13269, B1 => n14382, B2 => 
                           n13266, ZN => n3355);
   U2004 : OAI22_X1 port map( A1 => n14594, A2 => n13296, B1 => n14626, B2 => 
                           n13293, ZN => n3316);
   U2005 : OAI22_X1 port map( A1 => n14413, A2 => n13269, B1 => n14381, B2 => 
                           n13266, ZN => n3318);
   U2006 : OAI22_X1 port map( A1 => n14593, A2 => n13296, B1 => n14625, B2 => 
                           n13293, ZN => n3279);
   U2007 : OAI22_X1 port map( A1 => n14412, A2 => n13269, B1 => n14380, B2 => 
                           n13266, ZN => n3281);
   U2008 : OAI22_X1 port map( A1 => n14652, A2 => n13066, B1 => n14620, B2 => 
                           n13063, ZN => n5694);
   U2009 : OAI22_X1 port map( A1 => n14439, A2 => n13039, B1 => n14407, B2 => 
                           n13036, ZN => n5698);
   U2010 : OAI22_X1 port map( A1 => n14651, A2 => n13066, B1 => n14619, B2 => 
                           n13063, ZN => n5610);
   U2011 : OAI22_X1 port map( A1 => n14438, A2 => n13039, B1 => n14406, B2 => 
                           n13036, ZN => n5614);
   U2012 : OAI22_X1 port map( A1 => n14650, A2 => n13066, B1 => n14618, B2 => 
                           n13063, ZN => n5549);
   U2013 : OAI22_X1 port map( A1 => n14437, A2 => n13039, B1 => n14405, B2 => 
                           n13036, ZN => n5551);
   U2014 : OAI22_X1 port map( A1 => n14649, A2 => n13066, B1 => n14617, B2 => 
                           n13063, ZN => n5488);
   U2015 : OAI22_X1 port map( A1 => n14436, A2 => n13039, B1 => n14404, B2 => 
                           n13036, ZN => n5490);
   U2016 : OAI22_X1 port map( A1 => n14648, A2 => n13066, B1 => n14616, B2 => 
                           n13063, ZN => n5429);
   U2017 : OAI22_X1 port map( A1 => n14435, A2 => n13039, B1 => n14403, B2 => 
                           n13036, ZN => n5431);
   U2018 : OAI22_X1 port map( A1 => n14647, A2 => n13066, B1 => n14615, B2 => 
                           n13063, ZN => n5377);
   U2019 : OAI22_X1 port map( A1 => n14434, A2 => n13039, B1 => n14402, B2 => 
                           n13036, ZN => n5379);
   U2020 : OAI22_X1 port map( A1 => n14646, A2 => n13066, B1 => n14614, B2 => 
                           n13063, ZN => n5340);
   U2021 : OAI22_X1 port map( A1 => n14433, A2 => n13039, B1 => n14401, B2 => 
                           n13036, ZN => n5342);
   U2022 : OAI22_X1 port map( A1 => n14645, A2 => n13066, B1 => n14613, B2 => 
                           n13063, ZN => n5303);
   U2023 : OAI22_X1 port map( A1 => n14432, A2 => n13039, B1 => n14400, B2 => 
                           n13036, ZN => n5305);
   U2024 : OAI22_X1 port map( A1 => n14644, A2 => n13066, B1 => n14612, B2 => 
                           n13063, ZN => n5266);
   U2025 : OAI22_X1 port map( A1 => n14431, A2 => n13039, B1 => n14399, B2 => 
                           n13036, ZN => n5268);
   U2026 : OAI22_X1 port map( A1 => n14643, A2 => n13066, B1 => n14611, B2 => 
                           n13063, ZN => n5229);
   U2027 : OAI22_X1 port map( A1 => n14430, A2 => n13039, B1 => n14398, B2 => 
                           n13036, ZN => n5231);
   U2028 : OAI22_X1 port map( A1 => n14642, A2 => n13066, B1 => n14610, B2 => 
                           n13063, ZN => n5192);
   U2029 : OAI22_X1 port map( A1 => n14429, A2 => n13039, B1 => n14397, B2 => 
                           n13036, ZN => n5194);
   U2030 : OAI22_X1 port map( A1 => n14641, A2 => n13066, B1 => n14609, B2 => 
                           n13063, ZN => n5155);
   U2031 : OAI22_X1 port map( A1 => n14428, A2 => n13039, B1 => n14396, B2 => 
                           n13036, ZN => n5157);
   U2032 : OAI22_X1 port map( A1 => n14640, A2 => n13067, B1 => n14608, B2 => 
                           n13064, ZN => n5118);
   U2033 : OAI22_X1 port map( A1 => n14427, A2 => n13040, B1 => n14395, B2 => 
                           n13037, ZN => n5120);
   U2034 : OAI22_X1 port map( A1 => n14639, A2 => n13067, B1 => n14607, B2 => 
                           n13064, ZN => n5081);
   U2035 : OAI22_X1 port map( A1 => n14426, A2 => n13040, B1 => n14394, B2 => 
                           n13037, ZN => n5083);
   U2036 : OAI22_X1 port map( A1 => n14638, A2 => n13067, B1 => n14606, B2 => 
                           n13064, ZN => n5044);
   U2037 : OAI22_X1 port map( A1 => n14425, A2 => n13040, B1 => n14393, B2 => 
                           n13037, ZN => n5046);
   U2038 : OAI22_X1 port map( A1 => n14637, A2 => n13067, B1 => n14605, B2 => 
                           n13064, ZN => n5007);
   U2039 : OAI22_X1 port map( A1 => n14424, A2 => n13040, B1 => n14392, B2 => 
                           n13037, ZN => n5009);
   U2040 : OAI22_X1 port map( A1 => n14636, A2 => n13067, B1 => n14604, B2 => 
                           n13064, ZN => n4970);
   U2041 : OAI22_X1 port map( A1 => n14423, A2 => n13040, B1 => n14391, B2 => 
                           n13037, ZN => n4972);
   U2042 : OAI22_X1 port map( A1 => n14635, A2 => n13067, B1 => n14603, B2 => 
                           n13064, ZN => n4933);
   U2043 : OAI22_X1 port map( A1 => n14422, A2 => n13040, B1 => n14390, B2 => 
                           n13037, ZN => n4935);
   U2044 : OAI22_X1 port map( A1 => n14634, A2 => n13067, B1 => n14602, B2 => 
                           n13064, ZN => n4896);
   U2045 : OAI22_X1 port map( A1 => n14421, A2 => n13040, B1 => n14389, B2 => 
                           n13037, ZN => n4898);
   U2046 : OAI22_X1 port map( A1 => n14633, A2 => n13067, B1 => n14601, B2 => 
                           n13064, ZN => n4859);
   U2047 : OAI22_X1 port map( A1 => n14420, A2 => n13040, B1 => n14388, B2 => 
                           n13037, ZN => n4861);
   U2048 : OAI22_X1 port map( A1 => n14632, A2 => n13067, B1 => n14600, B2 => 
                           n13064, ZN => n4822);
   U2049 : OAI22_X1 port map( A1 => n14419, A2 => n13040, B1 => n14387, B2 => 
                           n13037, ZN => n4824);
   U2050 : OAI22_X1 port map( A1 => n14631, A2 => n13067, B1 => n14599, B2 => 
                           n13064, ZN => n4785);
   U2051 : OAI22_X1 port map( A1 => n14418, A2 => n13040, B1 => n14386, B2 => 
                           n13037, ZN => n4787);
   U2052 : OAI22_X1 port map( A1 => n14630, A2 => n13067, B1 => n14598, B2 => 
                           n13064, ZN => n4748);
   U2053 : OAI22_X1 port map( A1 => n14417, A2 => n13040, B1 => n14385, B2 => 
                           n13037, ZN => n4750);
   U2054 : OAI22_X1 port map( A1 => n14629, A2 => n13067, B1 => n14597, B2 => 
                           n13064, ZN => n4711);
   U2055 : OAI22_X1 port map( A1 => n14416, A2 => n13040, B1 => n14384, B2 => 
                           n13037, ZN => n4713);
   U2056 : OAI22_X1 port map( A1 => n14620, A2 => n13294, B1 => n14652, B2 => 
                           n13291, ZN => n4291);
   U2057 : OAI22_X1 port map( A1 => n14439, A2 => n13267, B1 => n14407, B2 => 
                           n13264, ZN => n4293);
   U2058 : OAI22_X1 port map( A1 => n14619, A2 => n13294, B1 => n14651, B2 => 
                           n13291, ZN => n4241);
   U2059 : OAI22_X1 port map( A1 => n14438, A2 => n13267, B1 => n14406, B2 => 
                           n13264, ZN => n4243);
   U2060 : OAI22_X1 port map( A1 => n14618, A2 => n13294, B1 => n14650, B2 => 
                           n13291, ZN => n4204);
   U2061 : OAI22_X1 port map( A1 => n14437, A2 => n13267, B1 => n14405, B2 => 
                           n13264, ZN => n4206);
   U2062 : OAI22_X1 port map( A1 => n14617, A2 => n13294, B1 => n14649, B2 => 
                           n13291, ZN => n4167);
   U2063 : OAI22_X1 port map( A1 => n14436, A2 => n13267, B1 => n14404, B2 => 
                           n13264, ZN => n4169);
   U2064 : OAI22_X1 port map( A1 => n14616, A2 => n13294, B1 => n14648, B2 => 
                           n13291, ZN => n4130);
   U2065 : OAI22_X1 port map( A1 => n14435, A2 => n13267, B1 => n14403, B2 => 
                           n13264, ZN => n4132);
   U2066 : OAI22_X1 port map( A1 => n14615, A2 => n13294, B1 => n14647, B2 => 
                           n13291, ZN => n4093);
   U2067 : OAI22_X1 port map( A1 => n14434, A2 => n13267, B1 => n14402, B2 => 
                           n13264, ZN => n4095);
   U2068 : OAI22_X1 port map( A1 => n14614, A2 => n13294, B1 => n14646, B2 => 
                           n13291, ZN => n4056);
   U2069 : OAI22_X1 port map( A1 => n14433, A2 => n13267, B1 => n14401, B2 => 
                           n13264, ZN => n4058);
   U2070 : OAI22_X1 port map( A1 => n14613, A2 => n13294, B1 => n14645, B2 => 
                           n13291, ZN => n4019);
   U2071 : OAI22_X1 port map( A1 => n14432, A2 => n13267, B1 => n14400, B2 => 
                           n13264, ZN => n4021);
   U2072 : OAI22_X1 port map( A1 => n14612, A2 => n13294, B1 => n14644, B2 => 
                           n13291, ZN => n3982);
   U2073 : OAI22_X1 port map( A1 => n14431, A2 => n13267, B1 => n14399, B2 => 
                           n13264, ZN => n3984);
   U2074 : OAI22_X1 port map( A1 => n14611, A2 => n13294, B1 => n14643, B2 => 
                           n13291, ZN => n3945);
   U2075 : OAI22_X1 port map( A1 => n14430, A2 => n13267, B1 => n14398, B2 => 
                           n13264, ZN => n3947);
   U2076 : OAI22_X1 port map( A1 => n14610, A2 => n13294, B1 => n14642, B2 => 
                           n13291, ZN => n3908);
   U2077 : OAI22_X1 port map( A1 => n14429, A2 => n13267, B1 => n14397, B2 => 
                           n13264, ZN => n3910);
   U2078 : OAI22_X1 port map( A1 => n14609, A2 => n13294, B1 => n14641, B2 => 
                           n13291, ZN => n3871);
   U2079 : OAI22_X1 port map( A1 => n14428, A2 => n13267, B1 => n14396, B2 => 
                           n13264, ZN => n3873);
   U2080 : OAI22_X1 port map( A1 => n14608, A2 => n13295, B1 => n14640, B2 => 
                           n13292, ZN => n3834);
   U2081 : OAI22_X1 port map( A1 => n14427, A2 => n13268, B1 => n14395, B2 => 
                           n13265, ZN => n3836);
   U2082 : OAI22_X1 port map( A1 => n14607, A2 => n13295, B1 => n14639, B2 => 
                           n13292, ZN => n3797);
   U2083 : OAI22_X1 port map( A1 => n14426, A2 => n13268, B1 => n14394, B2 => 
                           n13265, ZN => n3799);
   U2084 : OAI22_X1 port map( A1 => n14606, A2 => n13295, B1 => n14638, B2 => 
                           n13292, ZN => n3760);
   U2085 : OAI22_X1 port map( A1 => n14425, A2 => n13268, B1 => n14393, B2 => 
                           n13265, ZN => n3762);
   U2086 : OAI22_X1 port map( A1 => n14605, A2 => n13295, B1 => n14637, B2 => 
                           n13292, ZN => n3723);
   U2087 : OAI22_X1 port map( A1 => n14424, A2 => n13268, B1 => n14392, B2 => 
                           n13265, ZN => n3725);
   U2088 : OAI22_X1 port map( A1 => n14604, A2 => n13295, B1 => n14636, B2 => 
                           n13292, ZN => n3686);
   U2089 : OAI22_X1 port map( A1 => n14423, A2 => n13268, B1 => n14391, B2 => 
                           n13265, ZN => n3688);
   U2090 : OAI22_X1 port map( A1 => n14603, A2 => n13295, B1 => n14635, B2 => 
                           n13292, ZN => n3649);
   U2091 : OAI22_X1 port map( A1 => n14422, A2 => n13268, B1 => n14390, B2 => 
                           n13265, ZN => n3651);
   U2092 : OAI22_X1 port map( A1 => n14602, A2 => n13295, B1 => n14634, B2 => 
                           n13292, ZN => n3612);
   U2093 : OAI22_X1 port map( A1 => n14421, A2 => n13268, B1 => n14389, B2 => 
                           n13265, ZN => n3614);
   U2094 : OAI22_X1 port map( A1 => n14601, A2 => n13295, B1 => n14633, B2 => 
                           n13292, ZN => n3575);
   U2095 : OAI22_X1 port map( A1 => n14420, A2 => n13268, B1 => n14388, B2 => 
                           n13265, ZN => n3577);
   U2096 : OAI22_X1 port map( A1 => n14600, A2 => n13295, B1 => n14632, B2 => 
                           n13292, ZN => n3538);
   U2097 : OAI22_X1 port map( A1 => n14419, A2 => n13268, B1 => n14387, B2 => 
                           n13265, ZN => n3540);
   U2098 : OAI22_X1 port map( A1 => n14599, A2 => n13295, B1 => n14631, B2 => 
                           n13292, ZN => n3501);
   U2099 : OAI22_X1 port map( A1 => n14418, A2 => n13268, B1 => n14386, B2 => 
                           n13265, ZN => n3503);
   U2100 : OAI22_X1 port map( A1 => n14598, A2 => n13295, B1 => n14630, B2 => 
                           n13292, ZN => n3464);
   U2101 : OAI22_X1 port map( A1 => n14417, A2 => n13268, B1 => n14385, B2 => 
                           n13265, ZN => n3466);
   U2102 : OAI22_X1 port map( A1 => n14597, A2 => n13295, B1 => n14629, B2 => 
                           n13292, ZN => n3427);
   U2103 : OAI22_X1 port map( A1 => n14416, A2 => n13268, B1 => n14384, B2 => 
                           n13265, ZN => n3429);
   U2104 : AOI221_X1 port map( B1 => n12992, B2 => n15741, C1 => n12989, C2 => 
                           n15709, A => n4832, ZN => n4825);
   U2105 : OAI22_X1 port map( A1 => n14831, A2 => n12986, B1 => n14799, B2 => 
                           n12983, ZN => n4832);
   U2106 : AOI221_X1 port map( B1 => n12992, B2 => n15740, C1 => n12989, C2 => 
                           n15708, A => n4795, ZN => n4788);
   U2107 : OAI22_X1 port map( A1 => n14830, A2 => n12986, B1 => n14798, B2 => 
                           n12983, ZN => n4795);
   U2108 : AOI221_X1 port map( B1 => n12992, B2 => n15739, C1 => n12989, C2 => 
                           n15707, A => n4758, ZN => n4751);
   U2109 : OAI22_X1 port map( A1 => n14829, A2 => n12986, B1 => n14797, B2 => 
                           n12983, ZN => n4758);
   U2110 : AOI221_X1 port map( B1 => n12992, B2 => n15738, C1 => n12989, C2 => 
                           n15706, A => n4721, ZN => n4714);
   U2111 : OAI22_X1 port map( A1 => n14828, A2 => n12986, B1 => n14796, B2 => 
                           n12983, ZN => n4721);
   U2112 : AOI221_X1 port map( B1 => n13220, B2 => n15741, C1 => n13217, C2 => 
                           n15709, A => n3548, ZN => n3541);
   U2113 : OAI22_X1 port map( A1 => n14831, A2 => n13214, B1 => n14799, B2 => 
                           n13211, ZN => n3548);
   U2114 : AOI221_X1 port map( B1 => n13220, B2 => n15740, C1 => n13217, C2 => 
                           n15708, A => n3511, ZN => n3504);
   U2115 : OAI22_X1 port map( A1 => n14830, A2 => n13214, B1 => n14798, B2 => 
                           n13211, ZN => n3511);
   U2116 : AOI221_X1 port map( B1 => n13220, B2 => n15739, C1 => n13217, C2 => 
                           n15707, A => n3474, ZN => n3467);
   U2117 : OAI22_X1 port map( A1 => n14829, A2 => n13214, B1 => n14797, B2 => 
                           n13211, ZN => n3474);
   U2118 : AOI221_X1 port map( B1 => n13220, B2 => n15738, C1 => n13217, C2 => 
                           n15706, A => n3437, ZN => n3430);
   U2119 : OAI22_X1 port map( A1 => n14828, A2 => n13214, B1 => n14796, B2 => 
                           n13211, ZN => n3437);
   U2120 : OAI22_X1 port map( A1 => n13829, A2 => n13384, B1 => n13387, B2 => 
                           n15557, ZN => n7674);
   U2121 : OAI22_X1 port map( A1 => n13829, A2 => n13395, B1 => n13390, B2 => 
                           n15525, ZN => n7706);
   U2122 : OAI22_X1 port map( A1 => n13829, A2 => n13401, B1 => n13396, B2 => 
                           n15493, ZN => n7738);
   U2123 : OAI22_X1 port map( A1 => n13835, A2 => n13401, B1 => n13396, B2 => 
                           n15492, ZN => n7739);
   U2124 : OAI22_X1 port map( A1 => n13841, A2 => n13401, B1 => n13396, B2 => 
                           n15491, ZN => n7740);
   U2125 : OAI22_X1 port map( A1 => n13847, A2 => n13401, B1 => n13396, B2 => 
                           n15490, ZN => n7741);
   U2126 : OAI22_X1 port map( A1 => n13853, A2 => n13401, B1 => n13396, B2 => 
                           n15489, ZN => n7742);
   U2127 : OAI22_X1 port map( A1 => n13859, A2 => n13401, B1 => n13396, B2 => 
                           n15488, ZN => n7743);
   U2128 : OAI22_X1 port map( A1 => n13865, A2 => n13401, B1 => n13396, B2 => 
                           n15487, ZN => n7744);
   U2129 : OAI22_X1 port map( A1 => n13871, A2 => n13401, B1 => n13396, B2 => 
                           n15486, ZN => n7745);
   U2130 : OAI22_X1 port map( A1 => n13877, A2 => n13400, B1 => n13396, B2 => 
                           n15485, ZN => n7746);
   U2131 : OAI22_X1 port map( A1 => n13883, A2 => n13400, B1 => n13396, B2 => 
                           n15484, ZN => n7747);
   U2132 : OAI22_X1 port map( A1 => n13889, A2 => n13400, B1 => n13396, B2 => 
                           n15483, ZN => n7748);
   U2133 : OAI22_X1 port map( A1 => n13895, A2 => n13400, B1 => n13396, B2 => 
                           n15482, ZN => n7749);
   U2134 : OAI22_X1 port map( A1 => n13901, A2 => n13400, B1 => n13397, B2 => 
                           n15481, ZN => n7750);
   U2135 : OAI22_X1 port map( A1 => n13907, A2 => n13400, B1 => n13397, B2 => 
                           n15480, ZN => n7751);
   U2136 : OAI22_X1 port map( A1 => n13913, A2 => n13400, B1 => n13397, B2 => 
                           n15479, ZN => n7752);
   U2137 : OAI22_X1 port map( A1 => n13919, A2 => n13400, B1 => n13397, B2 => 
                           n15478, ZN => n7753);
   U2138 : OAI22_X1 port map( A1 => n13925, A2 => n13400, B1 => n13397, B2 => 
                           n15477, ZN => n7754);
   U2139 : OAI22_X1 port map( A1 => n13931, A2 => n13400, B1 => n13397, B2 => 
                           n15476, ZN => n7755);
   U2140 : OAI22_X1 port map( A1 => n13937, A2 => n13400, B1 => n13397, B2 => 
                           n15475, ZN => n7756);
   U2141 : OAI22_X1 port map( A1 => n13943, A2 => n13400, B1 => n13397, B2 => 
                           n15474, ZN => n7757);
   U2142 : OAI22_X1 port map( A1 => n13949, A2 => n13399, B1 => n13397, B2 => 
                           n15473, ZN => n7758);
   U2143 : OAI22_X1 port map( A1 => n13955, A2 => n13399, B1 => n13397, B2 => 
                           n15472, ZN => n7759);
   U2144 : OAI22_X1 port map( A1 => n13961, A2 => n13399, B1 => n13397, B2 => 
                           n15471, ZN => n7760);
   U2145 : OAI22_X1 port map( A1 => n13967, A2 => n13399, B1 => n13397, B2 => 
                           n15470, ZN => n7761);
   U2146 : OAI22_X1 port map( A1 => n13973, A2 => n13399, B1 => n13398, B2 => 
                           n15469, ZN => n7762);
   U2147 : OAI22_X1 port map( A1 => n13979, A2 => n13399, B1 => n13398, B2 => 
                           n15468, ZN => n7763);
   U2148 : OAI22_X1 port map( A1 => n13985, A2 => n13399, B1 => n13398, B2 => 
                           n15467, ZN => n7764);
   U2149 : OAI22_X1 port map( A1 => n13991, A2 => n13399, B1 => n13398, B2 => 
                           n15466, ZN => n7765);
   U2150 : OAI22_X1 port map( A1 => n13997, A2 => n13399, B1 => n13398, B2 => 
                           n15465, ZN => n7766);
   U2151 : OAI22_X1 port map( A1 => n14003, A2 => n13399, B1 => n13398, B2 => 
                           n15464, ZN => n7767);
   U2152 : OAI22_X1 port map( A1 => n14009, A2 => n13399, B1 => n13398, B2 => 
                           n15463, ZN => n7768);
   U2153 : OAI22_X1 port map( A1 => n14018, A2 => n13399, B1 => n13398, B2 => 
                           n15462, ZN => n7769);
   U2154 : OAI22_X1 port map( A1 => n13829, A2 => n13419, B1 => n13414, B2 => 
                           n15397, ZN => n7834);
   U2155 : OAI22_X1 port map( A1 => n13835, A2 => n13419, B1 => n13414, B2 => 
                           n15396, ZN => n7835);
   U2156 : OAI22_X1 port map( A1 => n13841, A2 => n13419, B1 => n13414, B2 => 
                           n15395, ZN => n7836);
   U2157 : OAI22_X1 port map( A1 => n13847, A2 => n13419, B1 => n13414, B2 => 
                           n15394, ZN => n7837);
   U2158 : OAI22_X1 port map( A1 => n13853, A2 => n13419, B1 => n13414, B2 => 
                           n15393, ZN => n7838);
   U2159 : OAI22_X1 port map( A1 => n13859, A2 => n13419, B1 => n13414, B2 => 
                           n15392, ZN => n7839);
   U2160 : OAI22_X1 port map( A1 => n13865, A2 => n13419, B1 => n13414, B2 => 
                           n15391, ZN => n7840);
   U2161 : OAI22_X1 port map( A1 => n13871, A2 => n13419, B1 => n13414, B2 => 
                           n15390, ZN => n7841);
   U2162 : OAI22_X1 port map( A1 => n13877, A2 => n13418, B1 => n13414, B2 => 
                           n15389, ZN => n7842);
   U2163 : OAI22_X1 port map( A1 => n13883, A2 => n13418, B1 => n13414, B2 => 
                           n15388, ZN => n7843);
   U2164 : OAI22_X1 port map( A1 => n13889, A2 => n13418, B1 => n13414, B2 => 
                           n15387, ZN => n7844);
   U2165 : OAI22_X1 port map( A1 => n13895, A2 => n13418, B1 => n13414, B2 => 
                           n15386, ZN => n7845);
   U2166 : OAI22_X1 port map( A1 => n13901, A2 => n13418, B1 => n13415, B2 => 
                           n15385, ZN => n7846);
   U2167 : OAI22_X1 port map( A1 => n13907, A2 => n13418, B1 => n13415, B2 => 
                           n15384, ZN => n7847);
   U2168 : OAI22_X1 port map( A1 => n13913, A2 => n13418, B1 => n13415, B2 => 
                           n15383, ZN => n7848);
   U2169 : OAI22_X1 port map( A1 => n13919, A2 => n13418, B1 => n13415, B2 => 
                           n15382, ZN => n7849);
   U2170 : OAI22_X1 port map( A1 => n13925, A2 => n13418, B1 => n13415, B2 => 
                           n15381, ZN => n7850);
   U2171 : OAI22_X1 port map( A1 => n13931, A2 => n13418, B1 => n13415, B2 => 
                           n15380, ZN => n7851);
   U2172 : OAI22_X1 port map( A1 => n13937, A2 => n13418, B1 => n13415, B2 => 
                           n15379, ZN => n7852);
   U2173 : OAI22_X1 port map( A1 => n13943, A2 => n13418, B1 => n13415, B2 => 
                           n15378, ZN => n7853);
   U2174 : OAI22_X1 port map( A1 => n13949, A2 => n13417, B1 => n13415, B2 => 
                           n15377, ZN => n7854);
   U2175 : OAI22_X1 port map( A1 => n13955, A2 => n13417, B1 => n13415, B2 => 
                           n15376, ZN => n7855);
   U2176 : OAI22_X1 port map( A1 => n13961, A2 => n13417, B1 => n13415, B2 => 
                           n15375, ZN => n7856);
   U2177 : OAI22_X1 port map( A1 => n13967, A2 => n13417, B1 => n13415, B2 => 
                           n15374, ZN => n7857);
   U2178 : OAI22_X1 port map( A1 => n13973, A2 => n13417, B1 => n13416, B2 => 
                           n15373, ZN => n7858);
   U2179 : OAI22_X1 port map( A1 => n13979, A2 => n13417, B1 => n13416, B2 => 
                           n15372, ZN => n7859);
   U2180 : OAI22_X1 port map( A1 => n13985, A2 => n13417, B1 => n13416, B2 => 
                           n15371, ZN => n7860);
   U2181 : OAI22_X1 port map( A1 => n13991, A2 => n13417, B1 => n13416, B2 => 
                           n15370, ZN => n7861);
   U2182 : OAI22_X1 port map( A1 => n13997, A2 => n13417, B1 => n13416, B2 => 
                           n15369, ZN => n7862);
   U2183 : OAI22_X1 port map( A1 => n14003, A2 => n13417, B1 => n13416, B2 => 
                           n15368, ZN => n7863);
   U2184 : OAI22_X1 port map( A1 => n14009, A2 => n13417, B1 => n13416, B2 => 
                           n15367, ZN => n7864);
   U2185 : OAI22_X1 port map( A1 => n14018, A2 => n13417, B1 => n13416, B2 => 
                           n15366, ZN => n7865);
   U2186 : OAI22_X1 port map( A1 => n13829, A2 => n13425, B1 => n13420, B2 => 
                           n15365, ZN => n7866);
   U2187 : OAI22_X1 port map( A1 => n13835, A2 => n13425, B1 => n13420, B2 => 
                           n15364, ZN => n7867);
   U2188 : OAI22_X1 port map( A1 => n13841, A2 => n13425, B1 => n13420, B2 => 
                           n15363, ZN => n7868);
   U2189 : OAI22_X1 port map( A1 => n13847, A2 => n13425, B1 => n13420, B2 => 
                           n15362, ZN => n7869);
   U2190 : OAI22_X1 port map( A1 => n13853, A2 => n13425, B1 => n13420, B2 => 
                           n15361, ZN => n7870);
   U2191 : OAI22_X1 port map( A1 => n13859, A2 => n13425, B1 => n13420, B2 => 
                           n15360, ZN => n7871);
   U2192 : OAI22_X1 port map( A1 => n13865, A2 => n13425, B1 => n13420, B2 => 
                           n15359, ZN => n7872);
   U2193 : OAI22_X1 port map( A1 => n13871, A2 => n13425, B1 => n13420, B2 => 
                           n15358, ZN => n7873);
   U2194 : OAI22_X1 port map( A1 => n13877, A2 => n13424, B1 => n13420, B2 => 
                           n15357, ZN => n7874);
   U2195 : OAI22_X1 port map( A1 => n13883, A2 => n13424, B1 => n13420, B2 => 
                           n15356, ZN => n7875);
   U2196 : OAI22_X1 port map( A1 => n13889, A2 => n13424, B1 => n13420, B2 => 
                           n15355, ZN => n7876);
   U2197 : OAI22_X1 port map( A1 => n13895, A2 => n13424, B1 => n13420, B2 => 
                           n15354, ZN => n7877);
   U2198 : OAI22_X1 port map( A1 => n13901, A2 => n13424, B1 => n13421, B2 => 
                           n15353, ZN => n7878);
   U2199 : OAI22_X1 port map( A1 => n13907, A2 => n13424, B1 => n13421, B2 => 
                           n15352, ZN => n7879);
   U2200 : OAI22_X1 port map( A1 => n13913, A2 => n13424, B1 => n13421, B2 => 
                           n15351, ZN => n7880);
   U2201 : OAI22_X1 port map( A1 => n13919, A2 => n13424, B1 => n13421, B2 => 
                           n15350, ZN => n7881);
   U2202 : OAI22_X1 port map( A1 => n13925, A2 => n13424, B1 => n13421, B2 => 
                           n15349, ZN => n7882);
   U2203 : OAI22_X1 port map( A1 => n13931, A2 => n13424, B1 => n13421, B2 => 
                           n15348, ZN => n7883);
   U2204 : OAI22_X1 port map( A1 => n13937, A2 => n13424, B1 => n13421, B2 => 
                           n15347, ZN => n7884);
   U2205 : OAI22_X1 port map( A1 => n13943, A2 => n13424, B1 => n13421, B2 => 
                           n15346, ZN => n7885);
   U2206 : OAI22_X1 port map( A1 => n13949, A2 => n13423, B1 => n13421, B2 => 
                           n15345, ZN => n7886);
   U2207 : OAI22_X1 port map( A1 => n13955, A2 => n13423, B1 => n13421, B2 => 
                           n15344, ZN => n7887);
   U2208 : OAI22_X1 port map( A1 => n13961, A2 => n13423, B1 => n13421, B2 => 
                           n15343, ZN => n7888);
   U2209 : OAI22_X1 port map( A1 => n13967, A2 => n13423, B1 => n13421, B2 => 
                           n15342, ZN => n7889);
   U2210 : OAI22_X1 port map( A1 => n13973, A2 => n13423, B1 => n13422, B2 => 
                           n15341, ZN => n7890);
   U2211 : OAI22_X1 port map( A1 => n13979, A2 => n13423, B1 => n13422, B2 => 
                           n15340, ZN => n7891);
   U2212 : OAI22_X1 port map( A1 => n13985, A2 => n13423, B1 => n13422, B2 => 
                           n15339, ZN => n7892);
   U2213 : OAI22_X1 port map( A1 => n13991, A2 => n13423, B1 => n13422, B2 => 
                           n15338, ZN => n7893);
   U2214 : OAI22_X1 port map( A1 => n13997, A2 => n13423, B1 => n13422, B2 => 
                           n15337, ZN => n7894);
   U2215 : OAI22_X1 port map( A1 => n14003, A2 => n13423, B1 => n13422, B2 => 
                           n15336, ZN => n7895);
   U2216 : OAI22_X1 port map( A1 => n14009, A2 => n13423, B1 => n13422, B2 => 
                           n15335, ZN => n7896);
   U2217 : OAI22_X1 port map( A1 => n14018, A2 => n13423, B1 => n13422, B2 => 
                           n15334, ZN => n7897);
   U2218 : OAI22_X1 port map( A1 => n13968, A2 => n13393, B1 => n13392, B2 => 
                           n15501, ZN => n7730);
   U2219 : OAI22_X1 port map( A1 => n13974, A2 => n13393, B1 => n13392, B2 => 
                           n15500, ZN => n7731);
   U2220 : OAI22_X1 port map( A1 => n13980, A2 => n13393, B1 => n13392, B2 => 
                           n15499, ZN => n7732);
   U2221 : OAI22_X1 port map( A1 => n13986, A2 => n13393, B1 => n13392, B2 => 
                           n15498, ZN => n7733);
   U2222 : OAI22_X1 port map( A1 => n13992, A2 => n13393, B1 => n13392, B2 => 
                           n15497, ZN => n7734);
   U2223 : OAI22_X1 port map( A1 => n13998, A2 => n13393, B1 => n13392, B2 => 
                           n15496, ZN => n7735);
   U2224 : OAI22_X1 port map( A1 => n14004, A2 => n13393, B1 => n13392, B2 => 
                           n15495, ZN => n7736);
   U2225 : OAI22_X1 port map( A1 => n14013, A2 => n13393, B1 => n13392, B2 => 
                           n15494, ZN => n7737);
   U2226 : OAI22_X1 port map( A1 => n13971, A2 => n13525, B1 => n13524, B2 => 
                           n15930, ZN => n8434);
   U2227 : OAI22_X1 port map( A1 => n13977, A2 => n13525, B1 => n13524, B2 => 
                           n15929, ZN => n8435);
   U2228 : OAI22_X1 port map( A1 => n13983, A2 => n13525, B1 => n13524, B2 => 
                           n15928, ZN => n8436);
   U2229 : OAI22_X1 port map( A1 => n13989, A2 => n13525, B1 => n13524, B2 => 
                           n15927, ZN => n8437);
   U2230 : OAI22_X1 port map( A1 => n13995, A2 => n13525, B1 => n13524, B2 => 
                           n15926, ZN => n8438);
   U2231 : OAI22_X1 port map( A1 => n14001, A2 => n13525, B1 => n13524, B2 => 
                           n15925, ZN => n8439);
   U2232 : OAI22_X1 port map( A1 => n14007, A2 => n13525, B1 => n13524, B2 => 
                           n15924, ZN => n8440);
   U2233 : OAI22_X1 port map( A1 => n14016, A2 => n13525, B1 => n13524, B2 => 
                           n15923, ZN => n8441);
   U2234 : OAI22_X1 port map( A1 => n13972, A2 => n13441, B1 => n13440, B2 => 
                           n15277, ZN => n7986);
   U2235 : OAI22_X1 port map( A1 => n13978, A2 => n13441, B1 => n13440, B2 => 
                           n15276, ZN => n7987);
   U2236 : OAI22_X1 port map( A1 => n13984, A2 => n13441, B1 => n13440, B2 => 
                           n15275, ZN => n7988);
   U2237 : OAI22_X1 port map( A1 => n13990, A2 => n13441, B1 => n13440, B2 => 
                           n15274, ZN => n7989);
   U2238 : OAI22_X1 port map( A1 => n13996, A2 => n13441, B1 => n13440, B2 => 
                           n15273, ZN => n7990);
   U2239 : OAI22_X1 port map( A1 => n14002, A2 => n13441, B1 => n13440, B2 => 
                           n15272, ZN => n7991);
   U2240 : OAI22_X1 port map( A1 => n14008, A2 => n13441, B1 => n13440, B2 => 
                           n15271, ZN => n7992);
   U2241 : OAI22_X1 port map( A1 => n14017, A2 => n13441, B1 => n13440, B2 => 
                           n15270, ZN => n7993);
   U2242 : OAI22_X1 port map( A1 => n13972, A2 => n13447, B1 => n13446, B2 => 
                           n15245, ZN => n8018);
   U2243 : OAI22_X1 port map( A1 => n13978, A2 => n13447, B1 => n13446, B2 => 
                           n15244, ZN => n8019);
   U2244 : OAI22_X1 port map( A1 => n13984, A2 => n13447, B1 => n13446, B2 => 
                           n15243, ZN => n8020);
   U2245 : OAI22_X1 port map( A1 => n13990, A2 => n13447, B1 => n13446, B2 => 
                           n15242, ZN => n8021);
   U2246 : OAI22_X1 port map( A1 => n13996, A2 => n13447, B1 => n13446, B2 => 
                           n15241, ZN => n8022);
   U2247 : OAI22_X1 port map( A1 => n14002, A2 => n13447, B1 => n13446, B2 => 
                           n15240, ZN => n8023);
   U2248 : OAI22_X1 port map( A1 => n14008, A2 => n13447, B1 => n13446, B2 => 
                           n15239, ZN => n8024);
   U2249 : OAI22_X1 port map( A1 => n14017, A2 => n13447, B1 => n13446, B2 => 
                           n15238, ZN => n8025);
   U2250 : OAI22_X1 port map( A1 => n13972, A2 => n13453, B1 => n13452, B2 => 
                           n15213, ZN => n8050);
   U2251 : OAI22_X1 port map( A1 => n13978, A2 => n13453, B1 => n13452, B2 => 
                           n15212, ZN => n8051);
   U2252 : OAI22_X1 port map( A1 => n13984, A2 => n13453, B1 => n13452, B2 => 
                           n15211, ZN => n8052);
   U2253 : OAI22_X1 port map( A1 => n13990, A2 => n13453, B1 => n13452, B2 => 
                           n15210, ZN => n8053);
   U2254 : OAI22_X1 port map( A1 => n13996, A2 => n13453, B1 => n13452, B2 => 
                           n15209, ZN => n8054);
   U2255 : OAI22_X1 port map( A1 => n14002, A2 => n13453, B1 => n13452, B2 => 
                           n15208, ZN => n8055);
   U2256 : OAI22_X1 port map( A1 => n14008, A2 => n13453, B1 => n13452, B2 => 
                           n15207, ZN => n8056);
   U2257 : OAI22_X1 port map( A1 => n14017, A2 => n13453, B1 => n13452, B2 => 
                           n15206, ZN => n8057);
   U2258 : OAI22_X1 port map( A1 => n13972, A2 => n13483, B1 => n13482, B2 => 
                           n15149, ZN => n8210);
   U2259 : OAI22_X1 port map( A1 => n13978, A2 => n13483, B1 => n13482, B2 => 
                           n15148, ZN => n8211);
   U2260 : OAI22_X1 port map( A1 => n13984, A2 => n13483, B1 => n13482, B2 => 
                           n15147, ZN => n8212);
   U2261 : OAI22_X1 port map( A1 => n13990, A2 => n13483, B1 => n13482, B2 => 
                           n15146, ZN => n8213);
   U2262 : OAI22_X1 port map( A1 => n13996, A2 => n13483, B1 => n13482, B2 => 
                           n15145, ZN => n8214);
   U2263 : OAI22_X1 port map( A1 => n14002, A2 => n13483, B1 => n13482, B2 => 
                           n15144, ZN => n8215);
   U2264 : OAI22_X1 port map( A1 => n14008, A2 => n13483, B1 => n13482, B2 => 
                           n15143, ZN => n8216);
   U2265 : OAI22_X1 port map( A1 => n14017, A2 => n13483, B1 => n13482, B2 => 
                           n15142, ZN => n8217);
   U2266 : OAI22_X1 port map( A1 => n13972, A2 => n13489, B1 => n13488, B2 => 
                           n15117, ZN => n8242);
   U2267 : OAI22_X1 port map( A1 => n13978, A2 => n13489, B1 => n13488, B2 => 
                           n15116, ZN => n8243);
   U2268 : OAI22_X1 port map( A1 => n13984, A2 => n13489, B1 => n13488, B2 => 
                           n15115, ZN => n8244);
   U2269 : OAI22_X1 port map( A1 => n13990, A2 => n13489, B1 => n13488, B2 => 
                           n15114, ZN => n8245);
   U2270 : OAI22_X1 port map( A1 => n13996, A2 => n13489, B1 => n13488, B2 => 
                           n15113, ZN => n8246);
   U2271 : OAI22_X1 port map( A1 => n14002, A2 => n13489, B1 => n13488, B2 => 
                           n15112, ZN => n8247);
   U2272 : OAI22_X1 port map( A1 => n14008, A2 => n13489, B1 => n13488, B2 => 
                           n15111, ZN => n8248);
   U2273 : OAI22_X1 port map( A1 => n14017, A2 => n13489, B1 => n13488, B2 => 
                           n15110, ZN => n8249);
   U2274 : OAI22_X1 port map( A1 => n13972, A2 => n13495, B1 => n13494, B2 => 
                           n15085, ZN => n8274);
   U2275 : OAI22_X1 port map( A1 => n13978, A2 => n13495, B1 => n13494, B2 => 
                           n15084, ZN => n8275);
   U2276 : OAI22_X1 port map( A1 => n13984, A2 => n13495, B1 => n13494, B2 => 
                           n15083, ZN => n8276);
   U2277 : OAI22_X1 port map( A1 => n13990, A2 => n13495, B1 => n13494, B2 => 
                           n15082, ZN => n8277);
   U2278 : OAI22_X1 port map( A1 => n13996, A2 => n13495, B1 => n13494, B2 => 
                           n15081, ZN => n8278);
   U2279 : OAI22_X1 port map( A1 => n14002, A2 => n13495, B1 => n13494, B2 => 
                           n15080, ZN => n8279);
   U2280 : OAI22_X1 port map( A1 => n14008, A2 => n13495, B1 => n13494, B2 => 
                           n15079, ZN => n8280);
   U2281 : OAI22_X1 port map( A1 => n14017, A2 => n13495, B1 => n13494, B2 => 
                           n15078, ZN => n8281);
   U2282 : OAI22_X1 port map( A1 => n13972, A2 => n13501, B1 => n13500, B2 => 
                           n15053, ZN => n8306);
   U2283 : OAI22_X1 port map( A1 => n13978, A2 => n13501, B1 => n13500, B2 => 
                           n15052, ZN => n8307);
   U2284 : OAI22_X1 port map( A1 => n13984, A2 => n13501, B1 => n13500, B2 => 
                           n15051, ZN => n8308);
   U2285 : OAI22_X1 port map( A1 => n13990, A2 => n13501, B1 => n13500, B2 => 
                           n15050, ZN => n8309);
   U2286 : OAI22_X1 port map( A1 => n13996, A2 => n13501, B1 => n13500, B2 => 
                           n15049, ZN => n8310);
   U2287 : OAI22_X1 port map( A1 => n14002, A2 => n13501, B1 => n13500, B2 => 
                           n15048, ZN => n8311);
   U2288 : OAI22_X1 port map( A1 => n14008, A2 => n13501, B1 => n13500, B2 => 
                           n15047, ZN => n8312);
   U2289 : OAI22_X1 port map( A1 => n14017, A2 => n13501, B1 => n13500, B2 => 
                           n15046, ZN => n8313);
   U2290 : OAI22_X1 port map( A1 => n13972, A2 => n13507, B1 => n13506, B2 => 
                           n15021, ZN => n8338);
   U2291 : OAI22_X1 port map( A1 => n13978, A2 => n13507, B1 => n13506, B2 => 
                           n15020, ZN => n8339);
   U2292 : OAI22_X1 port map( A1 => n13984, A2 => n13507, B1 => n13506, B2 => 
                           n15019, ZN => n8340);
   U2293 : OAI22_X1 port map( A1 => n13990, A2 => n13507, B1 => n13506, B2 => 
                           n15018, ZN => n8341);
   U2294 : OAI22_X1 port map( A1 => n13996, A2 => n13507, B1 => n13506, B2 => 
                           n15017, ZN => n8342);
   U2295 : OAI22_X1 port map( A1 => n14002, A2 => n13507, B1 => n13506, B2 => 
                           n15016, ZN => n8343);
   U2296 : OAI22_X1 port map( A1 => n14008, A2 => n13507, B1 => n13506, B2 => 
                           n15015, ZN => n8344);
   U2297 : OAI22_X1 port map( A1 => n14017, A2 => n13507, B1 => n13506, B2 => 
                           n15014, ZN => n8345);
   U2298 : OAI22_X1 port map( A1 => n13971, A2 => n13531, B1 => n13530, B2 => 
                           n14956, ZN => n8466);
   U2299 : OAI22_X1 port map( A1 => n13977, A2 => n13531, B1 => n13530, B2 => 
                           n14955, ZN => n8467);
   U2300 : OAI22_X1 port map( A1 => n13983, A2 => n13531, B1 => n13530, B2 => 
                           n14954, ZN => n8468);
   U2301 : OAI22_X1 port map( A1 => n13989, A2 => n13531, B1 => n13530, B2 => 
                           n14953, ZN => n8469);
   U2302 : OAI22_X1 port map( A1 => n13995, A2 => n13531, B1 => n13530, B2 => 
                           n14952, ZN => n8470);
   U2303 : OAI22_X1 port map( A1 => n14001, A2 => n13531, B1 => n13530, B2 => 
                           n14951, ZN => n8471);
   U2304 : OAI22_X1 port map( A1 => n14007, A2 => n13531, B1 => n13530, B2 => 
                           n14950, ZN => n8472);
   U2305 : OAI22_X1 port map( A1 => n14016, A2 => n13531, B1 => n13530, B2 => 
                           n14949, ZN => n8473);
   U2306 : OAI22_X1 port map( A1 => n13971, A2 => n13549, B1 => n13548, B2 => 
                           n14923, ZN => n8562);
   U2307 : OAI22_X1 port map( A1 => n13977, A2 => n13549, B1 => n13548, B2 => 
                           n14922, ZN => n8563);
   U2308 : OAI22_X1 port map( A1 => n13983, A2 => n13549, B1 => n13548, B2 => 
                           n14921, ZN => n8564);
   U2309 : OAI22_X1 port map( A1 => n13989, A2 => n13549, B1 => n13548, B2 => 
                           n14920, ZN => n8565);
   U2310 : OAI22_X1 port map( A1 => n13995, A2 => n13549, B1 => n13548, B2 => 
                           n14919, ZN => n8566);
   U2311 : OAI22_X1 port map( A1 => n14001, A2 => n13549, B1 => n13548, B2 => 
                           n14918, ZN => n8567);
   U2312 : OAI22_X1 port map( A1 => n14007, A2 => n13549, B1 => n13548, B2 => 
                           n14917, ZN => n8568);
   U2313 : OAI22_X1 port map( A1 => n14016, A2 => n13549, B1 => n13548, B2 => 
                           n14916, ZN => n8569);
   U2314 : OAI22_X1 port map( A1 => n13971, A2 => n13555, B1 => n13554, B2 => 
                           n14891, ZN => n8594);
   U2315 : OAI22_X1 port map( A1 => n13977, A2 => n13555, B1 => n13554, B2 => 
                           n14890, ZN => n8595);
   U2316 : OAI22_X1 port map( A1 => n13983, A2 => n13555, B1 => n13554, B2 => 
                           n14889, ZN => n8596);
   U2317 : OAI22_X1 port map( A1 => n13989, A2 => n13555, B1 => n13554, B2 => 
                           n14888, ZN => n8597);
   U2318 : OAI22_X1 port map( A1 => n13995, A2 => n13555, B1 => n13554, B2 => 
                           n14887, ZN => n8598);
   U2319 : OAI22_X1 port map( A1 => n14001, A2 => n13555, B1 => n13554, B2 => 
                           n14886, ZN => n8599);
   U2320 : OAI22_X1 port map( A1 => n14007, A2 => n13555, B1 => n13554, B2 => 
                           n14885, ZN => n8600);
   U2321 : OAI22_X1 port map( A1 => n14016, A2 => n13555, B1 => n13554, B2 => 
                           n14884, ZN => n8601);
   U2322 : OAI22_X1 port map( A1 => n13971, A2 => n13561, B1 => n13560, B2 => 
                           n14859, ZN => n8626);
   U2323 : OAI22_X1 port map( A1 => n13977, A2 => n13561, B1 => n13560, B2 => 
                           n14858, ZN => n8627);
   U2324 : OAI22_X1 port map( A1 => n13983, A2 => n13561, B1 => n13560, B2 => 
                           n14857, ZN => n8628);
   U2325 : OAI22_X1 port map( A1 => n13989, A2 => n13561, B1 => n13560, B2 => 
                           n14856, ZN => n8629);
   U2326 : OAI22_X1 port map( A1 => n13995, A2 => n13561, B1 => n13560, B2 => 
                           n14855, ZN => n8630);
   U2327 : OAI22_X1 port map( A1 => n14001, A2 => n13561, B1 => n13560, B2 => 
                           n14854, ZN => n8631);
   U2328 : OAI22_X1 port map( A1 => n14007, A2 => n13561, B1 => n13560, B2 => 
                           n14853, ZN => n8632);
   U2329 : OAI22_X1 port map( A1 => n14016, A2 => n13561, B1 => n13560, B2 => 
                           n14852, ZN => n8633);
   U2330 : OAI22_X1 port map( A1 => n13971, A2 => n13591, B1 => n13590, B2 => 
                           n14827, ZN => n8786);
   U2331 : OAI22_X1 port map( A1 => n13977, A2 => n13591, B1 => n13590, B2 => 
                           n14826, ZN => n8787);
   U2332 : OAI22_X1 port map( A1 => n13983, A2 => n13591, B1 => n13590, B2 => 
                           n14825, ZN => n8788);
   U2333 : OAI22_X1 port map( A1 => n13989, A2 => n13591, B1 => n13590, B2 => 
                           n14824, ZN => n8789);
   U2334 : OAI22_X1 port map( A1 => n13995, A2 => n13591, B1 => n13590, B2 => 
                           n14823, ZN => n8790);
   U2335 : OAI22_X1 port map( A1 => n14001, A2 => n13591, B1 => n13590, B2 => 
                           n14822, ZN => n8791);
   U2336 : OAI22_X1 port map( A1 => n14007, A2 => n13591, B1 => n13590, B2 => 
                           n14821, ZN => n8792);
   U2337 : OAI22_X1 port map( A1 => n14016, A2 => n13591, B1 => n13590, B2 => 
                           n14820, ZN => n8793);
   U2338 : OAI22_X1 port map( A1 => n13970, A2 => n13597, B1 => n13596, B2 => 
                           n14795, ZN => n8818);
   U2339 : OAI22_X1 port map( A1 => n13976, A2 => n13597, B1 => n13596, B2 => 
                           n14794, ZN => n8819);
   U2340 : OAI22_X1 port map( A1 => n13982, A2 => n13597, B1 => n13596, B2 => 
                           n14793, ZN => n8820);
   U2341 : OAI22_X1 port map( A1 => n13988, A2 => n13597, B1 => n13596, B2 => 
                           n14792, ZN => n8821);
   U2342 : OAI22_X1 port map( A1 => n13994, A2 => n13597, B1 => n13596, B2 => 
                           n14791, ZN => n8822);
   U2343 : OAI22_X1 port map( A1 => n14000, A2 => n13597, B1 => n13596, B2 => 
                           n14790, ZN => n8823);
   U2344 : OAI22_X1 port map( A1 => n14006, A2 => n13597, B1 => n13596, B2 => 
                           n14789, ZN => n8824);
   U2345 : OAI22_X1 port map( A1 => n14015, A2 => n13597, B1 => n13596, B2 => 
                           n14788, ZN => n8825);
   U2346 : OAI22_X1 port map( A1 => n13970, A2 => n13603, B1 => n13602, B2 => 
                           n14763, ZN => n8850);
   U2347 : OAI22_X1 port map( A1 => n13976, A2 => n13603, B1 => n13602, B2 => 
                           n14762, ZN => n8851);
   U2348 : OAI22_X1 port map( A1 => n13982, A2 => n13603, B1 => n13602, B2 => 
                           n14761, ZN => n8852);
   U2349 : OAI22_X1 port map( A1 => n13988, A2 => n13603, B1 => n13602, B2 => 
                           n14760, ZN => n8853);
   U2350 : OAI22_X1 port map( A1 => n13994, A2 => n13603, B1 => n13602, B2 => 
                           n14759, ZN => n8854);
   U2351 : OAI22_X1 port map( A1 => n14000, A2 => n13603, B1 => n13602, B2 => 
                           n14758, ZN => n8855);
   U2352 : OAI22_X1 port map( A1 => n14006, A2 => n13603, B1 => n13602, B2 => 
                           n14757, ZN => n8856);
   U2353 : OAI22_X1 port map( A1 => n14015, A2 => n13603, B1 => n13602, B2 => 
                           n14756, ZN => n8857);
   U2354 : OAI22_X1 port map( A1 => n13970, A2 => n13609, B1 => n13608, B2 => 
                           n14731, ZN => n8882);
   U2355 : OAI22_X1 port map( A1 => n13976, A2 => n13609, B1 => n13608, B2 => 
                           n14730, ZN => n8883);
   U2356 : OAI22_X1 port map( A1 => n13982, A2 => n13609, B1 => n13608, B2 => 
                           n14729, ZN => n8884);
   U2357 : OAI22_X1 port map( A1 => n13988, A2 => n13609, B1 => n13608, B2 => 
                           n14728, ZN => n8885);
   U2358 : OAI22_X1 port map( A1 => n13994, A2 => n13609, B1 => n13608, B2 => 
                           n14727, ZN => n8886);
   U2359 : OAI22_X1 port map( A1 => n14000, A2 => n13609, B1 => n13608, B2 => 
                           n14726, ZN => n8887);
   U2360 : OAI22_X1 port map( A1 => n14006, A2 => n13609, B1 => n13608, B2 => 
                           n14725, ZN => n8888);
   U2361 : OAI22_X1 port map( A1 => n14015, A2 => n13609, B1 => n13608, B2 => 
                           n14724, ZN => n8889);
   U2362 : OAI22_X1 port map( A1 => n13970, A2 => n13615, B1 => n13614, B2 => 
                           n14699, ZN => n8914);
   U2363 : OAI22_X1 port map( A1 => n13976, A2 => n13615, B1 => n13614, B2 => 
                           n14698, ZN => n8915);
   U2364 : OAI22_X1 port map( A1 => n13982, A2 => n13615, B1 => n13614, B2 => 
                           n14697, ZN => n8916);
   U2365 : OAI22_X1 port map( A1 => n13988, A2 => n13615, B1 => n13614, B2 => 
                           n14696, ZN => n8917);
   U2366 : OAI22_X1 port map( A1 => n13994, A2 => n13615, B1 => n13614, B2 => 
                           n14695, ZN => n8918);
   U2367 : OAI22_X1 port map( A1 => n14000, A2 => n13615, B1 => n13614, B2 => 
                           n14694, ZN => n8919);
   U2368 : OAI22_X1 port map( A1 => n14006, A2 => n13615, B1 => n13614, B2 => 
                           n14693, ZN => n8920);
   U2369 : OAI22_X1 port map( A1 => n14015, A2 => n13615, B1 => n13614, B2 => 
                           n14692, ZN => n8921);
   U2370 : OAI22_X1 port map( A1 => n13970, A2 => n13645, B1 => n13644, B2 => 
                           n14628, ZN => n9074);
   U2371 : OAI22_X1 port map( A1 => n13976, A2 => n13645, B1 => n13644, B2 => 
                           n14627, ZN => n9075);
   U2372 : OAI22_X1 port map( A1 => n13982, A2 => n13645, B1 => n13644, B2 => 
                           n14626, ZN => n9076);
   U2373 : OAI22_X1 port map( A1 => n13988, A2 => n13645, B1 => n13644, B2 => 
                           n14625, ZN => n9077);
   U2374 : OAI22_X1 port map( A1 => n13994, A2 => n13645, B1 => n13644, B2 => 
                           n14624, ZN => n9078);
   U2375 : OAI22_X1 port map( A1 => n14000, A2 => n13645, B1 => n13644, B2 => 
                           n14623, ZN => n9079);
   U2376 : OAI22_X1 port map( A1 => n14006, A2 => n13645, B1 => n13644, B2 => 
                           n14622, ZN => n9080);
   U2377 : OAI22_X1 port map( A1 => n14015, A2 => n13645, B1 => n13644, B2 => 
                           n14621, ZN => n9081);
   U2378 : OAI22_X1 port map( A1 => n13970, A2 => n13651, B1 => n13650, B2 => 
                           n14596, ZN => n9106);
   U2379 : OAI22_X1 port map( A1 => n13976, A2 => n13651, B1 => n13650, B2 => 
                           n14595, ZN => n9107);
   U2380 : OAI22_X1 port map( A1 => n13982, A2 => n13651, B1 => n13650, B2 => 
                           n14594, ZN => n9108);
   U2381 : OAI22_X1 port map( A1 => n13988, A2 => n13651, B1 => n13650, B2 => 
                           n14593, ZN => n9109);
   U2382 : OAI22_X1 port map( A1 => n13994, A2 => n13651, B1 => n13650, B2 => 
                           n14592, ZN => n9110);
   U2383 : OAI22_X1 port map( A1 => n14000, A2 => n13651, B1 => n13650, B2 => 
                           n14591, ZN => n9111);
   U2384 : OAI22_X1 port map( A1 => n14006, A2 => n13651, B1 => n13650, B2 => 
                           n14590, ZN => n9112);
   U2385 : OAI22_X1 port map( A1 => n14015, A2 => n13651, B1 => n13650, B2 => 
                           n14589, ZN => n9113);
   U2386 : OAI22_X1 port map( A1 => n13970, A2 => n13657, B1 => n13656, B2 => 
                           n14564, ZN => n9138);
   U2387 : OAI22_X1 port map( A1 => n13976, A2 => n13657, B1 => n13656, B2 => 
                           n14563, ZN => n9139);
   U2388 : OAI22_X1 port map( A1 => n13982, A2 => n13657, B1 => n13656, B2 => 
                           n14562, ZN => n9140);
   U2389 : OAI22_X1 port map( A1 => n13988, A2 => n13657, B1 => n13656, B2 => 
                           n14561, ZN => n9141);
   U2390 : OAI22_X1 port map( A1 => n13994, A2 => n13657, B1 => n13656, B2 => 
                           n14560, ZN => n9142);
   U2391 : OAI22_X1 port map( A1 => n14000, A2 => n13657, B1 => n13656, B2 => 
                           n14559, ZN => n9143);
   U2392 : OAI22_X1 port map( A1 => n14006, A2 => n13657, B1 => n13656, B2 => 
                           n14558, ZN => n9144);
   U2393 : OAI22_X1 port map( A1 => n14015, A2 => n13657, B1 => n13656, B2 => 
                           n14557, ZN => n9145);
   U2394 : OAI22_X1 port map( A1 => n13970, A2 => n13663, B1 => n13662, B2 => 
                           n14532, ZN => n9170);
   U2395 : OAI22_X1 port map( A1 => n13976, A2 => n13663, B1 => n13662, B2 => 
                           n14531, ZN => n9171);
   U2396 : OAI22_X1 port map( A1 => n13982, A2 => n13663, B1 => n13662, B2 => 
                           n14530, ZN => n9172);
   U2397 : OAI22_X1 port map( A1 => n13988, A2 => n13663, B1 => n13662, B2 => 
                           n14529, ZN => n9173);
   U2398 : OAI22_X1 port map( A1 => n13994, A2 => n13663, B1 => n13662, B2 => 
                           n14528, ZN => n9174);
   U2399 : OAI22_X1 port map( A1 => n14000, A2 => n13663, B1 => n13662, B2 => 
                           n14527, ZN => n9175);
   U2400 : OAI22_X1 port map( A1 => n14006, A2 => n13663, B1 => n13662, B2 => 
                           n14526, ZN => n9176);
   U2401 : OAI22_X1 port map( A1 => n14015, A2 => n13663, B1 => n13662, B2 => 
                           n14525, ZN => n9177);
   U2402 : OAI22_X1 port map( A1 => n13969, A2 => n13669, B1 => n13668, B2 => 
                           n14500, ZN => n9202);
   U2403 : OAI22_X1 port map( A1 => n13975, A2 => n13669, B1 => n13668, B2 => 
                           n14499, ZN => n9203);
   U2404 : OAI22_X1 port map( A1 => n13981, A2 => n13669, B1 => n13668, B2 => 
                           n14498, ZN => n9204);
   U2405 : OAI22_X1 port map( A1 => n13987, A2 => n13669, B1 => n13668, B2 => 
                           n14497, ZN => n9205);
   U2406 : OAI22_X1 port map( A1 => n13993, A2 => n13669, B1 => n13668, B2 => 
                           n14496, ZN => n9206);
   U2407 : OAI22_X1 port map( A1 => n13999, A2 => n13669, B1 => n13668, B2 => 
                           n14495, ZN => n9207);
   U2408 : OAI22_X1 port map( A1 => n14005, A2 => n13669, B1 => n13668, B2 => 
                           n14494, ZN => n9208);
   U2409 : OAI22_X1 port map( A1 => n14014, A2 => n13669, B1 => n13668, B2 => 
                           n14493, ZN => n9209);
   U2410 : OAI22_X1 port map( A1 => n13969, A2 => n13699, B1 => n13698, B2 => 
                           n14415, ZN => n9362);
   U2411 : OAI22_X1 port map( A1 => n13975, A2 => n13699, B1 => n13698, B2 => 
                           n14414, ZN => n9363);
   U2412 : OAI22_X1 port map( A1 => n13981, A2 => n13699, B1 => n13698, B2 => 
                           n14413, ZN => n9364);
   U2413 : OAI22_X1 port map( A1 => n13987, A2 => n13699, B1 => n13698, B2 => 
                           n14412, ZN => n9365);
   U2414 : OAI22_X1 port map( A1 => n13993, A2 => n13699, B1 => n13698, B2 => 
                           n14411, ZN => n9366);
   U2415 : OAI22_X1 port map( A1 => n13999, A2 => n13699, B1 => n13698, B2 => 
                           n14410, ZN => n9367);
   U2416 : OAI22_X1 port map( A1 => n14005, A2 => n13699, B1 => n13698, B2 => 
                           n14409, ZN => n9368);
   U2417 : OAI22_X1 port map( A1 => n14014, A2 => n13699, B1 => n13698, B2 => 
                           n14408, ZN => n9369);
   U2418 : OAI22_X1 port map( A1 => n13970, A2 => n13705, B1 => n13704, B2 => 
                           n14383, ZN => n9394);
   U2419 : OAI22_X1 port map( A1 => n13976, A2 => n13705, B1 => n13704, B2 => 
                           n14382, ZN => n9395);
   U2420 : OAI22_X1 port map( A1 => n13982, A2 => n13705, B1 => n13704, B2 => 
                           n14381, ZN => n9396);
   U2421 : OAI22_X1 port map( A1 => n13988, A2 => n13705, B1 => n13704, B2 => 
                           n14380, ZN => n9397);
   U2422 : OAI22_X1 port map( A1 => n13994, A2 => n13705, B1 => n13704, B2 => 
                           n14379, ZN => n9398);
   U2423 : OAI22_X1 port map( A1 => n14000, A2 => n13705, B1 => n13704, B2 => 
                           n14378, ZN => n9399);
   U2424 : OAI22_X1 port map( A1 => n14006, A2 => n13705, B1 => n13704, B2 => 
                           n14377, ZN => n9400);
   U2425 : OAI22_X1 port map( A1 => n14015, A2 => n13705, B1 => n13704, B2 => 
                           n14376, ZN => n9401);
   U2426 : OAI22_X1 port map( A1 => n13969, A2 => n13711, B1 => n13710, B2 => 
                           n14351, ZN => n9426);
   U2427 : OAI22_X1 port map( A1 => n13975, A2 => n13711, B1 => n13710, B2 => 
                           n14350, ZN => n9427);
   U2428 : OAI22_X1 port map( A1 => n13981, A2 => n13711, B1 => n13710, B2 => 
                           n14349, ZN => n9428);
   U2429 : OAI22_X1 port map( A1 => n13987, A2 => n13711, B1 => n13710, B2 => 
                           n14348, ZN => n9429);
   U2430 : OAI22_X1 port map( A1 => n13993, A2 => n13711, B1 => n13710, B2 => 
                           n14347, ZN => n9430);
   U2431 : OAI22_X1 port map( A1 => n13999, A2 => n13711, B1 => n13710, B2 => 
                           n14346, ZN => n9431);
   U2432 : OAI22_X1 port map( A1 => n14005, A2 => n13711, B1 => n13710, B2 => 
                           n14345, ZN => n9432);
   U2433 : OAI22_X1 port map( A1 => n14014, A2 => n13711, B1 => n13710, B2 => 
                           n14344, ZN => n9433);
   U2434 : OAI22_X1 port map( A1 => n13969, A2 => n13717, B1 => n13716, B2 => 
                           n14319, ZN => n9458);
   U2435 : OAI22_X1 port map( A1 => n13975, A2 => n13717, B1 => n13716, B2 => 
                           n14318, ZN => n9459);
   U2436 : OAI22_X1 port map( A1 => n13981, A2 => n13717, B1 => n13716, B2 => 
                           n14317, ZN => n9460);
   U2437 : OAI22_X1 port map( A1 => n13987, A2 => n13717, B1 => n13716, B2 => 
                           n14316, ZN => n9461);
   U2438 : OAI22_X1 port map( A1 => n13993, A2 => n13717, B1 => n13716, B2 => 
                           n14315, ZN => n9462);
   U2439 : OAI22_X1 port map( A1 => n13999, A2 => n13717, B1 => n13716, B2 => 
                           n14314, ZN => n9463);
   U2440 : OAI22_X1 port map( A1 => n14005, A2 => n13717, B1 => n13716, B2 => 
                           n14313, ZN => n9464);
   U2441 : OAI22_X1 port map( A1 => n14014, A2 => n13717, B1 => n13716, B2 => 
                           n14312, ZN => n9465);
   U2442 : OAI22_X1 port map( A1 => n13969, A2 => n13723, B1 => n13722, B2 => 
                           n14287, ZN => n9490);
   U2443 : OAI22_X1 port map( A1 => n13975, A2 => n13723, B1 => n13722, B2 => 
                           n14286, ZN => n9491);
   U2444 : OAI22_X1 port map( A1 => n13981, A2 => n13723, B1 => n13722, B2 => 
                           n14285, ZN => n9492);
   U2445 : OAI22_X1 port map( A1 => n13987, A2 => n13723, B1 => n13722, B2 => 
                           n14284, ZN => n9493);
   U2446 : OAI22_X1 port map( A1 => n13993, A2 => n13723, B1 => n13722, B2 => 
                           n14283, ZN => n9494);
   U2447 : OAI22_X1 port map( A1 => n13999, A2 => n13723, B1 => n13722, B2 => 
                           n14282, ZN => n9495);
   U2448 : OAI22_X1 port map( A1 => n14005, A2 => n13723, B1 => n13722, B2 => 
                           n14281, ZN => n9496);
   U2449 : OAI22_X1 port map( A1 => n14014, A2 => n13723, B1 => n13722, B2 => 
                           n14280, ZN => n9497);
   U2450 : OAI22_X1 port map( A1 => n13968, A2 => n13747, B1 => n13746, B2 => 
                           n12657, ZN => n9618);
   U2451 : OAI22_X1 port map( A1 => n13974, A2 => n13747, B1 => n13746, B2 => 
                           n12658, ZN => n9619);
   U2452 : OAI22_X1 port map( A1 => n13980, A2 => n13747, B1 => n13746, B2 => 
                           n12659, ZN => n9620);
   U2453 : OAI22_X1 port map( A1 => n13986, A2 => n13747, B1 => n13746, B2 => 
                           n12660, ZN => n9621);
   U2454 : OAI22_X1 port map( A1 => n13992, A2 => n13747, B1 => n13746, B2 => 
                           n12653, ZN => n9622);
   U2455 : OAI22_X1 port map( A1 => n13998, A2 => n13747, B1 => n13746, B2 => 
                           n12654, ZN => n9623);
   U2456 : OAI22_X1 port map( A1 => n14004, A2 => n13747, B1 => n13746, B2 => 
                           n12655, ZN => n9624);
   U2457 : OAI22_X1 port map( A1 => n14013, A2 => n13747, B1 => n13746, B2 => 
                           n12656, ZN => n9625);
   U2458 : OAI22_X1 port map( A1 => n13968, A2 => n13765, B1 => n13764, B2 => 
                           n14179, ZN => n9714);
   U2459 : OAI22_X1 port map( A1 => n13974, A2 => n13765, B1 => n13764, B2 => 
                           n14178, ZN => n9715);
   U2460 : OAI22_X1 port map( A1 => n13980, A2 => n13765, B1 => n13764, B2 => 
                           n14177, ZN => n9716);
   U2461 : OAI22_X1 port map( A1 => n13986, A2 => n13765, B1 => n13764, B2 => 
                           n14176, ZN => n9717);
   U2462 : OAI22_X1 port map( A1 => n13992, A2 => n13765, B1 => n13764, B2 => 
                           n14175, ZN => n9718);
   U2463 : OAI22_X1 port map( A1 => n13998, A2 => n13765, B1 => n13764, B2 => 
                           n14174, ZN => n9719);
   U2464 : OAI22_X1 port map( A1 => n14004, A2 => n13765, B1 => n13764, B2 => 
                           n14173, ZN => n9720);
   U2465 : OAI22_X1 port map( A1 => n14013, A2 => n13765, B1 => n13764, B2 => 
                           n14172, ZN => n9721);
   U2466 : OAI22_X1 port map( A1 => n13968, A2 => n13771, B1 => n13770, B2 => 
                           n14147, ZN => n9746);
   U2467 : OAI22_X1 port map( A1 => n13974, A2 => n13771, B1 => n13770, B2 => 
                           n14146, ZN => n9747);
   U2468 : OAI22_X1 port map( A1 => n13980, A2 => n13771, B1 => n13770, B2 => 
                           n14145, ZN => n9748);
   U2469 : OAI22_X1 port map( A1 => n13986, A2 => n13771, B1 => n13770, B2 => 
                           n14144, ZN => n9749);
   U2470 : OAI22_X1 port map( A1 => n13992, A2 => n13771, B1 => n13770, B2 => 
                           n14143, ZN => n9750);
   U2471 : OAI22_X1 port map( A1 => n13998, A2 => n13771, B1 => n13770, B2 => 
                           n14142, ZN => n9751);
   U2472 : OAI22_X1 port map( A1 => n14004, A2 => n13771, B1 => n13770, B2 => 
                           n14141, ZN => n9752);
   U2473 : OAI22_X1 port map( A1 => n14013, A2 => n13771, B1 => n13770, B2 => 
                           n14140, ZN => n9753);
   U2474 : OAI22_X1 port map( A1 => n13968, A2 => n13777, B1 => n13776, B2 => 
                           n14115, ZN => n9778);
   U2475 : OAI22_X1 port map( A1 => n13974, A2 => n13777, B1 => n13776, B2 => 
                           n14114, ZN => n9779);
   U2476 : OAI22_X1 port map( A1 => n13980, A2 => n13777, B1 => n13776, B2 => 
                           n14113, ZN => n9780);
   U2477 : OAI22_X1 port map( A1 => n13986, A2 => n13777, B1 => n13776, B2 => 
                           n14112, ZN => n9781);
   U2478 : OAI22_X1 port map( A1 => n13992, A2 => n13777, B1 => n13776, B2 => 
                           n14111, ZN => n9782);
   U2479 : OAI22_X1 port map( A1 => n13998, A2 => n13777, B1 => n13776, B2 => 
                           n14110, ZN => n9783);
   U2480 : OAI22_X1 port map( A1 => n14004, A2 => n13777, B1 => n13776, B2 => 
                           n14109, ZN => n9784);
   U2481 : OAI22_X1 port map( A1 => n14013, A2 => n13777, B1 => n13776, B2 => 
                           n14108, ZN => n9785);
   U2482 : OAI22_X1 port map( A1 => n13968, A2 => n13801, B1 => n13800, B2 => 
                           n12649, ZN => n9906);
   U2483 : OAI22_X1 port map( A1 => n13974, A2 => n13801, B1 => n13800, B2 => 
                           n12650, ZN => n9907);
   U2484 : OAI22_X1 port map( A1 => n13980, A2 => n13801, B1 => n13800, B2 => 
                           n12651, ZN => n9908);
   U2485 : OAI22_X1 port map( A1 => n13986, A2 => n13801, B1 => n13800, B2 => 
                           n12652, ZN => n9909);
   U2486 : OAI22_X1 port map( A1 => n13992, A2 => n13801, B1 => n13800, B2 => 
                           n12645, ZN => n9910);
   U2487 : OAI22_X1 port map( A1 => n13998, A2 => n13801, B1 => n13800, B2 => 
                           n12646, ZN => n9911);
   U2488 : OAI22_X1 port map( A1 => n14004, A2 => n13801, B1 => n13800, B2 => 
                           n12647, ZN => n9912);
   U2489 : OAI22_X1 port map( A1 => n14013, A2 => n13801, B1 => n13800, B2 => 
                           n12648, ZN => n9913);
   U2490 : OAI22_X1 port map( A1 => n13387, A2 => n15556, B1 => n13830, B2 => 
                           n13386, ZN => n7675);
   U2491 : OAI22_X1 port map( A1 => n13387, A2 => n15555, B1 => n13836, B2 => 
                           n13386, ZN => n7676);
   U2492 : OAI22_X1 port map( A1 => n13387, A2 => n15554, B1 => n13842, B2 => 
                           n13386, ZN => n7677);
   U2493 : OAI22_X1 port map( A1 => n13387, A2 => n15553, B1 => n13848, B2 => 
                           n13386, ZN => n7678);
   U2494 : OAI22_X1 port map( A1 => n13387, A2 => n15552, B1 => n13854, B2 => 
                           n13386, ZN => n7679);
   U2495 : OAI22_X1 port map( A1 => n13387, A2 => n15551, B1 => n13860, B2 => 
                           n13386, ZN => n7680);
   U2496 : OAI22_X1 port map( A1 => n13387, A2 => n15550, B1 => n13866, B2 => 
                           n13386, ZN => n7681);
   U2497 : OAI22_X1 port map( A1 => n13387, A2 => n15549, B1 => n13872, B2 => 
                           n13386, ZN => n7682);
   U2498 : OAI22_X1 port map( A1 => n13827, A2 => n13527, B1 => n13522, B2 => 
                           n15970, ZN => n8410);
   U2499 : OAI22_X1 port map( A1 => n13833, A2 => n13527, B1 => n13522, B2 => 
                           n15969, ZN => n8411);
   U2500 : OAI22_X1 port map( A1 => n13839, A2 => n13527, B1 => n13522, B2 => 
                           n15968, ZN => n8412);
   U2501 : OAI22_X1 port map( A1 => n13845, A2 => n13527, B1 => n13522, B2 => 
                           n15967, ZN => n8413);
   U2502 : OAI22_X1 port map( A1 => n13851, A2 => n13527, B1 => n13522, B2 => 
                           n15966, ZN => n8414);
   U2503 : OAI22_X1 port map( A1 => n13857, A2 => n13527, B1 => n13522, B2 => 
                           n15965, ZN => n8415);
   U2504 : OAI22_X1 port map( A1 => n13863, A2 => n13527, B1 => n13522, B2 => 
                           n15964, ZN => n8416);
   U2505 : OAI22_X1 port map( A1 => n13869, A2 => n13527, B1 => n13522, B2 => 
                           n15963, ZN => n8417);
   U2506 : OAI22_X1 port map( A1 => n13875, A2 => n13526, B1 => n13522, B2 => 
                           n15962, ZN => n8418);
   U2507 : OAI22_X1 port map( A1 => n13881, A2 => n13526, B1 => n13522, B2 => 
                           n15961, ZN => n8419);
   U2508 : OAI22_X1 port map( A1 => n13887, A2 => n13526, B1 => n13522, B2 => 
                           n15960, ZN => n8420);
   U2509 : OAI22_X1 port map( A1 => n13893, A2 => n13526, B1 => n13522, B2 => 
                           n15959, ZN => n8421);
   U2510 : OAI22_X1 port map( A1 => n13899, A2 => n13526, B1 => n13523, B2 => 
                           n15958, ZN => n8422);
   U2511 : OAI22_X1 port map( A1 => n13905, A2 => n13526, B1 => n13523, B2 => 
                           n15957, ZN => n8423);
   U2512 : OAI22_X1 port map( A1 => n13911, A2 => n13526, B1 => n13523, B2 => 
                           n15956, ZN => n8424);
   U2513 : OAI22_X1 port map( A1 => n13917, A2 => n13526, B1 => n13523, B2 => 
                           n15955, ZN => n8425);
   U2514 : OAI22_X1 port map( A1 => n13923, A2 => n13526, B1 => n13523, B2 => 
                           n15954, ZN => n8426);
   U2515 : OAI22_X1 port map( A1 => n13929, A2 => n13526, B1 => n13523, B2 => 
                           n15953, ZN => n8427);
   U2516 : OAI22_X1 port map( A1 => n13935, A2 => n13526, B1 => n13523, B2 => 
                           n15952, ZN => n8428);
   U2517 : OAI22_X1 port map( A1 => n13941, A2 => n13526, B1 => n13523, B2 => 
                           n15951, ZN => n8429);
   U2518 : OAI22_X1 port map( A1 => n13947, A2 => n13525, B1 => n13523, B2 => 
                           n15950, ZN => n8430);
   U2519 : OAI22_X1 port map( A1 => n13953, A2 => n13525, B1 => n13523, B2 => 
                           n15949, ZN => n8431);
   U2520 : OAI22_X1 port map( A1 => n13959, A2 => n13525, B1 => n13523, B2 => 
                           n15948, ZN => n8432);
   U2521 : OAI22_X1 port map( A1 => n13965, A2 => n13525, B1 => n13523, B2 => 
                           n15947, ZN => n8433);
   U2522 : OAI22_X1 port map( A1 => n13830, A2 => n13395, B1 => n13390, B2 => 
                           n15524, ZN => n7707);
   U2523 : OAI22_X1 port map( A1 => n13836, A2 => n13395, B1 => n13390, B2 => 
                           n15523, ZN => n7708);
   U2524 : OAI22_X1 port map( A1 => n13842, A2 => n13395, B1 => n13390, B2 => 
                           n15522, ZN => n7709);
   U2525 : OAI22_X1 port map( A1 => n13848, A2 => n13395, B1 => n13390, B2 => 
                           n15521, ZN => n7710);
   U2526 : OAI22_X1 port map( A1 => n13854, A2 => n13395, B1 => n13390, B2 => 
                           n15520, ZN => n7711);
   U2527 : OAI22_X1 port map( A1 => n13860, A2 => n13395, B1 => n13390, B2 => 
                           n15519, ZN => n7712);
   U2528 : OAI22_X1 port map( A1 => n13866, A2 => n13395, B1 => n13390, B2 => 
                           n15518, ZN => n7713);
   U2529 : OAI22_X1 port map( A1 => n13872, A2 => n13394, B1 => n13390, B2 => 
                           n15517, ZN => n7714);
   U2530 : OAI22_X1 port map( A1 => n13878, A2 => n13394, B1 => n13390, B2 => 
                           n15516, ZN => n7715);
   U2531 : OAI22_X1 port map( A1 => n13884, A2 => n13394, B1 => n13390, B2 => 
                           n15515, ZN => n7716);
   U2532 : OAI22_X1 port map( A1 => n13890, A2 => n13394, B1 => n13390, B2 => 
                           n15514, ZN => n7717);
   U2533 : OAI22_X1 port map( A1 => n13896, A2 => n13394, B1 => n13391, B2 => 
                           n15513, ZN => n7718);
   U2534 : OAI22_X1 port map( A1 => n13902, A2 => n13394, B1 => n13391, B2 => 
                           n15512, ZN => n7719);
   U2535 : OAI22_X1 port map( A1 => n13908, A2 => n13394, B1 => n13391, B2 => 
                           n15511, ZN => n7720);
   U2536 : OAI22_X1 port map( A1 => n13914, A2 => n13394, B1 => n13391, B2 => 
                           n15510, ZN => n7721);
   U2537 : OAI22_X1 port map( A1 => n13920, A2 => n13394, B1 => n13391, B2 => 
                           n15509, ZN => n7722);
   U2538 : OAI22_X1 port map( A1 => n13926, A2 => n13394, B1 => n13391, B2 => 
                           n15508, ZN => n7723);
   U2539 : OAI22_X1 port map( A1 => n13932, A2 => n13394, B1 => n13391, B2 => 
                           n15507, ZN => n7724);
   U2540 : OAI22_X1 port map( A1 => n13938, A2 => n13394, B1 => n13391, B2 => 
                           n15506, ZN => n7725);
   U2541 : OAI22_X1 port map( A1 => n13944, A2 => n13393, B1 => n13391, B2 => 
                           n15505, ZN => n7726);
   U2542 : OAI22_X1 port map( A1 => n13950, A2 => n13393, B1 => n13391, B2 => 
                           n15504, ZN => n7727);
   U2543 : OAI22_X1 port map( A1 => n13956, A2 => n13393, B1 => n13391, B2 => 
                           n15503, ZN => n7728);
   U2544 : OAI22_X1 port map( A1 => n13962, A2 => n13393, B1 => n13391, B2 => 
                           n15502, ZN => n7729);
   U2545 : OAI22_X1 port map( A1 => n13828, A2 => n13443, B1 => n13438, B2 => 
                           n15301, ZN => n7962);
   U2546 : OAI22_X1 port map( A1 => n13834, A2 => n13443, B1 => n13438, B2 => 
                           n15300, ZN => n7963);
   U2547 : OAI22_X1 port map( A1 => n13840, A2 => n13443, B1 => n13438, B2 => 
                           n15299, ZN => n7964);
   U2548 : OAI22_X1 port map( A1 => n13846, A2 => n13443, B1 => n13438, B2 => 
                           n15298, ZN => n7965);
   U2549 : OAI22_X1 port map( A1 => n13852, A2 => n13443, B1 => n13438, B2 => 
                           n15297, ZN => n7966);
   U2550 : OAI22_X1 port map( A1 => n13858, A2 => n13443, B1 => n13438, B2 => 
                           n15296, ZN => n7967);
   U2551 : OAI22_X1 port map( A1 => n13864, A2 => n13443, B1 => n13438, B2 => 
                           n15295, ZN => n7968);
   U2552 : OAI22_X1 port map( A1 => n13870, A2 => n13443, B1 => n13438, B2 => 
                           n15294, ZN => n7969);
   U2553 : OAI22_X1 port map( A1 => n13876, A2 => n13442, B1 => n13438, B2 => 
                           n15293, ZN => n7970);
   U2554 : OAI22_X1 port map( A1 => n13882, A2 => n13442, B1 => n13438, B2 => 
                           n15292, ZN => n7971);
   U2555 : OAI22_X1 port map( A1 => n13888, A2 => n13442, B1 => n13438, B2 => 
                           n15291, ZN => n7972);
   U2556 : OAI22_X1 port map( A1 => n13894, A2 => n13442, B1 => n13438, B2 => 
                           n15290, ZN => n7973);
   U2557 : OAI22_X1 port map( A1 => n13900, A2 => n13442, B1 => n13439, B2 => 
                           n15289, ZN => n7974);
   U2558 : OAI22_X1 port map( A1 => n13906, A2 => n13442, B1 => n13439, B2 => 
                           n15288, ZN => n7975);
   U2559 : OAI22_X1 port map( A1 => n13912, A2 => n13442, B1 => n13439, B2 => 
                           n15287, ZN => n7976);
   U2560 : OAI22_X1 port map( A1 => n13918, A2 => n13442, B1 => n13439, B2 => 
                           n15286, ZN => n7977);
   U2561 : OAI22_X1 port map( A1 => n13924, A2 => n13442, B1 => n13439, B2 => 
                           n15285, ZN => n7978);
   U2562 : OAI22_X1 port map( A1 => n13930, A2 => n13442, B1 => n13439, B2 => 
                           n15284, ZN => n7979);
   U2563 : OAI22_X1 port map( A1 => n13936, A2 => n13442, B1 => n13439, B2 => 
                           n15283, ZN => n7980);
   U2564 : OAI22_X1 port map( A1 => n13942, A2 => n13442, B1 => n13439, B2 => 
                           n15282, ZN => n7981);
   U2565 : OAI22_X1 port map( A1 => n13948, A2 => n13441, B1 => n13439, B2 => 
                           n15281, ZN => n7982);
   U2566 : OAI22_X1 port map( A1 => n13954, A2 => n13441, B1 => n13439, B2 => 
                           n15280, ZN => n7983);
   U2567 : OAI22_X1 port map( A1 => n13960, A2 => n13441, B1 => n13439, B2 => 
                           n15279, ZN => n7984);
   U2568 : OAI22_X1 port map( A1 => n13966, A2 => n13441, B1 => n13439, B2 => 
                           n15278, ZN => n7985);
   U2569 : OAI22_X1 port map( A1 => n13828, A2 => n13449, B1 => n13444, B2 => 
                           n15269, ZN => n7994);
   U2570 : OAI22_X1 port map( A1 => n13834, A2 => n13449, B1 => n13444, B2 => 
                           n15268, ZN => n7995);
   U2571 : OAI22_X1 port map( A1 => n13840, A2 => n13449, B1 => n13444, B2 => 
                           n15267, ZN => n7996);
   U2572 : OAI22_X1 port map( A1 => n13846, A2 => n13449, B1 => n13444, B2 => 
                           n15266, ZN => n7997);
   U2573 : OAI22_X1 port map( A1 => n13852, A2 => n13449, B1 => n13444, B2 => 
                           n15265, ZN => n7998);
   U2574 : OAI22_X1 port map( A1 => n13858, A2 => n13449, B1 => n13444, B2 => 
                           n15264, ZN => n7999);
   U2575 : OAI22_X1 port map( A1 => n13864, A2 => n13449, B1 => n13444, B2 => 
                           n15263, ZN => n8000);
   U2576 : OAI22_X1 port map( A1 => n13870, A2 => n13449, B1 => n13444, B2 => 
                           n15262, ZN => n8001);
   U2577 : OAI22_X1 port map( A1 => n13876, A2 => n13448, B1 => n13444, B2 => 
                           n15261, ZN => n8002);
   U2578 : OAI22_X1 port map( A1 => n13882, A2 => n13448, B1 => n13444, B2 => 
                           n15260, ZN => n8003);
   U2579 : OAI22_X1 port map( A1 => n13888, A2 => n13448, B1 => n13444, B2 => 
                           n15259, ZN => n8004);
   U2580 : OAI22_X1 port map( A1 => n13894, A2 => n13448, B1 => n13444, B2 => 
                           n15258, ZN => n8005);
   U2581 : OAI22_X1 port map( A1 => n13900, A2 => n13448, B1 => n13445, B2 => 
                           n15257, ZN => n8006);
   U2582 : OAI22_X1 port map( A1 => n13906, A2 => n13448, B1 => n13445, B2 => 
                           n15256, ZN => n8007);
   U2583 : OAI22_X1 port map( A1 => n13912, A2 => n13448, B1 => n13445, B2 => 
                           n15255, ZN => n8008);
   U2584 : OAI22_X1 port map( A1 => n13918, A2 => n13448, B1 => n13445, B2 => 
                           n15254, ZN => n8009);
   U2585 : OAI22_X1 port map( A1 => n13924, A2 => n13448, B1 => n13445, B2 => 
                           n15253, ZN => n8010);
   U2586 : OAI22_X1 port map( A1 => n13930, A2 => n13448, B1 => n13445, B2 => 
                           n15252, ZN => n8011);
   U2587 : OAI22_X1 port map( A1 => n13936, A2 => n13448, B1 => n13445, B2 => 
                           n15251, ZN => n8012);
   U2588 : OAI22_X1 port map( A1 => n13942, A2 => n13448, B1 => n13445, B2 => 
                           n15250, ZN => n8013);
   U2589 : OAI22_X1 port map( A1 => n13948, A2 => n13447, B1 => n13445, B2 => 
                           n15249, ZN => n8014);
   U2590 : OAI22_X1 port map( A1 => n13954, A2 => n13447, B1 => n13445, B2 => 
                           n15248, ZN => n8015);
   U2591 : OAI22_X1 port map( A1 => n13960, A2 => n13447, B1 => n13445, B2 => 
                           n15247, ZN => n8016);
   U2592 : OAI22_X1 port map( A1 => n13966, A2 => n13447, B1 => n13445, B2 => 
                           n15246, ZN => n8017);
   U2593 : OAI22_X1 port map( A1 => n13828, A2 => n13455, B1 => n13450, B2 => 
                           n15237, ZN => n8026);
   U2594 : OAI22_X1 port map( A1 => n13834, A2 => n13455, B1 => n13450, B2 => 
                           n15236, ZN => n8027);
   U2595 : OAI22_X1 port map( A1 => n13840, A2 => n13455, B1 => n13450, B2 => 
                           n15235, ZN => n8028);
   U2596 : OAI22_X1 port map( A1 => n13846, A2 => n13455, B1 => n13450, B2 => 
                           n15234, ZN => n8029);
   U2597 : OAI22_X1 port map( A1 => n13852, A2 => n13455, B1 => n13450, B2 => 
                           n15233, ZN => n8030);
   U2598 : OAI22_X1 port map( A1 => n13858, A2 => n13455, B1 => n13450, B2 => 
                           n15232, ZN => n8031);
   U2599 : OAI22_X1 port map( A1 => n13864, A2 => n13455, B1 => n13450, B2 => 
                           n15231, ZN => n8032);
   U2600 : OAI22_X1 port map( A1 => n13870, A2 => n13455, B1 => n13450, B2 => 
                           n15230, ZN => n8033);
   U2601 : OAI22_X1 port map( A1 => n13876, A2 => n13454, B1 => n13450, B2 => 
                           n15229, ZN => n8034);
   U2602 : OAI22_X1 port map( A1 => n13882, A2 => n13454, B1 => n13450, B2 => 
                           n15228, ZN => n8035);
   U2603 : OAI22_X1 port map( A1 => n13888, A2 => n13454, B1 => n13450, B2 => 
                           n15227, ZN => n8036);
   U2604 : OAI22_X1 port map( A1 => n13894, A2 => n13454, B1 => n13450, B2 => 
                           n15226, ZN => n8037);
   U2605 : OAI22_X1 port map( A1 => n13900, A2 => n13454, B1 => n13451, B2 => 
                           n15225, ZN => n8038);
   U2606 : OAI22_X1 port map( A1 => n13906, A2 => n13454, B1 => n13451, B2 => 
                           n15224, ZN => n8039);
   U2607 : OAI22_X1 port map( A1 => n13912, A2 => n13454, B1 => n13451, B2 => 
                           n15223, ZN => n8040);
   U2608 : OAI22_X1 port map( A1 => n13918, A2 => n13454, B1 => n13451, B2 => 
                           n15222, ZN => n8041);
   U2609 : OAI22_X1 port map( A1 => n13924, A2 => n13454, B1 => n13451, B2 => 
                           n15221, ZN => n8042);
   U2610 : OAI22_X1 port map( A1 => n13930, A2 => n13454, B1 => n13451, B2 => 
                           n15220, ZN => n8043);
   U2611 : OAI22_X1 port map( A1 => n13936, A2 => n13454, B1 => n13451, B2 => 
                           n15219, ZN => n8044);
   U2612 : OAI22_X1 port map( A1 => n13942, A2 => n13454, B1 => n13451, B2 => 
                           n15218, ZN => n8045);
   U2613 : OAI22_X1 port map( A1 => n13948, A2 => n13453, B1 => n13451, B2 => 
                           n15217, ZN => n8046);
   U2614 : OAI22_X1 port map( A1 => n13954, A2 => n13453, B1 => n13451, B2 => 
                           n15216, ZN => n8047);
   U2615 : OAI22_X1 port map( A1 => n13960, A2 => n13453, B1 => n13451, B2 => 
                           n15215, ZN => n8048);
   U2616 : OAI22_X1 port map( A1 => n13966, A2 => n13453, B1 => n13451, B2 => 
                           n15214, ZN => n8049);
   U2617 : OAI22_X1 port map( A1 => n13828, A2 => n13485, B1 => n13480, B2 => 
                           n15173, ZN => n8186);
   U2618 : OAI22_X1 port map( A1 => n13834, A2 => n13485, B1 => n13480, B2 => 
                           n15172, ZN => n8187);
   U2619 : OAI22_X1 port map( A1 => n13840, A2 => n13485, B1 => n13480, B2 => 
                           n15171, ZN => n8188);
   U2620 : OAI22_X1 port map( A1 => n13846, A2 => n13485, B1 => n13480, B2 => 
                           n15170, ZN => n8189);
   U2621 : OAI22_X1 port map( A1 => n13852, A2 => n13485, B1 => n13480, B2 => 
                           n15169, ZN => n8190);
   U2622 : OAI22_X1 port map( A1 => n13858, A2 => n13485, B1 => n13480, B2 => 
                           n15168, ZN => n8191);
   U2623 : OAI22_X1 port map( A1 => n13864, A2 => n13485, B1 => n13480, B2 => 
                           n15167, ZN => n8192);
   U2624 : OAI22_X1 port map( A1 => n13870, A2 => n13485, B1 => n13480, B2 => 
                           n15166, ZN => n8193);
   U2625 : OAI22_X1 port map( A1 => n13876, A2 => n13484, B1 => n13480, B2 => 
                           n15165, ZN => n8194);
   U2626 : OAI22_X1 port map( A1 => n13882, A2 => n13484, B1 => n13480, B2 => 
                           n15164, ZN => n8195);
   U2627 : OAI22_X1 port map( A1 => n13888, A2 => n13484, B1 => n13480, B2 => 
                           n15163, ZN => n8196);
   U2628 : OAI22_X1 port map( A1 => n13894, A2 => n13484, B1 => n13480, B2 => 
                           n15162, ZN => n8197);
   U2629 : OAI22_X1 port map( A1 => n13900, A2 => n13484, B1 => n13481, B2 => 
                           n15161, ZN => n8198);
   U2630 : OAI22_X1 port map( A1 => n13906, A2 => n13484, B1 => n13481, B2 => 
                           n15160, ZN => n8199);
   U2631 : OAI22_X1 port map( A1 => n13912, A2 => n13484, B1 => n13481, B2 => 
                           n15159, ZN => n8200);
   U2632 : OAI22_X1 port map( A1 => n13918, A2 => n13484, B1 => n13481, B2 => 
                           n15158, ZN => n8201);
   U2633 : OAI22_X1 port map( A1 => n13924, A2 => n13484, B1 => n13481, B2 => 
                           n15157, ZN => n8202);
   U2634 : OAI22_X1 port map( A1 => n13930, A2 => n13484, B1 => n13481, B2 => 
                           n15156, ZN => n8203);
   U2635 : OAI22_X1 port map( A1 => n13936, A2 => n13484, B1 => n13481, B2 => 
                           n15155, ZN => n8204);
   U2636 : OAI22_X1 port map( A1 => n13942, A2 => n13484, B1 => n13481, B2 => 
                           n15154, ZN => n8205);
   U2637 : OAI22_X1 port map( A1 => n13948, A2 => n13483, B1 => n13481, B2 => 
                           n15153, ZN => n8206);
   U2638 : OAI22_X1 port map( A1 => n13954, A2 => n13483, B1 => n13481, B2 => 
                           n15152, ZN => n8207);
   U2639 : OAI22_X1 port map( A1 => n13960, A2 => n13483, B1 => n13481, B2 => 
                           n15151, ZN => n8208);
   U2640 : OAI22_X1 port map( A1 => n13966, A2 => n13483, B1 => n13481, B2 => 
                           n15150, ZN => n8209);
   U2641 : OAI22_X1 port map( A1 => n13828, A2 => n13491, B1 => n13486, B2 => 
                           n15141, ZN => n8218);
   U2642 : OAI22_X1 port map( A1 => n13834, A2 => n13491, B1 => n13486, B2 => 
                           n15140, ZN => n8219);
   U2643 : OAI22_X1 port map( A1 => n13840, A2 => n13491, B1 => n13486, B2 => 
                           n15139, ZN => n8220);
   U2644 : OAI22_X1 port map( A1 => n13846, A2 => n13491, B1 => n13486, B2 => 
                           n15138, ZN => n8221);
   U2645 : OAI22_X1 port map( A1 => n13852, A2 => n13491, B1 => n13486, B2 => 
                           n15137, ZN => n8222);
   U2646 : OAI22_X1 port map( A1 => n13858, A2 => n13491, B1 => n13486, B2 => 
                           n15136, ZN => n8223);
   U2647 : OAI22_X1 port map( A1 => n13864, A2 => n13491, B1 => n13486, B2 => 
                           n15135, ZN => n8224);
   U2648 : OAI22_X1 port map( A1 => n13870, A2 => n13491, B1 => n13486, B2 => 
                           n15134, ZN => n8225);
   U2649 : OAI22_X1 port map( A1 => n13876, A2 => n13490, B1 => n13486, B2 => 
                           n15133, ZN => n8226);
   U2650 : OAI22_X1 port map( A1 => n13882, A2 => n13490, B1 => n13486, B2 => 
                           n15132, ZN => n8227);
   U2651 : OAI22_X1 port map( A1 => n13888, A2 => n13490, B1 => n13486, B2 => 
                           n15131, ZN => n8228);
   U2652 : OAI22_X1 port map( A1 => n13894, A2 => n13490, B1 => n13486, B2 => 
                           n15130, ZN => n8229);
   U2653 : OAI22_X1 port map( A1 => n13900, A2 => n13490, B1 => n13487, B2 => 
                           n15129, ZN => n8230);
   U2654 : OAI22_X1 port map( A1 => n13906, A2 => n13490, B1 => n13487, B2 => 
                           n15128, ZN => n8231);
   U2655 : OAI22_X1 port map( A1 => n13912, A2 => n13490, B1 => n13487, B2 => 
                           n15127, ZN => n8232);
   U2656 : OAI22_X1 port map( A1 => n13918, A2 => n13490, B1 => n13487, B2 => 
                           n15126, ZN => n8233);
   U2657 : OAI22_X1 port map( A1 => n13924, A2 => n13490, B1 => n13487, B2 => 
                           n15125, ZN => n8234);
   U2658 : OAI22_X1 port map( A1 => n13930, A2 => n13490, B1 => n13487, B2 => 
                           n15124, ZN => n8235);
   U2659 : OAI22_X1 port map( A1 => n13936, A2 => n13490, B1 => n13487, B2 => 
                           n15123, ZN => n8236);
   U2660 : OAI22_X1 port map( A1 => n13942, A2 => n13490, B1 => n13487, B2 => 
                           n15122, ZN => n8237);
   U2661 : OAI22_X1 port map( A1 => n13948, A2 => n13489, B1 => n13487, B2 => 
                           n15121, ZN => n8238);
   U2662 : OAI22_X1 port map( A1 => n13954, A2 => n13489, B1 => n13487, B2 => 
                           n15120, ZN => n8239);
   U2663 : OAI22_X1 port map( A1 => n13960, A2 => n13489, B1 => n13487, B2 => 
                           n15119, ZN => n8240);
   U2664 : OAI22_X1 port map( A1 => n13966, A2 => n13489, B1 => n13487, B2 => 
                           n15118, ZN => n8241);
   U2665 : OAI22_X1 port map( A1 => n13828, A2 => n13497, B1 => n13492, B2 => 
                           n15109, ZN => n8250);
   U2666 : OAI22_X1 port map( A1 => n13834, A2 => n13497, B1 => n13492, B2 => 
                           n15108, ZN => n8251);
   U2667 : OAI22_X1 port map( A1 => n13840, A2 => n13497, B1 => n13492, B2 => 
                           n15107, ZN => n8252);
   U2668 : OAI22_X1 port map( A1 => n13846, A2 => n13497, B1 => n13492, B2 => 
                           n15106, ZN => n8253);
   U2669 : OAI22_X1 port map( A1 => n13852, A2 => n13497, B1 => n13492, B2 => 
                           n15105, ZN => n8254);
   U2670 : OAI22_X1 port map( A1 => n13858, A2 => n13497, B1 => n13492, B2 => 
                           n15104, ZN => n8255);
   U2671 : OAI22_X1 port map( A1 => n13864, A2 => n13497, B1 => n13492, B2 => 
                           n15103, ZN => n8256);
   U2672 : OAI22_X1 port map( A1 => n13870, A2 => n13497, B1 => n13492, B2 => 
                           n15102, ZN => n8257);
   U2673 : OAI22_X1 port map( A1 => n13876, A2 => n13496, B1 => n13492, B2 => 
                           n15101, ZN => n8258);
   U2674 : OAI22_X1 port map( A1 => n13882, A2 => n13496, B1 => n13492, B2 => 
                           n15100, ZN => n8259);
   U2675 : OAI22_X1 port map( A1 => n13888, A2 => n13496, B1 => n13492, B2 => 
                           n15099, ZN => n8260);
   U2676 : OAI22_X1 port map( A1 => n13894, A2 => n13496, B1 => n13492, B2 => 
                           n15098, ZN => n8261);
   U2677 : OAI22_X1 port map( A1 => n13900, A2 => n13496, B1 => n13493, B2 => 
                           n15097, ZN => n8262);
   U2678 : OAI22_X1 port map( A1 => n13906, A2 => n13496, B1 => n13493, B2 => 
                           n15096, ZN => n8263);
   U2679 : OAI22_X1 port map( A1 => n13912, A2 => n13496, B1 => n13493, B2 => 
                           n15095, ZN => n8264);
   U2680 : OAI22_X1 port map( A1 => n13918, A2 => n13496, B1 => n13493, B2 => 
                           n15094, ZN => n8265);
   U2681 : OAI22_X1 port map( A1 => n13924, A2 => n13496, B1 => n13493, B2 => 
                           n15093, ZN => n8266);
   U2682 : OAI22_X1 port map( A1 => n13930, A2 => n13496, B1 => n13493, B2 => 
                           n15092, ZN => n8267);
   U2683 : OAI22_X1 port map( A1 => n13936, A2 => n13496, B1 => n13493, B2 => 
                           n15091, ZN => n8268);
   U2684 : OAI22_X1 port map( A1 => n13942, A2 => n13496, B1 => n13493, B2 => 
                           n15090, ZN => n8269);
   U2685 : OAI22_X1 port map( A1 => n13948, A2 => n13495, B1 => n13493, B2 => 
                           n15089, ZN => n8270);
   U2686 : OAI22_X1 port map( A1 => n13954, A2 => n13495, B1 => n13493, B2 => 
                           n15088, ZN => n8271);
   U2687 : OAI22_X1 port map( A1 => n13960, A2 => n13495, B1 => n13493, B2 => 
                           n15087, ZN => n8272);
   U2688 : OAI22_X1 port map( A1 => n13966, A2 => n13495, B1 => n13493, B2 => 
                           n15086, ZN => n8273);
   U2689 : OAI22_X1 port map( A1 => n13828, A2 => n13503, B1 => n13498, B2 => 
                           n15077, ZN => n8282);
   U2690 : OAI22_X1 port map( A1 => n13834, A2 => n13503, B1 => n13498, B2 => 
                           n15076, ZN => n8283);
   U2691 : OAI22_X1 port map( A1 => n13840, A2 => n13503, B1 => n13498, B2 => 
                           n15075, ZN => n8284);
   U2692 : OAI22_X1 port map( A1 => n13846, A2 => n13503, B1 => n13498, B2 => 
                           n15074, ZN => n8285);
   U2693 : OAI22_X1 port map( A1 => n13852, A2 => n13503, B1 => n13498, B2 => 
                           n15073, ZN => n8286);
   U2694 : OAI22_X1 port map( A1 => n13858, A2 => n13503, B1 => n13498, B2 => 
                           n15072, ZN => n8287);
   U2695 : OAI22_X1 port map( A1 => n13864, A2 => n13503, B1 => n13498, B2 => 
                           n15071, ZN => n8288);
   U2696 : OAI22_X1 port map( A1 => n13870, A2 => n13503, B1 => n13498, B2 => 
                           n15070, ZN => n8289);
   U2697 : OAI22_X1 port map( A1 => n13876, A2 => n13502, B1 => n13498, B2 => 
                           n15069, ZN => n8290);
   U2698 : OAI22_X1 port map( A1 => n13882, A2 => n13502, B1 => n13498, B2 => 
                           n15068, ZN => n8291);
   U2699 : OAI22_X1 port map( A1 => n13888, A2 => n13502, B1 => n13498, B2 => 
                           n15067, ZN => n8292);
   U2700 : OAI22_X1 port map( A1 => n13894, A2 => n13502, B1 => n13498, B2 => 
                           n15066, ZN => n8293);
   U2701 : OAI22_X1 port map( A1 => n13900, A2 => n13502, B1 => n13499, B2 => 
                           n15065, ZN => n8294);
   U2702 : OAI22_X1 port map( A1 => n13906, A2 => n13502, B1 => n13499, B2 => 
                           n15064, ZN => n8295);
   U2703 : OAI22_X1 port map( A1 => n13912, A2 => n13502, B1 => n13499, B2 => 
                           n15063, ZN => n8296);
   U2704 : OAI22_X1 port map( A1 => n13918, A2 => n13502, B1 => n13499, B2 => 
                           n15062, ZN => n8297);
   U2705 : OAI22_X1 port map( A1 => n13924, A2 => n13502, B1 => n13499, B2 => 
                           n15061, ZN => n8298);
   U2706 : OAI22_X1 port map( A1 => n13930, A2 => n13502, B1 => n13499, B2 => 
                           n15060, ZN => n8299);
   U2707 : OAI22_X1 port map( A1 => n13936, A2 => n13502, B1 => n13499, B2 => 
                           n15059, ZN => n8300);
   U2708 : OAI22_X1 port map( A1 => n13942, A2 => n13502, B1 => n13499, B2 => 
                           n15058, ZN => n8301);
   U2709 : OAI22_X1 port map( A1 => n13948, A2 => n13501, B1 => n13499, B2 => 
                           n15057, ZN => n8302);
   U2710 : OAI22_X1 port map( A1 => n13954, A2 => n13501, B1 => n13499, B2 => 
                           n15056, ZN => n8303);
   U2711 : OAI22_X1 port map( A1 => n13960, A2 => n13501, B1 => n13499, B2 => 
                           n15055, ZN => n8304);
   U2712 : OAI22_X1 port map( A1 => n13966, A2 => n13501, B1 => n13499, B2 => 
                           n15054, ZN => n8305);
   U2713 : OAI22_X1 port map( A1 => n13827, A2 => n13509, B1 => n13504, B2 => 
                           n15045, ZN => n8314);
   U2714 : OAI22_X1 port map( A1 => n13834, A2 => n13509, B1 => n13504, B2 => 
                           n15044, ZN => n8315);
   U2715 : OAI22_X1 port map( A1 => n13840, A2 => n13509, B1 => n13504, B2 => 
                           n15043, ZN => n8316);
   U2716 : OAI22_X1 port map( A1 => n13846, A2 => n13509, B1 => n13504, B2 => 
                           n15042, ZN => n8317);
   U2717 : OAI22_X1 port map( A1 => n13852, A2 => n13509, B1 => n13504, B2 => 
                           n15041, ZN => n8318);
   U2718 : OAI22_X1 port map( A1 => n13858, A2 => n13509, B1 => n13504, B2 => 
                           n15040, ZN => n8319);
   U2719 : OAI22_X1 port map( A1 => n13864, A2 => n13509, B1 => n13504, B2 => 
                           n15039, ZN => n8320);
   U2720 : OAI22_X1 port map( A1 => n13870, A2 => n13509, B1 => n13504, B2 => 
                           n15038, ZN => n8321);
   U2721 : OAI22_X1 port map( A1 => n13876, A2 => n13508, B1 => n13504, B2 => 
                           n15037, ZN => n8322);
   U2722 : OAI22_X1 port map( A1 => n13882, A2 => n13508, B1 => n13504, B2 => 
                           n15036, ZN => n8323);
   U2723 : OAI22_X1 port map( A1 => n13888, A2 => n13508, B1 => n13504, B2 => 
                           n15035, ZN => n8324);
   U2724 : OAI22_X1 port map( A1 => n13894, A2 => n13508, B1 => n13504, B2 => 
                           n15034, ZN => n8325);
   U2725 : OAI22_X1 port map( A1 => n13900, A2 => n13508, B1 => n13505, B2 => 
                           n15033, ZN => n8326);
   U2726 : OAI22_X1 port map( A1 => n13906, A2 => n13508, B1 => n13505, B2 => 
                           n15032, ZN => n8327);
   U2727 : OAI22_X1 port map( A1 => n13912, A2 => n13508, B1 => n13505, B2 => 
                           n15031, ZN => n8328);
   U2728 : OAI22_X1 port map( A1 => n13918, A2 => n13508, B1 => n13505, B2 => 
                           n15030, ZN => n8329);
   U2729 : OAI22_X1 port map( A1 => n13924, A2 => n13508, B1 => n13505, B2 => 
                           n15029, ZN => n8330);
   U2730 : OAI22_X1 port map( A1 => n13930, A2 => n13508, B1 => n13505, B2 => 
                           n15028, ZN => n8331);
   U2731 : OAI22_X1 port map( A1 => n13936, A2 => n13508, B1 => n13505, B2 => 
                           n15027, ZN => n8332);
   U2732 : OAI22_X1 port map( A1 => n13942, A2 => n13508, B1 => n13505, B2 => 
                           n15026, ZN => n8333);
   U2733 : OAI22_X1 port map( A1 => n13948, A2 => n13507, B1 => n13505, B2 => 
                           n15025, ZN => n8334);
   U2734 : OAI22_X1 port map( A1 => n13954, A2 => n13507, B1 => n13505, B2 => 
                           n15024, ZN => n8335);
   U2735 : OAI22_X1 port map( A1 => n13960, A2 => n13507, B1 => n13505, B2 => 
                           n15023, ZN => n8336);
   U2736 : OAI22_X1 port map( A1 => n13966, A2 => n13507, B1 => n13505, B2 => 
                           n15022, ZN => n8337);
   U2737 : OAI22_X1 port map( A1 => n13827, A2 => n13533, B1 => n13528, B2 => 
                           n14980, ZN => n8442);
   U2738 : OAI22_X1 port map( A1 => n13833, A2 => n13533, B1 => n13528, B2 => 
                           n14979, ZN => n8443);
   U2739 : OAI22_X1 port map( A1 => n13839, A2 => n13533, B1 => n13528, B2 => 
                           n14978, ZN => n8444);
   U2740 : OAI22_X1 port map( A1 => n13845, A2 => n13533, B1 => n13528, B2 => 
                           n14977, ZN => n8445);
   U2741 : OAI22_X1 port map( A1 => n13851, A2 => n13533, B1 => n13528, B2 => 
                           n14976, ZN => n8446);
   U2742 : OAI22_X1 port map( A1 => n13857, A2 => n13533, B1 => n13528, B2 => 
                           n14975, ZN => n8447);
   U2743 : OAI22_X1 port map( A1 => n13863, A2 => n13533, B1 => n13528, B2 => 
                           n14974, ZN => n8448);
   U2744 : OAI22_X1 port map( A1 => n13869, A2 => n13533, B1 => n13528, B2 => 
                           n14973, ZN => n8449);
   U2745 : OAI22_X1 port map( A1 => n13875, A2 => n13532, B1 => n13528, B2 => 
                           n14972, ZN => n8450);
   U2746 : OAI22_X1 port map( A1 => n13881, A2 => n13532, B1 => n13528, B2 => 
                           n14971, ZN => n8451);
   U2747 : OAI22_X1 port map( A1 => n13887, A2 => n13532, B1 => n13528, B2 => 
                           n14970, ZN => n8452);
   U2748 : OAI22_X1 port map( A1 => n13893, A2 => n13532, B1 => n13528, B2 => 
                           n14969, ZN => n8453);
   U2749 : OAI22_X1 port map( A1 => n13899, A2 => n13532, B1 => n13529, B2 => 
                           n14968, ZN => n8454);
   U2750 : OAI22_X1 port map( A1 => n13905, A2 => n13532, B1 => n13529, B2 => 
                           n14967, ZN => n8455);
   U2751 : OAI22_X1 port map( A1 => n13911, A2 => n13532, B1 => n13529, B2 => 
                           n14966, ZN => n8456);
   U2752 : OAI22_X1 port map( A1 => n13917, A2 => n13532, B1 => n13529, B2 => 
                           n14965, ZN => n8457);
   U2753 : OAI22_X1 port map( A1 => n13923, A2 => n13532, B1 => n13529, B2 => 
                           n14964, ZN => n8458);
   U2754 : OAI22_X1 port map( A1 => n13929, A2 => n13532, B1 => n13529, B2 => 
                           n14963, ZN => n8459);
   U2755 : OAI22_X1 port map( A1 => n13935, A2 => n13532, B1 => n13529, B2 => 
                           n14962, ZN => n8460);
   U2756 : OAI22_X1 port map( A1 => n13941, A2 => n13532, B1 => n13529, B2 => 
                           n14961, ZN => n8461);
   U2757 : OAI22_X1 port map( A1 => n13947, A2 => n13531, B1 => n13529, B2 => 
                           n14960, ZN => n8462);
   U2758 : OAI22_X1 port map( A1 => n13953, A2 => n13531, B1 => n13529, B2 => 
                           n14959, ZN => n8463);
   U2759 : OAI22_X1 port map( A1 => n13959, A2 => n13531, B1 => n13529, B2 => 
                           n14958, ZN => n8464);
   U2760 : OAI22_X1 port map( A1 => n13965, A2 => n13531, B1 => n13529, B2 => 
                           n14957, ZN => n8465);
   U2761 : OAI22_X1 port map( A1 => n13827, A2 => n13551, B1 => n13546, B2 => 
                           n14947, ZN => n8538);
   U2762 : OAI22_X1 port map( A1 => n13833, A2 => n13551, B1 => n13546, B2 => 
                           n14946, ZN => n8539);
   U2763 : OAI22_X1 port map( A1 => n13839, A2 => n13551, B1 => n13546, B2 => 
                           n14945, ZN => n8540);
   U2764 : OAI22_X1 port map( A1 => n13845, A2 => n13551, B1 => n13546, B2 => 
                           n14944, ZN => n8541);
   U2765 : OAI22_X1 port map( A1 => n13851, A2 => n13551, B1 => n13546, B2 => 
                           n14943, ZN => n8542);
   U2766 : OAI22_X1 port map( A1 => n13857, A2 => n13551, B1 => n13546, B2 => 
                           n14942, ZN => n8543);
   U2767 : OAI22_X1 port map( A1 => n13863, A2 => n13551, B1 => n13546, B2 => 
                           n14941, ZN => n8544);
   U2768 : OAI22_X1 port map( A1 => n13869, A2 => n13551, B1 => n13546, B2 => 
                           n14940, ZN => n8545);
   U2769 : OAI22_X1 port map( A1 => n13875, A2 => n13550, B1 => n13546, B2 => 
                           n14939, ZN => n8546);
   U2770 : OAI22_X1 port map( A1 => n13881, A2 => n13550, B1 => n13546, B2 => 
                           n14938, ZN => n8547);
   U2771 : OAI22_X1 port map( A1 => n13887, A2 => n13550, B1 => n13546, B2 => 
                           n14937, ZN => n8548);
   U2772 : OAI22_X1 port map( A1 => n13893, A2 => n13550, B1 => n13546, B2 => 
                           n14936, ZN => n8549);
   U2773 : OAI22_X1 port map( A1 => n13899, A2 => n13550, B1 => n13547, B2 => 
                           n14935, ZN => n8550);
   U2774 : OAI22_X1 port map( A1 => n13905, A2 => n13550, B1 => n13547, B2 => 
                           n14934, ZN => n8551);
   U2775 : OAI22_X1 port map( A1 => n13911, A2 => n13550, B1 => n13547, B2 => 
                           n14933, ZN => n8552);
   U2776 : OAI22_X1 port map( A1 => n13917, A2 => n13550, B1 => n13547, B2 => 
                           n14932, ZN => n8553);
   U2777 : OAI22_X1 port map( A1 => n13923, A2 => n13550, B1 => n13547, B2 => 
                           n14931, ZN => n8554);
   U2778 : OAI22_X1 port map( A1 => n13929, A2 => n13550, B1 => n13547, B2 => 
                           n14930, ZN => n8555);
   U2779 : OAI22_X1 port map( A1 => n13935, A2 => n13550, B1 => n13547, B2 => 
                           n14929, ZN => n8556);
   U2780 : OAI22_X1 port map( A1 => n13941, A2 => n13550, B1 => n13547, B2 => 
                           n14928, ZN => n8557);
   U2781 : OAI22_X1 port map( A1 => n13947, A2 => n13549, B1 => n13547, B2 => 
                           n14927, ZN => n8558);
   U2782 : OAI22_X1 port map( A1 => n13953, A2 => n13549, B1 => n13547, B2 => 
                           n14926, ZN => n8559);
   U2783 : OAI22_X1 port map( A1 => n13959, A2 => n13549, B1 => n13547, B2 => 
                           n14925, ZN => n8560);
   U2784 : OAI22_X1 port map( A1 => n13965, A2 => n13549, B1 => n13547, B2 => 
                           n14924, ZN => n8561);
   U2785 : OAI22_X1 port map( A1 => n13827, A2 => n13557, B1 => n13552, B2 => 
                           n14915, ZN => n8570);
   U2786 : OAI22_X1 port map( A1 => n13833, A2 => n13557, B1 => n13552, B2 => 
                           n14914, ZN => n8571);
   U2787 : OAI22_X1 port map( A1 => n13839, A2 => n13557, B1 => n13552, B2 => 
                           n14913, ZN => n8572);
   U2788 : OAI22_X1 port map( A1 => n13845, A2 => n13557, B1 => n13552, B2 => 
                           n14912, ZN => n8573);
   U2789 : OAI22_X1 port map( A1 => n13851, A2 => n13557, B1 => n13552, B2 => 
                           n14911, ZN => n8574);
   U2790 : OAI22_X1 port map( A1 => n13857, A2 => n13557, B1 => n13552, B2 => 
                           n14910, ZN => n8575);
   U2791 : OAI22_X1 port map( A1 => n13863, A2 => n13557, B1 => n13552, B2 => 
                           n14909, ZN => n8576);
   U2792 : OAI22_X1 port map( A1 => n13869, A2 => n13557, B1 => n13552, B2 => 
                           n14908, ZN => n8577);
   U2793 : OAI22_X1 port map( A1 => n13875, A2 => n13556, B1 => n13552, B2 => 
                           n14907, ZN => n8578);
   U2794 : OAI22_X1 port map( A1 => n13881, A2 => n13556, B1 => n13552, B2 => 
                           n14906, ZN => n8579);
   U2795 : OAI22_X1 port map( A1 => n13887, A2 => n13556, B1 => n13552, B2 => 
                           n14905, ZN => n8580);
   U2796 : OAI22_X1 port map( A1 => n13893, A2 => n13556, B1 => n13552, B2 => 
                           n14904, ZN => n8581);
   U2797 : OAI22_X1 port map( A1 => n13899, A2 => n13556, B1 => n13553, B2 => 
                           n14903, ZN => n8582);
   U2798 : OAI22_X1 port map( A1 => n13905, A2 => n13556, B1 => n13553, B2 => 
                           n14902, ZN => n8583);
   U2799 : OAI22_X1 port map( A1 => n13911, A2 => n13556, B1 => n13553, B2 => 
                           n14901, ZN => n8584);
   U2800 : OAI22_X1 port map( A1 => n13917, A2 => n13556, B1 => n13553, B2 => 
                           n14900, ZN => n8585);
   U2801 : OAI22_X1 port map( A1 => n13923, A2 => n13556, B1 => n13553, B2 => 
                           n14899, ZN => n8586);
   U2802 : OAI22_X1 port map( A1 => n13929, A2 => n13556, B1 => n13553, B2 => 
                           n14898, ZN => n8587);
   U2803 : OAI22_X1 port map( A1 => n13935, A2 => n13556, B1 => n13553, B2 => 
                           n14897, ZN => n8588);
   U2804 : OAI22_X1 port map( A1 => n13941, A2 => n13556, B1 => n13553, B2 => 
                           n14896, ZN => n8589);
   U2805 : OAI22_X1 port map( A1 => n13947, A2 => n13555, B1 => n13553, B2 => 
                           n14895, ZN => n8590);
   U2806 : OAI22_X1 port map( A1 => n13953, A2 => n13555, B1 => n13553, B2 => 
                           n14894, ZN => n8591);
   U2807 : OAI22_X1 port map( A1 => n13959, A2 => n13555, B1 => n13553, B2 => 
                           n14893, ZN => n8592);
   U2808 : OAI22_X1 port map( A1 => n13965, A2 => n13555, B1 => n13553, B2 => 
                           n14892, ZN => n8593);
   U2809 : OAI22_X1 port map( A1 => n13827, A2 => n13563, B1 => n13558, B2 => 
                           n14883, ZN => n8602);
   U2810 : OAI22_X1 port map( A1 => n13833, A2 => n13563, B1 => n13558, B2 => 
                           n14882, ZN => n8603);
   U2811 : OAI22_X1 port map( A1 => n13839, A2 => n13563, B1 => n13558, B2 => 
                           n14881, ZN => n8604);
   U2812 : OAI22_X1 port map( A1 => n13845, A2 => n13563, B1 => n13558, B2 => 
                           n14880, ZN => n8605);
   U2813 : OAI22_X1 port map( A1 => n13851, A2 => n13563, B1 => n13558, B2 => 
                           n14879, ZN => n8606);
   U2814 : OAI22_X1 port map( A1 => n13857, A2 => n13563, B1 => n13558, B2 => 
                           n14878, ZN => n8607);
   U2815 : OAI22_X1 port map( A1 => n13863, A2 => n13563, B1 => n13558, B2 => 
                           n14877, ZN => n8608);
   U2816 : OAI22_X1 port map( A1 => n13869, A2 => n13563, B1 => n13558, B2 => 
                           n14876, ZN => n8609);
   U2817 : OAI22_X1 port map( A1 => n13875, A2 => n13562, B1 => n13558, B2 => 
                           n14875, ZN => n8610);
   U2818 : OAI22_X1 port map( A1 => n13881, A2 => n13562, B1 => n13558, B2 => 
                           n14874, ZN => n8611);
   U2819 : OAI22_X1 port map( A1 => n13887, A2 => n13562, B1 => n13558, B2 => 
                           n14873, ZN => n8612);
   U2820 : OAI22_X1 port map( A1 => n13893, A2 => n13562, B1 => n13558, B2 => 
                           n14872, ZN => n8613);
   U2821 : OAI22_X1 port map( A1 => n13899, A2 => n13562, B1 => n13559, B2 => 
                           n14871, ZN => n8614);
   U2822 : OAI22_X1 port map( A1 => n13905, A2 => n13562, B1 => n13559, B2 => 
                           n14870, ZN => n8615);
   U2823 : OAI22_X1 port map( A1 => n13911, A2 => n13562, B1 => n13559, B2 => 
                           n14869, ZN => n8616);
   U2824 : OAI22_X1 port map( A1 => n13917, A2 => n13562, B1 => n13559, B2 => 
                           n14868, ZN => n8617);
   U2825 : OAI22_X1 port map( A1 => n13923, A2 => n13562, B1 => n13559, B2 => 
                           n14867, ZN => n8618);
   U2826 : OAI22_X1 port map( A1 => n13929, A2 => n13562, B1 => n13559, B2 => 
                           n14866, ZN => n8619);
   U2827 : OAI22_X1 port map( A1 => n13935, A2 => n13562, B1 => n13559, B2 => 
                           n14865, ZN => n8620);
   U2828 : OAI22_X1 port map( A1 => n13941, A2 => n13562, B1 => n13559, B2 => 
                           n14864, ZN => n8621);
   U2829 : OAI22_X1 port map( A1 => n13947, A2 => n13561, B1 => n13559, B2 => 
                           n14863, ZN => n8622);
   U2830 : OAI22_X1 port map( A1 => n13953, A2 => n13561, B1 => n13559, B2 => 
                           n14862, ZN => n8623);
   U2831 : OAI22_X1 port map( A1 => n13959, A2 => n13561, B1 => n13559, B2 => 
                           n14861, ZN => n8624);
   U2832 : OAI22_X1 port map( A1 => n13965, A2 => n13561, B1 => n13559, B2 => 
                           n14860, ZN => n8625);
   U2833 : OAI22_X1 port map( A1 => n13826, A2 => n13593, B1 => n13588, B2 => 
                           n14851, ZN => n8762);
   U2834 : OAI22_X1 port map( A1 => n13833, A2 => n13593, B1 => n13588, B2 => 
                           n14850, ZN => n8763);
   U2835 : OAI22_X1 port map( A1 => n13839, A2 => n13593, B1 => n13588, B2 => 
                           n14849, ZN => n8764);
   U2836 : OAI22_X1 port map( A1 => n13845, A2 => n13593, B1 => n13588, B2 => 
                           n14848, ZN => n8765);
   U2837 : OAI22_X1 port map( A1 => n13851, A2 => n13593, B1 => n13588, B2 => 
                           n14847, ZN => n8766);
   U2838 : OAI22_X1 port map( A1 => n13857, A2 => n13593, B1 => n13588, B2 => 
                           n14846, ZN => n8767);
   U2839 : OAI22_X1 port map( A1 => n13863, A2 => n13593, B1 => n13588, B2 => 
                           n14845, ZN => n8768);
   U2840 : OAI22_X1 port map( A1 => n13869, A2 => n13593, B1 => n13588, B2 => 
                           n14844, ZN => n8769);
   U2841 : OAI22_X1 port map( A1 => n13875, A2 => n13592, B1 => n13588, B2 => 
                           n14843, ZN => n8770);
   U2842 : OAI22_X1 port map( A1 => n13881, A2 => n13592, B1 => n13588, B2 => 
                           n14842, ZN => n8771);
   U2843 : OAI22_X1 port map( A1 => n13887, A2 => n13592, B1 => n13588, B2 => 
                           n14841, ZN => n8772);
   U2844 : OAI22_X1 port map( A1 => n13893, A2 => n13592, B1 => n13588, B2 => 
                           n14840, ZN => n8773);
   U2845 : OAI22_X1 port map( A1 => n13899, A2 => n13592, B1 => n13589, B2 => 
                           n14839, ZN => n8774);
   U2846 : OAI22_X1 port map( A1 => n13905, A2 => n13592, B1 => n13589, B2 => 
                           n14838, ZN => n8775);
   U2847 : OAI22_X1 port map( A1 => n13911, A2 => n13592, B1 => n13589, B2 => 
                           n14837, ZN => n8776);
   U2848 : OAI22_X1 port map( A1 => n13917, A2 => n13592, B1 => n13589, B2 => 
                           n14836, ZN => n8777);
   U2849 : OAI22_X1 port map( A1 => n13923, A2 => n13592, B1 => n13589, B2 => 
                           n14835, ZN => n8778);
   U2850 : OAI22_X1 port map( A1 => n13929, A2 => n13592, B1 => n13589, B2 => 
                           n14834, ZN => n8779);
   U2851 : OAI22_X1 port map( A1 => n13935, A2 => n13592, B1 => n13589, B2 => 
                           n14833, ZN => n8780);
   U2852 : OAI22_X1 port map( A1 => n13941, A2 => n13592, B1 => n13589, B2 => 
                           n14832, ZN => n8781);
   U2853 : OAI22_X1 port map( A1 => n13947, A2 => n13591, B1 => n13589, B2 => 
                           n14831, ZN => n8782);
   U2854 : OAI22_X1 port map( A1 => n13953, A2 => n13591, B1 => n13589, B2 => 
                           n14830, ZN => n8783);
   U2855 : OAI22_X1 port map( A1 => n13959, A2 => n13591, B1 => n13589, B2 => 
                           n14829, ZN => n8784);
   U2856 : OAI22_X1 port map( A1 => n13965, A2 => n13591, B1 => n13589, B2 => 
                           n14828, ZN => n8785);
   U2857 : OAI22_X1 port map( A1 => n13826, A2 => n13599, B1 => n13594, B2 => 
                           n14819, ZN => n8794);
   U2858 : OAI22_X1 port map( A1 => n13832, A2 => n13599, B1 => n13594, B2 => 
                           n14818, ZN => n8795);
   U2859 : OAI22_X1 port map( A1 => n13838, A2 => n13599, B1 => n13594, B2 => 
                           n14817, ZN => n8796);
   U2860 : OAI22_X1 port map( A1 => n13844, A2 => n13599, B1 => n13594, B2 => 
                           n14816, ZN => n8797);
   U2861 : OAI22_X1 port map( A1 => n13850, A2 => n13599, B1 => n13594, B2 => 
                           n14815, ZN => n8798);
   U2862 : OAI22_X1 port map( A1 => n13856, A2 => n13599, B1 => n13594, B2 => 
                           n14814, ZN => n8799);
   U2863 : OAI22_X1 port map( A1 => n13862, A2 => n13599, B1 => n13594, B2 => 
                           n14813, ZN => n8800);
   U2864 : OAI22_X1 port map( A1 => n13868, A2 => n13599, B1 => n13594, B2 => 
                           n14812, ZN => n8801);
   U2865 : OAI22_X1 port map( A1 => n13874, A2 => n13598, B1 => n13594, B2 => 
                           n14811, ZN => n8802);
   U2866 : OAI22_X1 port map( A1 => n13880, A2 => n13598, B1 => n13594, B2 => 
                           n14810, ZN => n8803);
   U2867 : OAI22_X1 port map( A1 => n13886, A2 => n13598, B1 => n13594, B2 => 
                           n14809, ZN => n8804);
   U2868 : OAI22_X1 port map( A1 => n13892, A2 => n13598, B1 => n13594, B2 => 
                           n14808, ZN => n8805);
   U2869 : OAI22_X1 port map( A1 => n13898, A2 => n13598, B1 => n13595, B2 => 
                           n14807, ZN => n8806);
   U2870 : OAI22_X1 port map( A1 => n13904, A2 => n13598, B1 => n13595, B2 => 
                           n14806, ZN => n8807);
   U2871 : OAI22_X1 port map( A1 => n13910, A2 => n13598, B1 => n13595, B2 => 
                           n14805, ZN => n8808);
   U2872 : OAI22_X1 port map( A1 => n13916, A2 => n13598, B1 => n13595, B2 => 
                           n14804, ZN => n8809);
   U2873 : OAI22_X1 port map( A1 => n13922, A2 => n13598, B1 => n13595, B2 => 
                           n14803, ZN => n8810);
   U2874 : OAI22_X1 port map( A1 => n13928, A2 => n13598, B1 => n13595, B2 => 
                           n14802, ZN => n8811);
   U2875 : OAI22_X1 port map( A1 => n13934, A2 => n13598, B1 => n13595, B2 => 
                           n14801, ZN => n8812);
   U2876 : OAI22_X1 port map( A1 => n13940, A2 => n13598, B1 => n13595, B2 => 
                           n14800, ZN => n8813);
   U2877 : OAI22_X1 port map( A1 => n13946, A2 => n13597, B1 => n13595, B2 => 
                           n14799, ZN => n8814);
   U2878 : OAI22_X1 port map( A1 => n13952, A2 => n13597, B1 => n13595, B2 => 
                           n14798, ZN => n8815);
   U2879 : OAI22_X1 port map( A1 => n13958, A2 => n13597, B1 => n13595, B2 => 
                           n14797, ZN => n8816);
   U2880 : OAI22_X1 port map( A1 => n13964, A2 => n13597, B1 => n13595, B2 => 
                           n14796, ZN => n8817);
   U2881 : OAI22_X1 port map( A1 => n13826, A2 => n13605, B1 => n13600, B2 => 
                           n14787, ZN => n8826);
   U2882 : OAI22_X1 port map( A1 => n13832, A2 => n13605, B1 => n13600, B2 => 
                           n14786, ZN => n8827);
   U2883 : OAI22_X1 port map( A1 => n13838, A2 => n13605, B1 => n13600, B2 => 
                           n14785, ZN => n8828);
   U2884 : OAI22_X1 port map( A1 => n13844, A2 => n13605, B1 => n13600, B2 => 
                           n14784, ZN => n8829);
   U2885 : OAI22_X1 port map( A1 => n13850, A2 => n13605, B1 => n13600, B2 => 
                           n14783, ZN => n8830);
   U2886 : OAI22_X1 port map( A1 => n13856, A2 => n13605, B1 => n13600, B2 => 
                           n14782, ZN => n8831);
   U2887 : OAI22_X1 port map( A1 => n13862, A2 => n13605, B1 => n13600, B2 => 
                           n14781, ZN => n8832);
   U2888 : OAI22_X1 port map( A1 => n13868, A2 => n13605, B1 => n13600, B2 => 
                           n14780, ZN => n8833);
   U2889 : OAI22_X1 port map( A1 => n13874, A2 => n13604, B1 => n13600, B2 => 
                           n14779, ZN => n8834);
   U2890 : OAI22_X1 port map( A1 => n13880, A2 => n13604, B1 => n13600, B2 => 
                           n14778, ZN => n8835);
   U2891 : OAI22_X1 port map( A1 => n13886, A2 => n13604, B1 => n13600, B2 => 
                           n14777, ZN => n8836);
   U2892 : OAI22_X1 port map( A1 => n13892, A2 => n13604, B1 => n13600, B2 => 
                           n14776, ZN => n8837);
   U2893 : OAI22_X1 port map( A1 => n13898, A2 => n13604, B1 => n13601, B2 => 
                           n14775, ZN => n8838);
   U2894 : OAI22_X1 port map( A1 => n13904, A2 => n13604, B1 => n13601, B2 => 
                           n14774, ZN => n8839);
   U2895 : OAI22_X1 port map( A1 => n13910, A2 => n13604, B1 => n13601, B2 => 
                           n14773, ZN => n8840);
   U2896 : OAI22_X1 port map( A1 => n13916, A2 => n13604, B1 => n13601, B2 => 
                           n14772, ZN => n8841);
   U2897 : OAI22_X1 port map( A1 => n13922, A2 => n13604, B1 => n13601, B2 => 
                           n14771, ZN => n8842);
   U2898 : OAI22_X1 port map( A1 => n13928, A2 => n13604, B1 => n13601, B2 => 
                           n14770, ZN => n8843);
   U2899 : OAI22_X1 port map( A1 => n13934, A2 => n13604, B1 => n13601, B2 => 
                           n14769, ZN => n8844);
   U2900 : OAI22_X1 port map( A1 => n13940, A2 => n13604, B1 => n13601, B2 => 
                           n14768, ZN => n8845);
   U2901 : OAI22_X1 port map( A1 => n13946, A2 => n13603, B1 => n13601, B2 => 
                           n14767, ZN => n8846);
   U2902 : OAI22_X1 port map( A1 => n13952, A2 => n13603, B1 => n13601, B2 => 
                           n14766, ZN => n8847);
   U2903 : OAI22_X1 port map( A1 => n13958, A2 => n13603, B1 => n13601, B2 => 
                           n14765, ZN => n8848);
   U2904 : OAI22_X1 port map( A1 => n13964, A2 => n13603, B1 => n13601, B2 => 
                           n14764, ZN => n8849);
   U2905 : OAI22_X1 port map( A1 => n13826, A2 => n13611, B1 => n13606, B2 => 
                           n14755, ZN => n8858);
   U2906 : OAI22_X1 port map( A1 => n13832, A2 => n13611, B1 => n13606, B2 => 
                           n14754, ZN => n8859);
   U2907 : OAI22_X1 port map( A1 => n13838, A2 => n13611, B1 => n13606, B2 => 
                           n14753, ZN => n8860);
   U2908 : OAI22_X1 port map( A1 => n13844, A2 => n13611, B1 => n13606, B2 => 
                           n14752, ZN => n8861);
   U2909 : OAI22_X1 port map( A1 => n13850, A2 => n13611, B1 => n13606, B2 => 
                           n14751, ZN => n8862);
   U2910 : OAI22_X1 port map( A1 => n13856, A2 => n13611, B1 => n13606, B2 => 
                           n14750, ZN => n8863);
   U2911 : OAI22_X1 port map( A1 => n13862, A2 => n13611, B1 => n13606, B2 => 
                           n14749, ZN => n8864);
   U2912 : OAI22_X1 port map( A1 => n13868, A2 => n13611, B1 => n13606, B2 => 
                           n14748, ZN => n8865);
   U2913 : OAI22_X1 port map( A1 => n13874, A2 => n13610, B1 => n13606, B2 => 
                           n14747, ZN => n8866);
   U2914 : OAI22_X1 port map( A1 => n13880, A2 => n13610, B1 => n13606, B2 => 
                           n14746, ZN => n8867);
   U2915 : OAI22_X1 port map( A1 => n13886, A2 => n13610, B1 => n13606, B2 => 
                           n14745, ZN => n8868);
   U2916 : OAI22_X1 port map( A1 => n13892, A2 => n13610, B1 => n13606, B2 => 
                           n14744, ZN => n8869);
   U2917 : OAI22_X1 port map( A1 => n13898, A2 => n13610, B1 => n13607, B2 => 
                           n14743, ZN => n8870);
   U2918 : OAI22_X1 port map( A1 => n13904, A2 => n13610, B1 => n13607, B2 => 
                           n14742, ZN => n8871);
   U2919 : OAI22_X1 port map( A1 => n13910, A2 => n13610, B1 => n13607, B2 => 
                           n14741, ZN => n8872);
   U2920 : OAI22_X1 port map( A1 => n13916, A2 => n13610, B1 => n13607, B2 => 
                           n14740, ZN => n8873);
   U2921 : OAI22_X1 port map( A1 => n13922, A2 => n13610, B1 => n13607, B2 => 
                           n14739, ZN => n8874);
   U2922 : OAI22_X1 port map( A1 => n13928, A2 => n13610, B1 => n13607, B2 => 
                           n14738, ZN => n8875);
   U2923 : OAI22_X1 port map( A1 => n13934, A2 => n13610, B1 => n13607, B2 => 
                           n14737, ZN => n8876);
   U2924 : OAI22_X1 port map( A1 => n13940, A2 => n13610, B1 => n13607, B2 => 
                           n14736, ZN => n8877);
   U2925 : OAI22_X1 port map( A1 => n13946, A2 => n13609, B1 => n13607, B2 => 
                           n14735, ZN => n8878);
   U2926 : OAI22_X1 port map( A1 => n13952, A2 => n13609, B1 => n13607, B2 => 
                           n14734, ZN => n8879);
   U2927 : OAI22_X1 port map( A1 => n13958, A2 => n13609, B1 => n13607, B2 => 
                           n14733, ZN => n8880);
   U2928 : OAI22_X1 port map( A1 => n13964, A2 => n13609, B1 => n13607, B2 => 
                           n14732, ZN => n8881);
   U2929 : OAI22_X1 port map( A1 => n13826, A2 => n13617, B1 => n13612, B2 => 
                           n14723, ZN => n8890);
   U2930 : OAI22_X1 port map( A1 => n13832, A2 => n13617, B1 => n13612, B2 => 
                           n14722, ZN => n8891);
   U2931 : OAI22_X1 port map( A1 => n13838, A2 => n13617, B1 => n13612, B2 => 
                           n14721, ZN => n8892);
   U2932 : OAI22_X1 port map( A1 => n13844, A2 => n13617, B1 => n13612, B2 => 
                           n14720, ZN => n8893);
   U2933 : OAI22_X1 port map( A1 => n13850, A2 => n13617, B1 => n13612, B2 => 
                           n14719, ZN => n8894);
   U2934 : OAI22_X1 port map( A1 => n13856, A2 => n13617, B1 => n13612, B2 => 
                           n14718, ZN => n8895);
   U2935 : OAI22_X1 port map( A1 => n13862, A2 => n13617, B1 => n13612, B2 => 
                           n14717, ZN => n8896);
   U2936 : OAI22_X1 port map( A1 => n13868, A2 => n13617, B1 => n13612, B2 => 
                           n14716, ZN => n8897);
   U2937 : OAI22_X1 port map( A1 => n13874, A2 => n13616, B1 => n13612, B2 => 
                           n14715, ZN => n8898);
   U2938 : OAI22_X1 port map( A1 => n13880, A2 => n13616, B1 => n13612, B2 => 
                           n14714, ZN => n8899);
   U2939 : OAI22_X1 port map( A1 => n13886, A2 => n13616, B1 => n13612, B2 => 
                           n14713, ZN => n8900);
   U2940 : OAI22_X1 port map( A1 => n13892, A2 => n13616, B1 => n13612, B2 => 
                           n14712, ZN => n8901);
   U2941 : OAI22_X1 port map( A1 => n13898, A2 => n13616, B1 => n13613, B2 => 
                           n14711, ZN => n8902);
   U2942 : OAI22_X1 port map( A1 => n13904, A2 => n13616, B1 => n13613, B2 => 
                           n14710, ZN => n8903);
   U2943 : OAI22_X1 port map( A1 => n13910, A2 => n13616, B1 => n13613, B2 => 
                           n14709, ZN => n8904);
   U2944 : OAI22_X1 port map( A1 => n13916, A2 => n13616, B1 => n13613, B2 => 
                           n14708, ZN => n8905);
   U2945 : OAI22_X1 port map( A1 => n13922, A2 => n13616, B1 => n13613, B2 => 
                           n14707, ZN => n8906);
   U2946 : OAI22_X1 port map( A1 => n13928, A2 => n13616, B1 => n13613, B2 => 
                           n14706, ZN => n8907);
   U2947 : OAI22_X1 port map( A1 => n13934, A2 => n13616, B1 => n13613, B2 => 
                           n14705, ZN => n8908);
   U2948 : OAI22_X1 port map( A1 => n13940, A2 => n13616, B1 => n13613, B2 => 
                           n14704, ZN => n8909);
   U2949 : OAI22_X1 port map( A1 => n13946, A2 => n13615, B1 => n13613, B2 => 
                           n14703, ZN => n8910);
   U2950 : OAI22_X1 port map( A1 => n13952, A2 => n13615, B1 => n13613, B2 => 
                           n14702, ZN => n8911);
   U2951 : OAI22_X1 port map( A1 => n13958, A2 => n13615, B1 => n13613, B2 => 
                           n14701, ZN => n8912);
   U2952 : OAI22_X1 port map( A1 => n13964, A2 => n13615, B1 => n13613, B2 => 
                           n14700, ZN => n8913);
   U2953 : OAI22_X1 port map( A1 => n13826, A2 => n13647, B1 => n13642, B2 => 
                           n14652, ZN => n9050);
   U2954 : OAI22_X1 port map( A1 => n13832, A2 => n13647, B1 => n13642, B2 => 
                           n14651, ZN => n9051);
   U2955 : OAI22_X1 port map( A1 => n13838, A2 => n13647, B1 => n13642, B2 => 
                           n14650, ZN => n9052);
   U2956 : OAI22_X1 port map( A1 => n13844, A2 => n13647, B1 => n13642, B2 => 
                           n14649, ZN => n9053);
   U2957 : OAI22_X1 port map( A1 => n13850, A2 => n13647, B1 => n13642, B2 => 
                           n14648, ZN => n9054);
   U2958 : OAI22_X1 port map( A1 => n13856, A2 => n13647, B1 => n13642, B2 => 
                           n14647, ZN => n9055);
   U2959 : OAI22_X1 port map( A1 => n13862, A2 => n13647, B1 => n13642, B2 => 
                           n14646, ZN => n9056);
   U2960 : OAI22_X1 port map( A1 => n13868, A2 => n13647, B1 => n13642, B2 => 
                           n14645, ZN => n9057);
   U2961 : OAI22_X1 port map( A1 => n13874, A2 => n13646, B1 => n13642, B2 => 
                           n14644, ZN => n9058);
   U2962 : OAI22_X1 port map( A1 => n13880, A2 => n13646, B1 => n13642, B2 => 
                           n14643, ZN => n9059);
   U2963 : OAI22_X1 port map( A1 => n13886, A2 => n13646, B1 => n13642, B2 => 
                           n14642, ZN => n9060);
   U2964 : OAI22_X1 port map( A1 => n13892, A2 => n13646, B1 => n13642, B2 => 
                           n14641, ZN => n9061);
   U2965 : OAI22_X1 port map( A1 => n13898, A2 => n13646, B1 => n13643, B2 => 
                           n14640, ZN => n9062);
   U2966 : OAI22_X1 port map( A1 => n13904, A2 => n13646, B1 => n13643, B2 => 
                           n14639, ZN => n9063);
   U2967 : OAI22_X1 port map( A1 => n13910, A2 => n13646, B1 => n13643, B2 => 
                           n14638, ZN => n9064);
   U2968 : OAI22_X1 port map( A1 => n13916, A2 => n13646, B1 => n13643, B2 => 
                           n14637, ZN => n9065);
   U2969 : OAI22_X1 port map( A1 => n13922, A2 => n13646, B1 => n13643, B2 => 
                           n14636, ZN => n9066);
   U2970 : OAI22_X1 port map( A1 => n13928, A2 => n13646, B1 => n13643, B2 => 
                           n14635, ZN => n9067);
   U2971 : OAI22_X1 port map( A1 => n13934, A2 => n13646, B1 => n13643, B2 => 
                           n14634, ZN => n9068);
   U2972 : OAI22_X1 port map( A1 => n13940, A2 => n13646, B1 => n13643, B2 => 
                           n14633, ZN => n9069);
   U2973 : OAI22_X1 port map( A1 => n13946, A2 => n13645, B1 => n13643, B2 => 
                           n14632, ZN => n9070);
   U2974 : OAI22_X1 port map( A1 => n13952, A2 => n13645, B1 => n13643, B2 => 
                           n14631, ZN => n9071);
   U2975 : OAI22_X1 port map( A1 => n13958, A2 => n13645, B1 => n13643, B2 => 
                           n14630, ZN => n9072);
   U2976 : OAI22_X1 port map( A1 => n13964, A2 => n13645, B1 => n13643, B2 => 
                           n14629, ZN => n9073);
   U2977 : OAI22_X1 port map( A1 => n13826, A2 => n13653, B1 => n13648, B2 => 
                           n14620, ZN => n9082);
   U2978 : OAI22_X1 port map( A1 => n13832, A2 => n13653, B1 => n13648, B2 => 
                           n14619, ZN => n9083);
   U2979 : OAI22_X1 port map( A1 => n13838, A2 => n13653, B1 => n13648, B2 => 
                           n14618, ZN => n9084);
   U2980 : OAI22_X1 port map( A1 => n13844, A2 => n13653, B1 => n13648, B2 => 
                           n14617, ZN => n9085);
   U2981 : OAI22_X1 port map( A1 => n13850, A2 => n13653, B1 => n13648, B2 => 
                           n14616, ZN => n9086);
   U2982 : OAI22_X1 port map( A1 => n13856, A2 => n13653, B1 => n13648, B2 => 
                           n14615, ZN => n9087);
   U2983 : OAI22_X1 port map( A1 => n13862, A2 => n13653, B1 => n13648, B2 => 
                           n14614, ZN => n9088);
   U2984 : OAI22_X1 port map( A1 => n13868, A2 => n13653, B1 => n13648, B2 => 
                           n14613, ZN => n9089);
   U2985 : OAI22_X1 port map( A1 => n13874, A2 => n13652, B1 => n13648, B2 => 
                           n14612, ZN => n9090);
   U2986 : OAI22_X1 port map( A1 => n13880, A2 => n13652, B1 => n13648, B2 => 
                           n14611, ZN => n9091);
   U2987 : OAI22_X1 port map( A1 => n13886, A2 => n13652, B1 => n13648, B2 => 
                           n14610, ZN => n9092);
   U2988 : OAI22_X1 port map( A1 => n13892, A2 => n13652, B1 => n13648, B2 => 
                           n14609, ZN => n9093);
   U2989 : OAI22_X1 port map( A1 => n13898, A2 => n13652, B1 => n13649, B2 => 
                           n14608, ZN => n9094);
   U2990 : OAI22_X1 port map( A1 => n13904, A2 => n13652, B1 => n13649, B2 => 
                           n14607, ZN => n9095);
   U2991 : OAI22_X1 port map( A1 => n13910, A2 => n13652, B1 => n13649, B2 => 
                           n14606, ZN => n9096);
   U2992 : OAI22_X1 port map( A1 => n13916, A2 => n13652, B1 => n13649, B2 => 
                           n14605, ZN => n9097);
   U2993 : OAI22_X1 port map( A1 => n13922, A2 => n13652, B1 => n13649, B2 => 
                           n14604, ZN => n9098);
   U2994 : OAI22_X1 port map( A1 => n13928, A2 => n13652, B1 => n13649, B2 => 
                           n14603, ZN => n9099);
   U2995 : OAI22_X1 port map( A1 => n13934, A2 => n13652, B1 => n13649, B2 => 
                           n14602, ZN => n9100);
   U2996 : OAI22_X1 port map( A1 => n13940, A2 => n13652, B1 => n13649, B2 => 
                           n14601, ZN => n9101);
   U2997 : OAI22_X1 port map( A1 => n13946, A2 => n13651, B1 => n13649, B2 => 
                           n14600, ZN => n9102);
   U2998 : OAI22_X1 port map( A1 => n13952, A2 => n13651, B1 => n13649, B2 => 
                           n14599, ZN => n9103);
   U2999 : OAI22_X1 port map( A1 => n13958, A2 => n13651, B1 => n13649, B2 => 
                           n14598, ZN => n9104);
   U3000 : OAI22_X1 port map( A1 => n13964, A2 => n13651, B1 => n13649, B2 => 
                           n14597, ZN => n9105);
   U3001 : OAI22_X1 port map( A1 => n13826, A2 => n13659, B1 => n13654, B2 => 
                           n14588, ZN => n9114);
   U3002 : OAI22_X1 port map( A1 => n13832, A2 => n13659, B1 => n13654, B2 => 
                           n14587, ZN => n9115);
   U3003 : OAI22_X1 port map( A1 => n13838, A2 => n13659, B1 => n13654, B2 => 
                           n14586, ZN => n9116);
   U3004 : OAI22_X1 port map( A1 => n13844, A2 => n13659, B1 => n13654, B2 => 
                           n14585, ZN => n9117);
   U3005 : OAI22_X1 port map( A1 => n13850, A2 => n13659, B1 => n13654, B2 => 
                           n14584, ZN => n9118);
   U3006 : OAI22_X1 port map( A1 => n13856, A2 => n13659, B1 => n13654, B2 => 
                           n14583, ZN => n9119);
   U3007 : OAI22_X1 port map( A1 => n13862, A2 => n13659, B1 => n13654, B2 => 
                           n14582, ZN => n9120);
   U3008 : OAI22_X1 port map( A1 => n13868, A2 => n13659, B1 => n13654, B2 => 
                           n14581, ZN => n9121);
   U3009 : OAI22_X1 port map( A1 => n13874, A2 => n13658, B1 => n13654, B2 => 
                           n14580, ZN => n9122);
   U3010 : OAI22_X1 port map( A1 => n13880, A2 => n13658, B1 => n13654, B2 => 
                           n14579, ZN => n9123);
   U3011 : OAI22_X1 port map( A1 => n13886, A2 => n13658, B1 => n13654, B2 => 
                           n14578, ZN => n9124);
   U3012 : OAI22_X1 port map( A1 => n13892, A2 => n13658, B1 => n13654, B2 => 
                           n14577, ZN => n9125);
   U3013 : OAI22_X1 port map( A1 => n13898, A2 => n13658, B1 => n13655, B2 => 
                           n14576, ZN => n9126);
   U3014 : OAI22_X1 port map( A1 => n13904, A2 => n13658, B1 => n13655, B2 => 
                           n14575, ZN => n9127);
   U3015 : OAI22_X1 port map( A1 => n13910, A2 => n13658, B1 => n13655, B2 => 
                           n14574, ZN => n9128);
   U3016 : OAI22_X1 port map( A1 => n13916, A2 => n13658, B1 => n13655, B2 => 
                           n14573, ZN => n9129);
   U3017 : OAI22_X1 port map( A1 => n13922, A2 => n13658, B1 => n13655, B2 => 
                           n14572, ZN => n9130);
   U3018 : OAI22_X1 port map( A1 => n13928, A2 => n13658, B1 => n13655, B2 => 
                           n14571, ZN => n9131);
   U3019 : OAI22_X1 port map( A1 => n13934, A2 => n13658, B1 => n13655, B2 => 
                           n14570, ZN => n9132);
   U3020 : OAI22_X1 port map( A1 => n13940, A2 => n13658, B1 => n13655, B2 => 
                           n14569, ZN => n9133);
   U3021 : OAI22_X1 port map( A1 => n13946, A2 => n13657, B1 => n13655, B2 => 
                           n14568, ZN => n9134);
   U3022 : OAI22_X1 port map( A1 => n13952, A2 => n13657, B1 => n13655, B2 => 
                           n14567, ZN => n9135);
   U3023 : OAI22_X1 port map( A1 => n13958, A2 => n13657, B1 => n13655, B2 => 
                           n14566, ZN => n9136);
   U3024 : OAI22_X1 port map( A1 => n13964, A2 => n13657, B1 => n13655, B2 => 
                           n14565, ZN => n9137);
   U3025 : OAI22_X1 port map( A1 => n13825, A2 => n13665, B1 => n13660, B2 => 
                           n14556, ZN => n9146);
   U3026 : OAI22_X1 port map( A1 => n13832, A2 => n13665, B1 => n13660, B2 => 
                           n14555, ZN => n9147);
   U3027 : OAI22_X1 port map( A1 => n13838, A2 => n13665, B1 => n13660, B2 => 
                           n14554, ZN => n9148);
   U3028 : OAI22_X1 port map( A1 => n13844, A2 => n13665, B1 => n13660, B2 => 
                           n14553, ZN => n9149);
   U3029 : OAI22_X1 port map( A1 => n13850, A2 => n13665, B1 => n13660, B2 => 
                           n14552, ZN => n9150);
   U3030 : OAI22_X1 port map( A1 => n13856, A2 => n13665, B1 => n13660, B2 => 
                           n14551, ZN => n9151);
   U3031 : OAI22_X1 port map( A1 => n13862, A2 => n13665, B1 => n13660, B2 => 
                           n14550, ZN => n9152);
   U3032 : OAI22_X1 port map( A1 => n13868, A2 => n13665, B1 => n13660, B2 => 
                           n14549, ZN => n9153);
   U3033 : OAI22_X1 port map( A1 => n13874, A2 => n13664, B1 => n13660, B2 => 
                           n14548, ZN => n9154);
   U3034 : OAI22_X1 port map( A1 => n13880, A2 => n13664, B1 => n13660, B2 => 
                           n14547, ZN => n9155);
   U3035 : OAI22_X1 port map( A1 => n13886, A2 => n13664, B1 => n13660, B2 => 
                           n14546, ZN => n9156);
   U3036 : OAI22_X1 port map( A1 => n13892, A2 => n13664, B1 => n13660, B2 => 
                           n14545, ZN => n9157);
   U3037 : OAI22_X1 port map( A1 => n13898, A2 => n13664, B1 => n13661, B2 => 
                           n14544, ZN => n9158);
   U3038 : OAI22_X1 port map( A1 => n13904, A2 => n13664, B1 => n13661, B2 => 
                           n14543, ZN => n9159);
   U3039 : OAI22_X1 port map( A1 => n13910, A2 => n13664, B1 => n13661, B2 => 
                           n14542, ZN => n9160);
   U3040 : OAI22_X1 port map( A1 => n13916, A2 => n13664, B1 => n13661, B2 => 
                           n14541, ZN => n9161);
   U3041 : OAI22_X1 port map( A1 => n13922, A2 => n13664, B1 => n13661, B2 => 
                           n14540, ZN => n9162);
   U3042 : OAI22_X1 port map( A1 => n13928, A2 => n13664, B1 => n13661, B2 => 
                           n14539, ZN => n9163);
   U3043 : OAI22_X1 port map( A1 => n13934, A2 => n13664, B1 => n13661, B2 => 
                           n14538, ZN => n9164);
   U3044 : OAI22_X1 port map( A1 => n13940, A2 => n13664, B1 => n13661, B2 => 
                           n14537, ZN => n9165);
   U3045 : OAI22_X1 port map( A1 => n13946, A2 => n13663, B1 => n13661, B2 => 
                           n14536, ZN => n9166);
   U3046 : OAI22_X1 port map( A1 => n13952, A2 => n13663, B1 => n13661, B2 => 
                           n14535, ZN => n9167);
   U3047 : OAI22_X1 port map( A1 => n13958, A2 => n13663, B1 => n13661, B2 => 
                           n14534, ZN => n9168);
   U3048 : OAI22_X1 port map( A1 => n13964, A2 => n13663, B1 => n13661, B2 => 
                           n14533, ZN => n9169);
   U3049 : OAI22_X1 port map( A1 => n13825, A2 => n13671, B1 => n13666, B2 => 
                           n14524, ZN => n9178);
   U3050 : OAI22_X1 port map( A1 => n13831, A2 => n13671, B1 => n13666, B2 => 
                           n14523, ZN => n9179);
   U3051 : OAI22_X1 port map( A1 => n13837, A2 => n13671, B1 => n13666, B2 => 
                           n14522, ZN => n9180);
   U3052 : OAI22_X1 port map( A1 => n13843, A2 => n13671, B1 => n13666, B2 => 
                           n14521, ZN => n9181);
   U3053 : OAI22_X1 port map( A1 => n13849, A2 => n13671, B1 => n13666, B2 => 
                           n14520, ZN => n9182);
   U3054 : OAI22_X1 port map( A1 => n13855, A2 => n13671, B1 => n13666, B2 => 
                           n14519, ZN => n9183);
   U3055 : OAI22_X1 port map( A1 => n13861, A2 => n13671, B1 => n13666, B2 => 
                           n14518, ZN => n9184);
   U3056 : OAI22_X1 port map( A1 => n13867, A2 => n13671, B1 => n13666, B2 => 
                           n14517, ZN => n9185);
   U3057 : OAI22_X1 port map( A1 => n13873, A2 => n13670, B1 => n13666, B2 => 
                           n14516, ZN => n9186);
   U3058 : OAI22_X1 port map( A1 => n13879, A2 => n13670, B1 => n13666, B2 => 
                           n14515, ZN => n9187);
   U3059 : OAI22_X1 port map( A1 => n13885, A2 => n13670, B1 => n13666, B2 => 
                           n14514, ZN => n9188);
   U3060 : OAI22_X1 port map( A1 => n13891, A2 => n13670, B1 => n13666, B2 => 
                           n14513, ZN => n9189);
   U3061 : OAI22_X1 port map( A1 => n13897, A2 => n13670, B1 => n13667, B2 => 
                           n14512, ZN => n9190);
   U3062 : OAI22_X1 port map( A1 => n13903, A2 => n13670, B1 => n13667, B2 => 
                           n14511, ZN => n9191);
   U3063 : OAI22_X1 port map( A1 => n13909, A2 => n13670, B1 => n13667, B2 => 
                           n14510, ZN => n9192);
   U3064 : OAI22_X1 port map( A1 => n13915, A2 => n13670, B1 => n13667, B2 => 
                           n14509, ZN => n9193);
   U3065 : OAI22_X1 port map( A1 => n13921, A2 => n13670, B1 => n13667, B2 => 
                           n14508, ZN => n9194);
   U3066 : OAI22_X1 port map( A1 => n13927, A2 => n13670, B1 => n13667, B2 => 
                           n14507, ZN => n9195);
   U3067 : OAI22_X1 port map( A1 => n13933, A2 => n13670, B1 => n13667, B2 => 
                           n14506, ZN => n9196);
   U3068 : OAI22_X1 port map( A1 => n13939, A2 => n13670, B1 => n13667, B2 => 
                           n14505, ZN => n9197);
   U3069 : OAI22_X1 port map( A1 => n13945, A2 => n13669, B1 => n13667, B2 => 
                           n14504, ZN => n9198);
   U3070 : OAI22_X1 port map( A1 => n13951, A2 => n13669, B1 => n13667, B2 => 
                           n14503, ZN => n9199);
   U3071 : OAI22_X1 port map( A1 => n13957, A2 => n13669, B1 => n13667, B2 => 
                           n14502, ZN => n9200);
   U3072 : OAI22_X1 port map( A1 => n13963, A2 => n13669, B1 => n13667, B2 => 
                           n14501, ZN => n9201);
   U3073 : OAI22_X1 port map( A1 => n13825, A2 => n13701, B1 => n13696, B2 => 
                           n14439, ZN => n9338);
   U3074 : OAI22_X1 port map( A1 => n13831, A2 => n13701, B1 => n13696, B2 => 
                           n14438, ZN => n9339);
   U3075 : OAI22_X1 port map( A1 => n13837, A2 => n13701, B1 => n13696, B2 => 
                           n14437, ZN => n9340);
   U3076 : OAI22_X1 port map( A1 => n13843, A2 => n13701, B1 => n13696, B2 => 
                           n14436, ZN => n9341);
   U3077 : OAI22_X1 port map( A1 => n13849, A2 => n13701, B1 => n13696, B2 => 
                           n14435, ZN => n9342);
   U3078 : OAI22_X1 port map( A1 => n13855, A2 => n13701, B1 => n13696, B2 => 
                           n14434, ZN => n9343);
   U3079 : OAI22_X1 port map( A1 => n13861, A2 => n13701, B1 => n13696, B2 => 
                           n14433, ZN => n9344);
   U3080 : OAI22_X1 port map( A1 => n13867, A2 => n13701, B1 => n13696, B2 => 
                           n14432, ZN => n9345);
   U3081 : OAI22_X1 port map( A1 => n13873, A2 => n13700, B1 => n13696, B2 => 
                           n14431, ZN => n9346);
   U3082 : OAI22_X1 port map( A1 => n13879, A2 => n13700, B1 => n13696, B2 => 
                           n14430, ZN => n9347);
   U3083 : OAI22_X1 port map( A1 => n13885, A2 => n13700, B1 => n13696, B2 => 
                           n14429, ZN => n9348);
   U3084 : OAI22_X1 port map( A1 => n13891, A2 => n13700, B1 => n13696, B2 => 
                           n14428, ZN => n9349);
   U3085 : OAI22_X1 port map( A1 => n13897, A2 => n13700, B1 => n13697, B2 => 
                           n14427, ZN => n9350);
   U3086 : OAI22_X1 port map( A1 => n13903, A2 => n13700, B1 => n13697, B2 => 
                           n14426, ZN => n9351);
   U3087 : OAI22_X1 port map( A1 => n13909, A2 => n13700, B1 => n13697, B2 => 
                           n14425, ZN => n9352);
   U3088 : OAI22_X1 port map( A1 => n13915, A2 => n13700, B1 => n13697, B2 => 
                           n14424, ZN => n9353);
   U3089 : OAI22_X1 port map( A1 => n13921, A2 => n13700, B1 => n13697, B2 => 
                           n14423, ZN => n9354);
   U3090 : OAI22_X1 port map( A1 => n13927, A2 => n13700, B1 => n13697, B2 => 
                           n14422, ZN => n9355);
   U3091 : OAI22_X1 port map( A1 => n13933, A2 => n13700, B1 => n13697, B2 => 
                           n14421, ZN => n9356);
   U3092 : OAI22_X1 port map( A1 => n13939, A2 => n13700, B1 => n13697, B2 => 
                           n14420, ZN => n9357);
   U3093 : OAI22_X1 port map( A1 => n13945, A2 => n13699, B1 => n13697, B2 => 
                           n14419, ZN => n9358);
   U3094 : OAI22_X1 port map( A1 => n13951, A2 => n13699, B1 => n13697, B2 => 
                           n14418, ZN => n9359);
   U3095 : OAI22_X1 port map( A1 => n13957, A2 => n13699, B1 => n13697, B2 => 
                           n14417, ZN => n9360);
   U3096 : OAI22_X1 port map( A1 => n13963, A2 => n13699, B1 => n13697, B2 => 
                           n14416, ZN => n9361);
   U3097 : OAI22_X1 port map( A1 => n13825, A2 => n13707, B1 => n13702, B2 => 
                           n14407, ZN => n9370);
   U3098 : OAI22_X1 port map( A1 => n13832, A2 => n13707, B1 => n13702, B2 => 
                           n14406, ZN => n9371);
   U3099 : OAI22_X1 port map( A1 => n13838, A2 => n13707, B1 => n13702, B2 => 
                           n14405, ZN => n9372);
   U3100 : OAI22_X1 port map( A1 => n13844, A2 => n13707, B1 => n13702, B2 => 
                           n14404, ZN => n9373);
   U3101 : OAI22_X1 port map( A1 => n13850, A2 => n13707, B1 => n13702, B2 => 
                           n14403, ZN => n9374);
   U3102 : OAI22_X1 port map( A1 => n13856, A2 => n13707, B1 => n13702, B2 => 
                           n14402, ZN => n9375);
   U3103 : OAI22_X1 port map( A1 => n13862, A2 => n13707, B1 => n13702, B2 => 
                           n14401, ZN => n9376);
   U3104 : OAI22_X1 port map( A1 => n13868, A2 => n13707, B1 => n13702, B2 => 
                           n14400, ZN => n9377);
   U3105 : OAI22_X1 port map( A1 => n13874, A2 => n13706, B1 => n13702, B2 => 
                           n14399, ZN => n9378);
   U3106 : OAI22_X1 port map( A1 => n13880, A2 => n13706, B1 => n13702, B2 => 
                           n14398, ZN => n9379);
   U3107 : OAI22_X1 port map( A1 => n13886, A2 => n13706, B1 => n13702, B2 => 
                           n14397, ZN => n9380);
   U3108 : OAI22_X1 port map( A1 => n13892, A2 => n13706, B1 => n13702, B2 => 
                           n14396, ZN => n9381);
   U3109 : OAI22_X1 port map( A1 => n13898, A2 => n13706, B1 => n13703, B2 => 
                           n14395, ZN => n9382);
   U3110 : OAI22_X1 port map( A1 => n13904, A2 => n13706, B1 => n13703, B2 => 
                           n14394, ZN => n9383);
   U3111 : OAI22_X1 port map( A1 => n13910, A2 => n13706, B1 => n13703, B2 => 
                           n14393, ZN => n9384);
   U3112 : OAI22_X1 port map( A1 => n13916, A2 => n13706, B1 => n13703, B2 => 
                           n14392, ZN => n9385);
   U3113 : OAI22_X1 port map( A1 => n13922, A2 => n13706, B1 => n13703, B2 => 
                           n14391, ZN => n9386);
   U3114 : OAI22_X1 port map( A1 => n13928, A2 => n13706, B1 => n13703, B2 => 
                           n14390, ZN => n9387);
   U3115 : OAI22_X1 port map( A1 => n13934, A2 => n13706, B1 => n13703, B2 => 
                           n14389, ZN => n9388);
   U3116 : OAI22_X1 port map( A1 => n13940, A2 => n13706, B1 => n13703, B2 => 
                           n14388, ZN => n9389);
   U3117 : OAI22_X1 port map( A1 => n13946, A2 => n13705, B1 => n13703, B2 => 
                           n14387, ZN => n9390);
   U3118 : OAI22_X1 port map( A1 => n13952, A2 => n13705, B1 => n13703, B2 => 
                           n14386, ZN => n9391);
   U3119 : OAI22_X1 port map( A1 => n13958, A2 => n13705, B1 => n13703, B2 => 
                           n14385, ZN => n9392);
   U3120 : OAI22_X1 port map( A1 => n13964, A2 => n13705, B1 => n13703, B2 => 
                           n14384, ZN => n9393);
   U3121 : OAI22_X1 port map( A1 => n13825, A2 => n13713, B1 => n13708, B2 => 
                           n14375, ZN => n9402);
   U3122 : OAI22_X1 port map( A1 => n13831, A2 => n13713, B1 => n13708, B2 => 
                           n14374, ZN => n9403);
   U3123 : OAI22_X1 port map( A1 => n13837, A2 => n13713, B1 => n13708, B2 => 
                           n14373, ZN => n9404);
   U3124 : OAI22_X1 port map( A1 => n13843, A2 => n13713, B1 => n13708, B2 => 
                           n14372, ZN => n9405);
   U3125 : OAI22_X1 port map( A1 => n13849, A2 => n13713, B1 => n13708, B2 => 
                           n14371, ZN => n9406);
   U3126 : OAI22_X1 port map( A1 => n13855, A2 => n13713, B1 => n13708, B2 => 
                           n14370, ZN => n9407);
   U3127 : OAI22_X1 port map( A1 => n13861, A2 => n13713, B1 => n13708, B2 => 
                           n14369, ZN => n9408);
   U3128 : OAI22_X1 port map( A1 => n13867, A2 => n13713, B1 => n13708, B2 => 
                           n14368, ZN => n9409);
   U3129 : OAI22_X1 port map( A1 => n13873, A2 => n13712, B1 => n13708, B2 => 
                           n14367, ZN => n9410);
   U3130 : OAI22_X1 port map( A1 => n13879, A2 => n13712, B1 => n13708, B2 => 
                           n14366, ZN => n9411);
   U3131 : OAI22_X1 port map( A1 => n13885, A2 => n13712, B1 => n13708, B2 => 
                           n14365, ZN => n9412);
   U3132 : OAI22_X1 port map( A1 => n13891, A2 => n13712, B1 => n13708, B2 => 
                           n14364, ZN => n9413);
   U3133 : OAI22_X1 port map( A1 => n13897, A2 => n13712, B1 => n13709, B2 => 
                           n14363, ZN => n9414);
   U3134 : OAI22_X1 port map( A1 => n13903, A2 => n13712, B1 => n13709, B2 => 
                           n14362, ZN => n9415);
   U3135 : OAI22_X1 port map( A1 => n13909, A2 => n13712, B1 => n13709, B2 => 
                           n14361, ZN => n9416);
   U3136 : OAI22_X1 port map( A1 => n13915, A2 => n13712, B1 => n13709, B2 => 
                           n14360, ZN => n9417);
   U3137 : OAI22_X1 port map( A1 => n13921, A2 => n13712, B1 => n13709, B2 => 
                           n14359, ZN => n9418);
   U3138 : OAI22_X1 port map( A1 => n13927, A2 => n13712, B1 => n13709, B2 => 
                           n14358, ZN => n9419);
   U3139 : OAI22_X1 port map( A1 => n13933, A2 => n13712, B1 => n13709, B2 => 
                           n14357, ZN => n9420);
   U3140 : OAI22_X1 port map( A1 => n13939, A2 => n13712, B1 => n13709, B2 => 
                           n14356, ZN => n9421);
   U3141 : OAI22_X1 port map( A1 => n13945, A2 => n13711, B1 => n13709, B2 => 
                           n14355, ZN => n9422);
   U3142 : OAI22_X1 port map( A1 => n13951, A2 => n13711, B1 => n13709, B2 => 
                           n14354, ZN => n9423);
   U3143 : OAI22_X1 port map( A1 => n13957, A2 => n13711, B1 => n13709, B2 => 
                           n14353, ZN => n9424);
   U3144 : OAI22_X1 port map( A1 => n13963, A2 => n13711, B1 => n13709, B2 => 
                           n14352, ZN => n9425);
   U3145 : OAI22_X1 port map( A1 => n13825, A2 => n13719, B1 => n13714, B2 => 
                           n14343, ZN => n9434);
   U3146 : OAI22_X1 port map( A1 => n13831, A2 => n13719, B1 => n13714, B2 => 
                           n14342, ZN => n9435);
   U3147 : OAI22_X1 port map( A1 => n13837, A2 => n13719, B1 => n13714, B2 => 
                           n14341, ZN => n9436);
   U3148 : OAI22_X1 port map( A1 => n13843, A2 => n13719, B1 => n13714, B2 => 
                           n14340, ZN => n9437);
   U3149 : OAI22_X1 port map( A1 => n13849, A2 => n13719, B1 => n13714, B2 => 
                           n14339, ZN => n9438);
   U3150 : OAI22_X1 port map( A1 => n13855, A2 => n13719, B1 => n13714, B2 => 
                           n14338, ZN => n9439);
   U3151 : OAI22_X1 port map( A1 => n13861, A2 => n13719, B1 => n13714, B2 => 
                           n14337, ZN => n9440);
   U3152 : OAI22_X1 port map( A1 => n13867, A2 => n13719, B1 => n13714, B2 => 
                           n14336, ZN => n9441);
   U3153 : OAI22_X1 port map( A1 => n13873, A2 => n13718, B1 => n13714, B2 => 
                           n14335, ZN => n9442);
   U3154 : OAI22_X1 port map( A1 => n13879, A2 => n13718, B1 => n13714, B2 => 
                           n14334, ZN => n9443);
   U3155 : OAI22_X1 port map( A1 => n13885, A2 => n13718, B1 => n13714, B2 => 
                           n14333, ZN => n9444);
   U3156 : OAI22_X1 port map( A1 => n13891, A2 => n13718, B1 => n13714, B2 => 
                           n14332, ZN => n9445);
   U3157 : OAI22_X1 port map( A1 => n13897, A2 => n13718, B1 => n13715, B2 => 
                           n14331, ZN => n9446);
   U3158 : OAI22_X1 port map( A1 => n13903, A2 => n13718, B1 => n13715, B2 => 
                           n14330, ZN => n9447);
   U3159 : OAI22_X1 port map( A1 => n13909, A2 => n13718, B1 => n13715, B2 => 
                           n14329, ZN => n9448);
   U3160 : OAI22_X1 port map( A1 => n13915, A2 => n13718, B1 => n13715, B2 => 
                           n14328, ZN => n9449);
   U3161 : OAI22_X1 port map( A1 => n13921, A2 => n13718, B1 => n13715, B2 => 
                           n14327, ZN => n9450);
   U3162 : OAI22_X1 port map( A1 => n13927, A2 => n13718, B1 => n13715, B2 => 
                           n14326, ZN => n9451);
   U3163 : OAI22_X1 port map( A1 => n13933, A2 => n13718, B1 => n13715, B2 => 
                           n14325, ZN => n9452);
   U3164 : OAI22_X1 port map( A1 => n13939, A2 => n13718, B1 => n13715, B2 => 
                           n14324, ZN => n9453);
   U3165 : OAI22_X1 port map( A1 => n13945, A2 => n13717, B1 => n13715, B2 => 
                           n14323, ZN => n9454);
   U3166 : OAI22_X1 port map( A1 => n13951, A2 => n13717, B1 => n13715, B2 => 
                           n14322, ZN => n9455);
   U3167 : OAI22_X1 port map( A1 => n13957, A2 => n13717, B1 => n13715, B2 => 
                           n14321, ZN => n9456);
   U3168 : OAI22_X1 port map( A1 => n13963, A2 => n13717, B1 => n13715, B2 => 
                           n14320, ZN => n9457);
   U3169 : OAI22_X1 port map( A1 => n13825, A2 => n13725, B1 => n13720, B2 => 
                           n14311, ZN => n9466);
   U3170 : OAI22_X1 port map( A1 => n13831, A2 => n13725, B1 => n13720, B2 => 
                           n14310, ZN => n9467);
   U3171 : OAI22_X1 port map( A1 => n13837, A2 => n13725, B1 => n13720, B2 => 
                           n14309, ZN => n9468);
   U3172 : OAI22_X1 port map( A1 => n13843, A2 => n13725, B1 => n13720, B2 => 
                           n14308, ZN => n9469);
   U3173 : OAI22_X1 port map( A1 => n13849, A2 => n13725, B1 => n13720, B2 => 
                           n14307, ZN => n9470);
   U3174 : OAI22_X1 port map( A1 => n13855, A2 => n13725, B1 => n13720, B2 => 
                           n14306, ZN => n9471);
   U3175 : OAI22_X1 port map( A1 => n13861, A2 => n13725, B1 => n13720, B2 => 
                           n14305, ZN => n9472);
   U3176 : OAI22_X1 port map( A1 => n13867, A2 => n13725, B1 => n13720, B2 => 
                           n14304, ZN => n9473);
   U3177 : OAI22_X1 port map( A1 => n13873, A2 => n13724, B1 => n13720, B2 => 
                           n14303, ZN => n9474);
   U3178 : OAI22_X1 port map( A1 => n13879, A2 => n13724, B1 => n13720, B2 => 
                           n14302, ZN => n9475);
   U3179 : OAI22_X1 port map( A1 => n13885, A2 => n13724, B1 => n13720, B2 => 
                           n14301, ZN => n9476);
   U3180 : OAI22_X1 port map( A1 => n13891, A2 => n13724, B1 => n13720, B2 => 
                           n14300, ZN => n9477);
   U3181 : OAI22_X1 port map( A1 => n13897, A2 => n13724, B1 => n13721, B2 => 
                           n14299, ZN => n9478);
   U3182 : OAI22_X1 port map( A1 => n13903, A2 => n13724, B1 => n13721, B2 => 
                           n14298, ZN => n9479);
   U3183 : OAI22_X1 port map( A1 => n13909, A2 => n13724, B1 => n13721, B2 => 
                           n14297, ZN => n9480);
   U3184 : OAI22_X1 port map( A1 => n13915, A2 => n13724, B1 => n13721, B2 => 
                           n14296, ZN => n9481);
   U3185 : OAI22_X1 port map( A1 => n13921, A2 => n13724, B1 => n13721, B2 => 
                           n14295, ZN => n9482);
   U3186 : OAI22_X1 port map( A1 => n13927, A2 => n13724, B1 => n13721, B2 => 
                           n14294, ZN => n9483);
   U3187 : OAI22_X1 port map( A1 => n13933, A2 => n13724, B1 => n13721, B2 => 
                           n14293, ZN => n9484);
   U3188 : OAI22_X1 port map( A1 => n13939, A2 => n13724, B1 => n13721, B2 => 
                           n14292, ZN => n9485);
   U3189 : OAI22_X1 port map( A1 => n13945, A2 => n13723, B1 => n13721, B2 => 
                           n14291, ZN => n9486);
   U3190 : OAI22_X1 port map( A1 => n13951, A2 => n13723, B1 => n13721, B2 => 
                           n14290, ZN => n9487);
   U3191 : OAI22_X1 port map( A1 => n13957, A2 => n13723, B1 => n13721, B2 => 
                           n14289, ZN => n9488);
   U3192 : OAI22_X1 port map( A1 => n13963, A2 => n13723, B1 => n13721, B2 => 
                           n14288, ZN => n9489);
   U3193 : OAI22_X1 port map( A1 => n13824, A2 => n13749, B1 => n13744, B2 => 
                           n12661, ZN => n9594);
   U3194 : OAI22_X1 port map( A1 => n13830, A2 => n13749, B1 => n13744, B2 => 
                           n12663, ZN => n9595);
   U3195 : OAI22_X1 port map( A1 => n13836, A2 => n13749, B1 => n13744, B2 => 
                           n12665, ZN => n9596);
   U3196 : OAI22_X1 port map( A1 => n13842, A2 => n13749, B1 => n13744, B2 => 
                           n12667, ZN => n9597);
   U3197 : OAI22_X1 port map( A1 => n13848, A2 => n13749, B1 => n13744, B2 => 
                           n12669, ZN => n9598);
   U3198 : OAI22_X1 port map( A1 => n13854, A2 => n13749, B1 => n13744, B2 => 
                           n12671, ZN => n9599);
   U3199 : OAI22_X1 port map( A1 => n13860, A2 => n13749, B1 => n13744, B2 => 
                           n12673, ZN => n9600);
   U3200 : OAI22_X1 port map( A1 => n13866, A2 => n13749, B1 => n13744, B2 => 
                           n12675, ZN => n9601);
   U3201 : OAI22_X1 port map( A1 => n13872, A2 => n13748, B1 => n13744, B2 => 
                           n12677, ZN => n9602);
   U3202 : OAI22_X1 port map( A1 => n13878, A2 => n13748, B1 => n13744, B2 => 
                           n12679, ZN => n9603);
   U3203 : OAI22_X1 port map( A1 => n13884, A2 => n13748, B1 => n13744, B2 => 
                           n12681, ZN => n9604);
   U3204 : OAI22_X1 port map( A1 => n13890, A2 => n13748, B1 => n13744, B2 => 
                           n12683, ZN => n9605);
   U3205 : OAI22_X1 port map( A1 => n13896, A2 => n13748, B1 => n13745, B2 => 
                           n12685, ZN => n9606);
   U3206 : OAI22_X1 port map( A1 => n13902, A2 => n13748, B1 => n13745, B2 => 
                           n12687, ZN => n9607);
   U3207 : OAI22_X1 port map( A1 => n13908, A2 => n13748, B1 => n13745, B2 => 
                           n12689, ZN => n9608);
   U3208 : OAI22_X1 port map( A1 => n13914, A2 => n13748, B1 => n13745, B2 => 
                           n12691, ZN => n9609);
   U3209 : OAI22_X1 port map( A1 => n13920, A2 => n13748, B1 => n13745, B2 => 
                           n12693, ZN => n9610);
   U3210 : OAI22_X1 port map( A1 => n13926, A2 => n13748, B1 => n13745, B2 => 
                           n12695, ZN => n9611);
   U3211 : OAI22_X1 port map( A1 => n13932, A2 => n13748, B1 => n13745, B2 => 
                           n12697, ZN => n9612);
   U3212 : OAI22_X1 port map( A1 => n13938, A2 => n13748, B1 => n13745, B2 => 
                           n12699, ZN => n9613);
   U3213 : OAI22_X1 port map( A1 => n13944, A2 => n13747, B1 => n13745, B2 => 
                           n12701, ZN => n9614);
   U3214 : OAI22_X1 port map( A1 => n13950, A2 => n13747, B1 => n13745, B2 => 
                           n12703, ZN => n9615);
   U3215 : OAI22_X1 port map( A1 => n13956, A2 => n13747, B1 => n13745, B2 => 
                           n12705, ZN => n9616);
   U3216 : OAI22_X1 port map( A1 => n13962, A2 => n13747, B1 => n13745, B2 => 
                           n12707, ZN => n9617);
   U3217 : OAI22_X1 port map( A1 => n13824, A2 => n13767, B1 => n13762, B2 => 
                           n14203, ZN => n9690);
   U3218 : OAI22_X1 port map( A1 => n13830, A2 => n13767, B1 => n13762, B2 => 
                           n14202, ZN => n9691);
   U3219 : OAI22_X1 port map( A1 => n13836, A2 => n13767, B1 => n13762, B2 => 
                           n14201, ZN => n9692);
   U3220 : OAI22_X1 port map( A1 => n13842, A2 => n13767, B1 => n13762, B2 => 
                           n14200, ZN => n9693);
   U3221 : OAI22_X1 port map( A1 => n13848, A2 => n13767, B1 => n13762, B2 => 
                           n14199, ZN => n9694);
   U3222 : OAI22_X1 port map( A1 => n13854, A2 => n13767, B1 => n13762, B2 => 
                           n14198, ZN => n9695);
   U3223 : OAI22_X1 port map( A1 => n13860, A2 => n13767, B1 => n13762, B2 => 
                           n14197, ZN => n9696);
   U3224 : OAI22_X1 port map( A1 => n13866, A2 => n13767, B1 => n13762, B2 => 
                           n14196, ZN => n9697);
   U3225 : OAI22_X1 port map( A1 => n13872, A2 => n13766, B1 => n13762, B2 => 
                           n14195, ZN => n9698);
   U3226 : OAI22_X1 port map( A1 => n13878, A2 => n13766, B1 => n13762, B2 => 
                           n14194, ZN => n9699);
   U3227 : OAI22_X1 port map( A1 => n13884, A2 => n13766, B1 => n13762, B2 => 
                           n14193, ZN => n9700);
   U3228 : OAI22_X1 port map( A1 => n13890, A2 => n13766, B1 => n13762, B2 => 
                           n14192, ZN => n9701);
   U3229 : OAI22_X1 port map( A1 => n13896, A2 => n13766, B1 => n13763, B2 => 
                           n14191, ZN => n9702);
   U3230 : OAI22_X1 port map( A1 => n13902, A2 => n13766, B1 => n13763, B2 => 
                           n14190, ZN => n9703);
   U3231 : OAI22_X1 port map( A1 => n13908, A2 => n13766, B1 => n13763, B2 => 
                           n14189, ZN => n9704);
   U3232 : OAI22_X1 port map( A1 => n13914, A2 => n13766, B1 => n13763, B2 => 
                           n14188, ZN => n9705);
   U3233 : OAI22_X1 port map( A1 => n13920, A2 => n13766, B1 => n13763, B2 => 
                           n14187, ZN => n9706);
   U3234 : OAI22_X1 port map( A1 => n13926, A2 => n13766, B1 => n13763, B2 => 
                           n14186, ZN => n9707);
   U3235 : OAI22_X1 port map( A1 => n13932, A2 => n13766, B1 => n13763, B2 => 
                           n14185, ZN => n9708);
   U3236 : OAI22_X1 port map( A1 => n13938, A2 => n13766, B1 => n13763, B2 => 
                           n14184, ZN => n9709);
   U3237 : OAI22_X1 port map( A1 => n13944, A2 => n13765, B1 => n13763, B2 => 
                           n14183, ZN => n9710);
   U3238 : OAI22_X1 port map( A1 => n13950, A2 => n13765, B1 => n13763, B2 => 
                           n14182, ZN => n9711);
   U3239 : OAI22_X1 port map( A1 => n13956, A2 => n13765, B1 => n13763, B2 => 
                           n14181, ZN => n9712);
   U3240 : OAI22_X1 port map( A1 => n13962, A2 => n13765, B1 => n13763, B2 => 
                           n14180, ZN => n9713);
   U3241 : OAI22_X1 port map( A1 => n13824, A2 => n13773, B1 => n13768, B2 => 
                           n14171, ZN => n9722);
   U3242 : OAI22_X1 port map( A1 => n13830, A2 => n13773, B1 => n13768, B2 => 
                           n14170, ZN => n9723);
   U3243 : OAI22_X1 port map( A1 => n13836, A2 => n13773, B1 => n13768, B2 => 
                           n14169, ZN => n9724);
   U3244 : OAI22_X1 port map( A1 => n13842, A2 => n13773, B1 => n13768, B2 => 
                           n14168, ZN => n9725);
   U3245 : OAI22_X1 port map( A1 => n13848, A2 => n13773, B1 => n13768, B2 => 
                           n14167, ZN => n9726);
   U3246 : OAI22_X1 port map( A1 => n13854, A2 => n13773, B1 => n13768, B2 => 
                           n14166, ZN => n9727);
   U3247 : OAI22_X1 port map( A1 => n13860, A2 => n13773, B1 => n13768, B2 => 
                           n14165, ZN => n9728);
   U3248 : OAI22_X1 port map( A1 => n13866, A2 => n13773, B1 => n13768, B2 => 
                           n14164, ZN => n9729);
   U3249 : OAI22_X1 port map( A1 => n13872, A2 => n13772, B1 => n13768, B2 => 
                           n14163, ZN => n9730);
   U3250 : OAI22_X1 port map( A1 => n13878, A2 => n13772, B1 => n13768, B2 => 
                           n14162, ZN => n9731);
   U3251 : OAI22_X1 port map( A1 => n13884, A2 => n13772, B1 => n13768, B2 => 
                           n14161, ZN => n9732);
   U3252 : OAI22_X1 port map( A1 => n13890, A2 => n13772, B1 => n13768, B2 => 
                           n14160, ZN => n9733);
   U3253 : OAI22_X1 port map( A1 => n13896, A2 => n13772, B1 => n13769, B2 => 
                           n14159, ZN => n9734);
   U3254 : OAI22_X1 port map( A1 => n13902, A2 => n13772, B1 => n13769, B2 => 
                           n14158, ZN => n9735);
   U3255 : OAI22_X1 port map( A1 => n13908, A2 => n13772, B1 => n13769, B2 => 
                           n14157, ZN => n9736);
   U3256 : OAI22_X1 port map( A1 => n13914, A2 => n13772, B1 => n13769, B2 => 
                           n14156, ZN => n9737);
   U3257 : OAI22_X1 port map( A1 => n13920, A2 => n13772, B1 => n13769, B2 => 
                           n14155, ZN => n9738);
   U3258 : OAI22_X1 port map( A1 => n13926, A2 => n13772, B1 => n13769, B2 => 
                           n14154, ZN => n9739);
   U3259 : OAI22_X1 port map( A1 => n13932, A2 => n13772, B1 => n13769, B2 => 
                           n14153, ZN => n9740);
   U3260 : OAI22_X1 port map( A1 => n13938, A2 => n13772, B1 => n13769, B2 => 
                           n14152, ZN => n9741);
   U3261 : OAI22_X1 port map( A1 => n13944, A2 => n13771, B1 => n13769, B2 => 
                           n14151, ZN => n9742);
   U3262 : OAI22_X1 port map( A1 => n13950, A2 => n13771, B1 => n13769, B2 => 
                           n14150, ZN => n9743);
   U3263 : OAI22_X1 port map( A1 => n13956, A2 => n13771, B1 => n13769, B2 => 
                           n14149, ZN => n9744);
   U3264 : OAI22_X1 port map( A1 => n13962, A2 => n13771, B1 => n13769, B2 => 
                           n14148, ZN => n9745);
   U3265 : OAI22_X1 port map( A1 => n13824, A2 => n13779, B1 => n13774, B2 => 
                           n14139, ZN => n9754);
   U3266 : OAI22_X1 port map( A1 => n13830, A2 => n13779, B1 => n13774, B2 => 
                           n14138, ZN => n9755);
   U3267 : OAI22_X1 port map( A1 => n13836, A2 => n13779, B1 => n13774, B2 => 
                           n14137, ZN => n9756);
   U3268 : OAI22_X1 port map( A1 => n13842, A2 => n13779, B1 => n13774, B2 => 
                           n14136, ZN => n9757);
   U3269 : OAI22_X1 port map( A1 => n13848, A2 => n13779, B1 => n13774, B2 => 
                           n14135, ZN => n9758);
   U3270 : OAI22_X1 port map( A1 => n13854, A2 => n13779, B1 => n13774, B2 => 
                           n14134, ZN => n9759);
   U3271 : OAI22_X1 port map( A1 => n13860, A2 => n13779, B1 => n13774, B2 => 
                           n14133, ZN => n9760);
   U3272 : OAI22_X1 port map( A1 => n13866, A2 => n13779, B1 => n13774, B2 => 
                           n14132, ZN => n9761);
   U3273 : OAI22_X1 port map( A1 => n13872, A2 => n13778, B1 => n13774, B2 => 
                           n14131, ZN => n9762);
   U3274 : OAI22_X1 port map( A1 => n13878, A2 => n13778, B1 => n13774, B2 => 
                           n14130, ZN => n9763);
   U3275 : OAI22_X1 port map( A1 => n13884, A2 => n13778, B1 => n13774, B2 => 
                           n14129, ZN => n9764);
   U3276 : OAI22_X1 port map( A1 => n13890, A2 => n13778, B1 => n13774, B2 => 
                           n14128, ZN => n9765);
   U3277 : OAI22_X1 port map( A1 => n13896, A2 => n13778, B1 => n13775, B2 => 
                           n14127, ZN => n9766);
   U3278 : OAI22_X1 port map( A1 => n13902, A2 => n13778, B1 => n13775, B2 => 
                           n14126, ZN => n9767);
   U3279 : OAI22_X1 port map( A1 => n13908, A2 => n13778, B1 => n13775, B2 => 
                           n14125, ZN => n9768);
   U3280 : OAI22_X1 port map( A1 => n13914, A2 => n13778, B1 => n13775, B2 => 
                           n14124, ZN => n9769);
   U3281 : OAI22_X1 port map( A1 => n13920, A2 => n13778, B1 => n13775, B2 => 
                           n14123, ZN => n9770);
   U3282 : OAI22_X1 port map( A1 => n13926, A2 => n13778, B1 => n13775, B2 => 
                           n14122, ZN => n9771);
   U3283 : OAI22_X1 port map( A1 => n13932, A2 => n13778, B1 => n13775, B2 => 
                           n14121, ZN => n9772);
   U3284 : OAI22_X1 port map( A1 => n13938, A2 => n13778, B1 => n13775, B2 => 
                           n14120, ZN => n9773);
   U3285 : OAI22_X1 port map( A1 => n13944, A2 => n13777, B1 => n13775, B2 => 
                           n14119, ZN => n9774);
   U3286 : OAI22_X1 port map( A1 => n13950, A2 => n13777, B1 => n13775, B2 => 
                           n14118, ZN => n9775);
   U3287 : OAI22_X1 port map( A1 => n13956, A2 => n13777, B1 => n13775, B2 => 
                           n14117, ZN => n9776);
   U3288 : OAI22_X1 port map( A1 => n13962, A2 => n13777, B1 => n13775, B2 => 
                           n14116, ZN => n9777);
   U3289 : OAI22_X1 port map( A1 => n13824, A2 => n13803, B1 => n13798, B2 => 
                           n12662, ZN => n9882);
   U3290 : OAI22_X1 port map( A1 => n13830, A2 => n13803, B1 => n13798, B2 => 
                           n12664, ZN => n9883);
   U3291 : OAI22_X1 port map( A1 => n13836, A2 => n13803, B1 => n13798, B2 => 
                           n12666, ZN => n9884);
   U3292 : OAI22_X1 port map( A1 => n13842, A2 => n13803, B1 => n13798, B2 => 
                           n12668, ZN => n9885);
   U3293 : OAI22_X1 port map( A1 => n13848, A2 => n13803, B1 => n13798, B2 => 
                           n12670, ZN => n9886);
   U3294 : OAI22_X1 port map( A1 => n13854, A2 => n13803, B1 => n13798, B2 => 
                           n12672, ZN => n9887);
   U3295 : OAI22_X1 port map( A1 => n13860, A2 => n13803, B1 => n13798, B2 => 
                           n12674, ZN => n9888);
   U3296 : OAI22_X1 port map( A1 => n13866, A2 => n13803, B1 => n13798, B2 => 
                           n12676, ZN => n9889);
   U3297 : OAI22_X1 port map( A1 => n13872, A2 => n13802, B1 => n13798, B2 => 
                           n12678, ZN => n9890);
   U3298 : OAI22_X1 port map( A1 => n13878, A2 => n13802, B1 => n13798, B2 => 
                           n12680, ZN => n9891);
   U3299 : OAI22_X1 port map( A1 => n13884, A2 => n13802, B1 => n13798, B2 => 
                           n12682, ZN => n9892);
   U3300 : OAI22_X1 port map( A1 => n13890, A2 => n13802, B1 => n13798, B2 => 
                           n12684, ZN => n9893);
   U3301 : OAI22_X1 port map( A1 => n13896, A2 => n13802, B1 => n13799, B2 => 
                           n12686, ZN => n9894);
   U3302 : OAI22_X1 port map( A1 => n13902, A2 => n13802, B1 => n13799, B2 => 
                           n12688, ZN => n9895);
   U3303 : OAI22_X1 port map( A1 => n13908, A2 => n13802, B1 => n13799, B2 => 
                           n12690, ZN => n9896);
   U3304 : OAI22_X1 port map( A1 => n13914, A2 => n13802, B1 => n13799, B2 => 
                           n12692, ZN => n9897);
   U3305 : OAI22_X1 port map( A1 => n13920, A2 => n13802, B1 => n13799, B2 => 
                           n12694, ZN => n9898);
   U3306 : OAI22_X1 port map( A1 => n13926, A2 => n13802, B1 => n13799, B2 => 
                           n12696, ZN => n9899);
   U3307 : OAI22_X1 port map( A1 => n13932, A2 => n13802, B1 => n13799, B2 => 
                           n12698, ZN => n9900);
   U3308 : OAI22_X1 port map( A1 => n13938, A2 => n13802, B1 => n13799, B2 => 
                           n12700, ZN => n9901);
   U3309 : OAI22_X1 port map( A1 => n13944, A2 => n13801, B1 => n13799, B2 => 
                           n12702, ZN => n9902);
   U3310 : OAI22_X1 port map( A1 => n13950, A2 => n13801, B1 => n13799, B2 => 
                           n12704, ZN => n9903);
   U3311 : OAI22_X1 port map( A1 => n13956, A2 => n13801, B1 => n13799, B2 => 
                           n12706, ZN => n9904);
   U3312 : OAI22_X1 port map( A1 => n13962, A2 => n13801, B1 => n13799, B2 => 
                           n12708, ZN => n9905);
   U3313 : OAI22_X1 port map( A1 => n13387, A2 => n15548, B1 => n13878, B2 => 
                           n13385, ZN => n7683);
   U3314 : OAI22_X1 port map( A1 => n13387, A2 => n15547, B1 => n13884, B2 => 
                           n13385, ZN => n7684);
   U3315 : OAI22_X1 port map( A1 => n13387, A2 => n15546, B1 => n13890, B2 => 
                           n13385, ZN => n7685);
   U3316 : OAI22_X1 port map( A1 => n13388, A2 => n15545, B1 => n13896, B2 => 
                           n13385, ZN => n7686);
   U3317 : OAI22_X1 port map( A1 => n13388, A2 => n15544, B1 => n13902, B2 => 
                           n13385, ZN => n7687);
   U3318 : OAI22_X1 port map( A1 => n13388, A2 => n15543, B1 => n13908, B2 => 
                           n13385, ZN => n7688);
   U3319 : OAI22_X1 port map( A1 => n13388, A2 => n15542, B1 => n13914, B2 => 
                           n13385, ZN => n7689);
   U3320 : OAI22_X1 port map( A1 => n13388, A2 => n15541, B1 => n13920, B2 => 
                           n13385, ZN => n7690);
   U3321 : OAI22_X1 port map( A1 => n13388, A2 => n15540, B1 => n13926, B2 => 
                           n13385, ZN => n7691);
   U3322 : OAI22_X1 port map( A1 => n13388, A2 => n15539, B1 => n13932, B2 => 
                           n13385, ZN => n7692);
   U3323 : OAI22_X1 port map( A1 => n13388, A2 => n15538, B1 => n13938, B2 => 
                           n13385, ZN => n7693);
   U3324 : OAI22_X1 port map( A1 => n13388, A2 => n15537, B1 => n13944, B2 => 
                           n13384, ZN => n7694);
   U3325 : OAI22_X1 port map( A1 => n13388, A2 => n15536, B1 => n13950, B2 => 
                           n13384, ZN => n7695);
   U3326 : OAI22_X1 port map( A1 => n13388, A2 => n15535, B1 => n13956, B2 => 
                           n13384, ZN => n7696);
   U3327 : OAI22_X1 port map( A1 => n13388, A2 => n15534, B1 => n13962, B2 => 
                           n13384, ZN => n7697);
   U3328 : OAI22_X1 port map( A1 => n13389, A2 => n15533, B1 => n13968, B2 => 
                           n13384, ZN => n7698);
   U3329 : OAI22_X1 port map( A1 => n13389, A2 => n15532, B1 => n13974, B2 => 
                           n13384, ZN => n7699);
   U3330 : OAI22_X1 port map( A1 => n13389, A2 => n15531, B1 => n13980, B2 => 
                           n13384, ZN => n7700);
   U3331 : OAI22_X1 port map( A1 => n13389, A2 => n15530, B1 => n13986, B2 => 
                           n13384, ZN => n7701);
   U3332 : OAI22_X1 port map( A1 => n13389, A2 => n15529, B1 => n13992, B2 => 
                           n13384, ZN => n7702);
   U3333 : OAI22_X1 port map( A1 => n13389, A2 => n15528, B1 => n13998, B2 => 
                           n13384, ZN => n7703);
   U3334 : OAI22_X1 port map( A1 => n13389, A2 => n15527, B1 => n14004, B2 => 
                           n13384, ZN => n7704);
   U3335 : OAI22_X1 port map( A1 => n13389, A2 => n15526, B1 => n14013, B2 => 
                           n13385, ZN => n7705);
   U3336 : NAND4_X1 port map( A1 => n3229, A2 => n3230, A3 => n3231, A4 => 
                           n3232, ZN => n3228);
   U3337 : AOI221_X1 port map( B1 => n13329, B2 => n14047, C1 => n13326, C2 => 
                           n14031, A => n3236, ZN => n3229);
   U3338 : AOI221_X1 port map( B1 => n13356, B2 => n14219, C1 => n13353, C2 => 
                           n14207, A => n3234, ZN => n3231);
   U3339 : AOI221_X1 port map( B1 => n13344, B2 => n14079, C1 => n13341, C2 => 
                           n15601, A => n3235, ZN => n3230);
   U3340 : NAND4_X1 port map( A1 => n3192, A2 => n3193, A3 => n3194, A4 => 
                           n3195, ZN => n3191);
   U3341 : AOI221_X1 port map( B1 => n13329, B2 => n14046, C1 => n13326, C2 => 
                           n14030, A => n3199, ZN => n3192);
   U3342 : AOI221_X1 port map( B1 => n13356, B2 => n14218, C1 => n13353, C2 => 
                           n14206, A => n3197, ZN => n3194);
   U3343 : AOI221_X1 port map( B1 => n13344, B2 => n14078, C1 => n13341, C2 => 
                           n15600, A => n3198, ZN => n3193);
   U3344 : NAND4_X1 port map( A1 => n3155, A2 => n3156, A3 => n3157, A4 => 
                           n3158, ZN => n3154);
   U3345 : AOI221_X1 port map( B1 => n13329, B2 => n14045, C1 => n13326, C2 => 
                           n14029, A => n3162, ZN => n3155);
   U3346 : AOI221_X1 port map( B1 => n13356, B2 => n14217, C1 => n13353, C2 => 
                           n14205, A => n3160, ZN => n3157);
   U3347 : AOI221_X1 port map( B1 => n13344, B2 => n14077, C1 => n13341, C2 => 
                           n15599, A => n3161, ZN => n3156);
   U3348 : NAND4_X1 port map( A1 => n3046, A2 => n3047, A3 => n3048, A4 => 
                           n3049, ZN => n3045);
   U3349 : AOI221_X1 port map( B1 => n13329, B2 => n14044, C1 => n13326, C2 => 
                           n14028, A => n3069, ZN => n3046);
   U3350 : AOI221_X1 port map( B1 => n13356, B2 => n14216, C1 => n13353, C2 => 
                           n14204, A => n3058, ZN => n3048);
   U3351 : AOI221_X1 port map( B1 => n13344, B2 => n14076, C1 => n13341, C2 => 
                           n15598, A => n3063, ZN => n3047);
   U3352 : NAND4_X1 port map( A1 => n4265, A2 => n4266, A3 => n4267, A4 => 
                           n4268, ZN => n4264);
   U3353 : AOI221_X1 port map( B1 => n13327, B2 => n14075, C1 => n13324, C2 => 
                           n16042, A => n4283, ZN => n4265);
   U3354 : AOI221_X1 port map( B1 => n13354, B2 => n14247, C1 => n13351, C2 => 
                           n16006, A => n4277, ZN => n4267);
   U3355 : AOI221_X1 port map( B1 => n13342, B2 => n14107, C1 => n13339, C2 => 
                           n15921, A => n4281, ZN => n4266);
   U3356 : NAND4_X1 port map( A1 => n4228, A2 => n4229, A3 => n4230, A4 => 
                           n4231, ZN => n4227);
   U3357 : AOI221_X1 port map( B1 => n13327, B2 => n14074, C1 => n13324, C2 => 
                           n16041, A => n4235, ZN => n4228);
   U3358 : AOI221_X1 port map( B1 => n13354, B2 => n14246, C1 => n13351, C2 => 
                           n16005, A => n4233, ZN => n4230);
   U3359 : AOI221_X1 port map( B1 => n13342, B2 => n14106, C1 => n13339, C2 => 
                           n15920, A => n4234, ZN => n4229);
   U3360 : NAND4_X1 port map( A1 => n4191, A2 => n4192, A3 => n4193, A4 => 
                           n4194, ZN => n4190);
   U3361 : AOI221_X1 port map( B1 => n13327, B2 => n14073, C1 => n13324, C2 => 
                           n16040, A => n4198, ZN => n4191);
   U3362 : AOI221_X1 port map( B1 => n13354, B2 => n14245, C1 => n13351, C2 => 
                           n16004, A => n4196, ZN => n4193);
   U3363 : AOI221_X1 port map( B1 => n13342, B2 => n14105, C1 => n13339, C2 => 
                           n15919, A => n4197, ZN => n4192);
   U3364 : NAND4_X1 port map( A1 => n4154, A2 => n4155, A3 => n4156, A4 => 
                           n4157, ZN => n4153);
   U3365 : AOI221_X1 port map( B1 => n13327, B2 => n14072, C1 => n13324, C2 => 
                           n16039, A => n4161, ZN => n4154);
   U3366 : AOI221_X1 port map( B1 => n13354, B2 => n14244, C1 => n13351, C2 => 
                           n16003, A => n4159, ZN => n4156);
   U3367 : AOI221_X1 port map( B1 => n13342, B2 => n14104, C1 => n13339, C2 => 
                           n15918, A => n4160, ZN => n4155);
   U3368 : NAND4_X1 port map( A1 => n4117, A2 => n4118, A3 => n4119, A4 => 
                           n4120, ZN => n4116);
   U3369 : AOI221_X1 port map( B1 => n13327, B2 => n14071, C1 => n13324, C2 => 
                           n16038, A => n4124, ZN => n4117);
   U3370 : AOI221_X1 port map( B1 => n13354, B2 => n14243, C1 => n13351, C2 => 
                           n16002, A => n4122, ZN => n4119);
   U3371 : AOI221_X1 port map( B1 => n13342, B2 => n14103, C1 => n13339, C2 => 
                           n15917, A => n4123, ZN => n4118);
   U3372 : NAND4_X1 port map( A1 => n4080, A2 => n4081, A3 => n4082, A4 => 
                           n4083, ZN => n4079);
   U3373 : AOI221_X1 port map( B1 => n13327, B2 => n14070, C1 => n13324, C2 => 
                           n16037, A => n4087, ZN => n4080);
   U3374 : AOI221_X1 port map( B1 => n13354, B2 => n14242, C1 => n13351, C2 => 
                           n16001, A => n4085, ZN => n4082);
   U3375 : AOI221_X1 port map( B1 => n13342, B2 => n14102, C1 => n13339, C2 => 
                           n15916, A => n4086, ZN => n4081);
   U3376 : NAND4_X1 port map( A1 => n4043, A2 => n4044, A3 => n4045, A4 => 
                           n4046, ZN => n4042);
   U3377 : AOI221_X1 port map( B1 => n13327, B2 => n14069, C1 => n13324, C2 => 
                           n16036, A => n4050, ZN => n4043);
   U3378 : AOI221_X1 port map( B1 => n13354, B2 => n14241, C1 => n13351, C2 => 
                           n16000, A => n4048, ZN => n4045);
   U3379 : AOI221_X1 port map( B1 => n13342, B2 => n14101, C1 => n13339, C2 => 
                           n15915, A => n4049, ZN => n4044);
   U3380 : NAND4_X1 port map( A1 => n4006, A2 => n4007, A3 => n4008, A4 => 
                           n4009, ZN => n4005);
   U3381 : AOI221_X1 port map( B1 => n13327, B2 => n14068, C1 => n13324, C2 => 
                           n16035, A => n4013, ZN => n4006);
   U3382 : AOI221_X1 port map( B1 => n13354, B2 => n14240, C1 => n13351, C2 => 
                           n15999, A => n4011, ZN => n4008);
   U3383 : AOI221_X1 port map( B1 => n13342, B2 => n14100, C1 => n13339, C2 => 
                           n15914, A => n4012, ZN => n4007);
   U3384 : NAND4_X1 port map( A1 => n3969, A2 => n3970, A3 => n3971, A4 => 
                           n3972, ZN => n3968);
   U3385 : AOI221_X1 port map( B1 => n13327, B2 => n14067, C1 => n13324, C2 => 
                           n16034, A => n3976, ZN => n3969);
   U3386 : AOI221_X1 port map( B1 => n13354, B2 => n14239, C1 => n13351, C2 => 
                           n15998, A => n3974, ZN => n3971);
   U3387 : AOI221_X1 port map( B1 => n13342, B2 => n14099, C1 => n13339, C2 => 
                           n15913, A => n3975, ZN => n3970);
   U3388 : NAND4_X1 port map( A1 => n3932, A2 => n3933, A3 => n3934, A4 => 
                           n3935, ZN => n3931);
   U3389 : AOI221_X1 port map( B1 => n13327, B2 => n14066, C1 => n13324, C2 => 
                           n16033, A => n3939, ZN => n3932);
   U3390 : AOI221_X1 port map( B1 => n13354, B2 => n14238, C1 => n13351, C2 => 
                           n15997, A => n3937, ZN => n3934);
   U3391 : AOI221_X1 port map( B1 => n13342, B2 => n14098, C1 => n13339, C2 => 
                           n15912, A => n3938, ZN => n3933);
   U3392 : NAND4_X1 port map( A1 => n3895, A2 => n3896, A3 => n3897, A4 => 
                           n3898, ZN => n3894);
   U3393 : AOI221_X1 port map( B1 => n13327, B2 => n14065, C1 => n13324, C2 => 
                           n16032, A => n3902, ZN => n3895);
   U3394 : AOI221_X1 port map( B1 => n13354, B2 => n14237, C1 => n13351, C2 => 
                           n15996, A => n3900, ZN => n3897);
   U3395 : AOI221_X1 port map( B1 => n13342, B2 => n14097, C1 => n13339, C2 => 
                           n15911, A => n3901, ZN => n3896);
   U3396 : NAND4_X1 port map( A1 => n3858, A2 => n3859, A3 => n3860, A4 => 
                           n3861, ZN => n3857);
   U3397 : AOI221_X1 port map( B1 => n13327, B2 => n14064, C1 => n13324, C2 => 
                           n16031, A => n3865, ZN => n3858);
   U3398 : AOI221_X1 port map( B1 => n13354, B2 => n14236, C1 => n13351, C2 => 
                           n15995, A => n3863, ZN => n3860);
   U3399 : AOI221_X1 port map( B1 => n13342, B2 => n14096, C1 => n13339, C2 => 
                           n15910, A => n3864, ZN => n3859);
   U3400 : NAND4_X1 port map( A1 => n3821, A2 => n3822, A3 => n3823, A4 => 
                           n3824, ZN => n3820);
   U3401 : AOI221_X1 port map( B1 => n13328, B2 => n14063, C1 => n13325, C2 => 
                           n16054, A => n3828, ZN => n3821);
   U3402 : AOI221_X1 port map( B1 => n13355, B2 => n14235, C1 => n13352, C2 => 
                           n16050, A => n3826, ZN => n3823);
   U3403 : AOI221_X1 port map( B1 => n13343, B2 => n14095, C1 => n13340, C2 => 
                           n15909, A => n3827, ZN => n3822);
   U3404 : NAND4_X1 port map( A1 => n3784, A2 => n3785, A3 => n3786, A4 => 
                           n3787, ZN => n3783);
   U3405 : AOI221_X1 port map( B1 => n13328, B2 => n14062, C1 => n13325, C2 => 
                           n16053, A => n3791, ZN => n3784);
   U3406 : AOI221_X1 port map( B1 => n13355, B2 => n14234, C1 => n13352, C2 => 
                           n16049, A => n3789, ZN => n3786);
   U3407 : AOI221_X1 port map( B1 => n13343, B2 => n14094, C1 => n13340, C2 => 
                           n15908, A => n3790, ZN => n3785);
   U3408 : NAND4_X1 port map( A1 => n3747, A2 => n3748, A3 => n3749, A4 => 
                           n3750, ZN => n3746);
   U3409 : AOI221_X1 port map( B1 => n13328, B2 => n14061, C1 => n13325, C2 => 
                           n16052, A => n3754, ZN => n3747);
   U3410 : AOI221_X1 port map( B1 => n13355, B2 => n14233, C1 => n13352, C2 => 
                           n16048, A => n3752, ZN => n3749);
   U3411 : AOI221_X1 port map( B1 => n13343, B2 => n14093, C1 => n13340, C2 => 
                           n15907, A => n3753, ZN => n3748);
   U3412 : NAND4_X1 port map( A1 => n3710, A2 => n3711, A3 => n3712, A4 => 
                           n3713, ZN => n3709);
   U3413 : AOI221_X1 port map( B1 => n13328, B2 => n14060, C1 => n13325, C2 => 
                           n16051, A => n3717, ZN => n3710);
   U3414 : AOI221_X1 port map( B1 => n13355, B2 => n14232, C1 => n13352, C2 => 
                           n16047, A => n3715, ZN => n3712);
   U3415 : AOI221_X1 port map( B1 => n13343, B2 => n14092, C1 => n13340, C2 => 
                           n15906, A => n3716, ZN => n3711);
   U3416 : NAND4_X1 port map( A1 => n3673, A2 => n3674, A3 => n3675, A4 => 
                           n3676, ZN => n3672);
   U3417 : AOI221_X1 port map( B1 => n13328, B2 => n14059, C1 => n13325, C2 => 
                           n14043, A => n3680, ZN => n3673);
   U3418 : AOI221_X1 port map( B1 => n13355, B2 => n14231, C1 => n13352, C2 => 
                           n16046, A => n3678, ZN => n3675);
   U3419 : AOI221_X1 port map( B1 => n13343, B2 => n14091, C1 => n13340, C2 => 
                           n15905, A => n3679, ZN => n3674);
   U3420 : NAND4_X1 port map( A1 => n3636, A2 => n3637, A3 => n3638, A4 => 
                           n3639, ZN => n3635);
   U3421 : AOI221_X1 port map( B1 => n13328, B2 => n14058, C1 => n13325, C2 => 
                           n14042, A => n3643, ZN => n3636);
   U3422 : AOI221_X1 port map( B1 => n13355, B2 => n14230, C1 => n13352, C2 => 
                           n16045, A => n3641, ZN => n3638);
   U3423 : AOI221_X1 port map( B1 => n13343, B2 => n14090, C1 => n13340, C2 => 
                           n15904, A => n3642, ZN => n3637);
   U3424 : NAND4_X1 port map( A1 => n3599, A2 => n3600, A3 => n3601, A4 => 
                           n3602, ZN => n3598);
   U3425 : AOI221_X1 port map( B1 => n13328, B2 => n14057, C1 => n13325, C2 => 
                           n14041, A => n3606, ZN => n3599);
   U3426 : AOI221_X1 port map( B1 => n13355, B2 => n14229, C1 => n13352, C2 => 
                           n16044, A => n3604, ZN => n3601);
   U3427 : AOI221_X1 port map( B1 => n13343, B2 => n14089, C1 => n13340, C2 => 
                           n15903, A => n3605, ZN => n3600);
   U3428 : NAND4_X1 port map( A1 => n3562, A2 => n3563, A3 => n3564, A4 => 
                           n3565, ZN => n3561);
   U3429 : AOI221_X1 port map( B1 => n13328, B2 => n14056, C1 => n13325, C2 => 
                           n14040, A => n3569, ZN => n3562);
   U3430 : AOI221_X1 port map( B1 => n13355, B2 => n14228, C1 => n13352, C2 => 
                           n16043, A => n3567, ZN => n3564);
   U3431 : AOI221_X1 port map( B1 => n13343, B2 => n14088, C1 => n13340, C2 => 
                           n15902, A => n3568, ZN => n3563);
   U3432 : NAND4_X1 port map( A1 => n3525, A2 => n3526, A3 => n3527, A4 => 
                           n3528, ZN => n3524);
   U3433 : AOI221_X1 port map( B1 => n13328, B2 => n14055, C1 => n13325, C2 => 
                           n14039, A => n3532, ZN => n3525);
   U3434 : AOI221_X1 port map( B1 => n13355, B2 => n14227, C1 => n13352, C2 => 
                           n14215, A => n3530, ZN => n3527);
   U3435 : AOI221_X1 port map( B1 => n13343, B2 => n14087, C1 => n13340, C2 => 
                           n15901, A => n3531, ZN => n3526);
   U3436 : NAND4_X1 port map( A1 => n3488, A2 => n3489, A3 => n3490, A4 => 
                           n3491, ZN => n3487);
   U3437 : AOI221_X1 port map( B1 => n13328, B2 => n14054, C1 => n13325, C2 => 
                           n14038, A => n3495, ZN => n3488);
   U3438 : AOI221_X1 port map( B1 => n13355, B2 => n14226, C1 => n13352, C2 => 
                           n14214, A => n3493, ZN => n3490);
   U3439 : AOI221_X1 port map( B1 => n13343, B2 => n14086, C1 => n13340, C2 => 
                           n15900, A => n3494, ZN => n3489);
   U3440 : NAND4_X1 port map( A1 => n3451, A2 => n3452, A3 => n3453, A4 => 
                           n3454, ZN => n3450);
   U3441 : AOI221_X1 port map( B1 => n13328, B2 => n14053, C1 => n13325, C2 => 
                           n14037, A => n3458, ZN => n3451);
   U3442 : AOI221_X1 port map( B1 => n13355, B2 => n14225, C1 => n13352, C2 => 
                           n14213, A => n3456, ZN => n3453);
   U3443 : AOI221_X1 port map( B1 => n13343, B2 => n14085, C1 => n13340, C2 => 
                           n15899, A => n3457, ZN => n3452);
   U3444 : NAND4_X1 port map( A1 => n3414, A2 => n3415, A3 => n3416, A4 => 
                           n3417, ZN => n3413);
   U3445 : AOI221_X1 port map( B1 => n13328, B2 => n14052, C1 => n13325, C2 => 
                           n14036, A => n3421, ZN => n3414);
   U3446 : AOI221_X1 port map( B1 => n13355, B2 => n14224, C1 => n13352, C2 => 
                           n14212, A => n3419, ZN => n3416);
   U3447 : AOI221_X1 port map( B1 => n13343, B2 => n14084, C1 => n13340, C2 => 
                           n15898, A => n3420, ZN => n3415);
   U3448 : NAND4_X1 port map( A1 => n3377, A2 => n3378, A3 => n3379, A4 => 
                           n3380, ZN => n3376);
   U3449 : AOI221_X1 port map( B1 => n13329, B2 => n14051, C1 => n13326, C2 => 
                           n14035, A => n3384, ZN => n3377);
   U3450 : AOI221_X1 port map( B1 => n13356, B2 => n14223, C1 => n13353, C2 => 
                           n14211, A => n3382, ZN => n3379);
   U3451 : AOI221_X1 port map( B1 => n13344, B2 => n14083, C1 => n13341, C2 => 
                           n15605, A => n3383, ZN => n3378);
   U3452 : NAND4_X1 port map( A1 => n3340, A2 => n3341, A3 => n3342, A4 => 
                           n3343, ZN => n3339);
   U3453 : AOI221_X1 port map( B1 => n13329, B2 => n14050, C1 => n13326, C2 => 
                           n14034, A => n3347, ZN => n3340);
   U3454 : AOI221_X1 port map( B1 => n13356, B2 => n14222, C1 => n13353, C2 => 
                           n14210, A => n3345, ZN => n3342);
   U3455 : AOI221_X1 port map( B1 => n13344, B2 => n14082, C1 => n13341, C2 => 
                           n15604, A => n3346, ZN => n3341);
   U3456 : NAND4_X1 port map( A1 => n3303, A2 => n3304, A3 => n3305, A4 => 
                           n3306, ZN => n3302);
   U3457 : AOI221_X1 port map( B1 => n13329, B2 => n14049, C1 => n13326, C2 => 
                           n14033, A => n3310, ZN => n3303);
   U3458 : AOI221_X1 port map( B1 => n13356, B2 => n14221, C1 => n13353, C2 => 
                           n14209, A => n3308, ZN => n3305);
   U3459 : AOI221_X1 port map( B1 => n13344, B2 => n14081, C1 => n13341, C2 => 
                           n15603, A => n3309, ZN => n3304);
   U3460 : NAND4_X1 port map( A1 => n3266, A2 => n3267, A3 => n3268, A4 => 
                           n3269, ZN => n3265);
   U3461 : AOI221_X1 port map( B1 => n13329, B2 => n14048, C1 => n13326, C2 => 
                           n14032, A => n3273, ZN => n3266);
   U3462 : AOI221_X1 port map( B1 => n13356, B2 => n14220, C1 => n13353, C2 => 
                           n14208, A => n3271, ZN => n3268);
   U3463 : AOI221_X1 port map( B1 => n13344, B2 => n14080, C1 => n13341, C2 => 
                           n15602, A => n3272, ZN => n3267);
   U3464 : NAND4_X1 port map( A1 => n3237, A2 => n3238, A3 => n3239, A4 => 
                           n3240, ZN => n3227);
   U3465 : AOI221_X1 port map( B1 => n13275, B2 => n15865, C1 => n13272, C2 => 
                           n15628, A => n3244, ZN => n3237);
   U3466 : AOI221_X1 port map( B1 => n13302, B2 => n15577, C1 => n13299, C2 => 
                           n15793, A => n3242, ZN => n3239);
   U3467 : AOI221_X1 port map( B1 => n13290, B2 => n14464, C1 => n13287, C2 => 
                           n15585, A => n3243, ZN => n3238);
   U3468 : NAND4_X1 port map( A1 => n3200, A2 => n3201, A3 => n3202, A4 => 
                           n3203, ZN => n3190);
   U3469 : AOI221_X1 port map( B1 => n13275, B2 => n15864, C1 => n13272, C2 => 
                           n15627, A => n3207, ZN => n3200);
   U3470 : AOI221_X1 port map( B1 => n13302, B2 => n15576, C1 => n13299, C2 => 
                           n15792, A => n3205, ZN => n3202);
   U3471 : AOI221_X1 port map( B1 => n13290, B2 => n14463, C1 => n13287, C2 => 
                           n15584, A => n3206, ZN => n3201);
   U3472 : NAND4_X1 port map( A1 => n4632, A2 => n4633, A3 => n4634, A4 => 
                           n4635, ZN => n4622);
   U3473 : AOI221_X1 port map( B1 => n13047, B2 => n15868, C1 => n13044, C2 => 
                           n15631, A => n4639, ZN => n4632);
   U3474 : AOI221_X1 port map( B1 => n13074, B2 => n15796, C1 => n13071, C2 => 
                           n15580, A => n4637, ZN => n4634);
   U3475 : AOI221_X1 port map( B1 => n13062, B2 => n14467, C1 => n13059, C2 => 
                           n15588, A => n4638, ZN => n4633);
   U3476 : NAND4_X1 port map( A1 => n4595, A2 => n4596, A3 => n4597, A4 => 
                           n4598, ZN => n4585);
   U3477 : AOI221_X1 port map( B1 => n13047, B2 => n15867, C1 => n13044, C2 => 
                           n15630, A => n4602, ZN => n4595);
   U3478 : AOI221_X1 port map( B1 => n13074, B2 => n15795, C1 => n13071, C2 => 
                           n15579, A => n4600, ZN => n4597);
   U3479 : AOI221_X1 port map( B1 => n13062, B2 => n14466, C1 => n13059, C2 => 
                           n15587, A => n4601, ZN => n4596);
   U3480 : NAND4_X1 port map( A1 => n4558, A2 => n4559, A3 => n4560, A4 => 
                           n4561, ZN => n4548);
   U3481 : AOI221_X1 port map( B1 => n13047, B2 => n15866, C1 => n13044, C2 => 
                           n15629, A => n4565, ZN => n4558);
   U3482 : AOI221_X1 port map( B1 => n13074, B2 => n15794, C1 => n13071, C2 => 
                           n15578, A => n4563, ZN => n4560);
   U3483 : AOI221_X1 port map( B1 => n13062, B2 => n14465, C1 => n13059, C2 => 
                           n15586, A => n4564, ZN => n4559);
   U3484 : NAND4_X1 port map( A1 => n4521, A2 => n4522, A3 => n4523, A4 => 
                           n4524, ZN => n4511);
   U3485 : AOI221_X1 port map( B1 => n13047, B2 => n15865, C1 => n13044, C2 => 
                           n15628, A => n4528, ZN => n4521);
   U3486 : AOI221_X1 port map( B1 => n13074, B2 => n15793, C1 => n13071, C2 => 
                           n15577, A => n4526, ZN => n4523);
   U3487 : AOI221_X1 port map( B1 => n13062, B2 => n14464, C1 => n13059, C2 => 
                           n15585, A => n4527, ZN => n4522);
   U3488 : NAND4_X1 port map( A1 => n4484, A2 => n4485, A3 => n4486, A4 => 
                           n4487, ZN => n4474);
   U3489 : AOI221_X1 port map( B1 => n13047, B2 => n15864, C1 => n13044, C2 => 
                           n15627, A => n4491, ZN => n4484);
   U3490 : AOI221_X1 port map( B1 => n13074, B2 => n15792, C1 => n13071, C2 => 
                           n15576, A => n4489, ZN => n4486);
   U3491 : AOI221_X1 port map( B1 => n13062, B2 => n14463, C1 => n13059, C2 => 
                           n15584, A => n4490, ZN => n4485);
   U3492 : NAND4_X1 port map( A1 => n5681, A2 => n5684, A3 => n5686, A4 => 
                           n5688, ZN => n5648);
   U3493 : AOI221_X1 port map( B1 => n13045, B2 => n14458, C1 => n13042, C2 => 
                           n15861, A => n5698, ZN => n5681);
   U3494 : AOI221_X1 port map( B1 => n13072, B2 => n14659, C1 => n13069, C2 => 
                           n15789, A => n5694, ZN => n5686);
   U3495 : AOI221_X1 port map( B1 => n13060, B2 => n14492, C1 => n13057, C2 => 
                           n15837, A => n5696, ZN => n5684);
   U3496 : NAND4_X1 port map( A1 => n5601, A2 => n5604, A3 => n5606, A4 => 
                           n5608, ZN => n5586);
   U3497 : AOI221_X1 port map( B1 => n13045, B2 => n14457, C1 => n13042, C2 => 
                           n15860, A => n5614, ZN => n5601);
   U3498 : AOI221_X1 port map( B1 => n13072, B2 => n14658, C1 => n13069, C2 => 
                           n15788, A => n5610, ZN => n5606);
   U3499 : AOI221_X1 port map( B1 => n13060, B2 => n14491, C1 => n13057, C2 => 
                           n15836, A => n5611, ZN => n5604);
   U3500 : NAND4_X1 port map( A1 => n5540, A2 => n5541, A3 => n5544, A4 => 
                           n5546, ZN => n5524);
   U3501 : AOI221_X1 port map( B1 => n13045, B2 => n14456, C1 => n13042, C2 => 
                           n15859, A => n5551, ZN => n5540);
   U3502 : AOI221_X1 port map( B1 => n13072, B2 => n14657, C1 => n13069, C2 => 
                           n15787, A => n5549, ZN => n5544);
   U3503 : AOI221_X1 port map( B1 => n13060, B2 => n14490, C1 => n13057, C2 => 
                           n15835, A => n5550, ZN => n5541);
   U3504 : NAND4_X1 port map( A1 => n5479, A2 => n5480, A3 => n5481, A4 => 
                           n5484, ZN => n5461);
   U3505 : AOI221_X1 port map( B1 => n13045, B2 => n14455, C1 => n13042, C2 => 
                           n15858, A => n5490, ZN => n5479);
   U3506 : AOI221_X1 port map( B1 => n13072, B2 => n14656, C1 => n13069, C2 => 
                           n15786, A => n5488, ZN => n5481);
   U3507 : AOI221_X1 port map( B1 => n13060, B2 => n14489, C1 => n13057, C2 => 
                           n15834, A => n5489, ZN => n5480);
   U3508 : NAND4_X1 port map( A1 => n5421, A2 => n5422, A3 => n5424, A4 => 
                           n5426, ZN => n5408);
   U3509 : AOI221_X1 port map( B1 => n13045, B2 => n14454, C1 => n13042, C2 => 
                           n15857, A => n5431, ZN => n5421);
   U3510 : AOI221_X1 port map( B1 => n13072, B2 => n14655, C1 => n13069, C2 => 
                           n15785, A => n5429, ZN => n5424);
   U3511 : AOI221_X1 port map( B1 => n13060, B2 => n14488, C1 => n13057, C2 => 
                           n15833, A => n5430, ZN => n5422);
   U3512 : NAND4_X1 port map( A1 => n5372, A2 => n5373, A3 => n5374, A4 => 
                           n5375, ZN => n5362);
   U3513 : AOI221_X1 port map( B1 => n13045, B2 => n14453, C1 => n13042, C2 => 
                           n15856, A => n5379, ZN => n5372);
   U3514 : AOI221_X1 port map( B1 => n13072, B2 => n14654, C1 => n13069, C2 => 
                           n15784, A => n5377, ZN => n5374);
   U3515 : AOI221_X1 port map( B1 => n13060, B2 => n14487, C1 => n13057, C2 => 
                           n15832, A => n5378, ZN => n5373);
   U3516 : NAND4_X1 port map( A1 => n5335, A2 => n5336, A3 => n5337, A4 => 
                           n5338, ZN => n5325);
   U3517 : AOI221_X1 port map( B1 => n13045, B2 => n14452, C1 => n13042, C2 => 
                           n15855, A => n5342, ZN => n5335);
   U3518 : AOI221_X1 port map( B1 => n13072, B2 => n14653, C1 => n13069, C2 => 
                           n15783, A => n5340, ZN => n5337);
   U3519 : AOI221_X1 port map( B1 => n13060, B2 => n14486, C1 => n13057, C2 => 
                           n15831, A => n5341, ZN => n5336);
   U3520 : NAND4_X1 port map( A1 => n5298, A2 => n5299, A3 => n5300, A4 => 
                           n5301, ZN => n5288);
   U3521 : AOI221_X1 port map( B1 => n13045, B2 => n14451, C1 => n13042, C2 => 
                           n15854, A => n5305, ZN => n5298);
   U3522 : AOI221_X1 port map( B1 => n13072, B2 => n15633, C1 => n13069, C2 => 
                           n15782, A => n5303, ZN => n5300);
   U3523 : AOI221_X1 port map( B1 => n13060, B2 => n14485, C1 => n13057, C2 => 
                           n15830, A => n5304, ZN => n5299);
   U3524 : NAND4_X1 port map( A1 => n5261, A2 => n5262, A3 => n5263, A4 => 
                           n5264, ZN => n5251);
   U3525 : AOI221_X1 port map( B1 => n13045, B2 => n14450, C1 => n13042, C2 => 
                           n15853, A => n5268, ZN => n5261);
   U3526 : AOI221_X1 port map( B1 => n13072, B2 => n15813, C1 => n13069, C2 => 
                           n15781, A => n5266, ZN => n5263);
   U3527 : AOI221_X1 port map( B1 => n13060, B2 => n14484, C1 => n13057, C2 => 
                           n15829, A => n5267, ZN => n5262);
   U3528 : NAND4_X1 port map( A1 => n5224, A2 => n5225, A3 => n5226, A4 => 
                           n5227, ZN => n5214);
   U3529 : AOI221_X1 port map( B1 => n13045, B2 => n14449, C1 => n13042, C2 => 
                           n15852, A => n5231, ZN => n5224);
   U3530 : AOI221_X1 port map( B1 => n13072, B2 => n15812, C1 => n13069, C2 => 
                           n15780, A => n5229, ZN => n5226);
   U3531 : AOI221_X1 port map( B1 => n13060, B2 => n14483, C1 => n13057, C2 => 
                           n15828, A => n5230, ZN => n5225);
   U3532 : NAND4_X1 port map( A1 => n5187, A2 => n5188, A3 => n5189, A4 => 
                           n5190, ZN => n5177);
   U3533 : AOI221_X1 port map( B1 => n13045, B2 => n14448, C1 => n13042, C2 => 
                           n15851, A => n5194, ZN => n5187);
   U3534 : AOI221_X1 port map( B1 => n13072, B2 => n15811, C1 => n13069, C2 => 
                           n15779, A => n5192, ZN => n5189);
   U3535 : AOI221_X1 port map( B1 => n13060, B2 => n14482, C1 => n13057, C2 => 
                           n15827, A => n5193, ZN => n5188);
   U3536 : NAND4_X1 port map( A1 => n5150, A2 => n5151, A3 => n5152, A4 => 
                           n5153, ZN => n5140);
   U3537 : AOI221_X1 port map( B1 => n13045, B2 => n14447, C1 => n13042, C2 => 
                           n15850, A => n5157, ZN => n5150);
   U3538 : AOI221_X1 port map( B1 => n13072, B2 => n15810, C1 => n13069, C2 => 
                           n15778, A => n5155, ZN => n5152);
   U3539 : AOI221_X1 port map( B1 => n13060, B2 => n14481, C1 => n13057, C2 => 
                           n15826, A => n5156, ZN => n5151);
   U3540 : NAND4_X1 port map( A1 => n5113, A2 => n5114, A3 => n5115, A4 => 
                           n5116, ZN => n5103);
   U3541 : AOI221_X1 port map( B1 => n13046, B2 => n14446, C1 => n13043, C2 => 
                           n15849, A => n5120, ZN => n5113);
   U3542 : AOI221_X1 port map( B1 => n13073, B2 => n15809, C1 => n13070, C2 => 
                           n15777, A => n5118, ZN => n5115);
   U3543 : AOI221_X1 port map( B1 => n13061, B2 => n14480, C1 => n13058, C2 => 
                           n15825, A => n5119, ZN => n5114);
   U3544 : NAND4_X1 port map( A1 => n5076, A2 => n5077, A3 => n5078, A4 => 
                           n5079, ZN => n5066);
   U3545 : AOI221_X1 port map( B1 => n13046, B2 => n14445, C1 => n13043, C2 => 
                           n15848, A => n5083, ZN => n5076);
   U3546 : AOI221_X1 port map( B1 => n13073, B2 => n15808, C1 => n13070, C2 => 
                           n15776, A => n5081, ZN => n5078);
   U3547 : AOI221_X1 port map( B1 => n13061, B2 => n14479, C1 => n13058, C2 => 
                           n15824, A => n5082, ZN => n5077);
   U3548 : NAND4_X1 port map( A1 => n5039, A2 => n5040, A3 => n5041, A4 => 
                           n5042, ZN => n5029);
   U3549 : AOI221_X1 port map( B1 => n13046, B2 => n14444, C1 => n13043, C2 => 
                           n15847, A => n5046, ZN => n5039);
   U3550 : AOI221_X1 port map( B1 => n13073, B2 => n15807, C1 => n13070, C2 => 
                           n15775, A => n5044, ZN => n5041);
   U3551 : AOI221_X1 port map( B1 => n13061, B2 => n14478, C1 => n13058, C2 => 
                           n15823, A => n5045, ZN => n5040);
   U3552 : NAND4_X1 port map( A1 => n5002, A2 => n5003, A3 => n5004, A4 => 
                           n5005, ZN => n4992);
   U3553 : AOI221_X1 port map( B1 => n13046, B2 => n14443, C1 => n13043, C2 => 
                           n15846, A => n5009, ZN => n5002);
   U3554 : AOI221_X1 port map( B1 => n13073, B2 => n15806, C1 => n13070, C2 => 
                           n15774, A => n5007, ZN => n5004);
   U3555 : AOI221_X1 port map( B1 => n13061, B2 => n14477, C1 => n13058, C2 => 
                           n15822, A => n5008, ZN => n5003);
   U3556 : NAND4_X1 port map( A1 => n4965, A2 => n4966, A3 => n4967, A4 => 
                           n4968, ZN => n4955);
   U3557 : AOI221_X1 port map( B1 => n13046, B2 => n14442, C1 => n13043, C2 => 
                           n15845, A => n4972, ZN => n4965);
   U3558 : AOI221_X1 port map( B1 => n13073, B2 => n15805, C1 => n13070, C2 => 
                           n15773, A => n4970, ZN => n4967);
   U3559 : AOI221_X1 port map( B1 => n13061, B2 => n14476, C1 => n13058, C2 => 
                           n15821, A => n4971, ZN => n4966);
   U3560 : NAND4_X1 port map( A1 => n4928, A2 => n4929, A3 => n4930, A4 => 
                           n4931, ZN => n4918);
   U3561 : AOI221_X1 port map( B1 => n13046, B2 => n14441, C1 => n13043, C2 => 
                           n15844, A => n4935, ZN => n4928);
   U3562 : AOI221_X1 port map( B1 => n13073, B2 => n15804, C1 => n13070, C2 => 
                           n15772, A => n4933, ZN => n4930);
   U3563 : AOI221_X1 port map( B1 => n13061, B2 => n14475, C1 => n13058, C2 => 
                           n15820, A => n4934, ZN => n4929);
   U3564 : NAND4_X1 port map( A1 => n4891, A2 => n4892, A3 => n4893, A4 => 
                           n4894, ZN => n4881);
   U3565 : AOI221_X1 port map( B1 => n13046, B2 => n14440, C1 => n13043, C2 => 
                           n15843, A => n4898, ZN => n4891);
   U3566 : AOI221_X1 port map( B1 => n13073, B2 => n15803, C1 => n13070, C2 => 
                           n15771, A => n4896, ZN => n4893);
   U3567 : AOI221_X1 port map( B1 => n13061, B2 => n14474, C1 => n13058, C2 => 
                           n15819, A => n4897, ZN => n4892);
   U3568 : NAND4_X1 port map( A1 => n4854, A2 => n4855, A3 => n4856, A4 => 
                           n4857, ZN => n4844);
   U3569 : AOI221_X1 port map( B1 => n13046, B2 => n15922, C1 => n13043, C2 => 
                           n15842, A => n4861, ZN => n4854);
   U3570 : AOI221_X1 port map( B1 => n13073, B2 => n15802, C1 => n13070, C2 => 
                           n15770, A => n4859, ZN => n4856);
   U3571 : AOI221_X1 port map( B1 => n13061, B2 => n14473, C1 => n13058, C2 => 
                           n15818, A => n4860, ZN => n4855);
   U3572 : NAND4_X1 port map( A1 => n4817, A2 => n4818, A3 => n4819, A4 => 
                           n4820, ZN => n4807);
   U3573 : AOI221_X1 port map( B1 => n13046, B2 => n15873, C1 => n13043, C2 => 
                           n15841, A => n4824, ZN => n4817);
   U3574 : AOI221_X1 port map( B1 => n13073, B2 => n15801, C1 => n13070, C2 => 
                           n15769, A => n4822, ZN => n4819);
   U3575 : AOI221_X1 port map( B1 => n13061, B2 => n14472, C1 => n13058, C2 => 
                           n15817, A => n4823, ZN => n4818);
   U3576 : NAND4_X1 port map( A1 => n4780, A2 => n4781, A3 => n4782, A4 => 
                           n4783, ZN => n4770);
   U3577 : AOI221_X1 port map( B1 => n13046, B2 => n15872, C1 => n13043, C2 => 
                           n15840, A => n4787, ZN => n4780);
   U3578 : AOI221_X1 port map( B1 => n13073, B2 => n15800, C1 => n13070, C2 => 
                           n15768, A => n4785, ZN => n4782);
   U3579 : AOI221_X1 port map( B1 => n13061, B2 => n14471, C1 => n13058, C2 => 
                           n15816, A => n4786, ZN => n4781);
   U3580 : NAND4_X1 port map( A1 => n4743, A2 => n4744, A3 => n4745, A4 => 
                           n4746, ZN => n4733);
   U3581 : AOI221_X1 port map( B1 => n13046, B2 => n15871, C1 => n13043, C2 => 
                           n15839, A => n4750, ZN => n4743);
   U3582 : AOI221_X1 port map( B1 => n13073, B2 => n15799, C1 => n13070, C2 => 
                           n15767, A => n4748, ZN => n4745);
   U3583 : AOI221_X1 port map( B1 => n13061, B2 => n14470, C1 => n13058, C2 => 
                           n15815, A => n4749, ZN => n4744);
   U3584 : NAND4_X1 port map( A1 => n4706, A2 => n4707, A3 => n4708, A4 => 
                           n4709, ZN => n4696);
   U3585 : AOI221_X1 port map( B1 => n13046, B2 => n15870, C1 => n13043, C2 => 
                           n15838, A => n4713, ZN => n4706);
   U3586 : AOI221_X1 port map( B1 => n13073, B2 => n15798, C1 => n13070, C2 => 
                           n15766, A => n4711, ZN => n4708);
   U3587 : AOI221_X1 port map( B1 => n13061, B2 => n14469, C1 => n13058, C2 => 
                           n15814, A => n4712, ZN => n4707);
   U3588 : NAND4_X1 port map( A1 => n4669, A2 => n4670, A3 => n4671, A4 => 
                           n4672, ZN => n4659);
   U3589 : AOI221_X1 port map( B1 => n13047, B2 => n15869, C1 => n13044, C2 => 
                           n15632, A => n4676, ZN => n4669);
   U3590 : AOI221_X1 port map( B1 => n13074, B2 => n15797, C1 => n13071, C2 => 
                           n15581, A => n4674, ZN => n4671);
   U3591 : AOI221_X1 port map( B1 => n13062, B2 => n14468, C1 => n13059, C2 => 
                           n15589, A => n4675, ZN => n4670);
   U3592 : NAND4_X1 port map( A1 => n4284, A2 => n4285, A3 => n4286, A4 => 
                           n4287, ZN => n4263);
   U3593 : AOI221_X1 port map( B1 => n13273, B2 => n14458, C1 => n13270, C2 => 
                           n15861, A => n4293, ZN => n4284);
   U3594 : AOI221_X1 port map( B1 => n13300, B2 => n15789, C1 => n13297, C2 => 
                           n14659, A => n4291, ZN => n4286);
   U3595 : AOI221_X1 port map( B1 => n13288, B2 => n14492, C1 => n13285, C2 => 
                           n15837, A => n4292, ZN => n4285);
   U3596 : NAND4_X1 port map( A1 => n4236, A2 => n4237, A3 => n4238, A4 => 
                           n4239, ZN => n4226);
   U3597 : AOI221_X1 port map( B1 => n13273, B2 => n14457, C1 => n13270, C2 => 
                           n15860, A => n4243, ZN => n4236);
   U3598 : AOI221_X1 port map( B1 => n13300, B2 => n15788, C1 => n13297, C2 => 
                           n14658, A => n4241, ZN => n4238);
   U3599 : AOI221_X1 port map( B1 => n13288, B2 => n14491, C1 => n13285, C2 => 
                           n15836, A => n4242, ZN => n4237);
   U3600 : NAND4_X1 port map( A1 => n4199, A2 => n4200, A3 => n4201, A4 => 
                           n4202, ZN => n4189);
   U3601 : AOI221_X1 port map( B1 => n13273, B2 => n14456, C1 => n13270, C2 => 
                           n15859, A => n4206, ZN => n4199);
   U3602 : AOI221_X1 port map( B1 => n13300, B2 => n15787, C1 => n13297, C2 => 
                           n14657, A => n4204, ZN => n4201);
   U3603 : AOI221_X1 port map( B1 => n13288, B2 => n14490, C1 => n13285, C2 => 
                           n15835, A => n4205, ZN => n4200);
   U3604 : NAND4_X1 port map( A1 => n4162, A2 => n4163, A3 => n4164, A4 => 
                           n4165, ZN => n4152);
   U3605 : AOI221_X1 port map( B1 => n13273, B2 => n14455, C1 => n13270, C2 => 
                           n15858, A => n4169, ZN => n4162);
   U3606 : AOI221_X1 port map( B1 => n13300, B2 => n15786, C1 => n13297, C2 => 
                           n14656, A => n4167, ZN => n4164);
   U3607 : AOI221_X1 port map( B1 => n13288, B2 => n14489, C1 => n13285, C2 => 
                           n15834, A => n4168, ZN => n4163);
   U3608 : NAND4_X1 port map( A1 => n4125, A2 => n4126, A3 => n4127, A4 => 
                           n4128, ZN => n4115);
   U3609 : AOI221_X1 port map( B1 => n13273, B2 => n14454, C1 => n13270, C2 => 
                           n15857, A => n4132, ZN => n4125);
   U3610 : AOI221_X1 port map( B1 => n13300, B2 => n15785, C1 => n13297, C2 => 
                           n14655, A => n4130, ZN => n4127);
   U3611 : AOI221_X1 port map( B1 => n13288, B2 => n14488, C1 => n13285, C2 => 
                           n15833, A => n4131, ZN => n4126);
   U3612 : NAND4_X1 port map( A1 => n4088, A2 => n4089, A3 => n4090, A4 => 
                           n4091, ZN => n4078);
   U3613 : AOI221_X1 port map( B1 => n13273, B2 => n14453, C1 => n13270, C2 => 
                           n15856, A => n4095, ZN => n4088);
   U3614 : AOI221_X1 port map( B1 => n13300, B2 => n15784, C1 => n13297, C2 => 
                           n14654, A => n4093, ZN => n4090);
   U3615 : AOI221_X1 port map( B1 => n13288, B2 => n14487, C1 => n13285, C2 => 
                           n15832, A => n4094, ZN => n4089);
   U3616 : NAND4_X1 port map( A1 => n4051, A2 => n4052, A3 => n4053, A4 => 
                           n4054, ZN => n4041);
   U3617 : AOI221_X1 port map( B1 => n13273, B2 => n14452, C1 => n13270, C2 => 
                           n15855, A => n4058, ZN => n4051);
   U3618 : AOI221_X1 port map( B1 => n13300, B2 => n15783, C1 => n13297, C2 => 
                           n14653, A => n4056, ZN => n4053);
   U3619 : AOI221_X1 port map( B1 => n13288, B2 => n14486, C1 => n13285, C2 => 
                           n15831, A => n4057, ZN => n4052);
   U3620 : NAND4_X1 port map( A1 => n4014, A2 => n4015, A3 => n4016, A4 => 
                           n4017, ZN => n4004);
   U3621 : AOI221_X1 port map( B1 => n13273, B2 => n14451, C1 => n13270, C2 => 
                           n15854, A => n4021, ZN => n4014);
   U3622 : AOI221_X1 port map( B1 => n13300, B2 => n15782, C1 => n13297, C2 => 
                           n15633, A => n4019, ZN => n4016);
   U3623 : AOI221_X1 port map( B1 => n13288, B2 => n14485, C1 => n13285, C2 => 
                           n15830, A => n4020, ZN => n4015);
   U3624 : NAND4_X1 port map( A1 => n3977, A2 => n3978, A3 => n3979, A4 => 
                           n3980, ZN => n3967);
   U3625 : AOI221_X1 port map( B1 => n13273, B2 => n14450, C1 => n13270, C2 => 
                           n15853, A => n3984, ZN => n3977);
   U3626 : AOI221_X1 port map( B1 => n13300, B2 => n15781, C1 => n13297, C2 => 
                           n15813, A => n3982, ZN => n3979);
   U3627 : AOI221_X1 port map( B1 => n13288, B2 => n14484, C1 => n13285, C2 => 
                           n15829, A => n3983, ZN => n3978);
   U3628 : NAND4_X1 port map( A1 => n3940, A2 => n3941, A3 => n3942, A4 => 
                           n3943, ZN => n3930);
   U3629 : AOI221_X1 port map( B1 => n13273, B2 => n14449, C1 => n13270, C2 => 
                           n15852, A => n3947, ZN => n3940);
   U3630 : AOI221_X1 port map( B1 => n13300, B2 => n15780, C1 => n13297, C2 => 
                           n15812, A => n3945, ZN => n3942);
   U3631 : AOI221_X1 port map( B1 => n13288, B2 => n14483, C1 => n13285, C2 => 
                           n15828, A => n3946, ZN => n3941);
   U3632 : NAND4_X1 port map( A1 => n3903, A2 => n3904, A3 => n3905, A4 => 
                           n3906, ZN => n3893);
   U3633 : AOI221_X1 port map( B1 => n13273, B2 => n14448, C1 => n13270, C2 => 
                           n15851, A => n3910, ZN => n3903);
   U3634 : AOI221_X1 port map( B1 => n13300, B2 => n15779, C1 => n13297, C2 => 
                           n15811, A => n3908, ZN => n3905);
   U3635 : AOI221_X1 port map( B1 => n13288, B2 => n14482, C1 => n13285, C2 => 
                           n15827, A => n3909, ZN => n3904);
   U3636 : NAND4_X1 port map( A1 => n3866, A2 => n3867, A3 => n3868, A4 => 
                           n3869, ZN => n3856);
   U3637 : AOI221_X1 port map( B1 => n13273, B2 => n14447, C1 => n13270, C2 => 
                           n15850, A => n3873, ZN => n3866);
   U3638 : AOI221_X1 port map( B1 => n13300, B2 => n15778, C1 => n13297, C2 => 
                           n15810, A => n3871, ZN => n3868);
   U3639 : AOI221_X1 port map( B1 => n13288, B2 => n14481, C1 => n13285, C2 => 
                           n15826, A => n3872, ZN => n3867);
   U3640 : NAND4_X1 port map( A1 => n3829, A2 => n3830, A3 => n3831, A4 => 
                           n3832, ZN => n3819);
   U3641 : AOI221_X1 port map( B1 => n13274, B2 => n14446, C1 => n13271, C2 => 
                           n15849, A => n3836, ZN => n3829);
   U3642 : AOI221_X1 port map( B1 => n13301, B2 => n15777, C1 => n13298, C2 => 
                           n15809, A => n3834, ZN => n3831);
   U3643 : AOI221_X1 port map( B1 => n13289, B2 => n14480, C1 => n13286, C2 => 
                           n15825, A => n3835, ZN => n3830);
   U3644 : NAND4_X1 port map( A1 => n3792, A2 => n3793, A3 => n3794, A4 => 
                           n3795, ZN => n3782);
   U3645 : AOI221_X1 port map( B1 => n13274, B2 => n14445, C1 => n13271, C2 => 
                           n15848, A => n3799, ZN => n3792);
   U3646 : AOI221_X1 port map( B1 => n13301, B2 => n15776, C1 => n13298, C2 => 
                           n15808, A => n3797, ZN => n3794);
   U3647 : AOI221_X1 port map( B1 => n13289, B2 => n14479, C1 => n13286, C2 => 
                           n15824, A => n3798, ZN => n3793);
   U3648 : NAND4_X1 port map( A1 => n3755, A2 => n3756, A3 => n3757, A4 => 
                           n3758, ZN => n3745);
   U3649 : AOI221_X1 port map( B1 => n13274, B2 => n14444, C1 => n13271, C2 => 
                           n15847, A => n3762, ZN => n3755);
   U3650 : AOI221_X1 port map( B1 => n13301, B2 => n15775, C1 => n13298, C2 => 
                           n15807, A => n3760, ZN => n3757);
   U3651 : AOI221_X1 port map( B1 => n13289, B2 => n14478, C1 => n13286, C2 => 
                           n15823, A => n3761, ZN => n3756);
   U3652 : NAND4_X1 port map( A1 => n3718, A2 => n3719, A3 => n3720, A4 => 
                           n3721, ZN => n3708);
   U3653 : AOI221_X1 port map( B1 => n13274, B2 => n14443, C1 => n13271, C2 => 
                           n15846, A => n3725, ZN => n3718);
   U3654 : AOI221_X1 port map( B1 => n13301, B2 => n15774, C1 => n13298, C2 => 
                           n15806, A => n3723, ZN => n3720);
   U3655 : AOI221_X1 port map( B1 => n13289, B2 => n14477, C1 => n13286, C2 => 
                           n15822, A => n3724, ZN => n3719);
   U3656 : NAND4_X1 port map( A1 => n3681, A2 => n3682, A3 => n3683, A4 => 
                           n3684, ZN => n3671);
   U3657 : AOI221_X1 port map( B1 => n13274, B2 => n14442, C1 => n13271, C2 => 
                           n15845, A => n3688, ZN => n3681);
   U3658 : AOI221_X1 port map( B1 => n13301, B2 => n15773, C1 => n13298, C2 => 
                           n15805, A => n3686, ZN => n3683);
   U3659 : AOI221_X1 port map( B1 => n13289, B2 => n14476, C1 => n13286, C2 => 
                           n15821, A => n3687, ZN => n3682);
   U3660 : NAND4_X1 port map( A1 => n3644, A2 => n3645, A3 => n3646, A4 => 
                           n3647, ZN => n3634);
   U3661 : AOI221_X1 port map( B1 => n13274, B2 => n14441, C1 => n13271, C2 => 
                           n15844, A => n3651, ZN => n3644);
   U3662 : AOI221_X1 port map( B1 => n13301, B2 => n15772, C1 => n13298, C2 => 
                           n15804, A => n3649, ZN => n3646);
   U3663 : AOI221_X1 port map( B1 => n13289, B2 => n14475, C1 => n13286, C2 => 
                           n15820, A => n3650, ZN => n3645);
   U3664 : NAND4_X1 port map( A1 => n3607, A2 => n3608, A3 => n3609, A4 => 
                           n3610, ZN => n3597);
   U3665 : AOI221_X1 port map( B1 => n13274, B2 => n14440, C1 => n13271, C2 => 
                           n15843, A => n3614, ZN => n3607);
   U3666 : AOI221_X1 port map( B1 => n13301, B2 => n15771, C1 => n13298, C2 => 
                           n15803, A => n3612, ZN => n3609);
   U3667 : AOI221_X1 port map( B1 => n13289, B2 => n14474, C1 => n13286, C2 => 
                           n15819, A => n3613, ZN => n3608);
   U3668 : NAND4_X1 port map( A1 => n3570, A2 => n3571, A3 => n3572, A4 => 
                           n3573, ZN => n3560);
   U3669 : AOI221_X1 port map( B1 => n13274, B2 => n15922, C1 => n13271, C2 => 
                           n15842, A => n3577, ZN => n3570);
   U3670 : AOI221_X1 port map( B1 => n13301, B2 => n15770, C1 => n13298, C2 => 
                           n15802, A => n3575, ZN => n3572);
   U3671 : AOI221_X1 port map( B1 => n13289, B2 => n14473, C1 => n13286, C2 => 
                           n15818, A => n3576, ZN => n3571);
   U3672 : NAND4_X1 port map( A1 => n3533, A2 => n3534, A3 => n3535, A4 => 
                           n3536, ZN => n3523);
   U3673 : AOI221_X1 port map( B1 => n13274, B2 => n15873, C1 => n13271, C2 => 
                           n15841, A => n3540, ZN => n3533);
   U3674 : AOI221_X1 port map( B1 => n13301, B2 => n15769, C1 => n13298, C2 => 
                           n15801, A => n3538, ZN => n3535);
   U3675 : AOI221_X1 port map( B1 => n13289, B2 => n14472, C1 => n13286, C2 => 
                           n15817, A => n3539, ZN => n3534);
   U3676 : NAND4_X1 port map( A1 => n3496, A2 => n3497, A3 => n3498, A4 => 
                           n3499, ZN => n3486);
   U3677 : AOI221_X1 port map( B1 => n13274, B2 => n15872, C1 => n13271, C2 => 
                           n15840, A => n3503, ZN => n3496);
   U3678 : AOI221_X1 port map( B1 => n13301, B2 => n15768, C1 => n13298, C2 => 
                           n15800, A => n3501, ZN => n3498);
   U3679 : AOI221_X1 port map( B1 => n13289, B2 => n14471, C1 => n13286, C2 => 
                           n15816, A => n3502, ZN => n3497);
   U3680 : NAND4_X1 port map( A1 => n3459, A2 => n3460, A3 => n3461, A4 => 
                           n3462, ZN => n3449);
   U3681 : AOI221_X1 port map( B1 => n13274, B2 => n15871, C1 => n13271, C2 => 
                           n15839, A => n3466, ZN => n3459);
   U3682 : AOI221_X1 port map( B1 => n13301, B2 => n15767, C1 => n13298, C2 => 
                           n15799, A => n3464, ZN => n3461);
   U3683 : AOI221_X1 port map( B1 => n13289, B2 => n14470, C1 => n13286, C2 => 
                           n15815, A => n3465, ZN => n3460);
   U3684 : NAND4_X1 port map( A1 => n3422, A2 => n3423, A3 => n3424, A4 => 
                           n3425, ZN => n3412);
   U3685 : AOI221_X1 port map( B1 => n13274, B2 => n15870, C1 => n13271, C2 => 
                           n15838, A => n3429, ZN => n3422);
   U3686 : AOI221_X1 port map( B1 => n13301, B2 => n15766, C1 => n13298, C2 => 
                           n15798, A => n3427, ZN => n3424);
   U3687 : AOI221_X1 port map( B1 => n13289, B2 => n14469, C1 => n13286, C2 => 
                           n15814, A => n3428, ZN => n3423);
   U3688 : NAND4_X1 port map( A1 => n3385, A2 => n3386, A3 => n3387, A4 => 
                           n3388, ZN => n3375);
   U3689 : AOI221_X1 port map( B1 => n13275, B2 => n15869, C1 => n13272, C2 => 
                           n15632, A => n3392, ZN => n3385);
   U3690 : AOI221_X1 port map( B1 => n13302, B2 => n15581, C1 => n13299, C2 => 
                           n15797, A => n3390, ZN => n3387);
   U3691 : AOI221_X1 port map( B1 => n13290, B2 => n14468, C1 => n13287, C2 => 
                           n15589, A => n3391, ZN => n3386);
   U3692 : NAND4_X1 port map( A1 => n3348, A2 => n3349, A3 => n3350, A4 => 
                           n3351, ZN => n3338);
   U3693 : AOI221_X1 port map( B1 => n13275, B2 => n15868, C1 => n13272, C2 => 
                           n15631, A => n3355, ZN => n3348);
   U3694 : AOI221_X1 port map( B1 => n13302, B2 => n15580, C1 => n13299, C2 => 
                           n15796, A => n3353, ZN => n3350);
   U3695 : AOI221_X1 port map( B1 => n13290, B2 => n14467, C1 => n13287, C2 => 
                           n15588, A => n3354, ZN => n3349);
   U3696 : NAND4_X1 port map( A1 => n3311, A2 => n3312, A3 => n3313, A4 => 
                           n3314, ZN => n3301);
   U3697 : AOI221_X1 port map( B1 => n13275, B2 => n15867, C1 => n13272, C2 => 
                           n15630, A => n3318, ZN => n3311);
   U3698 : AOI221_X1 port map( B1 => n13302, B2 => n15579, C1 => n13299, C2 => 
                           n15795, A => n3316, ZN => n3313);
   U3699 : AOI221_X1 port map( B1 => n13290, B2 => n14466, C1 => n13287, C2 => 
                           n15587, A => n3317, ZN => n3312);
   U3700 : NAND4_X1 port map( A1 => n3274, A2 => n3275, A3 => n3276, A4 => 
                           n3277, ZN => n3264);
   U3701 : AOI221_X1 port map( B1 => n13275, B2 => n15866, C1 => n13272, C2 => 
                           n15629, A => n3281, ZN => n3274);
   U3702 : AOI221_X1 port map( B1 => n13302, B2 => n15578, C1 => n13299, C2 => 
                           n15794, A => n3279, ZN => n3276);
   U3703 : AOI221_X1 port map( B1 => n13290, B2 => n14465, C1 => n13287, C2 => 
                           n15586, A => n3280, ZN => n3275);
   U3704 : NOR3_X2 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(1), A3 => n16066, 
                           ZN => n4278);
   U3705 : NOR3_X2 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(2), A3 => n16068, 
                           ZN => n5671);
   U3706 : NOR3_X2 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), A3 => n16067, 
                           ZN => n5666);
   U3707 : NOR3_X2 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(2), A3 => n16065, 
                           ZN => n4280);
   U3708 : NOR3_X2 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(1), A3 => n16069, 
                           ZN => n5674);
   U3709 : NOR3_X2 port map( A1 => n16067, A2 => ADD_RD2(2), A3 => n16068, ZN 
                           => n5676);
   U3710 : BUF_X1 port map( A => n16063, Z => n12922);
   U3711 : BUF_X1 port map( A => n16063, Z => n12923);
   U3712 : BUF_X1 port map( A => n16063, Z => n12924);
   U3713 : BUF_X1 port map( A => n16063, Z => n12925);
   U3714 : BUF_X1 port map( A => n16063, Z => n12926);
   U3715 : BUF_X1 port map( A => n16063, Z => n12927);
   U3716 : INV_X1 port map( A => ADD_RD2(0), ZN => n16067);
   U3717 : INV_X1 port map( A => ADD_RD1(0), ZN => n16064);
   U3718 : BUF_X1 port map( A => n2864, Z => n13830);
   U3719 : BUF_X1 port map( A => n2863, Z => n13836);
   U3720 : BUF_X1 port map( A => n2862, Z => n13842);
   U3721 : BUF_X1 port map( A => n2861, Z => n13848);
   U3722 : BUF_X1 port map( A => n2860, Z => n13854);
   U3723 : BUF_X1 port map( A => n2859, Z => n13860);
   U3724 : BUF_X1 port map( A => n2858, Z => n13866);
   U3725 : BUF_X1 port map( A => n2857, Z => n13872);
   U3726 : BUF_X1 port map( A => n2856, Z => n13878);
   U3727 : BUF_X1 port map( A => n2855, Z => n13884);
   U3728 : BUF_X1 port map( A => n2854, Z => n13890);
   U3729 : BUF_X1 port map( A => n2853, Z => n13896);
   U3730 : BUF_X1 port map( A => n2852, Z => n13902);
   U3731 : BUF_X1 port map( A => n2851, Z => n13908);
   U3732 : BUF_X1 port map( A => n2850, Z => n13914);
   U3733 : BUF_X1 port map( A => n2849, Z => n13920);
   U3734 : BUF_X1 port map( A => n2848, Z => n13926);
   U3735 : BUF_X1 port map( A => n2847, Z => n13932);
   U3736 : BUF_X1 port map( A => n2846, Z => n13938);
   U3737 : BUF_X1 port map( A => n2845, Z => n13944);
   U3738 : BUF_X1 port map( A => n2844, Z => n13950);
   U3739 : BUF_X1 port map( A => n2843, Z => n13956);
   U3740 : BUF_X1 port map( A => n2842, Z => n13962);
   U3741 : BUF_X1 port map( A => n2841, Z => n13968);
   U3742 : BUF_X1 port map( A => n2840, Z => n13974);
   U3743 : BUF_X1 port map( A => n2839, Z => n13980);
   U3744 : BUF_X1 port map( A => n2838, Z => n13986);
   U3745 : BUF_X1 port map( A => n2837, Z => n13992);
   U3746 : BUF_X1 port map( A => n2836, Z => n13998);
   U3747 : BUF_X1 port map( A => n2835, Z => n14004);
   U3748 : BUF_X1 port map( A => n2833, Z => n14013);
   U3749 : BUF_X1 port map( A => n2865, Z => n13824);
   U3750 : BUF_X1 port map( A => n2865, Z => n13828);
   U3751 : BUF_X1 port map( A => n2864, Z => n13834);
   U3752 : BUF_X1 port map( A => n2863, Z => n13840);
   U3753 : BUF_X1 port map( A => n2862, Z => n13846);
   U3754 : BUF_X1 port map( A => n2861, Z => n13852);
   U3755 : BUF_X1 port map( A => n2860, Z => n13858);
   U3756 : BUF_X1 port map( A => n2859, Z => n13864);
   U3757 : BUF_X1 port map( A => n2858, Z => n13870);
   U3758 : BUF_X1 port map( A => n2857, Z => n13876);
   U3759 : BUF_X1 port map( A => n2856, Z => n13882);
   U3760 : BUF_X1 port map( A => n2855, Z => n13888);
   U3761 : BUF_X1 port map( A => n2854, Z => n13894);
   U3762 : BUF_X1 port map( A => n2853, Z => n13900);
   U3763 : BUF_X1 port map( A => n2852, Z => n13906);
   U3764 : BUF_X1 port map( A => n2851, Z => n13912);
   U3765 : BUF_X1 port map( A => n2850, Z => n13918);
   U3766 : BUF_X1 port map( A => n2849, Z => n13924);
   U3767 : BUF_X1 port map( A => n2848, Z => n13930);
   U3768 : BUF_X1 port map( A => n2847, Z => n13936);
   U3769 : BUF_X1 port map( A => n2846, Z => n13942);
   U3770 : BUF_X1 port map( A => n2845, Z => n13948);
   U3771 : BUF_X1 port map( A => n2844, Z => n13954);
   U3772 : BUF_X1 port map( A => n2843, Z => n13960);
   U3773 : BUF_X1 port map( A => n2842, Z => n13966);
   U3774 : BUF_X1 port map( A => n2841, Z => n13972);
   U3775 : BUF_X1 port map( A => n2840, Z => n13978);
   U3776 : BUF_X1 port map( A => n2839, Z => n13984);
   U3777 : BUF_X1 port map( A => n2838, Z => n13990);
   U3778 : BUF_X1 port map( A => n2837, Z => n13996);
   U3779 : BUF_X1 port map( A => n2836, Z => n14002);
   U3780 : BUF_X1 port map( A => n2835, Z => n14008);
   U3781 : BUF_X1 port map( A => n2833, Z => n14017);
   U3782 : BUF_X1 port map( A => n2865, Z => n13827);
   U3783 : BUF_X1 port map( A => n2864, Z => n13833);
   U3784 : BUF_X1 port map( A => n2863, Z => n13839);
   U3785 : BUF_X1 port map( A => n2862, Z => n13845);
   U3786 : BUF_X1 port map( A => n2861, Z => n13851);
   U3787 : BUF_X1 port map( A => n2860, Z => n13857);
   U3788 : BUF_X1 port map( A => n2859, Z => n13863);
   U3789 : BUF_X1 port map( A => n2858, Z => n13869);
   U3790 : BUF_X1 port map( A => n2857, Z => n13875);
   U3791 : BUF_X1 port map( A => n2856, Z => n13881);
   U3792 : BUF_X1 port map( A => n2855, Z => n13887);
   U3793 : BUF_X1 port map( A => n2854, Z => n13893);
   U3794 : BUF_X1 port map( A => n2853, Z => n13899);
   U3795 : BUF_X1 port map( A => n2852, Z => n13905);
   U3796 : BUF_X1 port map( A => n2851, Z => n13911);
   U3797 : BUF_X1 port map( A => n2850, Z => n13917);
   U3798 : BUF_X1 port map( A => n2849, Z => n13923);
   U3799 : BUF_X1 port map( A => n2848, Z => n13929);
   U3800 : BUF_X1 port map( A => n2847, Z => n13935);
   U3801 : BUF_X1 port map( A => n2846, Z => n13941);
   U3802 : BUF_X1 port map( A => n2845, Z => n13947);
   U3803 : BUF_X1 port map( A => n2844, Z => n13953);
   U3804 : BUF_X1 port map( A => n2843, Z => n13959);
   U3805 : BUF_X1 port map( A => n2842, Z => n13965);
   U3806 : BUF_X1 port map( A => n2841, Z => n13971);
   U3807 : BUF_X1 port map( A => n2840, Z => n13977);
   U3808 : BUF_X1 port map( A => n2839, Z => n13983);
   U3809 : BUF_X1 port map( A => n2838, Z => n13989);
   U3810 : BUF_X1 port map( A => n2837, Z => n13995);
   U3811 : BUF_X1 port map( A => n2836, Z => n14001);
   U3812 : BUF_X1 port map( A => n2835, Z => n14007);
   U3813 : BUF_X1 port map( A => n2833, Z => n14016);
   U3814 : BUF_X1 port map( A => n2865, Z => n13826);
   U3815 : BUF_X1 port map( A => n2864, Z => n13832);
   U3816 : BUF_X1 port map( A => n2863, Z => n13838);
   U3818 : BUF_X1 port map( A => n2862, Z => n13844);
   U3819 : BUF_X1 port map( A => n2861, Z => n13850);
   U3820 : BUF_X1 port map( A => n2860, Z => n13856);
   U3821 : BUF_X1 port map( A => n2859, Z => n13862);
   U3822 : BUF_X1 port map( A => n2858, Z => n13868);
   U3823 : BUF_X1 port map( A => n2857, Z => n13874);
   U3824 : BUF_X1 port map( A => n2856, Z => n13880);
   U3825 : BUF_X1 port map( A => n2855, Z => n13886);
   U3826 : BUF_X1 port map( A => n2854, Z => n13892);
   U3827 : BUF_X1 port map( A => n2853, Z => n13898);
   U3828 : BUF_X1 port map( A => n2852, Z => n13904);
   U3829 : BUF_X1 port map( A => n2851, Z => n13910);
   U3830 : BUF_X1 port map( A => n2850, Z => n13916);
   U3831 : BUF_X1 port map( A => n2849, Z => n13922);
   U3832 : BUF_X1 port map( A => n2848, Z => n13928);
   U3833 : BUF_X1 port map( A => n2847, Z => n13934);
   U3834 : BUF_X1 port map( A => n2846, Z => n13940);
   U3835 : BUF_X1 port map( A => n2845, Z => n13946);
   U3836 : BUF_X1 port map( A => n2844, Z => n13952);
   U3837 : BUF_X1 port map( A => n2843, Z => n13958);
   U3838 : BUF_X1 port map( A => n2842, Z => n13964);
   U3839 : BUF_X1 port map( A => n2841, Z => n13970);
   U3840 : BUF_X1 port map( A => n2840, Z => n13976);
   U3841 : BUF_X1 port map( A => n2839, Z => n13982);
   U3842 : BUF_X1 port map( A => n2838, Z => n13988);
   U3843 : BUF_X1 port map( A => n2837, Z => n13994);
   U3844 : BUF_X1 port map( A => n2836, Z => n14000);
   U3845 : BUF_X1 port map( A => n2835, Z => n14006);
   U3846 : BUF_X1 port map( A => n2833, Z => n14015);
   U3847 : BUF_X1 port map( A => n2865, Z => n13825);
   U3848 : BUF_X1 port map( A => n2864, Z => n13831);
   U3849 : BUF_X1 port map( A => n2863, Z => n13837);
   U3850 : BUF_X1 port map( A => n2862, Z => n13843);
   U3851 : BUF_X1 port map( A => n2861, Z => n13849);
   U3852 : BUF_X1 port map( A => n2860, Z => n13855);
   U3853 : BUF_X1 port map( A => n2859, Z => n13861);
   U3854 : BUF_X1 port map( A => n2858, Z => n13867);
   U3855 : BUF_X1 port map( A => n2857, Z => n13873);
   U3856 : BUF_X1 port map( A => n2856, Z => n13879);
   U3857 : BUF_X1 port map( A => n2855, Z => n13885);
   U3858 : BUF_X1 port map( A => n2854, Z => n13891);
   U3859 : BUF_X1 port map( A => n2853, Z => n13897);
   U3860 : BUF_X1 port map( A => n2852, Z => n13903);
   U3861 : BUF_X1 port map( A => n2851, Z => n13909);
   U3862 : BUF_X1 port map( A => n2850, Z => n13915);
   U3863 : BUF_X1 port map( A => n2849, Z => n13921);
   U3864 : BUF_X1 port map( A => n2848, Z => n13927);
   U3865 : BUF_X1 port map( A => n2847, Z => n13933);
   U3866 : BUF_X1 port map( A => n2846, Z => n13939);
   U3867 : BUF_X1 port map( A => n2845, Z => n13945);
   U3868 : BUF_X1 port map( A => n2844, Z => n13951);
   U3869 : BUF_X1 port map( A => n2843, Z => n13957);
   U3870 : BUF_X1 port map( A => n2842, Z => n13963);
   U3871 : BUF_X1 port map( A => n2841, Z => n13969);
   U3872 : BUF_X1 port map( A => n2840, Z => n13975);
   U3873 : BUF_X1 port map( A => n2839, Z => n13981);
   U3874 : BUF_X1 port map( A => n2838, Z => n13987);
   U3875 : BUF_X1 port map( A => n2837, Z => n13993);
   U3876 : BUF_X1 port map( A => n2836, Z => n13999);
   U3877 : BUF_X1 port map( A => n2835, Z => n14005);
   U3878 : BUF_X1 port map( A => n2833, Z => n14014);
   U3879 : INV_X1 port map( A => ADD_RD2(1), ZN => n16068);
   U3880 : INV_X1 port map( A => ADD_RD1(1), ZN => n16065);
   U3881 : INV_X1 port map( A => ADD_RD2(2), ZN => n16069);
   U3882 : INV_X1 port map( A => ADD_RD1(2), ZN => n16066);
   U3883 : NAND2_X1 port map( A1 => n14027, A2 => n16074, ZN => n4325);
   U3884 : NAND2_X1 port map( A1 => n14027, A2 => n16073, ZN => n3041);
   U3885 : NAND4_X1 port map( A1 => n5738, A2 => n5740, A3 => n5742, A4 => 
                           n5744, ZN => n4322);
   U3886 : NOR3_X1 port map( A1 => n5754, A2 => n16075, A3 => n16074, ZN => 
                           n5742);
   U3887 : NAND4_X1 port map( A1 => n4313, A2 => n4314, A3 => n4315, A4 => 
                           n4316, ZN => n3038);
   U3888 : NOR3_X1 port map( A1 => n4321, A2 => n16075, A3 => n16073, ZN => 
                           n4315);
   U3889 : NOR2_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(1), ZN => n3000);
   U3890 : NOR2_X1 port map( A1 => n16070, A2 => ADD_WR(1), ZN => n3003);
   U3891 : NOR2_X1 port map( A1 => n16071, A2 => ADD_WR(0), ZN => n3006);
   U3892 : NOR2_X1 port map( A1 => ADD_WR(2), A2 => ADD_WR(3), ZN => n3022);
   U3893 : INV_X1 port map( A => ADD_WR(1), ZN => n16071);
   U3894 : INV_X1 port map( A => ADD_WR(2), ZN => n16072);
   U3895 : AND2_X1 port map( A1 => ADD_WR(3), A2 => ADD_WR(2), ZN => n3012);
   U3896 : INV_X1 port map( A => ADD_WR(0), ZN => n16070);
   U3897 : INV_X1 port map( A => n13810, ZN => n13823);
   U3898 : AOI221_X1 port map( B1 => n13182, B2 => n5982, C1 => n13179, C2 => 
                           n15177, A => n3259, ZN => n3254);
   U3899 : OAI222_X1 port map( A1 => n15273, A2 => n13176, B1 => n15209, B2 => 
                           n13173, C1 => n15241, C2 => n13170, ZN => n3259);
   U3900 : AOI221_X1 port map( B1 => n13182, B2 => n5983, C1 => n13179, C2 => 
                           n15176, A => n3222, ZN => n3217);
   U3901 : OAI222_X1 port map( A1 => n15272, A2 => n13176, B1 => n15208, B2 => 
                           n13173, C1 => n15240, C2 => n13170, ZN => n3222);
   U3902 : AOI221_X1 port map( B1 => n13182, B2 => n5984, C1 => n13179, C2 => 
                           n15175, A => n3185, ZN => n3180);
   U3903 : OAI222_X1 port map( A1 => n15271, A2 => n13176, B1 => n15207, B2 => 
                           n13173, C1 => n15239, C2 => n13170, ZN => n3185);
   U3904 : AOI221_X1 port map( B1 => n13182, B2 => n5985, C1 => n13179, C2 => 
                           n15174, A => n3141, ZN => n3125);
   U3905 : OAI222_X1 port map( A1 => n15270, A2 => n13176, B1 => n15206, B2 => 
                           n13173, C1 => n15238, C2 => n13170, ZN => n3141);
   U3906 : AOI221_X1 port map( B1 => n12954, B2 => n5979, C1 => n12951, C2 => 
                           n15180, A => n4654, ZN => n4649);
   U3907 : OAI222_X1 port map( A1 => n15276, A2 => n12948, B1 => n15212, B2 => 
                           n12945, C1 => n15244, C2 => n12942, ZN => n4654);
   U3908 : AOI221_X1 port map( B1 => n12954, B2 => n5980, C1 => n12951, C2 => 
                           n15179, A => n4617, ZN => n4612);
   U3909 : OAI222_X1 port map( A1 => n15275, A2 => n12948, B1 => n15211, B2 => 
                           n12945, C1 => n15243, C2 => n12942, ZN => n4617);
   U3910 : AOI221_X1 port map( B1 => n12954, B2 => n5981, C1 => n12951, C2 => 
                           n15178, A => n4580, ZN => n4575);
   U3911 : OAI222_X1 port map( A1 => n15274, A2 => n12948, B1 => n15210, B2 => 
                           n12945, C1 => n15242, C2 => n12942, ZN => n4580);
   U3912 : AOI221_X1 port map( B1 => n12954, B2 => n5982, C1 => n12951, C2 => 
                           n15177, A => n4543, ZN => n4538);
   U3913 : OAI222_X1 port map( A1 => n15273, A2 => n12948, B1 => n15209, B2 => 
                           n12945, C1 => n15241, C2 => n12942, ZN => n4543);
   U3914 : AOI221_X1 port map( B1 => n12954, B2 => n5983, C1 => n12951, C2 => 
                           n15176, A => n4506, ZN => n4501);
   U3915 : OAI222_X1 port map( A1 => n15272, A2 => n12948, B1 => n15208, B2 => 
                           n12945, C1 => n15240, C2 => n12942, ZN => n4506);
   U3916 : AOI221_X1 port map( B1 => n12954, B2 => n5984, C1 => n12951, C2 => 
                           n15175, A => n4469, ZN => n4464);
   U3917 : OAI222_X1 port map( A1 => n15271, A2 => n12948, B1 => n15207, B2 => 
                           n12945, C1 => n15239, C2 => n12942, ZN => n4469);
   U3918 : AOI221_X1 port map( B1 => n12954, B2 => n5985, C1 => n12951, C2 => 
                           n15174, A => n4425, ZN => n4409);
   U3919 : OAI222_X1 port map( A1 => n15270, A2 => n12948, B1 => n15206, B2 => 
                           n12945, C1 => n15238, C2 => n12942, ZN => n4425);
   U3920 : AOI221_X1 port map( B1 => n13008, B2 => n6234, C1 => n13005, C2 => 
                           n15565, A => n4683, ZN => n4678);
   U3921 : OAI222_X1 port map( A1 => n14923, A2 => n13002, B1 => n14859, B2 => 
                           n12999, C1 => n14891, C2 => n12996, ZN => n4683);
   U3922 : AOI221_X1 port map( B1 => n13236, B2 => n6234, C1 => n13233, C2 => 
                           n15565, A => n3399, ZN => n3394);
   U3923 : OAI222_X1 port map( A1 => n14923, A2 => n13230, B1 => n14859, B2 => 
                           n13227, C1 => n14891, C2 => n13224, ZN => n3399);
   U3924 : AOI221_X1 port map( B1 => n13182, B2 => n5979, C1 => n13179, C2 => 
                           n15180, A => n3370, ZN => n3365);
   U3925 : OAI222_X1 port map( A1 => n15276, A2 => n13176, B1 => n15212, B2 => 
                           n13173, C1 => n15244, C2 => n13170, ZN => n3370);
   U3926 : AOI221_X1 port map( B1 => n13182, B2 => n5980, C1 => n13179, C2 => 
                           n15179, A => n3333, ZN => n3328);
   U3927 : OAI222_X1 port map( A1 => n15275, A2 => n13176, B1 => n15211, B2 => 
                           n13173, C1 => n15243, C2 => n13170, ZN => n3333);
   U3928 : AOI221_X1 port map( B1 => n13182, B2 => n5981, C1 => n13179, C2 => 
                           n15178, A => n3296, ZN => n3291);
   U3929 : OAI222_X1 port map( A1 => n15274, A2 => n13176, B1 => n15210, B2 => 
                           n13173, C1 => n15242, C2 => n13170, ZN => n3296);
   U3930 : OAI222_X1 port map( A1 => n16082, A2 => n13155, B1 => n4619, B2 => 
                           n13152, C1 => n13144, C2 => n1487, ZN => n7597);
   U3931 : NOR4_X1 port map( A1 => n4620, A2 => n4621, A3 => n4622, A4 => n4623
                           , ZN => n4619);
   U3932 : NAND4_X1 port map( A1 => n4648, A2 => n4649, A3 => n4650, A4 => 
                           n4651, ZN => n4620);
   U3933 : NAND4_X1 port map( A1 => n4640, A2 => n4641, A3 => n4642, A4 => 
                           n4643, ZN => n4621);
   U3934 : OAI222_X1 port map( A1 => n16081, A2 => n13155, B1 => n4582, B2 => 
                           n13152, C1 => n13144, C2 => n1486, ZN => n7599);
   U3935 : NOR4_X1 port map( A1 => n4583, A2 => n4584, A3 => n4585, A4 => n4586
                           , ZN => n4582);
   U3936 : NAND4_X1 port map( A1 => n4611, A2 => n4612, A3 => n4613, A4 => 
                           n4614, ZN => n4583);
   U3937 : NAND4_X1 port map( A1 => n4603, A2 => n4604, A3 => n4605, A4 => 
                           n4606, ZN => n4584);
   U3938 : OAI222_X1 port map( A1 => n16080, A2 => n13155, B1 => n4545, B2 => 
                           n13152, C1 => n13144, C2 => n1485, ZN => n7601);
   U3939 : NOR4_X1 port map( A1 => n4546, A2 => n4547, A3 => n4548, A4 => n4549
                           , ZN => n4545);
   U3940 : NAND4_X1 port map( A1 => n4574, A2 => n4575, A3 => n4576, A4 => 
                           n4577, ZN => n4546);
   U3941 : NAND4_X1 port map( A1 => n4566, A2 => n4567, A3 => n4568, A4 => 
                           n4569, ZN => n4547);
   U3942 : OAI222_X1 port map( A1 => n16079, A2 => n13155, B1 => n4508, B2 => 
                           n13152, C1 => n13144, C2 => n1484, ZN => n7603);
   U3943 : NOR4_X1 port map( A1 => n4509, A2 => n4510, A3 => n4511, A4 => n4512
                           , ZN => n4508);
   U3944 : NAND4_X1 port map( A1 => n4537, A2 => n4538, A3 => n4539, A4 => 
                           n4540, ZN => n4509);
   U3945 : NAND4_X1 port map( A1 => n4529, A2 => n4530, A3 => n4531, A4 => 
                           n4532, ZN => n4510);
   U3946 : OAI222_X1 port map( A1 => n16078, A2 => n13155, B1 => n4471, B2 => 
                           n13152, C1 => n13144, C2 => n1483, ZN => n7605);
   U3947 : NOR4_X1 port map( A1 => n4472, A2 => n4473, A3 => n4474, A4 => n4475
                           , ZN => n4471);
   U3948 : NAND4_X1 port map( A1 => n4500, A2 => n4501, A3 => n4502, A4 => 
                           n4503, ZN => n4472);
   U3949 : NAND4_X1 port map( A1 => n4492, A2 => n4493, A3 => n4494, A4 => 
                           n4495, ZN => n4473);
   U3950 : OAI222_X1 port map( A1 => n16077, A2 => n13155, B1 => n4434, B2 => 
                           n13152, C1 => n13144, C2 => n1482, ZN => n7607);
   U3951 : NOR4_X1 port map( A1 => n4435, A2 => n4436, A3 => n4437, A4 => n4438
                           , ZN => n4434);
   U3952 : NAND4_X1 port map( A1 => n4463, A2 => n4464, A3 => n4465, A4 => 
                           n4466, ZN => n4435);
   U3953 : NAND4_X1 port map( A1 => n4455, A2 => n4456, A3 => n4457, A4 => 
                           n4458, ZN => n4436);
   U3954 : OAI222_X1 port map( A1 => n16076, A2 => n13155, B1 => n4323, B2 => 
                           n13152, C1 => n13145, C2 => n1481, ZN => n7609);
   U3955 : NOR4_X1 port map( A1 => n4326, A2 => n4327, A3 => n4328, A4 => n4329
                           , ZN => n4323);
   U3956 : NAND4_X1 port map( A1 => n4408, A2 => n4409, A3 => n4410, A4 => 
                           n4411, ZN => n4326);
   U3957 : NAND4_X1 port map( A1 => n4382, A2 => n4383, A3 => n4384, A4 => 
                           n4385, ZN => n4327);
   U3958 : AOI221_X1 port map( B1 => n13248, B2 => n6174, C1 => n13245, C2 => 
                           n15615, A => n3250, ZN => n3247);
   U3959 : OAI22_X1 port map( A1 => n14952, A2 => n13242, B1 => n15926, B2 => 
                           n13239, ZN => n3250);
   U3960 : AOI221_X1 port map( B1 => n13194, B2 => n5918, C1 => n13191, C2 => 
                           n15305, A => n3258, ZN => n3255);
   U3961 : OAI22_X1 port map( A1 => n15337, A2 => n13188, B1 => n15369, B2 => 
                           n13185, ZN => n3258);
   U3962 : AOI221_X1 port map( B1 => n13248, B2 => n6175, C1 => n13245, C2 => 
                           n15614, A => n3213, ZN => n3210);
   U3963 : OAI22_X1 port map( A1 => n14951, A2 => n13242, B1 => n15925, B2 => 
                           n13239, ZN => n3213);
   U3964 : AOI221_X1 port map( B1 => n13194, B2 => n5919, C1 => n13191, C2 => 
                           n15304, A => n3221, ZN => n3218);
   U3965 : OAI22_X1 port map( A1 => n15336, A2 => n13188, B1 => n15368, B2 => 
                           n13185, ZN => n3221);
   U3966 : AOI221_X1 port map( B1 => n13248, B2 => n6176, C1 => n13245, C2 => 
                           n15613, A => n3176, ZN => n3173);
   U3967 : OAI22_X1 port map( A1 => n14950, A2 => n13242, B1 => n15924, B2 => 
                           n13239, ZN => n3176);
   U3968 : AOI221_X1 port map( B1 => n13194, B2 => n5920, C1 => n13191, C2 => 
                           n15303, A => n3184, ZN => n3181);
   U3969 : OAI22_X1 port map( A1 => n15335, A2 => n13188, B1 => n15367, B2 => 
                           n13185, ZN => n3184);
   U3970 : AOI221_X1 port map( B1 => n13248, B2 => n6177, C1 => n13245, C2 => 
                           n14948, A => n3110, ZN => n3100);
   U3971 : OAI22_X1 port map( A1 => n14949, A2 => n13242, B1 => n15923, B2 => 
                           n13239, ZN => n3110);
   U3972 : AOI221_X1 port map( B1 => n13194, B2 => n5921, C1 => n13191, C2 => 
                           n15302, A => n3136, ZN => n3126);
   U3973 : OAI22_X1 port map( A1 => n15334, A2 => n13188, B1 => n15366, B2 => 
                           n13185, ZN => n3136);
   U3974 : AOI221_X1 port map( B1 => n13020, B2 => n6171, C1 => n13017, C2 => 
                           n15618, A => n4645, ZN => n4642);
   U3975 : OAI22_X1 port map( A1 => n14955, A2 => n13014, B1 => n15929, B2 => 
                           n13011, ZN => n4645);
   U3976 : AOI221_X1 port map( B1 => n12966, B2 => n5915, C1 => n12963, C2 => 
                           n15308, A => n4653, ZN => n4650);
   U3977 : OAI22_X1 port map( A1 => n15340, A2 => n12960, B1 => n15372, B2 => 
                           n12957, ZN => n4653);
   U3978 : AOI221_X1 port map( B1 => n13020, B2 => n6172, C1 => n13017, C2 => 
                           n15617, A => n4608, ZN => n4605);
   U3979 : OAI22_X1 port map( A1 => n14954, A2 => n13014, B1 => n15928, B2 => 
                           n13011, ZN => n4608);
   U3980 : AOI221_X1 port map( B1 => n12966, B2 => n5916, C1 => n12963, C2 => 
                           n15307, A => n4616, ZN => n4613);
   U3981 : OAI22_X1 port map( A1 => n15339, A2 => n12960, B1 => n15371, B2 => 
                           n12957, ZN => n4616);
   U3982 : AOI221_X1 port map( B1 => n13020, B2 => n6173, C1 => n13017, C2 => 
                           n15616, A => n4571, ZN => n4568);
   U3983 : OAI22_X1 port map( A1 => n14953, A2 => n13014, B1 => n15927, B2 => 
                           n13011, ZN => n4571);
   U3984 : AOI221_X1 port map( B1 => n12966, B2 => n5917, C1 => n12963, C2 => 
                           n15306, A => n4579, ZN => n4576);
   U3985 : OAI22_X1 port map( A1 => n15338, A2 => n12960, B1 => n15370, B2 => 
                           n12957, ZN => n4579);
   U3986 : AOI221_X1 port map( B1 => n13020, B2 => n6174, C1 => n13017, C2 => 
                           n15615, A => n4534, ZN => n4531);
   U3987 : OAI22_X1 port map( A1 => n14952, A2 => n13014, B1 => n15926, B2 => 
                           n13011, ZN => n4534);
   U3988 : AOI221_X1 port map( B1 => n12966, B2 => n5918, C1 => n12963, C2 => 
                           n15305, A => n4542, ZN => n4539);
   U3989 : OAI22_X1 port map( A1 => n15337, A2 => n12960, B1 => n15369, B2 => 
                           n12957, ZN => n4542);
   U3990 : AOI221_X1 port map( B1 => n13020, B2 => n6175, C1 => n13017, C2 => 
                           n15614, A => n4497, ZN => n4494);
   U3991 : OAI22_X1 port map( A1 => n14951, A2 => n13014, B1 => n15925, B2 => 
                           n13011, ZN => n4497);
   U3992 : AOI221_X1 port map( B1 => n12966, B2 => n5919, C1 => n12963, C2 => 
                           n15304, A => n4505, ZN => n4502);
   U3993 : OAI22_X1 port map( A1 => n15336, A2 => n12960, B1 => n15368, B2 => 
                           n12957, ZN => n4505);
   U3994 : AOI221_X1 port map( B1 => n13020, B2 => n6176, C1 => n13017, C2 => 
                           n15613, A => n4460, ZN => n4457);
   U3995 : OAI22_X1 port map( A1 => n14950, A2 => n13014, B1 => n15924, B2 => 
                           n13011, ZN => n4460);
   U3996 : AOI221_X1 port map( B1 => n12966, B2 => n5920, C1 => n12963, C2 => 
                           n15303, A => n4468, ZN => n4465);
   U3997 : OAI22_X1 port map( A1 => n15335, A2 => n12960, B1 => n15367, B2 => 
                           n12957, ZN => n4468);
   U3998 : AOI221_X1 port map( B1 => n13020, B2 => n6177, C1 => n13017, C2 => 
                           n14948, A => n4394, ZN => n4384);
   U3999 : OAI22_X1 port map( A1 => n14949, A2 => n13014, B1 => n15923, B2 => 
                           n13011, ZN => n4394);
   U4000 : AOI221_X1 port map( B1 => n12966, B2 => n5921, C1 => n12963, C2 => 
                           n15302, A => n4420, ZN => n4410);
   U4001 : OAI22_X1 port map( A1 => n15334, A2 => n12960, B1 => n15366, B2 => 
                           n12957, ZN => n4420);
   U4002 : AOI221_X1 port map( B1 => n13018, B2 => n6146, C1 => n13015, C2 => 
                           n15681, A => n5712, ZN => n5704);
   U4003 : OAI22_X1 port map( A1 => n14980, A2 => n13012, B1 => n15970, B2 => 
                           n13009, ZN => n5712);
   U4004 : AOI221_X1 port map( B1 => n12964, B2 => n5890, C1 => n12961, C2 => 
                           n15333, A => n5730, ZN => n5724);
   U4005 : OAI22_X1 port map( A1 => n15365, A2 => n12958, B1 => n15397, B2 => 
                           n12955, ZN => n5730);
   U4006 : AOI221_X1 port map( B1 => n13018, B2 => n6147, C1 => n13015, C2 => 
                           n15680, A => n5624, ZN => n5619);
   U4007 : OAI22_X1 port map( A1 => n14979, A2 => n13012, B1 => n15969, B2 => 
                           n13009, ZN => n5624);
   U4008 : AOI221_X1 port map( B1 => n12964, B2 => n5891, C1 => n12961, C2 => 
                           n15332, A => n5638, ZN => n5631);
   U4009 : OAI22_X1 port map( A1 => n15364, A2 => n12958, B1 => n15396, B2 => 
                           n12955, ZN => n5638);
   U4010 : AOI221_X1 port map( B1 => n13018, B2 => n6148, C1 => n13015, C2 => 
                           n15679, A => n5561, ZN => n5558);
   U4011 : OAI22_X1 port map( A1 => n14978, A2 => n13012, B1 => n15968, B2 => 
                           n13009, ZN => n5561);
   U4012 : AOI221_X1 port map( B1 => n12964, B2 => n5892, C1 => n12961, C2 => 
                           n15331, A => n5576, ZN => n5570);
   U4013 : OAI22_X1 port map( A1 => n15363, A2 => n12958, B1 => n15395, B2 => 
                           n12955, ZN => n5576);
   U4014 : AOI221_X1 port map( B1 => n13018, B2 => n6149, C1 => n13015, C2 => 
                           n15678, A => n5500, ZN => n5496);
   U4015 : OAI22_X1 port map( A1 => n14977, A2 => n13012, B1 => n15967, B2 => 
                           n13009, ZN => n5500);
   U4016 : AOI221_X1 port map( B1 => n12964, B2 => n5893, C1 => n12961, C2 => 
                           n15330, A => n5514, ZN => n5509);
   U4017 : OAI22_X1 port map( A1 => n15362, A2 => n12958, B1 => n15394, B2 => 
                           n12955, ZN => n5514);
   U4018 : AOI221_X1 port map( B1 => n13018, B2 => n6150, C1 => n13015, C2 => 
                           n15677, A => n5440, ZN => n5436);
   U4019 : OAI22_X1 port map( A1 => n14976, A2 => n13012, B1 => n15966, B2 => 
                           n13009, ZN => n5440);
   U4020 : AOI221_X1 port map( B1 => n12964, B2 => n5894, C1 => n12961, C2 => 
                           n15329, A => n5451, ZN => n5448);
   U4021 : OAI22_X1 port map( A1 => n15361, A2 => n12958, B1 => n15393, B2 => 
                           n12955, ZN => n5451);
   U4022 : AOI221_X1 port map( B1 => n13018, B2 => n6151, C1 => n13015, C2 => 
                           n15676, A => n5388, ZN => n5382);
   U4023 : OAI22_X1 port map( A1 => n14975, A2 => n13012, B1 => n15965, B2 => 
                           n13009, ZN => n5388);
   U4024 : AOI221_X1 port map( B1 => n12964, B2 => n5895, C1 => n12961, C2 => 
                           n15328, A => n5399, ZN => n5394);
   U4025 : OAI22_X1 port map( A1 => n15360, A2 => n12958, B1 => n15392, B2 => 
                           n12955, ZN => n5399);
   U4026 : AOI221_X1 port map( B1 => n13018, B2 => n6152, C1 => n13015, C2 => 
                           n15675, A => n5348, ZN => n5345);
   U4027 : OAI22_X1 port map( A1 => n14974, A2 => n13012, B1 => n15964, B2 => 
                           n13009, ZN => n5348);
   U4028 : AOI221_X1 port map( B1 => n12964, B2 => n5896, C1 => n12961, C2 => 
                           n15327, A => n5356, ZN => n5353);
   U4029 : OAI22_X1 port map( A1 => n15359, A2 => n12958, B1 => n15391, B2 => 
                           n12955, ZN => n5356);
   U4030 : AOI221_X1 port map( B1 => n13018, B2 => n6153, C1 => n13015, C2 => 
                           n15674, A => n5311, ZN => n5308);
   U4031 : OAI22_X1 port map( A1 => n14973, A2 => n13012, B1 => n15963, B2 => 
                           n13009, ZN => n5311);
   U4032 : AOI221_X1 port map( B1 => n12964, B2 => n5897, C1 => n12961, C2 => 
                           n15326, A => n5319, ZN => n5316);
   U4033 : OAI22_X1 port map( A1 => n15358, A2 => n12958, B1 => n15390, B2 => 
                           n12955, ZN => n5319);
   U4034 : AOI221_X1 port map( B1 => n13018, B2 => n6154, C1 => n13015, C2 => 
                           n15673, A => n5274, ZN => n5271);
   U4035 : OAI22_X1 port map( A1 => n14972, A2 => n13012, B1 => n15962, B2 => 
                           n13009, ZN => n5274);
   U4036 : AOI221_X1 port map( B1 => n12964, B2 => n5898, C1 => n12961, C2 => 
                           n15325, A => n5282, ZN => n5279);
   U4037 : OAI22_X1 port map( A1 => n15357, A2 => n12958, B1 => n15389, B2 => 
                           n12955, ZN => n5282);
   U4038 : AOI221_X1 port map( B1 => n13018, B2 => n6155, C1 => n13015, C2 => 
                           n15672, A => n5237, ZN => n5234);
   U4039 : OAI22_X1 port map( A1 => n14971, A2 => n13012, B1 => n15961, B2 => 
                           n13009, ZN => n5237);
   U4040 : AOI221_X1 port map( B1 => n12964, B2 => n5899, C1 => n12961, C2 => 
                           n15324, A => n5245, ZN => n5242);
   U4041 : OAI22_X1 port map( A1 => n15356, A2 => n12958, B1 => n15388, B2 => 
                           n12955, ZN => n5245);
   U4042 : AOI221_X1 port map( B1 => n13018, B2 => n6156, C1 => n13015, C2 => 
                           n15671, A => n5200, ZN => n5197);
   U4043 : OAI22_X1 port map( A1 => n14970, A2 => n13012, B1 => n15960, B2 => 
                           n13009, ZN => n5200);
   U4044 : AOI221_X1 port map( B1 => n12964, B2 => n5900, C1 => n12961, C2 => 
                           n15323, A => n5208, ZN => n5205);
   U4045 : OAI22_X1 port map( A1 => n15355, A2 => n12958, B1 => n15387, B2 => 
                           n12955, ZN => n5208);
   U4046 : AOI221_X1 port map( B1 => n13018, B2 => n6157, C1 => n13015, C2 => 
                           n15670, A => n5163, ZN => n5160);
   U4047 : OAI22_X1 port map( A1 => n14969, A2 => n13012, B1 => n15959, B2 => 
                           n13009, ZN => n5163);
   U4048 : AOI221_X1 port map( B1 => n12964, B2 => n5901, C1 => n12961, C2 => 
                           n15322, A => n5171, ZN => n5168);
   U4049 : OAI22_X1 port map( A1 => n15354, A2 => n12958, B1 => n15386, B2 => 
                           n12955, ZN => n5171);
   U4050 : AOI221_X1 port map( B1 => n13019, B2 => n6158, C1 => n13016, C2 => 
                           n15669, A => n5126, ZN => n5123);
   U4051 : OAI22_X1 port map( A1 => n14968, A2 => n13013, B1 => n15958, B2 => 
                           n13010, ZN => n5126);
   U4052 : AOI221_X1 port map( B1 => n12965, B2 => n5902, C1 => n12962, C2 => 
                           n15321, A => n5134, ZN => n5131);
   U4053 : OAI22_X1 port map( A1 => n15353, A2 => n12959, B1 => n15385, B2 => 
                           n12956, ZN => n5134);
   U4054 : AOI221_X1 port map( B1 => n13019, B2 => n6159, C1 => n13016, C2 => 
                           n15668, A => n5089, ZN => n5086);
   U4055 : OAI22_X1 port map( A1 => n14967, A2 => n13013, B1 => n15957, B2 => 
                           n13010, ZN => n5089);
   U4056 : AOI221_X1 port map( B1 => n12965, B2 => n5903, C1 => n12962, C2 => 
                           n15320, A => n5097, ZN => n5094);
   U4057 : OAI22_X1 port map( A1 => n15352, A2 => n12959, B1 => n15384, B2 => 
                           n12956, ZN => n5097);
   U4058 : AOI221_X1 port map( B1 => n13019, B2 => n6160, C1 => n13016, C2 => 
                           n15667, A => n5052, ZN => n5049);
   U4059 : OAI22_X1 port map( A1 => n14966, A2 => n13013, B1 => n15956, B2 => 
                           n13010, ZN => n5052);
   U4060 : AOI221_X1 port map( B1 => n12965, B2 => n5904, C1 => n12962, C2 => 
                           n15319, A => n5060, ZN => n5057);
   U4061 : OAI22_X1 port map( A1 => n15351, A2 => n12959, B1 => n15383, B2 => 
                           n12956, ZN => n5060);
   U4062 : AOI221_X1 port map( B1 => n13019, B2 => n6161, C1 => n13016, C2 => 
                           n15666, A => n5015, ZN => n5012);
   U4063 : OAI22_X1 port map( A1 => n14965, A2 => n13013, B1 => n15955, B2 => 
                           n13010, ZN => n5015);
   U4064 : AOI221_X1 port map( B1 => n12965, B2 => n5905, C1 => n12962, C2 => 
                           n15318, A => n5023, ZN => n5020);
   U4065 : OAI22_X1 port map( A1 => n15350, A2 => n12959, B1 => n15382, B2 => 
                           n12956, ZN => n5023);
   U4066 : AOI221_X1 port map( B1 => n13019, B2 => n6162, C1 => n13016, C2 => 
                           n15665, A => n4978, ZN => n4975);
   U4067 : OAI22_X1 port map( A1 => n14964, A2 => n13013, B1 => n15954, B2 => 
                           n13010, ZN => n4978);
   U4068 : AOI221_X1 port map( B1 => n12965, B2 => n5906, C1 => n12962, C2 => 
                           n15317, A => n4986, ZN => n4983);
   U4069 : OAI22_X1 port map( A1 => n15349, A2 => n12959, B1 => n15381, B2 => 
                           n12956, ZN => n4986);
   U4070 : AOI221_X1 port map( B1 => n13019, B2 => n6163, C1 => n13016, C2 => 
                           n15664, A => n4941, ZN => n4938);
   U4071 : OAI22_X1 port map( A1 => n14963, A2 => n13013, B1 => n15953, B2 => 
                           n13010, ZN => n4941);
   U4072 : AOI221_X1 port map( B1 => n12965, B2 => n5907, C1 => n12962, C2 => 
                           n15316, A => n4949, ZN => n4946);
   U4073 : OAI22_X1 port map( A1 => n15348, A2 => n12959, B1 => n15380, B2 => 
                           n12956, ZN => n4949);
   U4074 : AOI221_X1 port map( B1 => n13019, B2 => n6164, C1 => n13016, C2 => 
                           n15663, A => n4904, ZN => n4901);
   U4075 : OAI22_X1 port map( A1 => n14962, A2 => n13013, B1 => n15952, B2 => 
                           n13010, ZN => n4904);
   U4076 : AOI221_X1 port map( B1 => n12965, B2 => n5908, C1 => n12962, C2 => 
                           n15315, A => n4912, ZN => n4909);
   U4077 : OAI22_X1 port map( A1 => n15347, A2 => n12959, B1 => n15379, B2 => 
                           n12956, ZN => n4912);
   U4078 : AOI221_X1 port map( B1 => n13019, B2 => n6165, C1 => n13016, C2 => 
                           n15662, A => n4867, ZN => n4864);
   U4079 : OAI22_X1 port map( A1 => n14961, A2 => n13013, B1 => n15951, B2 => 
                           n13010, ZN => n4867);
   U4080 : AOI221_X1 port map( B1 => n12965, B2 => n5909, C1 => n12962, C2 => 
                           n15314, A => n4875, ZN => n4872);
   U4081 : OAI22_X1 port map( A1 => n15346, A2 => n12959, B1 => n15378, B2 => 
                           n12956, ZN => n4875);
   U4082 : AOI221_X1 port map( B1 => n13019, B2 => n6166, C1 => n13016, C2 => 
                           n15661, A => n4830, ZN => n4827);
   U4083 : OAI22_X1 port map( A1 => n14960, A2 => n13013, B1 => n15950, B2 => 
                           n13010, ZN => n4830);
   U4084 : AOI221_X1 port map( B1 => n12965, B2 => n5910, C1 => n12962, C2 => 
                           n15313, A => n4838, ZN => n4835);
   U4085 : OAI22_X1 port map( A1 => n15345, A2 => n12959, B1 => n15377, B2 => 
                           n12956, ZN => n4838);
   U4086 : AOI221_X1 port map( B1 => n13019, B2 => n6167, C1 => n13016, C2 => 
                           n15660, A => n4793, ZN => n4790);
   U4087 : OAI22_X1 port map( A1 => n14959, A2 => n13013, B1 => n15949, B2 => 
                           n13010, ZN => n4793);
   U4088 : AOI221_X1 port map( B1 => n12965, B2 => n5911, C1 => n12962, C2 => 
                           n15312, A => n4801, ZN => n4798);
   U4089 : OAI22_X1 port map( A1 => n15344, A2 => n12959, B1 => n15376, B2 => 
                           n12956, ZN => n4801);
   U4090 : AOI221_X1 port map( B1 => n13019, B2 => n6168, C1 => n13016, C2 => 
                           n15659, A => n4756, ZN => n4753);
   U4091 : OAI22_X1 port map( A1 => n14958, A2 => n13013, B1 => n15948, B2 => 
                           n13010, ZN => n4756);
   U4092 : AOI221_X1 port map( B1 => n12965, B2 => n5912, C1 => n12962, C2 => 
                           n15311, A => n4764, ZN => n4761);
   U4093 : OAI22_X1 port map( A1 => n15343, A2 => n12959, B1 => n15375, B2 => 
                           n12956, ZN => n4764);
   U4094 : AOI221_X1 port map( B1 => n13019, B2 => n6169, C1 => n13016, C2 => 
                           n15658, A => n4719, ZN => n4716);
   U4095 : OAI22_X1 port map( A1 => n14957, A2 => n13013, B1 => n15947, B2 => 
                           n13010, ZN => n4719);
   U4096 : AOI221_X1 port map( B1 => n12965, B2 => n5913, C1 => n12962, C2 => 
                           n15310, A => n4727, ZN => n4724);
   U4097 : OAI22_X1 port map( A1 => n15342, A2 => n12959, B1 => n15374, B2 => 
                           n12956, ZN => n4727);
   U4098 : AOI221_X1 port map( B1 => n12966, B2 => n5914, C1 => n12963, C2 => 
                           n15309, A => n4690, ZN => n4687);
   U4099 : OAI22_X1 port map( A1 => n15341, A2 => n12960, B1 => n15373, B2 => 
                           n12957, ZN => n4690);
   U4100 : AOI221_X1 port map( B1 => n13246, B2 => n6146, C1 => n13243, C2 => 
                           n15681, A => n4300, ZN => n4296);
   U4101 : OAI22_X1 port map( A1 => n14980, A2 => n13240, B1 => n15970, B2 => 
                           n13237, ZN => n4300);
   U4102 : AOI221_X1 port map( B1 => n13192, B2 => n5890, C1 => n13189, C2 => 
                           n15333, A => n4309, ZN => n4306);
   U4103 : OAI22_X1 port map( A1 => n15365, A2 => n13186, B1 => n15397, B2 => 
                           n13183, ZN => n4309);
   U4104 : AOI221_X1 port map( B1 => n13246, B2 => n6147, C1 => n13243, C2 => 
                           n15680, A => n4249, ZN => n4246);
   U4105 : OAI22_X1 port map( A1 => n14979, A2 => n13240, B1 => n15969, B2 => 
                           n13237, ZN => n4249);
   U4106 : AOI221_X1 port map( B1 => n13192, B2 => n5891, C1 => n13189, C2 => 
                           n15332, A => n4257, ZN => n4254);
   U4107 : OAI22_X1 port map( A1 => n15364, A2 => n13186, B1 => n15396, B2 => 
                           n13183, ZN => n4257);
   U4108 : AOI221_X1 port map( B1 => n13246, B2 => n6148, C1 => n13243, C2 => 
                           n15679, A => n4212, ZN => n4209);
   U4109 : OAI22_X1 port map( A1 => n14978, A2 => n13240, B1 => n15968, B2 => 
                           n13237, ZN => n4212);
   U4110 : AOI221_X1 port map( B1 => n13192, B2 => n5892, C1 => n13189, C2 => 
                           n15331, A => n4220, ZN => n4217);
   U4111 : OAI22_X1 port map( A1 => n15363, A2 => n13186, B1 => n15395, B2 => 
                           n13183, ZN => n4220);
   U4112 : AOI221_X1 port map( B1 => n13246, B2 => n6149, C1 => n13243, C2 => 
                           n15678, A => n4175, ZN => n4172);
   U4113 : OAI22_X1 port map( A1 => n14977, A2 => n13240, B1 => n15967, B2 => 
                           n13237, ZN => n4175);
   U4114 : AOI221_X1 port map( B1 => n13192, B2 => n5893, C1 => n13189, C2 => 
                           n15330, A => n4183, ZN => n4180);
   U4115 : OAI22_X1 port map( A1 => n15362, A2 => n13186, B1 => n15394, B2 => 
                           n13183, ZN => n4183);
   U4116 : AOI221_X1 port map( B1 => n13246, B2 => n6150, C1 => n13243, C2 => 
                           n15677, A => n4138, ZN => n4135);
   U4117 : OAI22_X1 port map( A1 => n14976, A2 => n13240, B1 => n15966, B2 => 
                           n13237, ZN => n4138);
   U4118 : AOI221_X1 port map( B1 => n13192, B2 => n5894, C1 => n13189, C2 => 
                           n15329, A => n4146, ZN => n4143);
   U4119 : OAI22_X1 port map( A1 => n15361, A2 => n13186, B1 => n15393, B2 => 
                           n13183, ZN => n4146);
   U4120 : AOI221_X1 port map( B1 => n13246, B2 => n6151, C1 => n13243, C2 => 
                           n15676, A => n4101, ZN => n4098);
   U4121 : OAI22_X1 port map( A1 => n14975, A2 => n13240, B1 => n15965, B2 => 
                           n13237, ZN => n4101);
   U4122 : AOI221_X1 port map( B1 => n13192, B2 => n5895, C1 => n13189, C2 => 
                           n15328, A => n4109, ZN => n4106);
   U4123 : OAI22_X1 port map( A1 => n15360, A2 => n13186, B1 => n15392, B2 => 
                           n13183, ZN => n4109);
   U4124 : AOI221_X1 port map( B1 => n13246, B2 => n6152, C1 => n13243, C2 => 
                           n15675, A => n4064, ZN => n4061);
   U4125 : OAI22_X1 port map( A1 => n14974, A2 => n13240, B1 => n15964, B2 => 
                           n13237, ZN => n4064);
   U4126 : AOI221_X1 port map( B1 => n13192, B2 => n5896, C1 => n13189, C2 => 
                           n15327, A => n4072, ZN => n4069);
   U4127 : OAI22_X1 port map( A1 => n15359, A2 => n13186, B1 => n15391, B2 => 
                           n13183, ZN => n4072);
   U4128 : AOI221_X1 port map( B1 => n13246, B2 => n6153, C1 => n13243, C2 => 
                           n15674, A => n4027, ZN => n4024);
   U4129 : OAI22_X1 port map( A1 => n14973, A2 => n13240, B1 => n15963, B2 => 
                           n13237, ZN => n4027);
   U4130 : AOI221_X1 port map( B1 => n13192, B2 => n5897, C1 => n13189, C2 => 
                           n15326, A => n4035, ZN => n4032);
   U4131 : OAI22_X1 port map( A1 => n15358, A2 => n13186, B1 => n15390, B2 => 
                           n13183, ZN => n4035);
   U4132 : AOI221_X1 port map( B1 => n13246, B2 => n6154, C1 => n13243, C2 => 
                           n15673, A => n3990, ZN => n3987);
   U4133 : OAI22_X1 port map( A1 => n14972, A2 => n13240, B1 => n15962, B2 => 
                           n13237, ZN => n3990);
   U4134 : AOI221_X1 port map( B1 => n13192, B2 => n5898, C1 => n13189, C2 => 
                           n15325, A => n3998, ZN => n3995);
   U4135 : OAI22_X1 port map( A1 => n15357, A2 => n13186, B1 => n15389, B2 => 
                           n13183, ZN => n3998);
   U4136 : AOI221_X1 port map( B1 => n13246, B2 => n6155, C1 => n13243, C2 => 
                           n15672, A => n3953, ZN => n3950);
   U4137 : OAI22_X1 port map( A1 => n14971, A2 => n13240, B1 => n15961, B2 => 
                           n13237, ZN => n3953);
   U4138 : AOI221_X1 port map( B1 => n13192, B2 => n5899, C1 => n13189, C2 => 
                           n15324, A => n3961, ZN => n3958);
   U4139 : OAI22_X1 port map( A1 => n15356, A2 => n13186, B1 => n15388, B2 => 
                           n13183, ZN => n3961);
   U4140 : AOI221_X1 port map( B1 => n13246, B2 => n6156, C1 => n13243, C2 => 
                           n15671, A => n3916, ZN => n3913);
   U4141 : OAI22_X1 port map( A1 => n14970, A2 => n13240, B1 => n15960, B2 => 
                           n13237, ZN => n3916);
   U4142 : AOI221_X1 port map( B1 => n13192, B2 => n5900, C1 => n13189, C2 => 
                           n15323, A => n3924, ZN => n3921);
   U4143 : OAI22_X1 port map( A1 => n15355, A2 => n13186, B1 => n15387, B2 => 
                           n13183, ZN => n3924);
   U4144 : AOI221_X1 port map( B1 => n13246, B2 => n6157, C1 => n13243, C2 => 
                           n15670, A => n3879, ZN => n3876);
   U4145 : OAI22_X1 port map( A1 => n14969, A2 => n13240, B1 => n15959, B2 => 
                           n13237, ZN => n3879);
   U4146 : AOI221_X1 port map( B1 => n13192, B2 => n5901, C1 => n13189, C2 => 
                           n15322, A => n3887, ZN => n3884);
   U4147 : OAI22_X1 port map( A1 => n15354, A2 => n13186, B1 => n15386, B2 => 
                           n13183, ZN => n3887);
   U4148 : AOI221_X1 port map( B1 => n13247, B2 => n6158, C1 => n13244, C2 => 
                           n15669, A => n3842, ZN => n3839);
   U4149 : OAI22_X1 port map( A1 => n14968, A2 => n13241, B1 => n15958, B2 => 
                           n13238, ZN => n3842);
   U4150 : AOI221_X1 port map( B1 => n13193, B2 => n5902, C1 => n13190, C2 => 
                           n15321, A => n3850, ZN => n3847);
   U4151 : OAI22_X1 port map( A1 => n15353, A2 => n13187, B1 => n15385, B2 => 
                           n13184, ZN => n3850);
   U4152 : AOI221_X1 port map( B1 => n13247, B2 => n6159, C1 => n13244, C2 => 
                           n15668, A => n3805, ZN => n3802);
   U4153 : OAI22_X1 port map( A1 => n14967, A2 => n13241, B1 => n15957, B2 => 
                           n13238, ZN => n3805);
   U4154 : AOI221_X1 port map( B1 => n13193, B2 => n5903, C1 => n13190, C2 => 
                           n15320, A => n3813, ZN => n3810);
   U4155 : OAI22_X1 port map( A1 => n15352, A2 => n13187, B1 => n15384, B2 => 
                           n13184, ZN => n3813);
   U4156 : AOI221_X1 port map( B1 => n13247, B2 => n6160, C1 => n13244, C2 => 
                           n15667, A => n3768, ZN => n3765);
   U4157 : OAI22_X1 port map( A1 => n14966, A2 => n13241, B1 => n15956, B2 => 
                           n13238, ZN => n3768);
   U4158 : AOI221_X1 port map( B1 => n13193, B2 => n5904, C1 => n13190, C2 => 
                           n15319, A => n3776, ZN => n3773);
   U4159 : OAI22_X1 port map( A1 => n15351, A2 => n13187, B1 => n15383, B2 => 
                           n13184, ZN => n3776);
   U4160 : AOI221_X1 port map( B1 => n13247, B2 => n6161, C1 => n13244, C2 => 
                           n15666, A => n3731, ZN => n3728);
   U4161 : OAI22_X1 port map( A1 => n14965, A2 => n13241, B1 => n15955, B2 => 
                           n13238, ZN => n3731);
   U4162 : AOI221_X1 port map( B1 => n13193, B2 => n5905, C1 => n13190, C2 => 
                           n15318, A => n3739, ZN => n3736);
   U4163 : OAI22_X1 port map( A1 => n15350, A2 => n13187, B1 => n15382, B2 => 
                           n13184, ZN => n3739);
   U4164 : AOI221_X1 port map( B1 => n13247, B2 => n6162, C1 => n13244, C2 => 
                           n15665, A => n3694, ZN => n3691);
   U4165 : OAI22_X1 port map( A1 => n14964, A2 => n13241, B1 => n15954, B2 => 
                           n13238, ZN => n3694);
   U4166 : AOI221_X1 port map( B1 => n13193, B2 => n5906, C1 => n13190, C2 => 
                           n15317, A => n3702, ZN => n3699);
   U4167 : OAI22_X1 port map( A1 => n15349, A2 => n13187, B1 => n15381, B2 => 
                           n13184, ZN => n3702);
   U4168 : AOI221_X1 port map( B1 => n13247, B2 => n6163, C1 => n13244, C2 => 
                           n15664, A => n3657, ZN => n3654);
   U4169 : OAI22_X1 port map( A1 => n14963, A2 => n13241, B1 => n15953, B2 => 
                           n13238, ZN => n3657);
   U4170 : AOI221_X1 port map( B1 => n13193, B2 => n5907, C1 => n13190, C2 => 
                           n15316, A => n3665, ZN => n3662);
   U4171 : OAI22_X1 port map( A1 => n15348, A2 => n13187, B1 => n15380, B2 => 
                           n13184, ZN => n3665);
   U4172 : AOI221_X1 port map( B1 => n13247, B2 => n6164, C1 => n13244, C2 => 
                           n15663, A => n3620, ZN => n3617);
   U4173 : OAI22_X1 port map( A1 => n14962, A2 => n13241, B1 => n15952, B2 => 
                           n13238, ZN => n3620);
   U4174 : AOI221_X1 port map( B1 => n13193, B2 => n5908, C1 => n13190, C2 => 
                           n15315, A => n3628, ZN => n3625);
   U4175 : OAI22_X1 port map( A1 => n15347, A2 => n13187, B1 => n15379, B2 => 
                           n13184, ZN => n3628);
   U4176 : AOI221_X1 port map( B1 => n13247, B2 => n6165, C1 => n13244, C2 => 
                           n15662, A => n3583, ZN => n3580);
   U4177 : OAI22_X1 port map( A1 => n14961, A2 => n13241, B1 => n15951, B2 => 
                           n13238, ZN => n3583);
   U4178 : AOI221_X1 port map( B1 => n13193, B2 => n5909, C1 => n13190, C2 => 
                           n15314, A => n3591, ZN => n3588);
   U4179 : OAI22_X1 port map( A1 => n15346, A2 => n13187, B1 => n15378, B2 => 
                           n13184, ZN => n3591);
   U4180 : AOI221_X1 port map( B1 => n13247, B2 => n6166, C1 => n13244, C2 => 
                           n15661, A => n3546, ZN => n3543);
   U4181 : OAI22_X1 port map( A1 => n14960, A2 => n13241, B1 => n15950, B2 => 
                           n13238, ZN => n3546);
   U4182 : AOI221_X1 port map( B1 => n13193, B2 => n5910, C1 => n13190, C2 => 
                           n15313, A => n3554, ZN => n3551);
   U4183 : OAI22_X1 port map( A1 => n15345, A2 => n13187, B1 => n15377, B2 => 
                           n13184, ZN => n3554);
   U4184 : AOI221_X1 port map( B1 => n13247, B2 => n6167, C1 => n13244, C2 => 
                           n15660, A => n3509, ZN => n3506);
   U4185 : OAI22_X1 port map( A1 => n14959, A2 => n13241, B1 => n15949, B2 => 
                           n13238, ZN => n3509);
   U4186 : AOI221_X1 port map( B1 => n13193, B2 => n5911, C1 => n13190, C2 => 
                           n15312, A => n3517, ZN => n3514);
   U4187 : OAI22_X1 port map( A1 => n15344, A2 => n13187, B1 => n15376, B2 => 
                           n13184, ZN => n3517);
   U4188 : AOI221_X1 port map( B1 => n13247, B2 => n6168, C1 => n13244, C2 => 
                           n15659, A => n3472, ZN => n3469);
   U4189 : OAI22_X1 port map( A1 => n14958, A2 => n13241, B1 => n15948, B2 => 
                           n13238, ZN => n3472);
   U4190 : AOI221_X1 port map( B1 => n13193, B2 => n5912, C1 => n13190, C2 => 
                           n15311, A => n3480, ZN => n3477);
   U4191 : OAI22_X1 port map( A1 => n15343, A2 => n13187, B1 => n15375, B2 => 
                           n13184, ZN => n3480);
   U4192 : AOI221_X1 port map( B1 => n13247, B2 => n6169, C1 => n13244, C2 => 
                           n15658, A => n3435, ZN => n3432);
   U4193 : OAI22_X1 port map( A1 => n14957, A2 => n13241, B1 => n15947, B2 => 
                           n13238, ZN => n3435);
   U4194 : AOI221_X1 port map( B1 => n13193, B2 => n5913, C1 => n13190, C2 => 
                           n15310, A => n3443, ZN => n3440);
   U4195 : OAI22_X1 port map( A1 => n15342, A2 => n13187, B1 => n15374, B2 => 
                           n13184, ZN => n3443);
   U4196 : AOI221_X1 port map( B1 => n13194, B2 => n5914, C1 => n13191, C2 => 
                           n15309, A => n3406, ZN => n3403);
   U4197 : OAI22_X1 port map( A1 => n15341, A2 => n13188, B1 => n15373, B2 => 
                           n13185, ZN => n3406);
   U4198 : AOI221_X1 port map( B1 => n13248, B2 => n6171, C1 => n13245, C2 => 
                           n15618, A => n3361, ZN => n3358);
   U4199 : OAI22_X1 port map( A1 => n14955, A2 => n13242, B1 => n15929, B2 => 
                           n13239, ZN => n3361);
   U4200 : AOI221_X1 port map( B1 => n13194, B2 => n5915, C1 => n13191, C2 => 
                           n15308, A => n3369, ZN => n3366);
   U4201 : OAI22_X1 port map( A1 => n15340, A2 => n13188, B1 => n15372, B2 => 
                           n13185, ZN => n3369);
   U4202 : AOI221_X1 port map( B1 => n13248, B2 => n6172, C1 => n13245, C2 => 
                           n15617, A => n3324, ZN => n3321);
   U4203 : OAI22_X1 port map( A1 => n14954, A2 => n13242, B1 => n15928, B2 => 
                           n13239, ZN => n3324);
   U4204 : AOI221_X1 port map( B1 => n13194, B2 => n5916, C1 => n13191, C2 => 
                           n15307, A => n3332, ZN => n3329);
   U4205 : OAI22_X1 port map( A1 => n15339, A2 => n13188, B1 => n15371, B2 => 
                           n13185, ZN => n3332);
   U4206 : AOI221_X1 port map( B1 => n13248, B2 => n6173, C1 => n13245, C2 => 
                           n15616, A => n3287, ZN => n3284);
   U4207 : OAI22_X1 port map( A1 => n14953, A2 => n13242, B1 => n15927, B2 => 
                           n13239, ZN => n3287);
   U4208 : AOI221_X1 port map( B1 => n13194, B2 => n5917, C1 => n13191, C2 => 
                           n15306, A => n3295, ZN => n3292);
   U4209 : OAI22_X1 port map( A1 => n15338, A2 => n13188, B1 => n15370, B2 => 
                           n13185, ZN => n3295);
   U4210 : OAI222_X1 port map( A1 => n16079, A2 => n13383, B1 => n3224, B2 => 
                           n13380, C1 => n13372, C2 => n1452, ZN => n7667);
   U4211 : NOR4_X1 port map( A1 => n3225, A2 => n3226, A3 => n3227, A4 => n3228
                           , ZN => n3224);
   U4212 : NAND4_X1 port map( A1 => n3253, A2 => n3254, A3 => n3255, A4 => 
                           n3256, ZN => n3225);
   U4213 : NAND4_X1 port map( A1 => n3245, A2 => n3246, A3 => n3247, A4 => 
                           n3248, ZN => n3226);
   U4214 : OAI222_X1 port map( A1 => n16078, A2 => n13383, B1 => n3187, B2 => 
                           n13380, C1 => n13372, C2 => n1451, ZN => n7669);
   U4215 : NOR4_X1 port map( A1 => n3188, A2 => n3189, A3 => n3190, A4 => n3191
                           , ZN => n3187);
   U4216 : NAND4_X1 port map( A1 => n3216, A2 => n3217, A3 => n3218, A4 => 
                           n3219, ZN => n3188);
   U4217 : NAND4_X1 port map( A1 => n3208, A2 => n3209, A3 => n3210, A4 => 
                           n3211, ZN => n3189);
   U4218 : OAI222_X1 port map( A1 => n16077, A2 => n13383, B1 => n3150, B2 => 
                           n13380, C1 => n13372, C2 => n1450, ZN => n7671);
   U4219 : NOR4_X1 port map( A1 => n3151, A2 => n3152, A3 => n3153, A4 => n3154
                           , ZN => n3150);
   U4220 : NAND4_X1 port map( A1 => n3179, A2 => n3180, A3 => n3181, A4 => 
                           n3182, ZN => n3151);
   U4221 : NAND4_X1 port map( A1 => n3171, A2 => n3172, A3 => n3173, A4 => 
                           n3174, ZN => n3152);
   U4222 : OAI222_X1 port map( A1 => n16076, A2 => n13383, B1 => n3039, B2 => 
                           n13380, C1 => n13373, C2 => n1449, ZN => n7673);
   U4223 : NOR4_X1 port map( A1 => n3042, A2 => n3043, A3 => n3044, A4 => n3045
                           , ZN => n3039);
   U4224 : NAND4_X1 port map( A1 => n3124, A2 => n3125, A3 => n3126, A4 => 
                           n3127, ZN => n3042);
   U4225 : NAND4_X1 port map( A1 => n3098, A2 => n3099, A3 => n3100, A4 => 
                           n3101, ZN => n3043);
   U4226 : OAI222_X1 port map( A1 => n16107, A2 => n13153, B1 => n5641, B2 => 
                           n13150, C1 => n13146, C2 => n1512, ZN => n7547);
   U4227 : NOR4_X1 port map( A1 => n5644, A2 => n5646, A3 => n5648, A4 => n5649
                           , ZN => n5641);
   U4228 : NAND4_X1 port map( A1 => n5720, A2 => n5722, A3 => n5724, A4 => 
                           n5726, ZN => n5644);
   U4229 : NAND4_X1 port map( A1 => n5700, A2 => n5702, A3 => n5704, A4 => 
                           n5706, ZN => n5646);
   U4230 : OAI222_X1 port map( A1 => n16106, A2 => n13153, B1 => n5580, B2 => 
                           n13150, C1 => n13146, C2 => n1511, ZN => n7549);
   U4231 : NOR4_X1 port map( A1 => n5581, A2 => n5584, A3 => n5586, A4 => n5588
                           , ZN => n5580);
   U4232 : NAND4_X1 port map( A1 => n5629, A2 => n5630, A3 => n5631, A4 => 
                           n5634, ZN => n5581);
   U4233 : NAND4_X1 port map( A1 => n5616, A2 => n5618, A3 => n5619, A4 => 
                           n5620, ZN => n5584);
   U4234 : OAI222_X1 port map( A1 => n16105, A2 => n13153, B1 => n5519, B2 => 
                           n13150, C1 => n13146, C2 => n1510, ZN => n7551);
   U4235 : NOR4_X1 port map( A1 => n5520, A2 => n5521, A3 => n5524, A4 => n5526
                           , ZN => n5519);
   U4236 : NAND4_X1 port map( A1 => n5568, A2 => n5569, A3 => n5570, A4 => 
                           n5571, ZN => n5520);
   U4237 : NAND4_X1 port map( A1 => n5554, A2 => n5556, A3 => n5558, A4 => 
                           n5559, ZN => n5521);
   U4238 : OAI222_X1 port map( A1 => n16104, A2 => n13153, B1 => n5458, B2 => 
                           n13150, C1 => n13146, C2 => n1509, ZN => n7553);
   U4239 : NOR4_X1 port map( A1 => n5459, A2 => n5460, A3 => n5461, A4 => n5464
                           , ZN => n5458);
   U4240 : NAND4_X1 port map( A1 => n5506, A2 => n5508, A3 => n5509, A4 => 
                           n5510, ZN => n5459);
   U4241 : NAND4_X1 port map( A1 => n5491, A2 => n5494, A3 => n5496, A4 => 
                           n5498, ZN => n5460);
   U4242 : OAI222_X1 port map( A1 => n16103, A2 => n13153, B1 => n5402, B2 => 
                           n13150, C1 => n13146, C2 => n1508, ZN => n7555);
   U4243 : NOR4_X1 port map( A1 => n5404, A2 => n5406, A3 => n5408, A4 => n5409
                           , ZN => n5402);
   U4244 : NAND4_X1 port map( A1 => n5444, A2 => n5446, A3 => n5448, A4 => 
                           n5449, ZN => n5404);
   U4245 : NAND4_X1 port map( A1 => n5432, A2 => n5434, A3 => n5436, A4 => 
                           n5438, ZN => n5406);
   U4246 : OAI222_X1 port map( A1 => n16102, A2 => n13153, B1 => n5359, B2 => 
                           n13150, C1 => n13146, C2 => n1507, ZN => n7557);
   U4247 : NOR4_X1 port map( A1 => n5360, A2 => n5361, A3 => n5362, A4 => n5363
                           , ZN => n5359);
   U4248 : NAND4_X1 port map( A1 => n5391, A2 => n5392, A3 => n5394, A4 => 
                           n5396, ZN => n5360);
   U4249 : NAND4_X1 port map( A1 => n5380, A2 => n5381, A3 => n5382, A4 => 
                           n5384, ZN => n5361);
   U4250 : OAI222_X1 port map( A1 => n16101, A2 => n13153, B1 => n5322, B2 => 
                           n13150, C1 => n13146, C2 => n1506, ZN => n7559);
   U4251 : NOR4_X1 port map( A1 => n5323, A2 => n5324, A3 => n5325, A4 => n5326
                           , ZN => n5322);
   U4252 : NAND4_X1 port map( A1 => n5351, A2 => n5352, A3 => n5353, A4 => 
                           n5354, ZN => n5323);
   U4253 : NAND4_X1 port map( A1 => n5343, A2 => n5344, A3 => n5345, A4 => 
                           n5346, ZN => n5324);
   U4254 : OAI222_X1 port map( A1 => n16100, A2 => n13153, B1 => n5285, B2 => 
                           n13150, C1 => n13146, C2 => n1505, ZN => n7561);
   U4255 : NOR4_X1 port map( A1 => n5286, A2 => n5287, A3 => n5288, A4 => n5289
                           , ZN => n5285);
   U4256 : NAND4_X1 port map( A1 => n5314, A2 => n5315, A3 => n5316, A4 => 
                           n5317, ZN => n5286);
   U4257 : NAND4_X1 port map( A1 => n5306, A2 => n5307, A3 => n5308, A4 => 
                           n5309, ZN => n5287);
   U4258 : OAI222_X1 port map( A1 => n16099, A2 => n13153, B1 => n5248, B2 => 
                           n13150, C1 => n13145, C2 => n1504, ZN => n7563);
   U4259 : NOR4_X1 port map( A1 => n5249, A2 => n5250, A3 => n5251, A4 => n5252
                           , ZN => n5248);
   U4260 : NAND4_X1 port map( A1 => n5277, A2 => n5278, A3 => n5279, A4 => 
                           n5280, ZN => n5249);
   U4261 : NAND4_X1 port map( A1 => n5269, A2 => n5270, A3 => n5271, A4 => 
                           n5272, ZN => n5250);
   U4262 : OAI222_X1 port map( A1 => n16098, A2 => n13153, B1 => n5211, B2 => 
                           n13150, C1 => n13145, C2 => n1503, ZN => n7565);
   U4263 : NOR4_X1 port map( A1 => n5212, A2 => n5213, A3 => n5214, A4 => n5215
                           , ZN => n5211);
   U4264 : NAND4_X1 port map( A1 => n5240, A2 => n5241, A3 => n5242, A4 => 
                           n5243, ZN => n5212);
   U4265 : NAND4_X1 port map( A1 => n5232, A2 => n5233, A3 => n5234, A4 => 
                           n5235, ZN => n5213);
   U4266 : OAI222_X1 port map( A1 => n16097, A2 => n13153, B1 => n5174, B2 => 
                           n13150, C1 => n13145, C2 => n1502, ZN => n7567);
   U4267 : NOR4_X1 port map( A1 => n5175, A2 => n5176, A3 => n5177, A4 => n5178
                           , ZN => n5174);
   U4268 : NAND4_X1 port map( A1 => n5203, A2 => n5204, A3 => n5205, A4 => 
                           n5206, ZN => n5175);
   U4269 : NAND4_X1 port map( A1 => n5195, A2 => n5196, A3 => n5197, A4 => 
                           n5198, ZN => n5176);
   U4270 : OAI222_X1 port map( A1 => n16096, A2 => n13153, B1 => n5137, B2 => 
                           n13150, C1 => n13145, C2 => n1501, ZN => n7569);
   U4271 : NOR4_X1 port map( A1 => n5138, A2 => n5139, A3 => n5140, A4 => n5141
                           , ZN => n5137);
   U4272 : NAND4_X1 port map( A1 => n5166, A2 => n5167, A3 => n5168, A4 => 
                           n5169, ZN => n5138);
   U4273 : NAND4_X1 port map( A1 => n5158, A2 => n5159, A3 => n5160, A4 => 
                           n5161, ZN => n5139);
   U4274 : OAI222_X1 port map( A1 => n16095, A2 => n13154, B1 => n5100, B2 => 
                           n13151, C1 => n13145, C2 => n1500, ZN => n7571);
   U4275 : NOR4_X1 port map( A1 => n5101, A2 => n5102, A3 => n5103, A4 => n5104
                           , ZN => n5100);
   U4276 : NAND4_X1 port map( A1 => n5129, A2 => n5130, A3 => n5131, A4 => 
                           n5132, ZN => n5101);
   U4277 : NAND4_X1 port map( A1 => n5121, A2 => n5122, A3 => n5123, A4 => 
                           n5124, ZN => n5102);
   U4278 : OAI222_X1 port map( A1 => n16094, A2 => n13154, B1 => n5063, B2 => 
                           n13151, C1 => n13145, C2 => n1499, ZN => n7573);
   U4279 : NOR4_X1 port map( A1 => n5064, A2 => n5065, A3 => n5066, A4 => n5067
                           , ZN => n5063);
   U4280 : NAND4_X1 port map( A1 => n5092, A2 => n5093, A3 => n5094, A4 => 
                           n5095, ZN => n5064);
   U4281 : NAND4_X1 port map( A1 => n5084, A2 => n5085, A3 => n5086, A4 => 
                           n5087, ZN => n5065);
   U4282 : OAI222_X1 port map( A1 => n16093, A2 => n13154, B1 => n5026, B2 => 
                           n13151, C1 => n13145, C2 => n1498, ZN => n7575);
   U4283 : NOR4_X1 port map( A1 => n5027, A2 => n5028, A3 => n5029, A4 => n5030
                           , ZN => n5026);
   U4284 : NAND4_X1 port map( A1 => n5055, A2 => n5056, A3 => n5057, A4 => 
                           n5058, ZN => n5027);
   U4285 : NAND4_X1 port map( A1 => n5047, A2 => n5048, A3 => n5049, A4 => 
                           n5050, ZN => n5028);
   U4286 : OAI222_X1 port map( A1 => n16092, A2 => n13154, B1 => n4989, B2 => 
                           n13151, C1 => n13145, C2 => n1497, ZN => n7577);
   U4287 : NOR4_X1 port map( A1 => n4990, A2 => n4991, A3 => n4992, A4 => n4993
                           , ZN => n4989);
   U4288 : NAND4_X1 port map( A1 => n5018, A2 => n5019, A3 => n5020, A4 => 
                           n5021, ZN => n4990);
   U4289 : NAND4_X1 port map( A1 => n5010, A2 => n5011, A3 => n5012, A4 => 
                           n5013, ZN => n4991);
   U4290 : OAI222_X1 port map( A1 => n16091, A2 => n13154, B1 => n4952, B2 => 
                           n13151, C1 => n13145, C2 => n1496, ZN => n7579);
   U4291 : NOR4_X1 port map( A1 => n4953, A2 => n4954, A3 => n4955, A4 => n4956
                           , ZN => n4952);
   U4292 : NAND4_X1 port map( A1 => n4981, A2 => n4982, A3 => n4983, A4 => 
                           n4984, ZN => n4953);
   U4293 : NAND4_X1 port map( A1 => n4973, A2 => n4974, A3 => n4975, A4 => 
                           n4976, ZN => n4954);
   U4294 : OAI222_X1 port map( A1 => n16090, A2 => n13154, B1 => n4915, B2 => 
                           n13151, C1 => n13145, C2 => n1495, ZN => n7581);
   U4295 : NOR4_X1 port map( A1 => n4916, A2 => n4917, A3 => n4918, A4 => n4919
                           , ZN => n4915);
   U4296 : NAND4_X1 port map( A1 => n4944, A2 => n4945, A3 => n4946, A4 => 
                           n4947, ZN => n4916);
   U4297 : NAND4_X1 port map( A1 => n4936, A2 => n4937, A3 => n4938, A4 => 
                           n4939, ZN => n4917);
   U4298 : OAI222_X1 port map( A1 => n16089, A2 => n13154, B1 => n4878, B2 => 
                           n13151, C1 => n13145, C2 => n1494, ZN => n7583);
   U4299 : NOR4_X1 port map( A1 => n4879, A2 => n4880, A3 => n4881, A4 => n4882
                           , ZN => n4878);
   U4300 : NAND4_X1 port map( A1 => n4907, A2 => n4908, A3 => n4909, A4 => 
                           n4910, ZN => n4879);
   U4301 : NAND4_X1 port map( A1 => n4899, A2 => n4900, A3 => n4901, A4 => 
                           n4902, ZN => n4880);
   U4302 : OAI222_X1 port map( A1 => n16088, A2 => n13154, B1 => n4841, B2 => 
                           n13151, C1 => n13144, C2 => n1493, ZN => n7585);
   U4303 : NOR4_X1 port map( A1 => n4842, A2 => n4843, A3 => n4844, A4 => n4845
                           , ZN => n4841);
   U4304 : NAND4_X1 port map( A1 => n4870, A2 => n4871, A3 => n4872, A4 => 
                           n4873, ZN => n4842);
   U4305 : NAND4_X1 port map( A1 => n4862, A2 => n4863, A3 => n4864, A4 => 
                           n4865, ZN => n4843);
   U4306 : OAI222_X1 port map( A1 => n16087, A2 => n13154, B1 => n4804, B2 => 
                           n13151, C1 => n13144, C2 => n1492, ZN => n7587);
   U4307 : NOR4_X1 port map( A1 => n4805, A2 => n4806, A3 => n4807, A4 => n4808
                           , ZN => n4804);
   U4308 : NAND4_X1 port map( A1 => n4833, A2 => n4834, A3 => n4835, A4 => 
                           n4836, ZN => n4805);
   U4309 : NAND4_X1 port map( A1 => n4825, A2 => n4826, A3 => n4827, A4 => 
                           n4828, ZN => n4806);
   U4310 : OAI222_X1 port map( A1 => n16086, A2 => n13154, B1 => n4767, B2 => 
                           n13151, C1 => n13144, C2 => n1491, ZN => n7589);
   U4311 : NOR4_X1 port map( A1 => n4768, A2 => n4769, A3 => n4770, A4 => n4771
                           , ZN => n4767);
   U4312 : NAND4_X1 port map( A1 => n4796, A2 => n4797, A3 => n4798, A4 => 
                           n4799, ZN => n4768);
   U4313 : NAND4_X1 port map( A1 => n4788, A2 => n4789, A3 => n4790, A4 => 
                           n4791, ZN => n4769);
   U4314 : OAI222_X1 port map( A1 => n16085, A2 => n13154, B1 => n4730, B2 => 
                           n13151, C1 => n13144, C2 => n1490, ZN => n7591);
   U4315 : NOR4_X1 port map( A1 => n4731, A2 => n4732, A3 => n4733, A4 => n4734
                           , ZN => n4730);
   U4316 : NAND4_X1 port map( A1 => n4759, A2 => n4760, A3 => n4761, A4 => 
                           n4762, ZN => n4731);
   U4317 : NAND4_X1 port map( A1 => n4751, A2 => n4752, A3 => n4753, A4 => 
                           n4754, ZN => n4732);
   U4318 : OAI222_X1 port map( A1 => n16084, A2 => n13154, B1 => n4693, B2 => 
                           n13151, C1 => n13144, C2 => n1489, ZN => n7593);
   U4319 : NOR4_X1 port map( A1 => n4694, A2 => n4695, A3 => n4696, A4 => n4697
                           , ZN => n4693);
   U4320 : NAND4_X1 port map( A1 => n4722, A2 => n4723, A3 => n4724, A4 => 
                           n4725, ZN => n4694);
   U4321 : NAND4_X1 port map( A1 => n4714, A2 => n4715, A3 => n4716, A4 => 
                           n4717, ZN => n4695);
   U4322 : OAI222_X1 port map( A1 => n16083, A2 => n13154, B1 => n4656, B2 => 
                           n13152, C1 => n13144, C2 => n1488, ZN => n7595);
   U4323 : NOR4_X1 port map( A1 => n4657, A2 => n4658, A3 => n4659, A4 => n4660
                           , ZN => n4656);
   U4324 : NAND4_X1 port map( A1 => n4685, A2 => n4686, A3 => n4687, A4 => 
                           n4688, ZN => n4657);
   U4325 : NAND4_X1 port map( A1 => n4677, A2 => n4678, A3 => n4679, A4 => 
                           n4680, ZN => n4658);
   U4326 : OAI222_X1 port map( A1 => n16107, A2 => n13381, B1 => n4260, B2 => 
                           n13378, C1 => n13374, C2 => n1480, ZN => n7611);
   U4327 : NOR4_X1 port map( A1 => n4261, A2 => n4262, A3 => n4263, A4 => n4264
                           , ZN => n4260);
   U4328 : NAND4_X1 port map( A1 => n4304, A2 => n4305, A3 => n4306, A4 => 
                           n4307, ZN => n4261);
   U4329 : NAND4_X1 port map( A1 => n4294, A2 => n4295, A3 => n4296, A4 => 
                           n4297, ZN => n4262);
   U4330 : OAI222_X1 port map( A1 => n16106, A2 => n13381, B1 => n4223, B2 => 
                           n13378, C1 => n13374, C2 => n1479, ZN => n7613);
   U4331 : NOR4_X1 port map( A1 => n4224, A2 => n4225, A3 => n4226, A4 => n4227
                           , ZN => n4223);
   U4332 : NAND4_X1 port map( A1 => n4252, A2 => n4253, A3 => n4254, A4 => 
                           n4255, ZN => n4224);
   U4333 : NAND4_X1 port map( A1 => n4244, A2 => n4245, A3 => n4246, A4 => 
                           n4247, ZN => n4225);
   U4334 : OAI222_X1 port map( A1 => n16105, A2 => n13381, B1 => n4186, B2 => 
                           n13378, C1 => n13374, C2 => n1478, ZN => n7615);
   U4335 : NOR4_X1 port map( A1 => n4187, A2 => n4188, A3 => n4189, A4 => n4190
                           , ZN => n4186);
   U4336 : NAND4_X1 port map( A1 => n4215, A2 => n4216, A3 => n4217, A4 => 
                           n4218, ZN => n4187);
   U4337 : NAND4_X1 port map( A1 => n4207, A2 => n4208, A3 => n4209, A4 => 
                           n4210, ZN => n4188);
   U4338 : OAI222_X1 port map( A1 => n16104, A2 => n13381, B1 => n4149, B2 => 
                           n13378, C1 => n13374, C2 => n1477, ZN => n7617);
   U4339 : NOR4_X1 port map( A1 => n4150, A2 => n4151, A3 => n4152, A4 => n4153
                           , ZN => n4149);
   U4340 : NAND4_X1 port map( A1 => n4178, A2 => n4179, A3 => n4180, A4 => 
                           n4181, ZN => n4150);
   U4341 : NAND4_X1 port map( A1 => n4170, A2 => n4171, A3 => n4172, A4 => 
                           n4173, ZN => n4151);
   U4342 : OAI222_X1 port map( A1 => n16103, A2 => n13381, B1 => n4112, B2 => 
                           n13378, C1 => n13374, C2 => n1476, ZN => n7619);
   U4343 : NOR4_X1 port map( A1 => n4113, A2 => n4114, A3 => n4115, A4 => n4116
                           , ZN => n4112);
   U4344 : NAND4_X1 port map( A1 => n4141, A2 => n4142, A3 => n4143, A4 => 
                           n4144, ZN => n4113);
   U4345 : NAND4_X1 port map( A1 => n4133, A2 => n4134, A3 => n4135, A4 => 
                           n4136, ZN => n4114);
   U4346 : OAI222_X1 port map( A1 => n16102, A2 => n13381, B1 => n4075, B2 => 
                           n13378, C1 => n13374, C2 => n1475, ZN => n7621);
   U4347 : NOR4_X1 port map( A1 => n4076, A2 => n4077, A3 => n4078, A4 => n4079
                           , ZN => n4075);
   U4348 : NAND4_X1 port map( A1 => n4104, A2 => n4105, A3 => n4106, A4 => 
                           n4107, ZN => n4076);
   U4349 : NAND4_X1 port map( A1 => n4096, A2 => n4097, A3 => n4098, A4 => 
                           n4099, ZN => n4077);
   U4350 : OAI222_X1 port map( A1 => n16101, A2 => n13381, B1 => n4038, B2 => 
                           n13378, C1 => n13374, C2 => n1474, ZN => n7623);
   U4351 : NOR4_X1 port map( A1 => n4039, A2 => n4040, A3 => n4041, A4 => n4042
                           , ZN => n4038);
   U4352 : NAND4_X1 port map( A1 => n4067, A2 => n4068, A3 => n4069, A4 => 
                           n4070, ZN => n4039);
   U4353 : NAND4_X1 port map( A1 => n4059, A2 => n4060, A3 => n4061, A4 => 
                           n4062, ZN => n4040);
   U4354 : OAI222_X1 port map( A1 => n16100, A2 => n13381, B1 => n4001, B2 => 
                           n13378, C1 => n13374, C2 => n1473, ZN => n7625);
   U4355 : NOR4_X1 port map( A1 => n4002, A2 => n4003, A3 => n4004, A4 => n4005
                           , ZN => n4001);
   U4356 : NAND4_X1 port map( A1 => n4030, A2 => n4031, A3 => n4032, A4 => 
                           n4033, ZN => n4002);
   U4357 : NAND4_X1 port map( A1 => n4022, A2 => n4023, A3 => n4024, A4 => 
                           n4025, ZN => n4003);
   U4358 : OAI222_X1 port map( A1 => n16099, A2 => n13381, B1 => n3964, B2 => 
                           n13378, C1 => n13373, C2 => n1472, ZN => n7627);
   U4359 : NOR4_X1 port map( A1 => n3965, A2 => n3966, A3 => n3967, A4 => n3968
                           , ZN => n3964);
   U4360 : NAND4_X1 port map( A1 => n3993, A2 => n3994, A3 => n3995, A4 => 
                           n3996, ZN => n3965);
   U4361 : NAND4_X1 port map( A1 => n3985, A2 => n3986, A3 => n3987, A4 => 
                           n3988, ZN => n3966);
   U4362 : OAI222_X1 port map( A1 => n16098, A2 => n13381, B1 => n3927, B2 => 
                           n13378, C1 => n13373, C2 => n1471, ZN => n7629);
   U4363 : NOR4_X1 port map( A1 => n3928, A2 => n3929, A3 => n3930, A4 => n3931
                           , ZN => n3927);
   U4364 : NAND4_X1 port map( A1 => n3956, A2 => n3957, A3 => n3958, A4 => 
                           n3959, ZN => n3928);
   U4365 : NAND4_X1 port map( A1 => n3948, A2 => n3949, A3 => n3950, A4 => 
                           n3951, ZN => n3929);
   U4366 : OAI222_X1 port map( A1 => n16097, A2 => n13381, B1 => n3890, B2 => 
                           n13378, C1 => n13373, C2 => n1470, ZN => n7631);
   U4367 : NOR4_X1 port map( A1 => n3891, A2 => n3892, A3 => n3893, A4 => n3894
                           , ZN => n3890);
   U4368 : NAND4_X1 port map( A1 => n3919, A2 => n3920, A3 => n3921, A4 => 
                           n3922, ZN => n3891);
   U4369 : NAND4_X1 port map( A1 => n3911, A2 => n3912, A3 => n3913, A4 => 
                           n3914, ZN => n3892);
   U4370 : OAI222_X1 port map( A1 => n16096, A2 => n13381, B1 => n3853, B2 => 
                           n13378, C1 => n13373, C2 => n1469, ZN => n7633);
   U4371 : NOR4_X1 port map( A1 => n3854, A2 => n3855, A3 => n3856, A4 => n3857
                           , ZN => n3853);
   U4372 : NAND4_X1 port map( A1 => n3882, A2 => n3883, A3 => n3884, A4 => 
                           n3885, ZN => n3854);
   U4373 : NAND4_X1 port map( A1 => n3874, A2 => n3875, A3 => n3876, A4 => 
                           n3877, ZN => n3855);
   U4374 : OAI222_X1 port map( A1 => n16095, A2 => n13382, B1 => n3816, B2 => 
                           n13379, C1 => n13373, C2 => n1468, ZN => n7635);
   U4375 : NOR4_X1 port map( A1 => n3817, A2 => n3818, A3 => n3819, A4 => n3820
                           , ZN => n3816);
   U4376 : NAND4_X1 port map( A1 => n3845, A2 => n3846, A3 => n3847, A4 => 
                           n3848, ZN => n3817);
   U4377 : NAND4_X1 port map( A1 => n3837, A2 => n3838, A3 => n3839, A4 => 
                           n3840, ZN => n3818);
   U4378 : OAI222_X1 port map( A1 => n16094, A2 => n13382, B1 => n3779, B2 => 
                           n13379, C1 => n13373, C2 => n1467, ZN => n7637);
   U4379 : NOR4_X1 port map( A1 => n3780, A2 => n3781, A3 => n3782, A4 => n3783
                           , ZN => n3779);
   U4380 : NAND4_X1 port map( A1 => n3808, A2 => n3809, A3 => n3810, A4 => 
                           n3811, ZN => n3780);
   U4381 : NAND4_X1 port map( A1 => n3800, A2 => n3801, A3 => n3802, A4 => 
                           n3803, ZN => n3781);
   U4382 : OAI222_X1 port map( A1 => n16093, A2 => n13382, B1 => n3742, B2 => 
                           n13379, C1 => n13373, C2 => n1466, ZN => n7639);
   U4383 : NOR4_X1 port map( A1 => n3743, A2 => n3744, A3 => n3745, A4 => n3746
                           , ZN => n3742);
   U4384 : NAND4_X1 port map( A1 => n3771, A2 => n3772, A3 => n3773, A4 => 
                           n3774, ZN => n3743);
   U4385 : NAND4_X1 port map( A1 => n3763, A2 => n3764, A3 => n3765, A4 => 
                           n3766, ZN => n3744);
   U4386 : OAI222_X1 port map( A1 => n16092, A2 => n13382, B1 => n3705, B2 => 
                           n13379, C1 => n13373, C2 => n1465, ZN => n7641);
   U4387 : NOR4_X1 port map( A1 => n3706, A2 => n3707, A3 => n3708, A4 => n3709
                           , ZN => n3705);
   U4388 : NAND4_X1 port map( A1 => n3734, A2 => n3735, A3 => n3736, A4 => 
                           n3737, ZN => n3706);
   U4389 : NAND4_X1 port map( A1 => n3726, A2 => n3727, A3 => n3728, A4 => 
                           n3729, ZN => n3707);
   U4390 : OAI222_X1 port map( A1 => n16091, A2 => n13382, B1 => n3668, B2 => 
                           n13379, C1 => n13373, C2 => n1464, ZN => n7643);
   U4391 : NOR4_X1 port map( A1 => n3669, A2 => n3670, A3 => n3671, A4 => n3672
                           , ZN => n3668);
   U4392 : NAND4_X1 port map( A1 => n3697, A2 => n3698, A3 => n3699, A4 => 
                           n3700, ZN => n3669);
   U4393 : NAND4_X1 port map( A1 => n3689, A2 => n3690, A3 => n3691, A4 => 
                           n3692, ZN => n3670);
   U4394 : OAI222_X1 port map( A1 => n16090, A2 => n13382, B1 => n3631, B2 => 
                           n13379, C1 => n13373, C2 => n1463, ZN => n7645);
   U4395 : NOR4_X1 port map( A1 => n3632, A2 => n3633, A3 => n3634, A4 => n3635
                           , ZN => n3631);
   U4396 : NAND4_X1 port map( A1 => n3660, A2 => n3661, A3 => n3662, A4 => 
                           n3663, ZN => n3632);
   U4397 : NAND4_X1 port map( A1 => n3652, A2 => n3653, A3 => n3654, A4 => 
                           n3655, ZN => n3633);
   U4398 : OAI222_X1 port map( A1 => n16089, A2 => n13382, B1 => n3594, B2 => 
                           n13379, C1 => n13373, C2 => n1462, ZN => n7647);
   U4399 : NOR4_X1 port map( A1 => n3595, A2 => n3596, A3 => n3597, A4 => n3598
                           , ZN => n3594);
   U4400 : NAND4_X1 port map( A1 => n3623, A2 => n3624, A3 => n3625, A4 => 
                           n3626, ZN => n3595);
   U4401 : NAND4_X1 port map( A1 => n3615, A2 => n3616, A3 => n3617, A4 => 
                           n3618, ZN => n3596);
   U4402 : OAI222_X1 port map( A1 => n16088, A2 => n13382, B1 => n3557, B2 => 
                           n13379, C1 => n13372, C2 => n1461, ZN => n7649);
   U4403 : NOR4_X1 port map( A1 => n3558, A2 => n3559, A3 => n3560, A4 => n3561
                           , ZN => n3557);
   U4404 : NAND4_X1 port map( A1 => n3586, A2 => n3587, A3 => n3588, A4 => 
                           n3589, ZN => n3558);
   U4405 : NAND4_X1 port map( A1 => n3578, A2 => n3579, A3 => n3580, A4 => 
                           n3581, ZN => n3559);
   U4406 : OAI222_X1 port map( A1 => n16087, A2 => n13382, B1 => n3520, B2 => 
                           n13379, C1 => n13372, C2 => n1460, ZN => n7651);
   U4407 : NOR4_X1 port map( A1 => n3521, A2 => n3522, A3 => n3523, A4 => n3524
                           , ZN => n3520);
   U4408 : NAND4_X1 port map( A1 => n3549, A2 => n3550, A3 => n3551, A4 => 
                           n3552, ZN => n3521);
   U4409 : NAND4_X1 port map( A1 => n3541, A2 => n3542, A3 => n3543, A4 => 
                           n3544, ZN => n3522);
   U4410 : OAI222_X1 port map( A1 => n16086, A2 => n13382, B1 => n3483, B2 => 
                           n13379, C1 => n13372, C2 => n1459, ZN => n7653);
   U4411 : NOR4_X1 port map( A1 => n3484, A2 => n3485, A3 => n3486, A4 => n3487
                           , ZN => n3483);
   U4412 : NAND4_X1 port map( A1 => n3512, A2 => n3513, A3 => n3514, A4 => 
                           n3515, ZN => n3484);
   U4413 : NAND4_X1 port map( A1 => n3504, A2 => n3505, A3 => n3506, A4 => 
                           n3507, ZN => n3485);
   U4414 : OAI222_X1 port map( A1 => n16085, A2 => n13382, B1 => n3446, B2 => 
                           n13379, C1 => n13372, C2 => n1458, ZN => n7655);
   U4415 : NOR4_X1 port map( A1 => n3447, A2 => n3448, A3 => n3449, A4 => n3450
                           , ZN => n3446);
   U4416 : NAND4_X1 port map( A1 => n3475, A2 => n3476, A3 => n3477, A4 => 
                           n3478, ZN => n3447);
   U4417 : NAND4_X1 port map( A1 => n3467, A2 => n3468, A3 => n3469, A4 => 
                           n3470, ZN => n3448);
   U4418 : OAI222_X1 port map( A1 => n16084, A2 => n13382, B1 => n3409, B2 => 
                           n13379, C1 => n13372, C2 => n1457, ZN => n7657);
   U4419 : NOR4_X1 port map( A1 => n3410, A2 => n3411, A3 => n3412, A4 => n3413
                           , ZN => n3409);
   U4420 : NAND4_X1 port map( A1 => n3438, A2 => n3439, A3 => n3440, A4 => 
                           n3441, ZN => n3410);
   U4421 : NAND4_X1 port map( A1 => n3430, A2 => n3431, A3 => n3432, A4 => 
                           n3433, ZN => n3411);
   U4422 : OAI222_X1 port map( A1 => n16083, A2 => n13382, B1 => n3372, B2 => 
                           n13380, C1 => n13372, C2 => n1456, ZN => n7659);
   U4423 : NOR4_X1 port map( A1 => n3373, A2 => n3374, A3 => n3375, A4 => n3376
                           , ZN => n3372);
   U4424 : NAND4_X1 port map( A1 => n3401, A2 => n3402, A3 => n3403, A4 => 
                           n3404, ZN => n3373);
   U4425 : NAND4_X1 port map( A1 => n3393, A2 => n3394, A3 => n3395, A4 => 
                           n3396, ZN => n3374);
   U4426 : OAI222_X1 port map( A1 => n16082, A2 => n13383, B1 => n3335, B2 => 
                           n13380, C1 => n13372, C2 => n1455, ZN => n7661);
   U4427 : NOR4_X1 port map( A1 => n3336, A2 => n3337, A3 => n3338, A4 => n3339
                           , ZN => n3335);
   U4428 : NAND4_X1 port map( A1 => n3364, A2 => n3365, A3 => n3366, A4 => 
                           n3367, ZN => n3336);
   U4429 : NAND4_X1 port map( A1 => n3356, A2 => n3357, A3 => n3358, A4 => 
                           n3359, ZN => n3337);
   U4430 : OAI222_X1 port map( A1 => n16081, A2 => n13383, B1 => n3298, B2 => 
                           n13380, C1 => n13372, C2 => n1454, ZN => n7663);
   U4431 : NOR4_X1 port map( A1 => n3299, A2 => n3300, A3 => n3301, A4 => n3302
                           , ZN => n3298);
   U4432 : NAND4_X1 port map( A1 => n3327, A2 => n3328, A3 => n3329, A4 => 
                           n3330, ZN => n3299);
   U4433 : NAND4_X1 port map( A1 => n3319, A2 => n3320, A3 => n3321, A4 => 
                           n3322, ZN => n3300);
   U4434 : OAI222_X1 port map( A1 => n16080, A2 => n13383, B1 => n3261, B2 => 
                           n13380, C1 => n13372, C2 => n1453, ZN => n7665);
   U4435 : NOR4_X1 port map( A1 => n3262, A2 => n3263, A3 => n3264, A4 => n3265
                           , ZN => n3261);
   U4436 : NAND4_X1 port map( A1 => n3290, A2 => n3291, A3 => n3292, A4 => 
                           n3293, ZN => n3262);
   U4437 : NAND4_X1 port map( A1 => n3282, A2 => n3283, A3 => n3284, A4 => 
                           n3285, ZN => n3263);
   U4438 : AOI221_X1 port map( B1 => n13236, B2 => n6238, C1 => n13233, C2 => 
                           n15561, A => n3251, ZN => n3246);
   U4439 : OAI222_X1 port map( A1 => n14919, A2 => n13230, B1 => n14855, B2 => 
                           n13227, C1 => n14887, C2 => n13224, ZN => n3251);
   U4440 : AOI221_X1 port map( B1 => n13236, B2 => n6239, C1 => n13233, C2 => 
                           n15560, A => n3214, ZN => n3209);
   U4441 : OAI222_X1 port map( A1 => n14918, A2 => n13230, B1 => n14854, B2 => 
                           n13227, C1 => n14886, C2 => n13224, ZN => n3214);
   U4442 : AOI221_X1 port map( B1 => n13236, B2 => n6240, C1 => n13233, C2 => 
                           n15559, A => n3177, ZN => n3172);
   U4443 : OAI222_X1 port map( A1 => n14917, A2 => n13230, B1 => n14853, B2 => 
                           n13227, C1 => n14885, C2 => n13224, ZN => n3177);
   U4444 : AOI221_X1 port map( B1 => n13236, B2 => n6241, C1 => n13233, C2 => 
                           n15558, A => n3115, ZN => n3099);
   U4445 : OAI222_X1 port map( A1 => n14916, A2 => n13230, B1 => n14852, B2 => 
                           n13227, C1 => n14884, C2 => n13224, ZN => n3115);
   U4446 : AOI221_X1 port map( B1 => n13008, B2 => n6235, C1 => n13005, C2 => 
                           n15564, A => n4646, ZN => n4641);
   U4447 : OAI222_X1 port map( A1 => n14922, A2 => n13002, B1 => n14858, B2 => 
                           n12999, C1 => n14890, C2 => n12996, ZN => n4646);
   U4448 : AOI221_X1 port map( B1 => n13008, B2 => n6236, C1 => n13005, C2 => 
                           n15563, A => n4609, ZN => n4604);
   U4449 : OAI222_X1 port map( A1 => n14921, A2 => n13002, B1 => n14857, B2 => 
                           n12999, C1 => n14889, C2 => n12996, ZN => n4609);
   U4450 : AOI221_X1 port map( B1 => n13008, B2 => n6237, C1 => n13005, C2 => 
                           n15562, A => n4572, ZN => n4567);
   U4451 : OAI222_X1 port map( A1 => n14920, A2 => n13002, B1 => n14856, B2 => 
                           n12999, C1 => n14888, C2 => n12996, ZN => n4572);
   U4452 : AOI221_X1 port map( B1 => n13008, B2 => n6238, C1 => n13005, C2 => 
                           n15561, A => n4535, ZN => n4530);
   U4453 : OAI222_X1 port map( A1 => n14919, A2 => n13002, B1 => n14855, B2 => 
                           n12999, C1 => n14887, C2 => n12996, ZN => n4535);
   U4454 : AOI221_X1 port map( B1 => n13008, B2 => n6239, C1 => n13005, C2 => 
                           n15560, A => n4498, ZN => n4493);
   U4455 : OAI222_X1 port map( A1 => n14918, A2 => n13002, B1 => n14854, B2 => 
                           n12999, C1 => n14886, C2 => n12996, ZN => n4498);
   U4456 : AOI221_X1 port map( B1 => n13008, B2 => n6240, C1 => n13005, C2 => 
                           n15559, A => n4461, ZN => n4456);
   U4457 : OAI222_X1 port map( A1 => n14917, A2 => n13002, B1 => n14853, B2 => 
                           n12999, C1 => n14885, C2 => n12996, ZN => n4461);
   U4458 : AOI221_X1 port map( B1 => n13008, B2 => n6241, C1 => n13005, C2 => 
                           n15558, A => n4399, ZN => n4383);
   U4459 : OAI222_X1 port map( A1 => n14916, A2 => n13002, B1 => n14852, B2 => 
                           n12999, C1 => n14884, C2 => n12996, ZN => n4399);
   U4460 : AOI221_X1 port map( B1 => n13006, B2 => n6210, C1 => n13003, C2 => 
                           n15705, A => n5716, ZN => n5702);
   U4461 : OAI222_X1 port map( A1 => n14947, A2 => n13000, B1 => n14883, B2 => 
                           n12997, C1 => n14915, C2 => n12994, ZN => n5716);
   U4462 : AOI221_X1 port map( B1 => n12952, B2 => n5954, C1 => n12949, C2 => 
                           n15205, A => n5734, ZN => n5722);
   U4463 : OAI222_X1 port map( A1 => n15301, A2 => n12946, B1 => n15237, B2 => 
                           n12943, C1 => n15269, C2 => n12940, ZN => n5734);
   U4464 : AOI221_X1 port map( B1 => n13006, B2 => n6211, C1 => n13003, C2 => 
                           n15704, A => n5626, ZN => n5618);
   U4465 : OAI222_X1 port map( A1 => n14946, A2 => n13000, B1 => n14882, B2 => 
                           n12997, C1 => n14914, C2 => n12994, ZN => n5626);
   U4466 : AOI221_X1 port map( B1 => n12952, B2 => n5955, C1 => n12949, C2 => 
                           n15204, A => n5639, ZN => n5630);
   U4467 : OAI222_X1 port map( A1 => n15300, A2 => n12946, B1 => n15236, B2 => 
                           n12943, C1 => n15268, C2 => n12940, ZN => n5639);
   U4468 : AOI221_X1 port map( B1 => n13006, B2 => n6212, C1 => n13003, C2 => 
                           n15703, A => n5564, ZN => n5556);
   U4469 : OAI222_X1 port map( A1 => n14945, A2 => n13000, B1 => n14881, B2 => 
                           n12997, C1 => n14913, C2 => n12994, ZN => n5564);
   U4470 : AOI221_X1 port map( B1 => n12952, B2 => n5956, C1 => n12949, C2 => 
                           n15203, A => n5578, ZN => n5569);
   U4471 : OAI222_X1 port map( A1 => n15299, A2 => n12946, B1 => n15235, B2 => 
                           n12943, C1 => n15267, C2 => n12940, ZN => n5578);
   U4472 : AOI221_X1 port map( B1 => n13006, B2 => n6213, C1 => n13003, C2 => 
                           n15702, A => n5501, ZN => n5494);
   U4473 : OAI222_X1 port map( A1 => n14944, A2 => n13000, B1 => n14880, B2 => 
                           n12997, C1 => n14912, C2 => n12994, ZN => n5501);
   U4474 : AOI221_X1 port map( B1 => n12952, B2 => n5957, C1 => n12949, C2 => 
                           n15202, A => n5516, ZN => n5508);
   U4475 : OAI222_X1 port map( A1 => n15298, A2 => n12946, B1 => n15234, B2 => 
                           n12943, C1 => n15266, C2 => n12940, ZN => n5516);
   U4476 : AOI221_X1 port map( B1 => n13006, B2 => n6214, C1 => n13003, C2 => 
                           n15701, A => n5441, ZN => n5434);
   U4477 : OAI222_X1 port map( A1 => n14943, A2 => n13000, B1 => n14879, B2 => 
                           n12997, C1 => n14911, C2 => n12994, ZN => n5441);
   U4478 : AOI221_X1 port map( B1 => n12952, B2 => n5958, C1 => n12949, C2 => 
                           n15201, A => n5454, ZN => n5446);
   U4479 : OAI222_X1 port map( A1 => n15297, A2 => n12946, B1 => n15233, B2 => 
                           n12943, C1 => n15265, C2 => n12940, ZN => n5454);
   U4480 : AOI221_X1 port map( B1 => n13006, B2 => n6215, C1 => n13003, C2 => 
                           n15700, A => n5389, ZN => n5381);
   U4481 : OAI222_X1 port map( A1 => n14942, A2 => n13000, B1 => n14878, B2 => 
                           n12997, C1 => n14910, C2 => n12994, ZN => n5389);
   U4482 : AOI221_X1 port map( B1 => n12952, B2 => n5959, C1 => n12949, C2 => 
                           n15200, A => n5400, ZN => n5392);
   U4483 : OAI222_X1 port map( A1 => n15296, A2 => n12946, B1 => n15232, B2 => 
                           n12943, C1 => n15264, C2 => n12940, ZN => n5400);
   U4484 : AOI221_X1 port map( B1 => n13006, B2 => n6216, C1 => n13003, C2 => 
                           n15699, A => n5349, ZN => n5344);
   U4485 : OAI222_X1 port map( A1 => n14941, A2 => n13000, B1 => n14877, B2 => 
                           n12997, C1 => n14909, C2 => n12994, ZN => n5349);
   U4486 : AOI221_X1 port map( B1 => n12952, B2 => n5960, C1 => n12949, C2 => 
                           n15199, A => n5357, ZN => n5352);
   U4487 : OAI222_X1 port map( A1 => n15295, A2 => n12946, B1 => n15231, B2 => 
                           n12943, C1 => n15263, C2 => n12940, ZN => n5357);
   U4488 : AOI221_X1 port map( B1 => n13006, B2 => n6217, C1 => n13003, C2 => 
                           n15698, A => n5312, ZN => n5307);
   U4489 : OAI222_X1 port map( A1 => n14940, A2 => n13000, B1 => n14876, B2 => 
                           n12997, C1 => n14908, C2 => n12994, ZN => n5312);
   U4490 : AOI221_X1 port map( B1 => n12952, B2 => n5961, C1 => n12949, C2 => 
                           n15198, A => n5320, ZN => n5315);
   U4491 : OAI222_X1 port map( A1 => n15294, A2 => n12946, B1 => n15230, B2 => 
                           n12943, C1 => n15262, C2 => n12940, ZN => n5320);
   U4492 : AOI221_X1 port map( B1 => n13006, B2 => n6218, C1 => n13003, C2 => 
                           n15697, A => n5275, ZN => n5270);
   U4493 : OAI222_X1 port map( A1 => n14939, A2 => n13000, B1 => n14875, B2 => 
                           n12997, C1 => n14907, C2 => n12994, ZN => n5275);
   U4494 : AOI221_X1 port map( B1 => n12952, B2 => n5962, C1 => n12949, C2 => 
                           n15197, A => n5283, ZN => n5278);
   U4495 : OAI222_X1 port map( A1 => n15293, A2 => n12946, B1 => n15229, B2 => 
                           n12943, C1 => n15261, C2 => n12940, ZN => n5283);
   U4496 : AOI221_X1 port map( B1 => n13006, B2 => n6219, C1 => n13003, C2 => 
                           n15696, A => n5238, ZN => n5233);
   U4497 : OAI222_X1 port map( A1 => n14938, A2 => n13000, B1 => n14874, B2 => 
                           n12997, C1 => n14906, C2 => n12994, ZN => n5238);
   U4498 : AOI221_X1 port map( B1 => n12952, B2 => n5963, C1 => n12949, C2 => 
                           n15196, A => n5246, ZN => n5241);
   U4499 : OAI222_X1 port map( A1 => n15292, A2 => n12946, B1 => n15228, B2 => 
                           n12943, C1 => n15260, C2 => n12940, ZN => n5246);
   U4500 : AOI221_X1 port map( B1 => n13006, B2 => n6220, C1 => n13003, C2 => 
                           n15695, A => n5201, ZN => n5196);
   U4501 : OAI222_X1 port map( A1 => n14937, A2 => n13000, B1 => n14873, B2 => 
                           n12997, C1 => n14905, C2 => n12994, ZN => n5201);
   U4502 : AOI221_X1 port map( B1 => n12952, B2 => n5964, C1 => n12949, C2 => 
                           n15195, A => n5209, ZN => n5204);
   U4503 : OAI222_X1 port map( A1 => n15291, A2 => n12946, B1 => n15227, B2 => 
                           n12943, C1 => n15259, C2 => n12940, ZN => n5209);
   U4504 : AOI221_X1 port map( B1 => n13006, B2 => n6221, C1 => n13003, C2 => 
                           n15694, A => n5164, ZN => n5159);
   U4505 : OAI222_X1 port map( A1 => n14936, A2 => n13000, B1 => n14872, B2 => 
                           n12997, C1 => n14904, C2 => n12994, ZN => n5164);
   U4506 : AOI221_X1 port map( B1 => n12952, B2 => n5965, C1 => n12949, C2 => 
                           n15194, A => n5172, ZN => n5167);
   U4507 : OAI222_X1 port map( A1 => n15290, A2 => n12946, B1 => n15226, B2 => 
                           n12943, C1 => n15258, C2 => n12940, ZN => n5172);
   U4508 : AOI221_X1 port map( B1 => n13007, B2 => n6222, C1 => n13004, C2 => 
                           n15693, A => n5127, ZN => n5122);
   U4509 : OAI222_X1 port map( A1 => n14935, A2 => n13001, B1 => n14871, B2 => 
                           n12998, C1 => n14903, C2 => n12995, ZN => n5127);
   U4510 : AOI221_X1 port map( B1 => n12953, B2 => n5966, C1 => n12950, C2 => 
                           n15193, A => n5135, ZN => n5130);
   U4511 : OAI222_X1 port map( A1 => n15289, A2 => n12947, B1 => n15225, B2 => 
                           n12944, C1 => n15257, C2 => n12941, ZN => n5135);
   U4512 : AOI221_X1 port map( B1 => n13007, B2 => n6223, C1 => n13004, C2 => 
                           n15692, A => n5090, ZN => n5085);
   U4513 : OAI222_X1 port map( A1 => n14934, A2 => n13001, B1 => n14870, B2 => 
                           n12998, C1 => n14902, C2 => n12995, ZN => n5090);
   U4514 : AOI221_X1 port map( B1 => n12953, B2 => n5967, C1 => n12950, C2 => 
                           n15192, A => n5098, ZN => n5093);
   U4515 : OAI222_X1 port map( A1 => n15288, A2 => n12947, B1 => n15224, B2 => 
                           n12944, C1 => n15256, C2 => n12941, ZN => n5098);
   U4516 : AOI221_X1 port map( B1 => n13007, B2 => n6224, C1 => n13004, C2 => 
                           n15691, A => n5053, ZN => n5048);
   U4517 : OAI222_X1 port map( A1 => n14933, A2 => n13001, B1 => n14869, B2 => 
                           n12998, C1 => n14901, C2 => n12995, ZN => n5053);
   U4518 : AOI221_X1 port map( B1 => n12953, B2 => n5968, C1 => n12950, C2 => 
                           n15191, A => n5061, ZN => n5056);
   U4519 : OAI222_X1 port map( A1 => n15287, A2 => n12947, B1 => n15223, B2 => 
                           n12944, C1 => n15255, C2 => n12941, ZN => n5061);
   U4520 : AOI221_X1 port map( B1 => n13007, B2 => n6225, C1 => n13004, C2 => 
                           n15690, A => n5016, ZN => n5011);
   U4521 : OAI222_X1 port map( A1 => n14932, A2 => n13001, B1 => n14868, B2 => 
                           n12998, C1 => n14900, C2 => n12995, ZN => n5016);
   U4522 : AOI221_X1 port map( B1 => n12953, B2 => n5969, C1 => n12950, C2 => 
                           n15190, A => n5024, ZN => n5019);
   U4523 : OAI222_X1 port map( A1 => n15286, A2 => n12947, B1 => n15222, B2 => 
                           n12944, C1 => n15254, C2 => n12941, ZN => n5024);
   U4524 : AOI221_X1 port map( B1 => n13007, B2 => n6226, C1 => n13004, C2 => 
                           n15689, A => n4979, ZN => n4974);
   U4525 : OAI222_X1 port map( A1 => n14931, A2 => n13001, B1 => n14867, B2 => 
                           n12998, C1 => n14899, C2 => n12995, ZN => n4979);
   U4526 : AOI221_X1 port map( B1 => n12953, B2 => n5970, C1 => n12950, C2 => 
                           n15189, A => n4987, ZN => n4982);
   U4527 : OAI222_X1 port map( A1 => n15285, A2 => n12947, B1 => n15221, B2 => 
                           n12944, C1 => n15253, C2 => n12941, ZN => n4987);
   U4528 : AOI221_X1 port map( B1 => n13007, B2 => n6227, C1 => n13004, C2 => 
                           n15688, A => n4942, ZN => n4937);
   U4529 : OAI222_X1 port map( A1 => n14930, A2 => n13001, B1 => n14866, B2 => 
                           n12998, C1 => n14898, C2 => n12995, ZN => n4942);
   U4530 : AOI221_X1 port map( B1 => n12953, B2 => n5971, C1 => n12950, C2 => 
                           n15188, A => n4950, ZN => n4945);
   U4531 : OAI222_X1 port map( A1 => n15284, A2 => n12947, B1 => n15220, B2 => 
                           n12944, C1 => n15252, C2 => n12941, ZN => n4950);
   U4532 : AOI221_X1 port map( B1 => n13007, B2 => n6228, C1 => n13004, C2 => 
                           n15687, A => n4905, ZN => n4900);
   U4533 : OAI222_X1 port map( A1 => n14929, A2 => n13001, B1 => n14865, B2 => 
                           n12998, C1 => n14897, C2 => n12995, ZN => n4905);
   U4534 : AOI221_X1 port map( B1 => n12953, B2 => n5972, C1 => n12950, C2 => 
                           n15187, A => n4913, ZN => n4908);
   U4535 : OAI222_X1 port map( A1 => n15283, A2 => n12947, B1 => n15219, B2 => 
                           n12944, C1 => n15251, C2 => n12941, ZN => n4913);
   U4536 : AOI221_X1 port map( B1 => n13007, B2 => n6229, C1 => n13004, C2 => 
                           n15686, A => n4868, ZN => n4863);
   U4537 : OAI222_X1 port map( A1 => n14928, A2 => n13001, B1 => n14864, B2 => 
                           n12998, C1 => n14896, C2 => n12995, ZN => n4868);
   U4538 : AOI221_X1 port map( B1 => n12953, B2 => n5973, C1 => n12950, C2 => 
                           n15186, A => n4876, ZN => n4871);
   U4539 : OAI222_X1 port map( A1 => n15282, A2 => n12947, B1 => n15218, B2 => 
                           n12944, C1 => n15250, C2 => n12941, ZN => n4876);
   U4540 : AOI221_X1 port map( B1 => n13007, B2 => n6230, C1 => n13004, C2 => 
                           n15685, A => n4831, ZN => n4826);
   U4541 : OAI222_X1 port map( A1 => n14927, A2 => n13001, B1 => n14863, B2 => 
                           n12998, C1 => n14895, C2 => n12995, ZN => n4831);
   U4542 : AOI221_X1 port map( B1 => n12953, B2 => n5974, C1 => n12950, C2 => 
                           n15185, A => n4839, ZN => n4834);
   U4543 : OAI222_X1 port map( A1 => n15281, A2 => n12947, B1 => n15217, B2 => 
                           n12944, C1 => n15249, C2 => n12941, ZN => n4839);
   U4544 : AOI221_X1 port map( B1 => n13007, B2 => n6231, C1 => n13004, C2 => 
                           n15684, A => n4794, ZN => n4789);
   U4545 : OAI222_X1 port map( A1 => n14926, A2 => n13001, B1 => n14862, B2 => 
                           n12998, C1 => n14894, C2 => n12995, ZN => n4794);
   U4546 : AOI221_X1 port map( B1 => n12953, B2 => n5975, C1 => n12950, C2 => 
                           n15184, A => n4802, ZN => n4797);
   U4547 : OAI222_X1 port map( A1 => n15280, A2 => n12947, B1 => n15216, B2 => 
                           n12944, C1 => n15248, C2 => n12941, ZN => n4802);
   U4548 : AOI221_X1 port map( B1 => n13007, B2 => n6232, C1 => n13004, C2 => 
                           n15683, A => n4757, ZN => n4752);
   U4549 : OAI222_X1 port map( A1 => n14925, A2 => n13001, B1 => n14861, B2 => 
                           n12998, C1 => n14893, C2 => n12995, ZN => n4757);
   U4550 : AOI221_X1 port map( B1 => n12953, B2 => n5976, C1 => n12950, C2 => 
                           n15183, A => n4765, ZN => n4760);
   U4551 : OAI222_X1 port map( A1 => n15279, A2 => n12947, B1 => n15215, B2 => 
                           n12944, C1 => n15247, C2 => n12941, ZN => n4765);
   U4552 : AOI221_X1 port map( B1 => n13007, B2 => n6233, C1 => n13004, C2 => 
                           n15682, A => n4720, ZN => n4715);
   U4553 : OAI222_X1 port map( A1 => n14924, A2 => n13001, B1 => n14860, B2 => 
                           n12998, C1 => n14892, C2 => n12995, ZN => n4720);
   U4554 : AOI221_X1 port map( B1 => n12953, B2 => n5977, C1 => n12950, C2 => 
                           n15182, A => n4728, ZN => n4723);
   U4555 : OAI222_X1 port map( A1 => n15278, A2 => n12947, B1 => n15214, B2 => 
                           n12944, C1 => n15246, C2 => n12941, ZN => n4728);
   U4556 : AOI221_X1 port map( B1 => n12954, B2 => n5978, C1 => n12951, C2 => 
                           n15181, A => n4691, ZN => n4686);
   U4557 : OAI222_X1 port map( A1 => n15277, A2 => n12948, B1 => n15213, B2 => 
                           n12945, C1 => n15245, C2 => n12942, ZN => n4691);
   U4558 : AOI221_X1 port map( B1 => n13234, B2 => n6210, C1 => n13231, C2 => 
                           n15705, A => n4302, ZN => n4295);
   U4559 : OAI222_X1 port map( A1 => n14947, A2 => n13228, B1 => n14883, B2 => 
                           n13225, C1 => n14915, C2 => n13222, ZN => n4302);
   U4560 : AOI221_X1 port map( B1 => n13180, B2 => n5954, C1 => n13177, C2 => 
                           n15205, A => n4311, ZN => n4305);
   U4561 : OAI222_X1 port map( A1 => n15301, A2 => n13174, B1 => n15237, B2 => 
                           n13171, C1 => n15269, C2 => n13168, ZN => n4311);
   U4562 : AOI221_X1 port map( B1 => n13234, B2 => n6211, C1 => n13231, C2 => 
                           n15704, A => n4250, ZN => n4245);
   U4563 : OAI222_X1 port map( A1 => n14946, A2 => n13228, B1 => n14882, B2 => 
                           n13225, C1 => n14914, C2 => n13222, ZN => n4250);
   U4564 : AOI221_X1 port map( B1 => n13180, B2 => n5955, C1 => n13177, C2 => 
                           n15204, A => n4258, ZN => n4253);
   U4565 : OAI222_X1 port map( A1 => n15300, A2 => n13174, B1 => n15236, B2 => 
                           n13171, C1 => n15268, C2 => n13168, ZN => n4258);
   U4566 : AOI221_X1 port map( B1 => n13234, B2 => n6212, C1 => n13231, C2 => 
                           n15703, A => n4213, ZN => n4208);
   U4567 : OAI222_X1 port map( A1 => n14945, A2 => n13228, B1 => n14881, B2 => 
                           n13225, C1 => n14913, C2 => n13222, ZN => n4213);
   U4568 : AOI221_X1 port map( B1 => n13180, B2 => n5956, C1 => n13177, C2 => 
                           n15203, A => n4221, ZN => n4216);
   U4569 : OAI222_X1 port map( A1 => n15299, A2 => n13174, B1 => n15235, B2 => 
                           n13171, C1 => n15267, C2 => n13168, ZN => n4221);
   U4570 : AOI221_X1 port map( B1 => n13234, B2 => n6213, C1 => n13231, C2 => 
                           n15702, A => n4176, ZN => n4171);
   U4571 : OAI222_X1 port map( A1 => n14944, A2 => n13228, B1 => n14880, B2 => 
                           n13225, C1 => n14912, C2 => n13222, ZN => n4176);
   U4572 : AOI221_X1 port map( B1 => n13180, B2 => n5957, C1 => n13177, C2 => 
                           n15202, A => n4184, ZN => n4179);
   U4573 : OAI222_X1 port map( A1 => n15298, A2 => n13174, B1 => n15234, B2 => 
                           n13171, C1 => n15266, C2 => n13168, ZN => n4184);
   U4574 : AOI221_X1 port map( B1 => n13234, B2 => n6214, C1 => n13231, C2 => 
                           n15701, A => n4139, ZN => n4134);
   U4575 : OAI222_X1 port map( A1 => n14943, A2 => n13228, B1 => n14879, B2 => 
                           n13225, C1 => n14911, C2 => n13222, ZN => n4139);
   U4576 : AOI221_X1 port map( B1 => n13180, B2 => n5958, C1 => n13177, C2 => 
                           n15201, A => n4147, ZN => n4142);
   U4577 : OAI222_X1 port map( A1 => n15297, A2 => n13174, B1 => n15233, B2 => 
                           n13171, C1 => n15265, C2 => n13168, ZN => n4147);
   U4578 : AOI221_X1 port map( B1 => n13234, B2 => n6215, C1 => n13231, C2 => 
                           n15700, A => n4102, ZN => n4097);
   U4579 : OAI222_X1 port map( A1 => n14942, A2 => n13228, B1 => n14878, B2 => 
                           n13225, C1 => n14910, C2 => n13222, ZN => n4102);
   U4580 : AOI221_X1 port map( B1 => n13180, B2 => n5959, C1 => n13177, C2 => 
                           n15200, A => n4110, ZN => n4105);
   U4581 : OAI222_X1 port map( A1 => n15296, A2 => n13174, B1 => n15232, B2 => 
                           n13171, C1 => n15264, C2 => n13168, ZN => n4110);
   U4582 : AOI221_X1 port map( B1 => n13234, B2 => n6216, C1 => n13231, C2 => 
                           n15699, A => n4065, ZN => n4060);
   U4583 : OAI222_X1 port map( A1 => n14941, A2 => n13228, B1 => n14877, B2 => 
                           n13225, C1 => n14909, C2 => n13222, ZN => n4065);
   U4584 : AOI221_X1 port map( B1 => n13180, B2 => n5960, C1 => n13177, C2 => 
                           n15199, A => n4073, ZN => n4068);
   U4585 : OAI222_X1 port map( A1 => n15295, A2 => n13174, B1 => n15231, B2 => 
                           n13171, C1 => n15263, C2 => n13168, ZN => n4073);
   U4586 : AOI221_X1 port map( B1 => n13234, B2 => n6217, C1 => n13231, C2 => 
                           n15698, A => n4028, ZN => n4023);
   U4587 : OAI222_X1 port map( A1 => n14940, A2 => n13228, B1 => n14876, B2 => 
                           n13225, C1 => n14908, C2 => n13222, ZN => n4028);
   U4588 : AOI221_X1 port map( B1 => n13180, B2 => n5961, C1 => n13177, C2 => 
                           n15198, A => n4036, ZN => n4031);
   U4589 : OAI222_X1 port map( A1 => n15294, A2 => n13174, B1 => n15230, B2 => 
                           n13171, C1 => n15262, C2 => n13168, ZN => n4036);
   U4590 : AOI221_X1 port map( B1 => n13234, B2 => n6218, C1 => n13231, C2 => 
                           n15697, A => n3991, ZN => n3986);
   U4591 : OAI222_X1 port map( A1 => n14939, A2 => n13228, B1 => n14875, B2 => 
                           n13225, C1 => n14907, C2 => n13222, ZN => n3991);
   U4592 : AOI221_X1 port map( B1 => n13180, B2 => n5962, C1 => n13177, C2 => 
                           n15197, A => n3999, ZN => n3994);
   U4593 : OAI222_X1 port map( A1 => n15293, A2 => n13174, B1 => n15229, B2 => 
                           n13171, C1 => n15261, C2 => n13168, ZN => n3999);
   U4594 : AOI221_X1 port map( B1 => n13234, B2 => n6219, C1 => n13231, C2 => 
                           n15696, A => n3954, ZN => n3949);
   U4595 : OAI222_X1 port map( A1 => n14938, A2 => n13228, B1 => n14874, B2 => 
                           n13225, C1 => n14906, C2 => n13222, ZN => n3954);
   U4596 : AOI221_X1 port map( B1 => n13180, B2 => n5963, C1 => n13177, C2 => 
                           n15196, A => n3962, ZN => n3957);
   U4597 : OAI222_X1 port map( A1 => n15292, A2 => n13174, B1 => n15228, B2 => 
                           n13171, C1 => n15260, C2 => n13168, ZN => n3962);
   U4598 : AOI221_X1 port map( B1 => n13234, B2 => n6220, C1 => n13231, C2 => 
                           n15695, A => n3917, ZN => n3912);
   U4599 : OAI222_X1 port map( A1 => n14937, A2 => n13228, B1 => n14873, B2 => 
                           n13225, C1 => n14905, C2 => n13222, ZN => n3917);
   U4600 : AOI221_X1 port map( B1 => n13180, B2 => n5964, C1 => n13177, C2 => 
                           n15195, A => n3925, ZN => n3920);
   U4601 : OAI222_X1 port map( A1 => n15291, A2 => n13174, B1 => n15227, B2 => 
                           n13171, C1 => n15259, C2 => n13168, ZN => n3925);
   U4602 : AOI221_X1 port map( B1 => n13234, B2 => n6221, C1 => n13231, C2 => 
                           n15694, A => n3880, ZN => n3875);
   U4603 : OAI222_X1 port map( A1 => n14936, A2 => n13228, B1 => n14872, B2 => 
                           n13225, C1 => n14904, C2 => n13222, ZN => n3880);
   U4604 : AOI221_X1 port map( B1 => n13180, B2 => n5965, C1 => n13177, C2 => 
                           n15194, A => n3888, ZN => n3883);
   U4605 : OAI222_X1 port map( A1 => n15290, A2 => n13174, B1 => n15226, B2 => 
                           n13171, C1 => n15258, C2 => n13168, ZN => n3888);
   U4606 : AOI221_X1 port map( B1 => n13235, B2 => n6222, C1 => n13232, C2 => 
                           n15693, A => n3843, ZN => n3838);
   U4607 : OAI222_X1 port map( A1 => n14935, A2 => n13229, B1 => n14871, B2 => 
                           n13226, C1 => n14903, C2 => n13223, ZN => n3843);
   U4608 : AOI221_X1 port map( B1 => n13181, B2 => n5966, C1 => n13178, C2 => 
                           n15193, A => n3851, ZN => n3846);
   U4609 : OAI222_X1 port map( A1 => n15289, A2 => n13175, B1 => n15225, B2 => 
                           n13172, C1 => n15257, C2 => n13169, ZN => n3851);
   U4610 : AOI221_X1 port map( B1 => n13235, B2 => n6223, C1 => n13232, C2 => 
                           n15692, A => n3806, ZN => n3801);
   U4611 : OAI222_X1 port map( A1 => n14934, A2 => n13229, B1 => n14870, B2 => 
                           n13226, C1 => n14902, C2 => n13223, ZN => n3806);
   U4612 : AOI221_X1 port map( B1 => n13181, B2 => n5967, C1 => n13178, C2 => 
                           n15192, A => n3814, ZN => n3809);
   U4613 : OAI222_X1 port map( A1 => n15288, A2 => n13175, B1 => n15224, B2 => 
                           n13172, C1 => n15256, C2 => n13169, ZN => n3814);
   U4614 : AOI221_X1 port map( B1 => n13235, B2 => n6224, C1 => n13232, C2 => 
                           n15691, A => n3769, ZN => n3764);
   U4615 : OAI222_X1 port map( A1 => n14933, A2 => n13229, B1 => n14869, B2 => 
                           n13226, C1 => n14901, C2 => n13223, ZN => n3769);
   U4616 : AOI221_X1 port map( B1 => n13181, B2 => n5968, C1 => n13178, C2 => 
                           n15191, A => n3777, ZN => n3772);
   U4617 : OAI222_X1 port map( A1 => n15287, A2 => n13175, B1 => n15223, B2 => 
                           n13172, C1 => n15255, C2 => n13169, ZN => n3777);
   U4618 : AOI221_X1 port map( B1 => n13235, B2 => n6225, C1 => n13232, C2 => 
                           n15690, A => n3732, ZN => n3727);
   U4619 : OAI222_X1 port map( A1 => n14932, A2 => n13229, B1 => n14868, B2 => 
                           n13226, C1 => n14900, C2 => n13223, ZN => n3732);
   U4620 : AOI221_X1 port map( B1 => n13181, B2 => n5969, C1 => n13178, C2 => 
                           n15190, A => n3740, ZN => n3735);
   U4621 : OAI222_X1 port map( A1 => n15286, A2 => n13175, B1 => n15222, B2 => 
                           n13172, C1 => n15254, C2 => n13169, ZN => n3740);
   U4622 : AOI221_X1 port map( B1 => n13235, B2 => n6226, C1 => n13232, C2 => 
                           n15689, A => n3695, ZN => n3690);
   U4623 : OAI222_X1 port map( A1 => n14931, A2 => n13229, B1 => n14867, B2 => 
                           n13226, C1 => n14899, C2 => n13223, ZN => n3695);
   U4624 : AOI221_X1 port map( B1 => n13181, B2 => n5970, C1 => n13178, C2 => 
                           n15189, A => n3703, ZN => n3698);
   U4625 : OAI222_X1 port map( A1 => n15285, A2 => n13175, B1 => n15221, B2 => 
                           n13172, C1 => n15253, C2 => n13169, ZN => n3703);
   U4626 : AOI221_X1 port map( B1 => n13235, B2 => n6227, C1 => n13232, C2 => 
                           n15688, A => n3658, ZN => n3653);
   U4627 : OAI222_X1 port map( A1 => n14930, A2 => n13229, B1 => n14866, B2 => 
                           n13226, C1 => n14898, C2 => n13223, ZN => n3658);
   U4628 : AOI221_X1 port map( B1 => n13181, B2 => n5971, C1 => n13178, C2 => 
                           n15188, A => n3666, ZN => n3661);
   U4629 : OAI222_X1 port map( A1 => n15284, A2 => n13175, B1 => n15220, B2 => 
                           n13172, C1 => n15252, C2 => n13169, ZN => n3666);
   U4630 : AOI221_X1 port map( B1 => n13235, B2 => n6228, C1 => n13232, C2 => 
                           n15687, A => n3621, ZN => n3616);
   U4631 : OAI222_X1 port map( A1 => n14929, A2 => n13229, B1 => n14865, B2 => 
                           n13226, C1 => n14897, C2 => n13223, ZN => n3621);
   U4632 : AOI221_X1 port map( B1 => n13181, B2 => n5972, C1 => n13178, C2 => 
                           n15187, A => n3629, ZN => n3624);
   U4633 : OAI222_X1 port map( A1 => n15283, A2 => n13175, B1 => n15219, B2 => 
                           n13172, C1 => n15251, C2 => n13169, ZN => n3629);
   U4634 : AOI221_X1 port map( B1 => n13235, B2 => n6229, C1 => n13232, C2 => 
                           n15686, A => n3584, ZN => n3579);
   U4635 : OAI222_X1 port map( A1 => n14928, A2 => n13229, B1 => n14864, B2 => 
                           n13226, C1 => n14896, C2 => n13223, ZN => n3584);
   U4636 : AOI221_X1 port map( B1 => n13181, B2 => n5973, C1 => n13178, C2 => 
                           n15186, A => n3592, ZN => n3587);
   U4637 : OAI222_X1 port map( A1 => n15282, A2 => n13175, B1 => n15218, B2 => 
                           n13172, C1 => n15250, C2 => n13169, ZN => n3592);
   U4638 : AOI221_X1 port map( B1 => n13235, B2 => n6230, C1 => n13232, C2 => 
                           n15685, A => n3547, ZN => n3542);
   U4639 : OAI222_X1 port map( A1 => n14927, A2 => n13229, B1 => n14863, B2 => 
                           n13226, C1 => n14895, C2 => n13223, ZN => n3547);
   U4640 : AOI221_X1 port map( B1 => n13181, B2 => n5974, C1 => n13178, C2 => 
                           n15185, A => n3555, ZN => n3550);
   U4641 : OAI222_X1 port map( A1 => n15281, A2 => n13175, B1 => n15217, B2 => 
                           n13172, C1 => n15249, C2 => n13169, ZN => n3555);
   U4642 : AOI221_X1 port map( B1 => n13235, B2 => n6231, C1 => n13232, C2 => 
                           n15684, A => n3510, ZN => n3505);
   U4643 : OAI222_X1 port map( A1 => n14926, A2 => n13229, B1 => n14862, B2 => 
                           n13226, C1 => n14894, C2 => n13223, ZN => n3510);
   U4644 : AOI221_X1 port map( B1 => n13181, B2 => n5975, C1 => n13178, C2 => 
                           n15184, A => n3518, ZN => n3513);
   U4645 : OAI222_X1 port map( A1 => n15280, A2 => n13175, B1 => n15216, B2 => 
                           n13172, C1 => n15248, C2 => n13169, ZN => n3518);
   U4646 : AOI221_X1 port map( B1 => n13235, B2 => n6232, C1 => n13232, C2 => 
                           n15683, A => n3473, ZN => n3468);
   U4647 : OAI222_X1 port map( A1 => n14925, A2 => n13229, B1 => n14861, B2 => 
                           n13226, C1 => n14893, C2 => n13223, ZN => n3473);
   U4648 : AOI221_X1 port map( B1 => n13181, B2 => n5976, C1 => n13178, C2 => 
                           n15183, A => n3481, ZN => n3476);
   U4649 : OAI222_X1 port map( A1 => n15279, A2 => n13175, B1 => n15215, B2 => 
                           n13172, C1 => n15247, C2 => n13169, ZN => n3481);
   U4650 : AOI221_X1 port map( B1 => n13235, B2 => n6233, C1 => n13232, C2 => 
                           n15682, A => n3436, ZN => n3431);
   U4651 : OAI222_X1 port map( A1 => n14924, A2 => n13229, B1 => n14860, B2 => 
                           n13226, C1 => n14892, C2 => n13223, ZN => n3436);
   U4652 : AOI221_X1 port map( B1 => n13181, B2 => n5977, C1 => n13178, C2 => 
                           n15182, A => n3444, ZN => n3439);
   U4653 : OAI222_X1 port map( A1 => n15278, A2 => n13175, B1 => n15214, B2 => 
                           n13172, C1 => n15246, C2 => n13169, ZN => n3444);
   U4654 : AOI221_X1 port map( B1 => n13182, B2 => n5978, C1 => n13179, C2 => 
                           n15181, A => n3407, ZN => n3402);
   U4655 : OAI222_X1 port map( A1 => n15277, A2 => n13176, B1 => n15213, B2 => 
                           n13173, C1 => n15245, C2 => n13170, ZN => n3407);
   U4656 : AOI221_X1 port map( B1 => n13236, B2 => n6235, C1 => n13233, C2 => 
                           n15564, A => n3362, ZN => n3357);
   U4657 : OAI222_X1 port map( A1 => n14922, A2 => n13230, B1 => n14858, B2 => 
                           n13227, C1 => n14890, C2 => n13224, ZN => n3362);
   U4658 : AOI221_X1 port map( B1 => n13236, B2 => n6236, C1 => n13233, C2 => 
                           n15563, A => n3325, ZN => n3320);
   U4659 : OAI222_X1 port map( A1 => n14921, A2 => n13230, B1 => n14857, B2 => 
                           n13227, C1 => n14889, C2 => n13224, ZN => n3325);
   U4660 : AOI221_X1 port map( B1 => n13236, B2 => n6237, C1 => n13233, C2 => 
                           n15562, A => n3288, ZN => n3283);
   U4661 : OAI222_X1 port map( A1 => n14920, A2 => n13230, B1 => n14856, B2 => 
                           n13227, C1 => n14888, C2 => n13224, ZN => n3288);
   U4662 : AOI221_X1 port map( B1 => n13167, B2 => n6046, C1 => n13164, C2 => 
                           n6078, A => n3260, ZN => n3253);
   U4663 : OAI22_X1 port map( A1 => n15113, A2 => n13161, B1 => n15145, B2 => 
                           n13158, ZN => n3260);
   U4664 : AOI221_X1 port map( B1 => n13167, B2 => n6047, C1 => n13164, C2 => 
                           n6079, A => n3223, ZN => n3216);
   U4665 : OAI22_X1 port map( A1 => n15112, A2 => n13161, B1 => n15144, B2 => 
                           n13158, ZN => n3223);
   U4666 : AOI221_X1 port map( B1 => n13167, B2 => n6048, C1 => n13164, C2 => 
                           n6080, A => n3186, ZN => n3179);
   U4667 : OAI22_X1 port map( A1 => n15111, A2 => n13161, B1 => n15143, B2 => 
                           n13158, ZN => n3186);
   U4668 : AOI221_X1 port map( B1 => n13167, B2 => n6049, C1 => n13164, C2 => 
                           n6081, A => n3147, ZN => n3124);
   U4669 : OAI22_X1 port map( A1 => n15110, A2 => n13161, B1 => n15142, B2 => 
                           n13158, ZN => n3147);
   U4670 : AOI221_X1 port map( B1 => n12939, B2 => n6075, C1 => n12936, C2 => 
                           n6043, A => n4655, ZN => n4648);
   U4671 : OAI22_X1 port map( A1 => n15148, A2 => n12933, B1 => n15116, B2 => 
                           n12930, ZN => n4655);
   U4672 : AOI221_X1 port map( B1 => n12939, B2 => n6076, C1 => n12936, C2 => 
                           n6044, A => n4618, ZN => n4611);
   U4673 : OAI22_X1 port map( A1 => n15147, A2 => n12933, B1 => n15115, B2 => 
                           n12930, ZN => n4618);
   U4674 : AOI221_X1 port map( B1 => n12939, B2 => n6077, C1 => n12936, C2 => 
                           n6045, A => n4581, ZN => n4574);
   U4675 : OAI22_X1 port map( A1 => n15146, A2 => n12933, B1 => n15114, B2 => 
                           n12930, ZN => n4581);
   U4676 : AOI221_X1 port map( B1 => n12939, B2 => n6078, C1 => n12936, C2 => 
                           n6046, A => n4544, ZN => n4537);
   U4677 : OAI22_X1 port map( A1 => n15145, A2 => n12933, B1 => n15113, B2 => 
                           n12930, ZN => n4544);
   U4678 : AOI221_X1 port map( B1 => n12939, B2 => n6079, C1 => n12936, C2 => 
                           n6047, A => n4507, ZN => n4500);
   U4679 : OAI22_X1 port map( A1 => n15144, A2 => n12933, B1 => n15112, B2 => 
                           n12930, ZN => n4507);
   U4680 : AOI221_X1 port map( B1 => n12939, B2 => n6080, C1 => n12936, C2 => 
                           n6048, A => n4470, ZN => n4463);
   U4681 : OAI22_X1 port map( A1 => n15143, A2 => n12933, B1 => n15111, B2 => 
                           n12930, ZN => n4470);
   U4682 : AOI221_X1 port map( B1 => n12939, B2 => n6081, C1 => n12936, C2 => 
                           n6049, A => n4431, ZN => n4408);
   U4683 : OAI22_X1 port map( A1 => n15142, A2 => n12933, B1 => n15110, B2 => 
                           n12930, ZN => n4431);
   U4684 : AOI221_X1 port map( B1 => n12992, B2 => n592, C1 => n12989, C2 => 
                           n15717, A => n5128, ZN => n5121);
   U4685 : OAI22_X1 port map( A1 => n14839, A2 => n12986, B1 => n14807, B2 => 
                           n12983, ZN => n5128);
   U4686 : AOI221_X1 port map( B1 => n12992, B2 => n590, C1 => n12989, C2 => 
                           n15716, A => n5091, ZN => n5084);
   U4687 : OAI22_X1 port map( A1 => n14838, A2 => n12986, B1 => n14806, B2 => 
                           n12983, ZN => n5091);
   U4688 : AOI221_X1 port map( B1 => n12992, B2 => n588, C1 => n12989, C2 => 
                           n15715, A => n5054, ZN => n5047);
   U4689 : OAI22_X1 port map( A1 => n14837, A2 => n12986, B1 => n14805, B2 => 
                           n12983, ZN => n5054);
   U4690 : AOI221_X1 port map( B1 => n12992, B2 => n586, C1 => n12989, C2 => 
                           n15714, A => n5017, ZN => n5010);
   U4691 : OAI22_X1 port map( A1 => n14836, A2 => n12986, B1 => n14804, B2 => 
                           n12983, ZN => n5017);
   U4692 : AOI221_X1 port map( B1 => n12992, B2 => n584, C1 => n12989, C2 => 
                           n15713, A => n4980, ZN => n4973);
   U4693 : OAI22_X1 port map( A1 => n14835, A2 => n12986, B1 => n14803, B2 => 
                           n12983, ZN => n4980);
   U4694 : AOI221_X1 port map( B1 => n12992, B2 => n582, C1 => n12989, C2 => 
                           n15712, A => n4943, ZN => n4936);
   U4695 : OAI22_X1 port map( A1 => n14834, A2 => n12986, B1 => n14802, B2 => 
                           n12983, ZN => n4943);
   U4696 : AOI221_X1 port map( B1 => n12992, B2 => n580, C1 => n12989, C2 => 
                           n15711, A => n4906, ZN => n4899);
   U4697 : OAI22_X1 port map( A1 => n14833, A2 => n12986, B1 => n14801, B2 => 
                           n12983, ZN => n4906);
   U4698 : AOI221_X1 port map( B1 => n12992, B2 => n578, C1 => n12989, C2 => 
                           n15710, A => n4869, ZN => n4862);
   U4699 : OAI22_X1 port map( A1 => n14832, A2 => n12986, B1 => n14800, B2 => 
                           n12983, ZN => n4869);
   U4700 : AOI221_X1 port map( B1 => n12939, B2 => n6074, C1 => n12936, C2 => 
                           n6042, A => n4692, ZN => n4685);
   U4701 : OAI22_X1 port map( A1 => n15149, A2 => n12933, B1 => n15117, B2 => 
                           n12930, ZN => n4692);
   U4702 : AOI221_X1 port map( B1 => n13220, B2 => n592, C1 => n13217, C2 => 
                           n15717, A => n3844, ZN => n3837);
   U4703 : OAI22_X1 port map( A1 => n14839, A2 => n13214, B1 => n14807, B2 => 
                           n13211, ZN => n3844);
   U4704 : AOI221_X1 port map( B1 => n13166, B2 => n6030, C1 => n13163, C2 => 
                           n6062, A => n3852, ZN => n3845);
   U4705 : OAI22_X1 port map( A1 => n15129, A2 => n13160, B1 => n15161, B2 => 
                           n13157, ZN => n3852);
   U4706 : AOI221_X1 port map( B1 => n13220, B2 => n590, C1 => n13217, C2 => 
                           n15716, A => n3807, ZN => n3800);
   U4707 : OAI22_X1 port map( A1 => n14838, A2 => n13214, B1 => n14806, B2 => 
                           n13211, ZN => n3807);
   U4708 : AOI221_X1 port map( B1 => n13166, B2 => n6031, C1 => n13163, C2 => 
                           n6063, A => n3815, ZN => n3808);
   U4709 : OAI22_X1 port map( A1 => n15128, A2 => n13160, B1 => n15160, B2 => 
                           n13157, ZN => n3815);
   U4710 : AOI221_X1 port map( B1 => n13220, B2 => n588, C1 => n13217, C2 => 
                           n15715, A => n3770, ZN => n3763);
   U4711 : OAI22_X1 port map( A1 => n14837, A2 => n13214, B1 => n14805, B2 => 
                           n13211, ZN => n3770);
   U4712 : AOI221_X1 port map( B1 => n13166, B2 => n6032, C1 => n13163, C2 => 
                           n6064, A => n3778, ZN => n3771);
   U4713 : OAI22_X1 port map( A1 => n15127, A2 => n13160, B1 => n15159, B2 => 
                           n13157, ZN => n3778);
   U4714 : AOI221_X1 port map( B1 => n13220, B2 => n586, C1 => n13217, C2 => 
                           n15714, A => n3733, ZN => n3726);
   U4715 : OAI22_X1 port map( A1 => n14836, A2 => n13214, B1 => n14804, B2 => 
                           n13211, ZN => n3733);
   U4716 : AOI221_X1 port map( B1 => n13166, B2 => n6033, C1 => n13163, C2 => 
                           n6065, A => n3741, ZN => n3734);
   U4717 : OAI22_X1 port map( A1 => n15126, A2 => n13160, B1 => n15158, B2 => 
                           n13157, ZN => n3741);
   U4718 : AOI221_X1 port map( B1 => n13220, B2 => n584, C1 => n13217, C2 => 
                           n15713, A => n3696, ZN => n3689);
   U4719 : OAI22_X1 port map( A1 => n14835, A2 => n13214, B1 => n14803, B2 => 
                           n13211, ZN => n3696);
   U4720 : AOI221_X1 port map( B1 => n13166, B2 => n6034, C1 => n13163, C2 => 
                           n6066, A => n3704, ZN => n3697);
   U4721 : OAI22_X1 port map( A1 => n15125, A2 => n13160, B1 => n15157, B2 => 
                           n13157, ZN => n3704);
   U4722 : AOI221_X1 port map( B1 => n13220, B2 => n582, C1 => n13217, C2 => 
                           n15712, A => n3659, ZN => n3652);
   U4723 : OAI22_X1 port map( A1 => n14834, A2 => n13214, B1 => n14802, B2 => 
                           n13211, ZN => n3659);
   U4724 : AOI221_X1 port map( B1 => n13166, B2 => n6035, C1 => n13163, C2 => 
                           n6067, A => n3667, ZN => n3660);
   U4725 : OAI22_X1 port map( A1 => n15124, A2 => n13160, B1 => n15156, B2 => 
                           n13157, ZN => n3667);
   U4726 : AOI221_X1 port map( B1 => n13220, B2 => n580, C1 => n13217, C2 => 
                           n15711, A => n3622, ZN => n3615);
   U4727 : OAI22_X1 port map( A1 => n14833, A2 => n13214, B1 => n14801, B2 => 
                           n13211, ZN => n3622);
   U4728 : AOI221_X1 port map( B1 => n13166, B2 => n6036, C1 => n13163, C2 => 
                           n6068, A => n3630, ZN => n3623);
   U4729 : OAI22_X1 port map( A1 => n15123, A2 => n13160, B1 => n15155, B2 => 
                           n13157, ZN => n3630);
   U4730 : AOI221_X1 port map( B1 => n13220, B2 => n578, C1 => n13217, C2 => 
                           n15710, A => n3585, ZN => n3578);
   U4731 : OAI22_X1 port map( A1 => n14832, A2 => n13214, B1 => n14800, B2 => 
                           n13211, ZN => n3585);
   U4732 : AOI221_X1 port map( B1 => n13166, B2 => n6037, C1 => n13163, C2 => 
                           n6069, A => n3593, ZN => n3586);
   U4733 : OAI22_X1 port map( A1 => n15122, A2 => n13160, B1 => n15154, B2 => 
                           n13157, ZN => n3593);
   U4734 : AOI221_X1 port map( B1 => n13166, B2 => n6038, C1 => n13163, C2 => 
                           n6070, A => n3556, ZN => n3549);
   U4735 : OAI22_X1 port map( A1 => n15121, A2 => n13160, B1 => n15153, B2 => 
                           n13157, ZN => n3556);
   U4736 : AOI221_X1 port map( B1 => n13166, B2 => n6039, C1 => n13163, C2 => 
                           n6071, A => n3519, ZN => n3512);
   U4737 : OAI22_X1 port map( A1 => n15120, A2 => n13160, B1 => n15152, B2 => 
                           n13157, ZN => n3519);
   U4738 : AOI221_X1 port map( B1 => n13166, B2 => n6040, C1 => n13163, C2 => 
                           n6072, A => n3482, ZN => n3475);
   U4739 : OAI22_X1 port map( A1 => n15119, A2 => n13160, B1 => n15151, B2 => 
                           n13157, ZN => n3482);
   U4740 : AOI221_X1 port map( B1 => n13166, B2 => n6041, C1 => n13163, C2 => 
                           n6073, A => n3445, ZN => n3438);
   U4741 : OAI22_X1 port map( A1 => n15118, A2 => n13160, B1 => n15150, B2 => 
                           n13157, ZN => n3445);
   U4742 : AOI221_X1 port map( B1 => n13167, B2 => n6043, C1 => n13164, C2 => 
                           n6075, A => n3371, ZN => n3364);
   U4743 : OAI22_X1 port map( A1 => n15116, A2 => n13161, B1 => n15148, B2 => 
                           n13158, ZN => n3371);
   U4744 : AOI221_X1 port map( B1 => n13167, B2 => n6044, C1 => n13164, C2 => 
                           n6076, A => n3334, ZN => n3327);
   U4745 : OAI22_X1 port map( A1 => n15115, A2 => n13161, B1 => n15147, B2 => 
                           n13158, ZN => n3334);
   U4746 : AOI221_X1 port map( B1 => n13167, B2 => n6045, C1 => n13164, C2 => 
                           n6077, A => n3297, ZN => n3290);
   U4747 : OAI22_X1 port map( A1 => n15114, A2 => n13161, B1 => n15146, B2 => 
                           n13158, ZN => n3297);
   U4748 : AOI221_X1 port map( B1 => n13221, B2 => n15730, C1 => n13218, C2 => 
                           n98, A => n3121, ZN => n3098);
   U4749 : OAI22_X1 port map( A1 => n14820, A2 => n13215, B1 => n14788, B2 => 
                           n13212, ZN => n3121);
   U4750 : AOI221_X1 port map( B1 => n12993, B2 => n15730, C1 => n12990, C2 => 
                           n98, A => n4405, ZN => n4382);
   U4751 : OAI22_X1 port map( A1 => n14820, A2 => n12987, B1 => n14788, B2 => 
                           n12984, ZN => n4405);
   U4752 : OAI22_X1 port map( A1 => n12645, A2 => n13323, B1 => n5667, B2 => 
                           n13320, ZN => n3236);
   U4753 : OAI22_X1 port map( A1 => n12646, A2 => n13323, B1 => n5677, B2 => 
                           n13320, ZN => n3199);
   U4754 : OAI22_X1 port map( A1 => n12647, A2 => n13323, B1 => n5687, B2 => 
                           n13320, ZN => n3162);
   U4755 : OAI22_X1 port map( A1 => n12648, A2 => n13323, B1 => n5697, B2 => 
                           n13320, ZN => n3069);
   U4756 : OAI22_X1 port map( A1 => n6803, A2 => n13095, B1 => n6931, B2 => 
                           n13092, ZN => n4631);
   U4757 : OAI22_X1 port map( A1 => n6804, A2 => n13095, B1 => n6932, B2 => 
                           n13092, ZN => n4594);
   U4758 : OAI22_X1 port map( A1 => n6805, A2 => n13095, B1 => n6933, B2 => 
                           n13092, ZN => n4557);
   U4759 : OAI22_X1 port map( A1 => n6806, A2 => n13095, B1 => n6934, B2 => 
                           n13092, ZN => n4520);
   U4760 : OAI22_X1 port map( A1 => n6807, A2 => n13095, B1 => n6935, B2 => 
                           n13092, ZN => n4483);
   U4761 : OAI22_X1 port map( A1 => n6808, A2 => n13095, B1 => n6936, B2 => 
                           n13092, ZN => n4446);
   U4762 : OAI22_X1 port map( A1 => n6809, A2 => n13095, B1 => n6937, B2 => 
                           n13092, ZN => n4353);
   U4763 : OAI22_X1 port map( A1 => n6802, A2 => n13095, B1 => n6930, B2 => 
                           n13092, ZN => n4668);
   U4764 : OAI22_X1 port map( A1 => n12649, A2 => n13323, B1 => n5627, B2 => 
                           n13320, ZN => n3384);
   U4765 : OAI22_X1 port map( A1 => n12650, A2 => n13323, B1 => n5637, B2 => 
                           n13320, ZN => n3347);
   U4766 : OAI22_X1 port map( A1 => n12651, A2 => n13323, B1 => n5647, B2 => 
                           n13320, ZN => n3310);
   U4767 : OAI22_X1 port map( A1 => n12652, A2 => n13323, B1 => n5657, B2 => 
                           n13320, ZN => n3273);
   U4768 : OAI22_X1 port map( A1 => n12653, A2 => n13350, B1 => n5665, B2 => 
                           n13347, ZN => n3234);
   U4769 : OAI22_X1 port map( A1 => n12654, A2 => n13350, B1 => n5675, B2 => 
                           n13347, ZN => n3197);
   U4770 : OAI22_X1 port map( A1 => n12655, A2 => n13350, B1 => n5685, B2 => 
                           n13347, ZN => n3160);
   U4771 : OAI22_X1 port map( A1 => n12656, A2 => n13350, B1 => n5695, B2 => 
                           n13347, ZN => n3058);
   U4772 : OAI22_X1 port map( A1 => n6787, A2 => n13122, B1 => n6915, B2 => 
                           n13119, ZN => n4629);
   U4773 : OAI22_X1 port map( A1 => n6788, A2 => n13122, B1 => n6916, B2 => 
                           n13119, ZN => n4592);
   U4774 : OAI22_X1 port map( A1 => n6789, A2 => n13122, B1 => n6917, B2 => 
                           n13119, ZN => n4555);
   U4775 : OAI22_X1 port map( A1 => n6790, A2 => n13122, B1 => n6918, B2 => 
                           n13119, ZN => n4518);
   U4776 : OAI22_X1 port map( A1 => n6791, A2 => n13122, B1 => n6919, B2 => 
                           n13119, ZN => n4481);
   U4777 : OAI22_X1 port map( A1 => n6792, A2 => n13122, B1 => n6920, B2 => 
                           n13119, ZN => n4444);
   U4778 : OAI22_X1 port map( A1 => n6793, A2 => n13122, B1 => n6921, B2 => 
                           n13119, ZN => n4342);
   U4779 : OAI22_X1 port map( A1 => n6786, A2 => n13122, B1 => n6914, B2 => 
                           n13119, ZN => n4666);
   U4780 : OAI22_X1 port map( A1 => n12657, A2 => n13350, B1 => n5625, B2 => 
                           n13347, ZN => n3382);
   U4781 : OAI22_X1 port map( A1 => n12658, A2 => n13350, B1 => n5635, B2 => 
                           n13347, ZN => n3345);
   U4782 : OAI22_X1 port map( A1 => n12659, A2 => n13350, B1 => n5645, B2 => 
                           n13347, ZN => n3308);
   U4783 : OAI22_X1 port map( A1 => n12660, A2 => n13350, B1 => n5655, B2 => 
                           n13347, ZN => n3271);
   U4784 : AOI221_X1 port map( B1 => n13020, B2 => n6170, C1 => n13017, C2 => 
                           n15619, A => n4682, ZN => n4679);
   U4785 : OAI22_X1 port map( A1 => n14956, A2 => n13014, B1 => n15930, B2 => 
                           n13011, ZN => n4682);
   U4786 : AOI221_X1 port map( B1 => n13248, B2 => n6170, C1 => n13245, C2 => 
                           n15619, A => n3398, ZN => n3395);
   U4787 : OAI22_X1 port map( A1 => n14956, A2 => n13242, B1 => n15930, B2 => 
                           n13239, ZN => n3398);
   U4788 : AOI221_X1 port map( B1 => n13167, B2 => n6042, C1 => n13164, C2 => 
                           n6074, A => n3408, ZN => n3401);
   U4789 : OAI22_X1 port map( A1 => n15117, A2 => n13161, B1 => n15149, B2 => 
                           n13158, ZN => n3408);
   U4790 : OAI22_X1 port map( A1 => n6870, A2 => n13120, B1 => n710, B2 => 
                           n13117, ZN => n5670);
   U4791 : OAI22_X1 port map( A1 => n6830, A2 => n13093, B1 => n711, B2 => 
                           n13090, ZN => n5680);
   U4792 : OAI22_X1 port map( A1 => n6871, A2 => n13120, B1 => n707, B2 => 
                           n13117, ZN => n5598);
   U4793 : OAI22_X1 port map( A1 => n6831, A2 => n13093, B1 => n708, B2 => 
                           n13090, ZN => n5600);
   U4794 : OAI22_X1 port map( A1 => n6872, A2 => n13120, B1 => n704, B2 => 
                           n13117, ZN => n5536);
   U4795 : OAI22_X1 port map( A1 => n6832, A2 => n13093, B1 => n705, B2 => 
                           n13090, ZN => n5539);
   U4796 : OAI22_X1 port map( A1 => n6873, A2 => n13120, B1 => n701, B2 => 
                           n13117, ZN => n5474);
   U4797 : OAI22_X1 port map( A1 => n6833, A2 => n13093, B1 => n702, B2 => 
                           n13090, ZN => n5478);
   U4798 : OAI22_X1 port map( A1 => n6874, A2 => n13120, B1 => n698, B2 => 
                           n13117, ZN => n5418);
   U4799 : OAI22_X1 port map( A1 => n6834, A2 => n13093, B1 => n699, B2 => 
                           n13090, ZN => n5420);
   U4800 : OAI22_X1 port map( A1 => n6875, A2 => n13120, B1 => n695, B2 => 
                           n13117, ZN => n5369);
   U4801 : OAI22_X1 port map( A1 => n6835, A2 => n13093, B1 => n696, B2 => 
                           n13090, ZN => n5371);
   U4802 : OAI22_X1 port map( A1 => n6876, A2 => n13120, B1 => n692, B2 => 
                           n13117, ZN => n5332);
   U4803 : OAI22_X1 port map( A1 => n6836, A2 => n13093, B1 => n693, B2 => 
                           n13090, ZN => n5334);
   U4804 : OAI22_X1 port map( A1 => n6877, A2 => n13120, B1 => n689, B2 => 
                           n13117, ZN => n5295);
   U4805 : OAI22_X1 port map( A1 => n6837, A2 => n13093, B1 => n690, B2 => 
                           n13090, ZN => n5297);
   U4806 : OAI22_X1 port map( A1 => n6878, A2 => n13120, B1 => n686, B2 => 
                           n13117, ZN => n5258);
   U4807 : OAI22_X1 port map( A1 => n6838, A2 => n13093, B1 => n687, B2 => 
                           n13090, ZN => n5260);
   U4808 : OAI22_X1 port map( A1 => n6879, A2 => n13120, B1 => n683, B2 => 
                           n13117, ZN => n5221);
   U4809 : OAI22_X1 port map( A1 => n6839, A2 => n13093, B1 => n684, B2 => 
                           n13090, ZN => n5223);
   U4810 : OAI22_X1 port map( A1 => n6880, A2 => n13120, B1 => n680, B2 => 
                           n13117, ZN => n5184);
   U4811 : OAI22_X1 port map( A1 => n6840, A2 => n13093, B1 => n681, B2 => 
                           n13090, ZN => n5186);
   U4812 : OAI22_X1 port map( A1 => n6881, A2 => n13120, B1 => n677, B2 => 
                           n13117, ZN => n5147);
   U4813 : OAI22_X1 port map( A1 => n6841, A2 => n13093, B1 => n678, B2 => 
                           n13090, ZN => n5149);
   U4814 : OAI22_X1 port map( A1 => n6882, A2 => n13121, B1 => n674, B2 => 
                           n13118, ZN => n5110);
   U4815 : OAI22_X1 port map( A1 => n6883, A2 => n13094, B1 => n675, B2 => 
                           n13091, ZN => n5112);
   U4816 : OAI22_X1 port map( A1 => n6884, A2 => n13121, B1 => n671, B2 => 
                           n13118, ZN => n5073);
   U4817 : OAI22_X1 port map( A1 => n6885, A2 => n13094, B1 => n672, B2 => 
                           n13091, ZN => n5075);
   U4818 : OAI22_X1 port map( A1 => n6886, A2 => n13121, B1 => n668, B2 => 
                           n13118, ZN => n5036);
   U4819 : OAI22_X1 port map( A1 => n6887, A2 => n13094, B1 => n669, B2 => 
                           n13091, ZN => n5038);
   U4820 : OAI22_X1 port map( A1 => n6888, A2 => n13121, B1 => n665, B2 => 
                           n13118, ZN => n4999);
   U4821 : OAI22_X1 port map( A1 => n6889, A2 => n13094, B1 => n666, B2 => 
                           n13091, ZN => n5001);
   U4822 : OAI22_X1 port map( A1 => n6890, A2 => n13121, B1 => n662, B2 => 
                           n13118, ZN => n4962);
   U4823 : OAI22_X1 port map( A1 => n6794, A2 => n13094, B1 => n6922, B2 => 
                           n13091, ZN => n4964);
   U4824 : OAI22_X1 port map( A1 => n6891, A2 => n13121, B1 => n659, B2 => 
                           n13118, ZN => n4925);
   U4825 : OAI22_X1 port map( A1 => n6795, A2 => n13094, B1 => n6923, B2 => 
                           n13091, ZN => n4927);
   U4826 : OAI22_X1 port map( A1 => n6892, A2 => n13121, B1 => n656, B2 => 
                           n13118, ZN => n4888);
   U4827 : OAI22_X1 port map( A1 => n6796, A2 => n13094, B1 => n6924, B2 => 
                           n13091, ZN => n4890);
   U4828 : OAI22_X1 port map( A1 => n6893, A2 => n13121, B1 => n653, B2 => 
                           n13118, ZN => n4851);
   U4829 : OAI22_X1 port map( A1 => n6797, A2 => n13094, B1 => n6925, B2 => 
                           n13091, ZN => n4853);
   U4830 : OAI22_X1 port map( A1 => n6810, A2 => n13121, B1 => n6938, B2 => 
                           n13118, ZN => n4814);
   U4831 : OAI22_X1 port map( A1 => n6798, A2 => n13094, B1 => n6926, B2 => 
                           n13091, ZN => n4816);
   U4832 : OAI22_X1 port map( A1 => n6811, A2 => n13121, B1 => n6939, B2 => 
                           n13118, ZN => n4777);
   U4833 : OAI22_X1 port map( A1 => n6799, A2 => n13094, B1 => n6927, B2 => 
                           n13091, ZN => n4779);
   U4834 : OAI22_X1 port map( A1 => n6812, A2 => n13121, B1 => n6940, B2 => 
                           n13118, ZN => n4740);
   U4835 : OAI22_X1 port map( A1 => n6800, A2 => n13094, B1 => n6928, B2 => 
                           n13091, ZN => n4742);
   U4836 : OAI22_X1 port map( A1 => n6813, A2 => n13121, B1 => n6941, B2 => 
                           n13118, ZN => n4703);
   U4837 : OAI22_X1 port map( A1 => n6801, A2 => n13094, B1 => n6929, B2 => 
                           n13091, ZN => n4705);
   U4838 : OAI22_X1 port map( A1 => n12661, A2 => n13348, B1 => n5385, B2 => 
                           n13345, ZN => n4277);
   U4839 : OAI22_X1 port map( A1 => n12662, A2 => n13321, B1 => n5387, B2 => 
                           n13318, ZN => n4283);
   U4840 : OAI22_X1 port map( A1 => n12663, A2 => n13348, B1 => n5395, B2 => 
                           n13345, ZN => n4233);
   U4841 : OAI22_X1 port map( A1 => n12664, A2 => n13321, B1 => n5397, B2 => 
                           n13318, ZN => n4235);
   U4842 : OAI22_X1 port map( A1 => n12665, A2 => n13348, B1 => n5405, B2 => 
                           n13345, ZN => n4196);
   U4843 : OAI22_X1 port map( A1 => n12666, A2 => n13321, B1 => n5407, B2 => 
                           n13318, ZN => n4198);
   U4844 : OAI22_X1 port map( A1 => n12667, A2 => n13348, B1 => n5415, B2 => 
                           n13345, ZN => n4159);
   U4845 : OAI22_X1 port map( A1 => n12668, A2 => n13321, B1 => n5417, B2 => 
                           n13318, ZN => n4161);
   U4846 : OAI22_X1 port map( A1 => n12669, A2 => n13348, B1 => n5425, B2 => 
                           n13345, ZN => n4122);
   U4847 : OAI22_X1 port map( A1 => n12670, A2 => n13321, B1 => n5427, B2 => 
                           n13318, ZN => n4124);
   U4848 : OAI22_X1 port map( A1 => n12671, A2 => n13348, B1 => n5435, B2 => 
                           n13345, ZN => n4085);
   U4849 : OAI22_X1 port map( A1 => n12672, A2 => n13321, B1 => n5437, B2 => 
                           n13318, ZN => n4087);
   U4850 : OAI22_X1 port map( A1 => n12673, A2 => n13348, B1 => n5445, B2 => 
                           n13345, ZN => n4048);
   U4851 : OAI22_X1 port map( A1 => n12674, A2 => n13321, B1 => n5447, B2 => 
                           n13318, ZN => n4050);
   U4852 : OAI22_X1 port map( A1 => n12675, A2 => n13348, B1 => n5455, B2 => 
                           n13345, ZN => n4011);
   U4853 : OAI22_X1 port map( A1 => n12676, A2 => n13321, B1 => n5457, B2 => 
                           n13318, ZN => n4013);
   U4854 : OAI22_X1 port map( A1 => n12677, A2 => n13348, B1 => n5465, B2 => 
                           n13345, ZN => n3974);
   U4855 : OAI22_X1 port map( A1 => n12678, A2 => n13321, B1 => n5467, B2 => 
                           n13318, ZN => n3976);
   U4856 : OAI22_X1 port map( A1 => n12679, A2 => n13348, B1 => n5475, B2 => 
                           n13345, ZN => n3937);
   U4857 : OAI22_X1 port map( A1 => n12680, A2 => n13321, B1 => n5477, B2 => 
                           n13318, ZN => n3939);
   U4858 : OAI22_X1 port map( A1 => n12681, A2 => n13348, B1 => n5485, B2 => 
                           n13345, ZN => n3900);
   U4859 : OAI22_X1 port map( A1 => n12682, A2 => n13321, B1 => n5487, B2 => 
                           n13318, ZN => n3902);
   U4860 : OAI22_X1 port map( A1 => n12683, A2 => n13348, B1 => n5495, B2 => 
                           n13345, ZN => n3863);
   U4861 : OAI22_X1 port map( A1 => n12684, A2 => n13321, B1 => n5497, B2 => 
                           n13318, ZN => n3865);
   U4862 : OAI22_X1 port map( A1 => n12685, A2 => n13349, B1 => n5505, B2 => 
                           n13346, ZN => n3826);
   U4863 : OAI22_X1 port map( A1 => n12686, A2 => n13322, B1 => n5507, B2 => 
                           n13319, ZN => n3828);
   U4864 : OAI22_X1 port map( A1 => n12687, A2 => n13349, B1 => n5515, B2 => 
                           n13346, ZN => n3789);
   U4865 : OAI22_X1 port map( A1 => n12688, A2 => n13322, B1 => n5517, B2 => 
                           n13319, ZN => n3791);
   U4866 : OAI22_X1 port map( A1 => n12689, A2 => n13349, B1 => n5525, B2 => 
                           n13346, ZN => n3752);
   U4867 : OAI22_X1 port map( A1 => n12690, A2 => n13322, B1 => n5527, B2 => 
                           n13319, ZN => n3754);
   U4868 : OAI22_X1 port map( A1 => n12691, A2 => n13349, B1 => n5535, B2 => 
                           n13346, ZN => n3715);
   U4869 : OAI22_X1 port map( A1 => n12692, A2 => n13322, B1 => n5537, B2 => 
                           n13319, ZN => n3717);
   U4870 : OAI22_X1 port map( A1 => n12693, A2 => n13349, B1 => n5545, B2 => 
                           n13346, ZN => n3678);
   U4871 : OAI22_X1 port map( A1 => n12694, A2 => n13322, B1 => n5547, B2 => 
                           n13319, ZN => n3680);
   U4872 : OAI22_X1 port map( A1 => n12695, A2 => n13349, B1 => n5555, B2 => 
                           n13346, ZN => n3641);
   U4873 : OAI22_X1 port map( A1 => n12696, A2 => n13322, B1 => n5557, B2 => 
                           n13319, ZN => n3643);
   U4874 : OAI22_X1 port map( A1 => n12697, A2 => n13349, B1 => n5565, B2 => 
                           n13346, ZN => n3604);
   U4875 : OAI22_X1 port map( A1 => n12698, A2 => n13322, B1 => n5567, B2 => 
                           n13319, ZN => n3606);
   U4876 : OAI22_X1 port map( A1 => n12699, A2 => n13349, B1 => n5575, B2 => 
                           n13346, ZN => n3567);
   U4877 : OAI22_X1 port map( A1 => n12700, A2 => n13322, B1 => n5577, B2 => 
                           n13319, ZN => n3569);
   U4878 : OAI22_X1 port map( A1 => n12701, A2 => n13349, B1 => n5585, B2 => 
                           n13346, ZN => n3530);
   U4879 : OAI22_X1 port map( A1 => n12702, A2 => n13322, B1 => n5587, B2 => 
                           n13319, ZN => n3532);
   U4880 : OAI22_X1 port map( A1 => n12703, A2 => n13349, B1 => n5595, B2 => 
                           n13346, ZN => n3493);
   U4881 : OAI22_X1 port map( A1 => n12704, A2 => n13322, B1 => n5597, B2 => 
                           n13319, ZN => n3495);
   U4882 : OAI22_X1 port map( A1 => n12705, A2 => n13349, B1 => n5605, B2 => 
                           n13346, ZN => n3456);
   U4883 : OAI22_X1 port map( A1 => n12706, A2 => n13322, B1 => n5607, B2 => 
                           n13319, ZN => n3458);
   U4884 : OAI22_X1 port map( A1 => n12707, A2 => n13349, B1 => n5615, B2 => 
                           n13346, ZN => n3419);
   U4885 : OAI22_X1 port map( A1 => n12708, A2 => n13322, B1 => n5617, B2 => 
                           n13319, ZN => n3421);
   U4886 : AOI221_X1 port map( B1 => n12991, B2 => n616, C1 => n12988, C2 => 
                           n15729, A => n5718, ZN => n5700);
   U4887 : OAI22_X1 port map( A1 => n14851, A2 => n12985, B1 => n14819, B2 => 
                           n12982, ZN => n5718);
   U4888 : AOI221_X1 port map( B1 => n12937, B2 => n6050, C1 => n12934, C2 => 
                           n6018, A => n5736, ZN => n5720);
   U4889 : OAI22_X1 port map( A1 => n15173, A2 => n12931, B1 => n15141, B2 => 
                           n12928, ZN => n5736);
   U4890 : AOI221_X1 port map( B1 => n12991, B2 => n614, C1 => n12988, C2 => 
                           n15728, A => n5628, ZN => n5616);
   U4891 : OAI22_X1 port map( A1 => n14850, A2 => n12985, B1 => n14818, B2 => 
                           n12982, ZN => n5628);
   U4892 : AOI221_X1 port map( B1 => n12937, B2 => n6051, C1 => n12934, C2 => 
                           n6019, A => n5640, ZN => n5629);
   U4893 : OAI22_X1 port map( A1 => n15172, A2 => n12931, B1 => n15140, B2 => 
                           n12928, ZN => n5640);
   U4894 : AOI221_X1 port map( B1 => n12991, B2 => n612, C1 => n12988, C2 => 
                           n15727, A => n5566, ZN => n5554);
   U4895 : OAI22_X1 port map( A1 => n14849, A2 => n12985, B1 => n14817, B2 => 
                           n12982, ZN => n5566);
   U4896 : AOI221_X1 port map( B1 => n12937, B2 => n6052, C1 => n12934, C2 => 
                           n6020, A => n5579, ZN => n5568);
   U4897 : OAI22_X1 port map( A1 => n15171, A2 => n12931, B1 => n15139, B2 => 
                           n12928, ZN => n5579);
   U4898 : AOI221_X1 port map( B1 => n12991, B2 => n610, C1 => n12988, C2 => 
                           n15726, A => n5504, ZN => n5491);
   U4899 : OAI22_X1 port map( A1 => n14848, A2 => n12985, B1 => n14816, B2 => 
                           n12982, ZN => n5504);
   U4900 : AOI221_X1 port map( B1 => n12937, B2 => n6053, C1 => n12934, C2 => 
                           n6021, A => n5518, ZN => n5506);
   U4901 : OAI22_X1 port map( A1 => n15170, A2 => n12931, B1 => n15138, B2 => 
                           n12928, ZN => n5518);
   U4902 : AOI221_X1 port map( B1 => n12991, B2 => n608, C1 => n12988, C2 => 
                           n15725, A => n5442, ZN => n5432);
   U4903 : OAI22_X1 port map( A1 => n14847, A2 => n12985, B1 => n14815, B2 => 
                           n12982, ZN => n5442);
   U4904 : AOI221_X1 port map( B1 => n12937, B2 => n6054, C1 => n12934, C2 => 
                           n6022, A => n5456, ZN => n5444);
   U4905 : OAI22_X1 port map( A1 => n15169, A2 => n12931, B1 => n15137, B2 => 
                           n12928, ZN => n5456);
   U4906 : AOI221_X1 port map( B1 => n12991, B2 => n606, C1 => n12988, C2 => 
                           n15724, A => n5390, ZN => n5380);
   U4907 : OAI22_X1 port map( A1 => n14846, A2 => n12985, B1 => n14814, B2 => 
                           n12982, ZN => n5390);
   U4908 : AOI221_X1 port map( B1 => n12937, B2 => n6055, C1 => n12934, C2 => 
                           n6023, A => n5401, ZN => n5391);
   U4909 : OAI22_X1 port map( A1 => n15168, A2 => n12931, B1 => n15136, B2 => 
                           n12928, ZN => n5401);
   U4910 : AOI221_X1 port map( B1 => n12991, B2 => n604, C1 => n12988, C2 => 
                           n15723, A => n5350, ZN => n5343);
   U4911 : OAI22_X1 port map( A1 => n14845, A2 => n12985, B1 => n14813, B2 => 
                           n12982, ZN => n5350);
   U4912 : AOI221_X1 port map( B1 => n12937, B2 => n6056, C1 => n12934, C2 => 
                           n6024, A => n5358, ZN => n5351);
   U4913 : OAI22_X1 port map( A1 => n15167, A2 => n12931, B1 => n15135, B2 => 
                           n12928, ZN => n5358);
   U4914 : AOI221_X1 port map( B1 => n12991, B2 => n602, C1 => n12988, C2 => 
                           n15722, A => n5313, ZN => n5306);
   U4915 : OAI22_X1 port map( A1 => n14844, A2 => n12985, B1 => n14812, B2 => 
                           n12982, ZN => n5313);
   U4916 : AOI221_X1 port map( B1 => n12937, B2 => n6057, C1 => n12934, C2 => 
                           n6025, A => n5321, ZN => n5314);
   U4917 : OAI22_X1 port map( A1 => n15166, A2 => n12931, B1 => n15134, B2 => 
                           n12928, ZN => n5321);
   U4918 : AOI221_X1 port map( B1 => n12991, B2 => n600, C1 => n12988, C2 => 
                           n15721, A => n5276, ZN => n5269);
   U4919 : OAI22_X1 port map( A1 => n14843, A2 => n12985, B1 => n14811, B2 => 
                           n12982, ZN => n5276);
   U4920 : AOI221_X1 port map( B1 => n12937, B2 => n6058, C1 => n12934, C2 => 
                           n6026, A => n5284, ZN => n5277);
   U4921 : OAI22_X1 port map( A1 => n15165, A2 => n12931, B1 => n15133, B2 => 
                           n12928, ZN => n5284);
   U4922 : AOI221_X1 port map( B1 => n12991, B2 => n598, C1 => n12988, C2 => 
                           n15720, A => n5239, ZN => n5232);
   U4923 : OAI22_X1 port map( A1 => n14842, A2 => n12985, B1 => n14810, B2 => 
                           n12982, ZN => n5239);
   U4924 : AOI221_X1 port map( B1 => n12937, B2 => n6059, C1 => n12934, C2 => 
                           n6027, A => n5247, ZN => n5240);
   U4925 : OAI22_X1 port map( A1 => n15164, A2 => n12931, B1 => n15132, B2 => 
                           n12928, ZN => n5247);
   U4926 : AOI221_X1 port map( B1 => n12991, B2 => n596, C1 => n12988, C2 => 
                           n15719, A => n5202, ZN => n5195);
   U4927 : OAI22_X1 port map( A1 => n14841, A2 => n12985, B1 => n14809, B2 => 
                           n12982, ZN => n5202);
   U4928 : AOI221_X1 port map( B1 => n12937, B2 => n6060, C1 => n12934, C2 => 
                           n6028, A => n5210, ZN => n5203);
   U4929 : OAI22_X1 port map( A1 => n15163, A2 => n12931, B1 => n15131, B2 => 
                           n12928, ZN => n5210);
   U4930 : AOI221_X1 port map( B1 => n12991, B2 => n594, C1 => n12988, C2 => 
                           n15718, A => n5165, ZN => n5158);
   U4931 : OAI22_X1 port map( A1 => n14840, A2 => n12985, B1 => n14808, B2 => 
                           n12982, ZN => n5165);
   U4932 : AOI221_X1 port map( B1 => n12937, B2 => n6061, C1 => n12934, C2 => 
                           n6029, A => n5173, ZN => n5166);
   U4933 : OAI22_X1 port map( A1 => n15162, A2 => n12931, B1 => n15130, B2 => 
                           n12928, ZN => n5173);
   U4934 : AOI221_X1 port map( B1 => n12938, B2 => n6062, C1 => n12935, C2 => 
                           n6030, A => n5136, ZN => n5129);
   U4935 : OAI22_X1 port map( A1 => n15161, A2 => n12932, B1 => n15129, B2 => 
                           n12929, ZN => n5136);
   U4936 : AOI221_X1 port map( B1 => n12938, B2 => n6063, C1 => n12935, C2 => 
                           n6031, A => n5099, ZN => n5092);
   U4937 : OAI22_X1 port map( A1 => n15160, A2 => n12932, B1 => n15128, B2 => 
                           n12929, ZN => n5099);
   U4938 : AOI221_X1 port map( B1 => n12938, B2 => n6064, C1 => n12935, C2 => 
                           n6032, A => n5062, ZN => n5055);
   U4939 : OAI22_X1 port map( A1 => n15159, A2 => n12932, B1 => n15127, B2 => 
                           n12929, ZN => n5062);
   U4940 : AOI221_X1 port map( B1 => n12938, B2 => n6065, C1 => n12935, C2 => 
                           n6033, A => n5025, ZN => n5018);
   U4941 : OAI22_X1 port map( A1 => n15158, A2 => n12932, B1 => n15126, B2 => 
                           n12929, ZN => n5025);
   U4942 : AOI221_X1 port map( B1 => n12938, B2 => n6066, C1 => n12935, C2 => 
                           n6034, A => n4988, ZN => n4981);
   U4943 : OAI22_X1 port map( A1 => n15157, A2 => n12932, B1 => n15125, B2 => 
                           n12929, ZN => n4988);
   U4944 : AOI221_X1 port map( B1 => n12938, B2 => n6067, C1 => n12935, C2 => 
                           n6035, A => n4951, ZN => n4944);
   U4945 : OAI22_X1 port map( A1 => n15156, A2 => n12932, B1 => n15124, B2 => 
                           n12929, ZN => n4951);
   U4946 : AOI221_X1 port map( B1 => n12938, B2 => n6068, C1 => n12935, C2 => 
                           n6036, A => n4914, ZN => n4907);
   U4947 : OAI22_X1 port map( A1 => n15155, A2 => n12932, B1 => n15123, B2 => 
                           n12929, ZN => n4914);
   U4948 : AOI221_X1 port map( B1 => n12938, B2 => n6069, C1 => n12935, C2 => 
                           n6037, A => n4877, ZN => n4870);
   U4949 : OAI22_X1 port map( A1 => n15154, A2 => n12932, B1 => n15122, B2 => 
                           n12929, ZN => n4877);
   U4950 : AOI221_X1 port map( B1 => n12938, B2 => n6070, C1 => n12935, C2 => 
                           n6038, A => n4840, ZN => n4833);
   U4951 : OAI22_X1 port map( A1 => n15153, A2 => n12932, B1 => n15121, B2 => 
                           n12929, ZN => n4840);
   U4952 : AOI221_X1 port map( B1 => n12938, B2 => n6071, C1 => n12935, C2 => 
                           n6039, A => n4803, ZN => n4796);
   U4953 : OAI22_X1 port map( A1 => n15152, A2 => n12932, B1 => n15120, B2 => 
                           n12929, ZN => n4803);
   U4954 : AOI221_X1 port map( B1 => n12938, B2 => n6072, C1 => n12935, C2 => 
                           n6040, A => n4766, ZN => n4759);
   U4955 : OAI22_X1 port map( A1 => n15151, A2 => n12932, B1 => n15119, B2 => 
                           n12929, ZN => n4766);
   U4956 : AOI221_X1 port map( B1 => n12938, B2 => n6073, C1 => n12935, C2 => 
                           n6041, A => n4729, ZN => n4722);
   U4957 : OAI22_X1 port map( A1 => n15150, A2 => n12932, B1 => n15118, B2 => 
                           n12929, ZN => n4729);
   U4958 : AOI221_X1 port map( B1 => n13219, B2 => n616, C1 => n13216, C2 => 
                           n15729, A => n4303, ZN => n4294);
   U4959 : OAI22_X1 port map( A1 => n14851, A2 => n13213, B1 => n14819, B2 => 
                           n13210, ZN => n4303);
   U4960 : AOI221_X1 port map( B1 => n13165, B2 => n6018, C1 => n13162, C2 => 
                           n6050, A => n4312, ZN => n4304);
   U4961 : OAI22_X1 port map( A1 => n15141, A2 => n13159, B1 => n15173, B2 => 
                           n13156, ZN => n4312);
   U4962 : AOI221_X1 port map( B1 => n13219, B2 => n614, C1 => n13216, C2 => 
                           n15728, A => n4251, ZN => n4244);
   U4963 : OAI22_X1 port map( A1 => n14850, A2 => n13213, B1 => n14818, B2 => 
                           n13210, ZN => n4251);
   U4964 : AOI221_X1 port map( B1 => n13165, B2 => n6019, C1 => n13162, C2 => 
                           n6051, A => n4259, ZN => n4252);
   U4965 : OAI22_X1 port map( A1 => n15140, A2 => n13159, B1 => n15172, B2 => 
                           n13156, ZN => n4259);
   U4966 : AOI221_X1 port map( B1 => n13219, B2 => n612, C1 => n13216, C2 => 
                           n15727, A => n4214, ZN => n4207);
   U4967 : OAI22_X1 port map( A1 => n14849, A2 => n13213, B1 => n14817, B2 => 
                           n13210, ZN => n4214);
   U4968 : AOI221_X1 port map( B1 => n13165, B2 => n6020, C1 => n13162, C2 => 
                           n6052, A => n4222, ZN => n4215);
   U4969 : OAI22_X1 port map( A1 => n15139, A2 => n13159, B1 => n15171, B2 => 
                           n13156, ZN => n4222);
   U4970 : AOI221_X1 port map( B1 => n13219, B2 => n610, C1 => n13216, C2 => 
                           n15726, A => n4177, ZN => n4170);
   U4971 : OAI22_X1 port map( A1 => n14848, A2 => n13213, B1 => n14816, B2 => 
                           n13210, ZN => n4177);
   U4972 : AOI221_X1 port map( B1 => n13165, B2 => n6021, C1 => n13162, C2 => 
                           n6053, A => n4185, ZN => n4178);
   U4973 : OAI22_X1 port map( A1 => n15138, A2 => n13159, B1 => n15170, B2 => 
                           n13156, ZN => n4185);
   U4974 : AOI221_X1 port map( B1 => n13219, B2 => n608, C1 => n13216, C2 => 
                           n15725, A => n4140, ZN => n4133);
   U4975 : OAI22_X1 port map( A1 => n14847, A2 => n13213, B1 => n14815, B2 => 
                           n13210, ZN => n4140);
   U4976 : AOI221_X1 port map( B1 => n13165, B2 => n6022, C1 => n13162, C2 => 
                           n6054, A => n4148, ZN => n4141);
   U4977 : OAI22_X1 port map( A1 => n15137, A2 => n13159, B1 => n15169, B2 => 
                           n13156, ZN => n4148);
   U4978 : AOI221_X1 port map( B1 => n13219, B2 => n606, C1 => n13216, C2 => 
                           n15724, A => n4103, ZN => n4096);
   U4979 : OAI22_X1 port map( A1 => n14846, A2 => n13213, B1 => n14814, B2 => 
                           n13210, ZN => n4103);
   U4980 : AOI221_X1 port map( B1 => n13165, B2 => n6023, C1 => n13162, C2 => 
                           n6055, A => n4111, ZN => n4104);
   U4981 : OAI22_X1 port map( A1 => n15136, A2 => n13159, B1 => n15168, B2 => 
                           n13156, ZN => n4111);
   U4982 : AOI221_X1 port map( B1 => n13219, B2 => n604, C1 => n13216, C2 => 
                           n15723, A => n4066, ZN => n4059);
   U4983 : OAI22_X1 port map( A1 => n14845, A2 => n13213, B1 => n14813, B2 => 
                           n13210, ZN => n4066);
   U4984 : AOI221_X1 port map( B1 => n13165, B2 => n6024, C1 => n13162, C2 => 
                           n6056, A => n4074, ZN => n4067);
   U4985 : OAI22_X1 port map( A1 => n15135, A2 => n13159, B1 => n15167, B2 => 
                           n13156, ZN => n4074);
   U4986 : AOI221_X1 port map( B1 => n13219, B2 => n602, C1 => n13216, C2 => 
                           n15722, A => n4029, ZN => n4022);
   U4987 : OAI22_X1 port map( A1 => n14844, A2 => n13213, B1 => n14812, B2 => 
                           n13210, ZN => n4029);
   U4988 : AOI221_X1 port map( B1 => n13165, B2 => n6025, C1 => n13162, C2 => 
                           n6057, A => n4037, ZN => n4030);
   U4989 : OAI22_X1 port map( A1 => n15134, A2 => n13159, B1 => n15166, B2 => 
                           n13156, ZN => n4037);
   U4990 : AOI221_X1 port map( B1 => n13219, B2 => n600, C1 => n13216, C2 => 
                           n15721, A => n3992, ZN => n3985);
   U4991 : OAI22_X1 port map( A1 => n14843, A2 => n13213, B1 => n14811, B2 => 
                           n13210, ZN => n3992);
   U4992 : AOI221_X1 port map( B1 => n13165, B2 => n6026, C1 => n13162, C2 => 
                           n6058, A => n4000, ZN => n3993);
   U4993 : OAI22_X1 port map( A1 => n15133, A2 => n13159, B1 => n15165, B2 => 
                           n13156, ZN => n4000);
   U4994 : AOI221_X1 port map( B1 => n13219, B2 => n598, C1 => n13216, C2 => 
                           n15720, A => n3955, ZN => n3948);
   U4995 : OAI22_X1 port map( A1 => n14842, A2 => n13213, B1 => n14810, B2 => 
                           n13210, ZN => n3955);
   U4996 : AOI221_X1 port map( B1 => n13165, B2 => n6027, C1 => n13162, C2 => 
                           n6059, A => n3963, ZN => n3956);
   U4997 : OAI22_X1 port map( A1 => n15132, A2 => n13159, B1 => n15164, B2 => 
                           n13156, ZN => n3963);
   U4998 : AOI221_X1 port map( B1 => n13219, B2 => n596, C1 => n13216, C2 => 
                           n15719, A => n3918, ZN => n3911);
   U4999 : OAI22_X1 port map( A1 => n14841, A2 => n13213, B1 => n14809, B2 => 
                           n13210, ZN => n3918);
   U5000 : AOI221_X1 port map( B1 => n13165, B2 => n6028, C1 => n13162, C2 => 
                           n6060, A => n3926, ZN => n3919);
   U5001 : OAI22_X1 port map( A1 => n15131, A2 => n13159, B1 => n15163, B2 => 
                           n13156, ZN => n3926);
   U5002 : AOI221_X1 port map( B1 => n13219, B2 => n594, C1 => n13216, C2 => 
                           n15718, A => n3881, ZN => n3874);
   U5003 : OAI22_X1 port map( A1 => n14840, A2 => n13213, B1 => n14808, B2 => 
                           n13210, ZN => n3881);
   U5004 : AOI221_X1 port map( B1 => n13165, B2 => n6029, C1 => n13162, C2 => 
                           n6061, A => n3889, ZN => n3882);
   U5005 : OAI22_X1 port map( A1 => n15130, A2 => n13159, B1 => n15162, B2 => 
                           n13156, ZN => n3889);
   U5006 : OAI22_X1 port map( A1 => n13829, A2 => n13407, B1 => n6942, B2 => 
                           n13402, ZN => n7770);
   U5007 : OAI22_X1 port map( A1 => n13835, A2 => n13407, B1 => n6943, B2 => 
                           n13402, ZN => n7771);
   U5008 : OAI22_X1 port map( A1 => n13841, A2 => n13407, B1 => n6944, B2 => 
                           n13402, ZN => n7772);
   U5009 : OAI22_X1 port map( A1 => n13847, A2 => n13407, B1 => n6945, B2 => 
                           n13402, ZN => n7773);
   U5010 : OAI22_X1 port map( A1 => n13853, A2 => n13407, B1 => n6946, B2 => 
                           n13402, ZN => n7774);
   U5011 : OAI22_X1 port map( A1 => n13859, A2 => n13407, B1 => n6947, B2 => 
                           n13402, ZN => n7775);
   U5012 : OAI22_X1 port map( A1 => n13865, A2 => n13407, B1 => n6948, B2 => 
                           n13402, ZN => n7776);
   U5013 : OAI22_X1 port map( A1 => n13871, A2 => n13407, B1 => n6949, B2 => 
                           n13402, ZN => n7777);
   U5014 : OAI22_X1 port map( A1 => n13877, A2 => n13406, B1 => n6950, B2 => 
                           n13402, ZN => n7778);
   U5015 : OAI22_X1 port map( A1 => n13883, A2 => n13406, B1 => n6951, B2 => 
                           n13402, ZN => n7779);
   U5016 : OAI22_X1 port map( A1 => n13889, A2 => n13406, B1 => n6952, B2 => 
                           n13402, ZN => n7780);
   U5017 : OAI22_X1 port map( A1 => n13895, A2 => n13406, B1 => n6953, B2 => 
                           n13402, ZN => n7781);
   U5018 : OAI22_X1 port map( A1 => n13901, A2 => n13406, B1 => n6954, B2 => 
                           n13403, ZN => n7782);
   U5019 : OAI22_X1 port map( A1 => n13907, A2 => n13406, B1 => n6955, B2 => 
                           n13403, ZN => n7783);
   U5020 : OAI22_X1 port map( A1 => n13913, A2 => n13406, B1 => n6956, B2 => 
                           n13403, ZN => n7784);
   U5021 : OAI22_X1 port map( A1 => n13919, A2 => n13406, B1 => n6957, B2 => 
                           n13403, ZN => n7785);
   U5022 : OAI22_X1 port map( A1 => n13925, A2 => n13406, B1 => n6958, B2 => 
                           n13403, ZN => n7786);
   U5023 : OAI22_X1 port map( A1 => n13931, A2 => n13406, B1 => n6959, B2 => 
                           n13403, ZN => n7787);
   U5024 : OAI22_X1 port map( A1 => n13937, A2 => n13406, B1 => n6960, B2 => 
                           n13403, ZN => n7788);
   U5025 : OAI22_X1 port map( A1 => n13943, A2 => n13406, B1 => n6961, B2 => 
                           n13403, ZN => n7789);
   U5026 : OAI22_X1 port map( A1 => n13949, A2 => n13405, B1 => n6962, B2 => 
                           n13403, ZN => n7790);
   U5027 : OAI22_X1 port map( A1 => n13955, A2 => n13405, B1 => n6963, B2 => 
                           n13403, ZN => n7791);
   U5028 : OAI22_X1 port map( A1 => n13961, A2 => n13405, B1 => n6964, B2 => 
                           n13403, ZN => n7792);
   U5029 : OAI22_X1 port map( A1 => n13967, A2 => n13405, B1 => n6965, B2 => 
                           n13403, ZN => n7793);
   U5030 : OAI22_X1 port map( A1 => n13973, A2 => n13405, B1 => n6966, B2 => 
                           n13404, ZN => n7794);
   U5031 : OAI22_X1 port map( A1 => n13979, A2 => n13405, B1 => n6967, B2 => 
                           n13404, ZN => n7795);
   U5032 : OAI22_X1 port map( A1 => n13985, A2 => n13405, B1 => n6968, B2 => 
                           n13404, ZN => n7796);
   U5033 : OAI22_X1 port map( A1 => n13991, A2 => n13405, B1 => n6969, B2 => 
                           n13404, ZN => n7797);
   U5034 : OAI22_X1 port map( A1 => n13997, A2 => n13405, B1 => n6970, B2 => 
                           n13404, ZN => n7798);
   U5035 : OAI22_X1 port map( A1 => n14003, A2 => n13405, B1 => n6971, B2 => 
                           n13404, ZN => n7799);
   U5036 : OAI22_X1 port map( A1 => n14009, A2 => n13405, B1 => n6972, B2 => 
                           n13404, ZN => n7800);
   U5037 : OAI22_X1 port map( A1 => n14018, A2 => n13405, B1 => n6973, B2 => 
                           n13404, ZN => n7801);
   U5038 : OAI22_X1 port map( A1 => n13829, A2 => n13413, B1 => n7160, B2 => 
                           n13408, ZN => n7802);
   U5039 : OAI22_X1 port map( A1 => n13835, A2 => n13413, B1 => n7161, B2 => 
                           n13408, ZN => n7803);
   U5040 : OAI22_X1 port map( A1 => n13841, A2 => n13413, B1 => n7162, B2 => 
                           n13408, ZN => n7804);
   U5041 : OAI22_X1 port map( A1 => n13847, A2 => n13413, B1 => n7163, B2 => 
                           n13408, ZN => n7805);
   U5042 : OAI22_X1 port map( A1 => n13853, A2 => n13413, B1 => n7164, B2 => 
                           n13408, ZN => n7806);
   U5043 : OAI22_X1 port map( A1 => n13859, A2 => n13413, B1 => n7165, B2 => 
                           n13408, ZN => n7807);
   U5044 : OAI22_X1 port map( A1 => n13865, A2 => n13413, B1 => n7166, B2 => 
                           n13408, ZN => n7808);
   U5045 : OAI22_X1 port map( A1 => n13871, A2 => n13413, B1 => n7167, B2 => 
                           n13408, ZN => n7809);
   U5046 : OAI22_X1 port map( A1 => n13877, A2 => n13412, B1 => n7168, B2 => 
                           n13408, ZN => n7810);
   U5047 : OAI22_X1 port map( A1 => n13883, A2 => n13412, B1 => n7169, B2 => 
                           n13408, ZN => n7811);
   U5048 : OAI22_X1 port map( A1 => n13889, A2 => n13412, B1 => n7170, B2 => 
                           n13408, ZN => n7812);
   U5049 : OAI22_X1 port map( A1 => n13895, A2 => n13412, B1 => n7171, B2 => 
                           n13408, ZN => n7813);
   U5050 : OAI22_X1 port map( A1 => n13901, A2 => n13412, B1 => n7172, B2 => 
                           n13409, ZN => n7814);
   U5051 : OAI22_X1 port map( A1 => n13907, A2 => n13412, B1 => n7173, B2 => 
                           n13409, ZN => n7815);
   U5052 : OAI22_X1 port map( A1 => n13913, A2 => n13412, B1 => n7174, B2 => 
                           n13409, ZN => n7816);
   U5053 : OAI22_X1 port map( A1 => n13919, A2 => n13412, B1 => n7175, B2 => 
                           n13409, ZN => n7817);
   U5054 : OAI22_X1 port map( A1 => n13925, A2 => n13412, B1 => n7176, B2 => 
                           n13409, ZN => n7818);
   U5055 : OAI22_X1 port map( A1 => n13931, A2 => n13412, B1 => n7177, B2 => 
                           n13409, ZN => n7819);
   U5056 : OAI22_X1 port map( A1 => n13937, A2 => n13412, B1 => n7178, B2 => 
                           n13409, ZN => n7820);
   U5057 : OAI22_X1 port map( A1 => n13943, A2 => n13412, B1 => n7179, B2 => 
                           n13409, ZN => n7821);
   U5058 : OAI22_X1 port map( A1 => n13949, A2 => n13411, B1 => n7180, B2 => 
                           n13409, ZN => n7822);
   U5059 : OAI22_X1 port map( A1 => n13955, A2 => n13411, B1 => n7181, B2 => 
                           n13409, ZN => n7823);
   U5060 : OAI22_X1 port map( A1 => n13961, A2 => n13411, B1 => n7182, B2 => 
                           n13409, ZN => n7824);
   U5061 : OAI22_X1 port map( A1 => n13967, A2 => n13411, B1 => n7183, B2 => 
                           n13409, ZN => n7825);
   U5062 : OAI22_X1 port map( A1 => n13973, A2 => n13411, B1 => n7184, B2 => 
                           n13410, ZN => n7826);
   U5063 : OAI22_X1 port map( A1 => n13979, A2 => n13411, B1 => n7185, B2 => 
                           n13410, ZN => n7827);
   U5064 : OAI22_X1 port map( A1 => n13985, A2 => n13411, B1 => n7186, B2 => 
                           n13410, ZN => n7828);
   U5065 : OAI22_X1 port map( A1 => n13991, A2 => n13411, B1 => n7187, B2 => 
                           n13410, ZN => n7829);
   U5066 : OAI22_X1 port map( A1 => n13997, A2 => n13411, B1 => n7188, B2 => 
                           n13410, ZN => n7830);
   U5067 : OAI22_X1 port map( A1 => n14003, A2 => n13411, B1 => n7189, B2 => 
                           n13410, ZN => n7831);
   U5068 : OAI22_X1 port map( A1 => n14009, A2 => n13411, B1 => n7190, B2 => 
                           n13410, ZN => n7832);
   U5069 : OAI22_X1 port map( A1 => n14018, A2 => n13411, B1 => n7191, B2 => 
                           n13410, ZN => n7833);
   U5070 : OAI22_X1 port map( A1 => n13835, A2 => n13437, B1 => n7193, B2 => 
                           n13432, ZN => n7931);
   U5071 : OAI22_X1 port map( A1 => n13841, A2 => n13437, B1 => n7194, B2 => 
                           n13432, ZN => n7932);
   U5072 : OAI22_X1 port map( A1 => n13847, A2 => n13437, B1 => n7195, B2 => 
                           n13432, ZN => n7933);
   U5073 : OAI22_X1 port map( A1 => n13853, A2 => n13437, B1 => n7196, B2 => 
                           n13432, ZN => n7934);
   U5074 : OAI22_X1 port map( A1 => n13859, A2 => n13437, B1 => n7197, B2 => 
                           n13432, ZN => n7935);
   U5075 : OAI22_X1 port map( A1 => n13865, A2 => n13437, B1 => n7198, B2 => 
                           n13432, ZN => n7936);
   U5076 : OAI22_X1 port map( A1 => n13871, A2 => n13437, B1 => n7199, B2 => 
                           n13432, ZN => n7937);
   U5077 : OAI22_X1 port map( A1 => n13877, A2 => n13436, B1 => n7200, B2 => 
                           n13432, ZN => n7938);
   U5078 : OAI22_X1 port map( A1 => n13883, A2 => n13436, B1 => n7201, B2 => 
                           n13432, ZN => n7939);
   U5079 : OAI22_X1 port map( A1 => n13889, A2 => n13436, B1 => n7202, B2 => 
                           n13432, ZN => n7940);
   U5080 : OAI22_X1 port map( A1 => n13895, A2 => n13436, B1 => n7203, B2 => 
                           n13432, ZN => n7941);
   U5081 : OAI22_X1 port map( A1 => n13901, A2 => n13436, B1 => n7204, B2 => 
                           n13433, ZN => n7942);
   U5082 : OAI22_X1 port map( A1 => n13907, A2 => n13436, B1 => n7205, B2 => 
                           n13433, ZN => n7943);
   U5083 : OAI22_X1 port map( A1 => n13913, A2 => n13436, B1 => n7206, B2 => 
                           n13433, ZN => n7944);
   U5084 : OAI22_X1 port map( A1 => n13919, A2 => n13436, B1 => n7207, B2 => 
                           n13433, ZN => n7945);
   U5085 : OAI22_X1 port map( A1 => n13925, A2 => n13436, B1 => n7208, B2 => 
                           n13433, ZN => n7946);
   U5086 : OAI22_X1 port map( A1 => n13931, A2 => n13436, B1 => n7209, B2 => 
                           n13433, ZN => n7947);
   U5087 : OAI22_X1 port map( A1 => n13937, A2 => n13436, B1 => n7210, B2 => 
                           n13433, ZN => n7948);
   U5088 : OAI22_X1 port map( A1 => n13943, A2 => n13436, B1 => n7211, B2 => 
                           n13433, ZN => n7949);
   U5089 : OAI22_X1 port map( A1 => n13949, A2 => n13435, B1 => n7212, B2 => 
                           n13433, ZN => n7950);
   U5090 : OAI22_X1 port map( A1 => n13955, A2 => n13435, B1 => n7213, B2 => 
                           n13433, ZN => n7951);
   U5091 : OAI22_X1 port map( A1 => n13961, A2 => n13435, B1 => n7214, B2 => 
                           n13433, ZN => n7952);
   U5092 : OAI22_X1 port map( A1 => n13967, A2 => n13435, B1 => n7215, B2 => 
                           n13433, ZN => n7953);
   U5093 : OAI22_X1 port map( A1 => n13973, A2 => n13435, B1 => n7216, B2 => 
                           n13434, ZN => n7954);
   U5094 : OAI22_X1 port map( A1 => n13979, A2 => n13435, B1 => n7217, B2 => 
                           n13434, ZN => n7955);
   U5095 : OAI22_X1 port map( A1 => n13985, A2 => n13435, B1 => n7218, B2 => 
                           n13434, ZN => n7956);
   U5096 : OAI22_X1 port map( A1 => n13991, A2 => n13435, B1 => n7219, B2 => 
                           n13434, ZN => n7957);
   U5097 : OAI22_X1 port map( A1 => n13997, A2 => n13435, B1 => n7220, B2 => 
                           n13434, ZN => n7958);
   U5098 : OAI22_X1 port map( A1 => n14003, A2 => n13435, B1 => n7221, B2 => 
                           n13434, ZN => n7959);
   U5099 : OAI22_X1 port map( A1 => n14009, A2 => n13435, B1 => n7222, B2 => 
                           n13434, ZN => n7960);
   U5100 : OAI22_X1 port map( A1 => n14018, A2 => n13435, B1 => n7223, B2 => 
                           n13434, ZN => n7961);
   U5101 : OAI22_X1 port map( A1 => n14016, A2 => n13579, B1 => n13578, B2 => 
                           n12709, ZN => n8729);
   U5102 : OAI22_X1 port map( A1 => n14005, A2 => n13687, B1 => n13686, B2 => 
                           n14460, ZN => n9304);
   U5103 : OAI22_X1 port map( A1 => n14014, A2 => n13687, B1 => n13686, B2 => 
                           n14459, ZN => n9305);
   U5104 : OAI22_X1 port map( A1 => n13972, A2 => n13471, B1 => n13470, B2 => 
                           n12710, ZN => n8146);
   U5105 : OAI22_X1 port map( A1 => n13978, A2 => n13471, B1 => n13470, B2 => 
                           n12711, ZN => n8147);
   U5106 : OAI22_X1 port map( A1 => n13984, A2 => n13471, B1 => n13470, B2 => 
                           n12712, ZN => n8148);
   U5107 : OAI22_X1 port map( A1 => n13990, A2 => n13471, B1 => n13470, B2 => 
                           n12713, ZN => n8149);
   U5108 : OAI22_X1 port map( A1 => n13996, A2 => n13471, B1 => n13470, B2 => 
                           n12714, ZN => n8150);
   U5109 : OAI22_X1 port map( A1 => n14002, A2 => n13471, B1 => n13470, B2 => 
                           n12715, ZN => n8151);
   U5110 : OAI22_X1 port map( A1 => n14008, A2 => n13471, B1 => n13470, B2 => 
                           n12716, ZN => n8152);
   U5111 : OAI22_X1 port map( A1 => n14017, A2 => n13471, B1 => n13470, B2 => 
                           n12717, ZN => n8153);
   U5112 : OAI22_X1 port map( A1 => n13972, A2 => n13477, B1 => n13476, B2 => 
                           n12718, ZN => n8178);
   U5113 : OAI22_X1 port map( A1 => n13978, A2 => n13477, B1 => n13476, B2 => 
                           n12719, ZN => n8179);
   U5114 : OAI22_X1 port map( A1 => n13984, A2 => n13477, B1 => n13476, B2 => 
                           n12720, ZN => n8180);
   U5115 : OAI22_X1 port map( A1 => n13990, A2 => n13477, B1 => n13476, B2 => 
                           n12721, ZN => n8181);
   U5116 : OAI22_X1 port map( A1 => n13996, A2 => n13477, B1 => n13476, B2 => 
                           n12722, ZN => n8182);
   U5117 : OAI22_X1 port map( A1 => n14002, A2 => n13477, B1 => n13476, B2 => 
                           n12723, ZN => n8183);
   U5118 : OAI22_X1 port map( A1 => n14008, A2 => n13477, B1 => n13476, B2 => 
                           n12724, ZN => n8184);
   U5119 : OAI22_X1 port map( A1 => n14017, A2 => n13477, B1 => n13476, B2 => 
                           n12725, ZN => n8185);
   U5120 : OAI22_X1 port map( A1 => n14019, A2 => n13968, B1 => n6930, B2 => 
                           n14012, ZN => n9970);
   U5121 : OAI22_X1 port map( A1 => n14019, A2 => n13974, B1 => n6931, B2 => 
                           n14012, ZN => n9971);
   U5122 : OAI22_X1 port map( A1 => n14019, A2 => n13980, B1 => n6932, B2 => 
                           n14012, ZN => n9972);
   U5123 : OAI22_X1 port map( A1 => n14019, A2 => n13986, B1 => n6933, B2 => 
                           n14012, ZN => n9973);
   U5124 : OAI22_X1 port map( A1 => n14019, A2 => n13992, B1 => n6934, B2 => 
                           n14012, ZN => n9974);
   U5125 : OAI22_X1 port map( A1 => n14019, A2 => n13998, B1 => n6935, B2 => 
                           n14012, ZN => n9975);
   U5126 : OAI22_X1 port map( A1 => n14019, A2 => n14004, B1 => n6936, B2 => 
                           n14012, ZN => n9976);
   U5127 : OAI22_X1 port map( A1 => n14019, A2 => n14013, B1 => n6937, B2 => 
                           n14012, ZN => n9977);
   U5128 : OAI22_X1 port map( A1 => n13968, A2 => n13795, B1 => n5627, B2 => 
                           n13794, ZN => n9874);
   U5129 : OAI22_X1 port map( A1 => n13974, A2 => n13795, B1 => n5637, B2 => 
                           n13794, ZN => n9875);
   U5130 : OAI22_X1 port map( A1 => n13980, A2 => n13795, B1 => n5647, B2 => 
                           n13794, ZN => n9876);
   U5131 : OAI22_X1 port map( A1 => n13986, A2 => n13795, B1 => n5657, B2 => 
                           n13794, ZN => n9877);
   U5132 : OAI22_X1 port map( A1 => n13992, A2 => n13795, B1 => n5667, B2 => 
                           n13794, ZN => n9878);
   U5133 : OAI22_X1 port map( A1 => n13998, A2 => n13795, B1 => n5677, B2 => 
                           n13794, ZN => n9879);
   U5134 : OAI22_X1 port map( A1 => n14004, A2 => n13795, B1 => n5687, B2 => 
                           n13794, ZN => n9880);
   U5135 : OAI22_X1 port map( A1 => n14013, A2 => n13795, B1 => n5697, B2 => 
                           n13794, ZN => n9881);
   U5136 : OAI22_X1 port map( A1 => n13969, A2 => n13741, B1 => n5625, B2 => 
                           n13740, ZN => n9586);
   U5137 : OAI22_X1 port map( A1 => n13975, A2 => n13741, B1 => n5635, B2 => 
                           n13740, ZN => n9587);
   U5138 : OAI22_X1 port map( A1 => n13981, A2 => n13741, B1 => n5645, B2 => 
                           n13740, ZN => n9588);
   U5139 : OAI22_X1 port map( A1 => n13987, A2 => n13741, B1 => n5655, B2 => 
                           n13740, ZN => n9589);
   U5140 : OAI22_X1 port map( A1 => n13993, A2 => n13741, B1 => n5665, B2 => 
                           n13740, ZN => n9590);
   U5141 : OAI22_X1 port map( A1 => n13999, A2 => n13741, B1 => n5675, B2 => 
                           n13740, ZN => n9591);
   U5142 : OAI22_X1 port map( A1 => n14005, A2 => n13741, B1 => n5685, B2 => 
                           n13740, ZN => n9592);
   U5143 : OAI22_X1 port map( A1 => n14014, A2 => n13741, B1 => n5695, B2 => 
                           n13740, ZN => n9593);
   U5144 : OAI22_X1 port map( A1 => n13969, A2 => n13693, B1 => n5796, B2 => 
                           n13692, ZN => n9330);
   U5145 : OAI22_X1 port map( A1 => n13975, A2 => n13693, B1 => n5800, B2 => 
                           n13692, ZN => n9331);
   U5146 : OAI22_X1 port map( A1 => n13981, A2 => n13693, B1 => n5804, B2 => 
                           n13692, ZN => n9332);
   U5147 : OAI22_X1 port map( A1 => n13987, A2 => n13693, B1 => n5808, B2 => 
                           n13692, ZN => n9333);
   U5148 : OAI22_X1 port map( A1 => n13993, A2 => n13693, B1 => n5812, B2 => 
                           n13692, ZN => n9334);
   U5149 : OAI22_X1 port map( A1 => n13999, A2 => n13693, B1 => n5816, B2 => 
                           n13692, ZN => n9335);
   U5150 : OAI22_X1 port map( A1 => n14005, A2 => n13693, B1 => n5820, B2 => 
                           n13692, ZN => n9336);
   U5151 : OAI22_X1 port map( A1 => n14014, A2 => n13693, B1 => n5824, B2 => 
                           n13692, ZN => n9337);
   U5152 : OAI22_X1 port map( A1 => n13970, A2 => n13639, B1 => n5622, B2 => 
                           n13638, ZN => n9042);
   U5153 : OAI22_X1 port map( A1 => n13976, A2 => n13639, B1 => n5632, B2 => 
                           n13638, ZN => n9043);
   U5154 : OAI22_X1 port map( A1 => n13982, A2 => n13639, B1 => n5642, B2 => 
                           n13638, ZN => n9044);
   U5155 : OAI22_X1 port map( A1 => n13988, A2 => n13639, B1 => n5652, B2 => 
                           n13638, ZN => n9045);
   U5156 : OAI22_X1 port map( A1 => n13994, A2 => n13639, B1 => n5662, B2 => 
                           n13638, ZN => n9046);
   U5157 : OAI22_X1 port map( A1 => n14000, A2 => n13639, B1 => n5672, B2 => 
                           n13638, ZN => n9047);
   U5159 : OAI22_X1 port map( A1 => n14006, A2 => n13639, B1 => n5682, B2 => 
                           n13638, ZN => n9048);
   U5160 : OAI22_X1 port map( A1 => n14015, A2 => n13639, B1 => n5692, B2 => 
                           n13638, ZN => n9049);
   U5161 : OAI22_X1 port map( A1 => n13971, A2 => n13519, B1 => n976, B2 => 
                           n13518, ZN => n8402);
   U5162 : OAI22_X1 port map( A1 => n13977, A2 => n13519, B1 => n975, B2 => 
                           n13518, ZN => n8403);
   U5163 : OAI22_X1 port map( A1 => n13983, A2 => n13519, B1 => n974, B2 => 
                           n13518, ZN => n8404);
   U5164 : OAI22_X1 port map( A1 => n13989, A2 => n13519, B1 => n973, B2 => 
                           n13518, ZN => n8405);
   U5165 : OAI22_X1 port map( A1 => n13995, A2 => n13519, B1 => n972, B2 => 
                           n13518, ZN => n8406);
   U5166 : OAI22_X1 port map( A1 => n14001, A2 => n13519, B1 => n971, B2 => 
                           n13518, ZN => n8407);
   U5167 : OAI22_X1 port map( A1 => n14007, A2 => n13519, B1 => n970, B2 => 
                           n13518, ZN => n8408);
   U5168 : OAI22_X1 port map( A1 => n14016, A2 => n13519, B1 => n969, B2 => 
                           n13518, ZN => n8409);
   U5169 : OAI22_X1 port map( A1 => n13971, A2 => n13543, B1 => n640, B2 => 
                           n13542, ZN => n8530);
   U5170 : OAI22_X1 port map( A1 => n13977, A2 => n13543, B1 => n637, B2 => 
                           n13542, ZN => n8531);
   U5171 : OAI22_X1 port map( A1 => n13983, A2 => n13543, B1 => n634, B2 => 
                           n13542, ZN => n8532);
   U5172 : OAI22_X1 port map( A1 => n13989, A2 => n13543, B1 => n631, B2 => 
                           n13542, ZN => n8533);
   U5173 : OAI22_X1 port map( A1 => n13995, A2 => n13543, B1 => n628, B2 => 
                           n13542, ZN => n8534);
   U5174 : OAI22_X1 port map( A1 => n14001, A2 => n13543, B1 => n625, B2 => 
                           n13542, ZN => n8535);
   U5175 : OAI22_X1 port map( A1 => n14007, A2 => n13543, B1 => n622, B2 => 
                           n13542, ZN => n8536);
   U5176 : OAI22_X1 port map( A1 => n13968, A2 => n13789, B1 => n816, B2 => 
                           n13788, ZN => n9842);
   U5177 : OAI22_X1 port map( A1 => n13974, A2 => n13789, B1 => n815, B2 => 
                           n13788, ZN => n9843);
   U5178 : OAI22_X1 port map( A1 => n13980, A2 => n13789, B1 => n814, B2 => 
                           n13788, ZN => n9844);
   U5179 : OAI22_X1 port map( A1 => n13986, A2 => n13789, B1 => n813, B2 => 
                           n13788, ZN => n9845);
   U5180 : OAI22_X1 port map( A1 => n13992, A2 => n13789, B1 => n812, B2 => 
                           n13788, ZN => n9846);
   U5181 : OAI22_X1 port map( A1 => n13998, A2 => n13789, B1 => n811, B2 => 
                           n13788, ZN => n9847);
   U5182 : OAI22_X1 port map( A1 => n14004, A2 => n13789, B1 => n810, B2 => 
                           n13788, ZN => n9848);
   U5183 : OAI22_X1 port map( A1 => n14013, A2 => n13789, B1 => n809, B2 => 
                           n13788, ZN => n9849);
   U5184 : OAI22_X1 port map( A1 => n13969, A2 => n13735, B1 => n848, B2 => 
                           n13734, ZN => n9554);
   U5185 : OAI22_X1 port map( A1 => n13975, A2 => n13735, B1 => n847, B2 => 
                           n13734, ZN => n9555);
   U5186 : OAI22_X1 port map( A1 => n13981, A2 => n13735, B1 => n846, B2 => 
                           n13734, ZN => n9556);
   U5187 : OAI22_X1 port map( A1 => n13987, A2 => n13735, B1 => n845, B2 => 
                           n13734, ZN => n9557);
   U5188 : OAI22_X1 port map( A1 => n13993, A2 => n13735, B1 => n844, B2 => 
                           n13734, ZN => n9558);
   U5189 : OAI22_X1 port map( A1 => n13999, A2 => n13735, B1 => n843, B2 => 
                           n13734, ZN => n9559);
   U5190 : OAI22_X1 port map( A1 => n14005, A2 => n13735, B1 => n842, B2 => 
                           n13734, ZN => n9560);
   U5191 : OAI22_X1 port map( A1 => n14014, A2 => n13735, B1 => n841, B2 => 
                           n13734, ZN => n9561);
   U5192 : OAI22_X1 port map( A1 => n13969, A2 => n13681, B1 => n880, B2 => 
                           n13680, ZN => n9266);
   U5193 : OAI22_X1 port map( A1 => n13975, A2 => n13681, B1 => n879, B2 => 
                           n13680, ZN => n9267);
   U5194 : OAI22_X1 port map( A1 => n13981, A2 => n13681, B1 => n878, B2 => 
                           n13680, ZN => n9268);
   U5195 : OAI22_X1 port map( A1 => n13987, A2 => n13681, B1 => n877, B2 => 
                           n13680, ZN => n9269);
   U5196 : OAI22_X1 port map( A1 => n13993, A2 => n13681, B1 => n876, B2 => 
                           n13680, ZN => n9270);
   U5197 : OAI22_X1 port map( A1 => n13999, A2 => n13681, B1 => n875, B2 => 
                           n13680, ZN => n9271);
   U5198 : OAI22_X1 port map( A1 => n14005, A2 => n13681, B1 => n874, B2 => 
                           n13680, ZN => n9272);
   U5199 : OAI22_X1 port map( A1 => n14014, A2 => n13681, B1 => n873, B2 => 
                           n13680, ZN => n9273);
   U5200 : OAI22_X1 port map( A1 => n13970, A2 => n13633, B1 => n5623, B2 => 
                           n13632, ZN => n9010);
   U5201 : OAI22_X1 port map( A1 => n13976, A2 => n13633, B1 => n5633, B2 => 
                           n13632, ZN => n9011);
   U5202 : OAI22_X1 port map( A1 => n13982, A2 => n13633, B1 => n5643, B2 => 
                           n13632, ZN => n9012);
   U5203 : OAI22_X1 port map( A1 => n13988, A2 => n13633, B1 => n5653, B2 => 
                           n13632, ZN => n9013);
   U5204 : OAI22_X1 port map( A1 => n13994, A2 => n13633, B1 => n5663, B2 => 
                           n13632, ZN => n9014);
   U5205 : OAI22_X1 port map( A1 => n14000, A2 => n13633, B1 => n5673, B2 => 
                           n13632, ZN => n9015);
   U5206 : OAI22_X1 port map( A1 => n14006, A2 => n13633, B1 => n5683, B2 => 
                           n13632, ZN => n9016);
   U5207 : OAI22_X1 port map( A1 => n14015, A2 => n13633, B1 => n5693, B2 => 
                           n13632, ZN => n9017);
   U5208 : OAI22_X1 port map( A1 => n13970, A2 => n13627, B1 => n912, B2 => 
                           n13626, ZN => n8978);
   U5209 : OAI22_X1 port map( A1 => n13976, A2 => n13627, B1 => n911, B2 => 
                           n13626, ZN => n8979);
   U5210 : OAI22_X1 port map( A1 => n13982, A2 => n13627, B1 => n910, B2 => 
                           n13626, ZN => n8980);
   U5211 : OAI22_X1 port map( A1 => n13988, A2 => n13627, B1 => n909, B2 => 
                           n13626, ZN => n8981);
   U5212 : OAI22_X1 port map( A1 => n13994, A2 => n13627, B1 => n908, B2 => 
                           n13626, ZN => n8982);
   U5213 : OAI22_X1 port map( A1 => n14000, A2 => n13627, B1 => n907, B2 => 
                           n13626, ZN => n8983);
   U5214 : OAI22_X1 port map( A1 => n14006, A2 => n13627, B1 => n906, B2 => 
                           n13626, ZN => n8984);
   U5215 : OAI22_X1 port map( A1 => n14015, A2 => n13627, B1 => n905, B2 => 
                           n13626, ZN => n8985);
   U5216 : OAI22_X1 port map( A1 => n13971, A2 => n13573, B1 => n944, B2 => 
                           n13572, ZN => n8690);
   U5217 : OAI22_X1 port map( A1 => n13977, A2 => n13573, B1 => n943, B2 => 
                           n13572, ZN => n8691);
   U5218 : OAI22_X1 port map( A1 => n13983, A2 => n13573, B1 => n942, B2 => 
                           n13572, ZN => n8692);
   U5219 : OAI22_X1 port map( A1 => n13989, A2 => n13573, B1 => n941, B2 => 
                           n13572, ZN => n8693);
   U5220 : OAI22_X1 port map( A1 => n13995, A2 => n13573, B1 => n940, B2 => 
                           n13572, ZN => n8694);
   U5221 : OAI22_X1 port map( A1 => n14001, A2 => n13573, B1 => n939, B2 => 
                           n13572, ZN => n8695);
   U5222 : OAI22_X1 port map( A1 => n14007, A2 => n13573, B1 => n938, B2 => 
                           n13572, ZN => n8696);
   U5223 : OAI22_X1 port map( A1 => n14016, A2 => n13573, B1 => n937, B2 => 
                           n13572, ZN => n8697);
   U5224 : OAI22_X1 port map( A1 => n13972, A2 => n13465, B1 => n7248, B2 => 
                           n13464, ZN => n8114);
   U5225 : OAI22_X1 port map( A1 => n13978, A2 => n13465, B1 => n7249, B2 => 
                           n13464, ZN => n8115);
   U5226 : OAI22_X1 port map( A1 => n13984, A2 => n13465, B1 => n7250, B2 => 
                           n13464, ZN => n8116);
   U5227 : OAI22_X1 port map( A1 => n13990, A2 => n13465, B1 => n7251, B2 => 
                           n13464, ZN => n8117);
   U5228 : OAI22_X1 port map( A1 => n13996, A2 => n13465, B1 => n7252, B2 => 
                           n13464, ZN => n8118);
   U5229 : OAI22_X1 port map( A1 => n14002, A2 => n13465, B1 => n7253, B2 => 
                           n13464, ZN => n8119);
   U5230 : OAI22_X1 port map( A1 => n14008, A2 => n13465, B1 => n7254, B2 => 
                           n13464, ZN => n8120);
   U5231 : OAI22_X1 port map( A1 => n14017, A2 => n13465, B1 => n7255, B2 => 
                           n13464, ZN => n8121);
   U5232 : OAI22_X1 port map( A1 => n13972, A2 => n13513, B1 => n6974, B2 => 
                           n13512, ZN => n8370);
   U5233 : OAI22_X1 port map( A1 => n13978, A2 => n13513, B1 => n6975, B2 => 
                           n13512, ZN => n8371);
   U5234 : OAI22_X1 port map( A1 => n13984, A2 => n13513, B1 => n6976, B2 => 
                           n13512, ZN => n8372);
   U5235 : OAI22_X1 port map( A1 => n13990, A2 => n13513, B1 => n6977, B2 => 
                           n13512, ZN => n8373);
   U5236 : OAI22_X1 port map( A1 => n13996, A2 => n13513, B1 => n6978, B2 => 
                           n13512, ZN => n8374);
   U5237 : OAI22_X1 port map( A1 => n14002, A2 => n13513, B1 => n6979, B2 => 
                           n13512, ZN => n8375);
   U5238 : OAI22_X1 port map( A1 => n14008, A2 => n13513, B1 => n6980, B2 => 
                           n13512, ZN => n8376);
   U5239 : OAI22_X1 port map( A1 => n14017, A2 => n13513, B1 => n6981, B2 => 
                           n13512, ZN => n8377);
   U5240 : OAI22_X1 port map( A1 => n14016, A2 => n13543, B1 => n7257, B2 => 
                           n13542, ZN => n8537);
   U5241 : OAI22_X1 port map( A1 => n13970, A2 => n13621, B1 => n6982, B2 => 
                           n13620, ZN => n8946);
   U5242 : OAI22_X1 port map( A1 => n13976, A2 => n13621, B1 => n6983, B2 => 
                           n13620, ZN => n8947);
   U5243 : OAI22_X1 port map( A1 => n13982, A2 => n13621, B1 => n6984, B2 => 
                           n13620, ZN => n8948);
   U5244 : OAI22_X1 port map( A1 => n13988, A2 => n13621, B1 => n6985, B2 => 
                           n13620, ZN => n8949);
   U5245 : OAI22_X1 port map( A1 => n13994, A2 => n13621, B1 => n6986, B2 => 
                           n13620, ZN => n8950);
   U5246 : OAI22_X1 port map( A1 => n14000, A2 => n13621, B1 => n6987, B2 => 
                           n13620, ZN => n8951);
   U5247 : OAI22_X1 port map( A1 => n14006, A2 => n13621, B1 => n6988, B2 => 
                           n13620, ZN => n8952);
   U5248 : OAI22_X1 port map( A1 => n14015, A2 => n13621, B1 => n6989, B2 => 
                           n13620, ZN => n8953);
   U5249 : OAI22_X1 port map( A1 => n13969, A2 => n13675, B1 => n6990, B2 => 
                           n13674, ZN => n9234);
   U5250 : OAI22_X1 port map( A1 => n13975, A2 => n13675, B1 => n6991, B2 => 
                           n13674, ZN => n9235);
   U5251 : OAI22_X1 port map( A1 => n13981, A2 => n13675, B1 => n6992, B2 => 
                           n13674, ZN => n9236);
   U5253 : OAI22_X1 port map( A1 => n13987, A2 => n13675, B1 => n6993, B2 => 
                           n13674, ZN => n9237);
   U5254 : OAI22_X1 port map( A1 => n13993, A2 => n13675, B1 => n6994, B2 => 
                           n13674, ZN => n9238);
   U5255 : OAI22_X1 port map( A1 => n13999, A2 => n13675, B1 => n6995, B2 => 
                           n13674, ZN => n9239);
   U5256 : OAI22_X1 port map( A1 => n14005, A2 => n13675, B1 => n6996, B2 => 
                           n13674, ZN => n9240);
   U5257 : OAI22_X1 port map( A1 => n14014, A2 => n13675, B1 => n6997, B2 => 
                           n13674, ZN => n9241);
   U5258 : OAI22_X1 port map( A1 => n13969, A2 => n13729, B1 => n7006, B2 => 
                           n13728, ZN => n9522);
   U5259 : OAI22_X1 port map( A1 => n13975, A2 => n13729, B1 => n7007, B2 => 
                           n13728, ZN => n9523);
   U5260 : OAI22_X1 port map( A1 => n13981, A2 => n13729, B1 => n7008, B2 => 
                           n13728, ZN => n9524);
   U5261 : OAI22_X1 port map( A1 => n13987, A2 => n13729, B1 => n7009, B2 => 
                           n13728, ZN => n9525);
   U5262 : OAI22_X1 port map( A1 => n13993, A2 => n13729, B1 => n7010, B2 => 
                           n13728, ZN => n9526);
   U5263 : OAI22_X1 port map( A1 => n13999, A2 => n13729, B1 => n7011, B2 => 
                           n13728, ZN => n9527);
   U5264 : OAI22_X1 port map( A1 => n14005, A2 => n13729, B1 => n7012, B2 => 
                           n13728, ZN => n9528);
   U5265 : OAI22_X1 port map( A1 => n14014, A2 => n13729, B1 => n7013, B2 => 
                           n13728, ZN => n9529);
   U5266 : OAI22_X1 port map( A1 => n13969, A2 => n13753, B1 => n6786, B2 => 
                           n13752, ZN => n9650);
   U5267 : OAI22_X1 port map( A1 => n13975, A2 => n13753, B1 => n6787, B2 => 
                           n13752, ZN => n9651);
   U5268 : OAI22_X1 port map( A1 => n13981, A2 => n13753, B1 => n6788, B2 => 
                           n13752, ZN => n9652);
   U5269 : OAI22_X1 port map( A1 => n13987, A2 => n13753, B1 => n6789, B2 => 
                           n13752, ZN => n9653);
   U5270 : OAI22_X1 port map( A1 => n13993, A2 => n13753, B1 => n6790, B2 => 
                           n13752, ZN => n9654);
   U5271 : OAI22_X1 port map( A1 => n13999, A2 => n13753, B1 => n6791, B2 => 
                           n13752, ZN => n9655);
   U5272 : OAI22_X1 port map( A1 => n14005, A2 => n13753, B1 => n6792, B2 => 
                           n13752, ZN => n9656);
   U5273 : OAI22_X1 port map( A1 => n14014, A2 => n13753, B1 => n6793, B2 => 
                           n13752, ZN => n9657);
   U5274 : OAI22_X1 port map( A1 => n13968, A2 => n13759, B1 => n6914, B2 => 
                           n13758, ZN => n9682);
   U5275 : OAI22_X1 port map( A1 => n13974, A2 => n13759, B1 => n6915, B2 => 
                           n13758, ZN => n9683);
   U5276 : OAI22_X1 port map( A1 => n13980, A2 => n13759, B1 => n6916, B2 => 
                           n13758, ZN => n9684);
   U5277 : OAI22_X1 port map( A1 => n13986, A2 => n13759, B1 => n6917, B2 => 
                           n13758, ZN => n9685);
   U5278 : OAI22_X1 port map( A1 => n13992, A2 => n13759, B1 => n6918, B2 => 
                           n13758, ZN => n9686);
   U5279 : OAI22_X1 port map( A1 => n13998, A2 => n13759, B1 => n6919, B2 => 
                           n13758, ZN => n9687);
   U5280 : OAI22_X1 port map( A1 => n14004, A2 => n13759, B1 => n6920, B2 => 
                           n13758, ZN => n9688);
   U5281 : OAI22_X1 port map( A1 => n14013, A2 => n13759, B1 => n6921, B2 => 
                           n13758, ZN => n9689);
   U5282 : OAI22_X1 port map( A1 => n13968, A2 => n13783, B1 => n7014, B2 => 
                           n13782, ZN => n9810);
   U5283 : OAI22_X1 port map( A1 => n13974, A2 => n13783, B1 => n7015, B2 => 
                           n13782, ZN => n9811);
   U5284 : OAI22_X1 port map( A1 => n13980, A2 => n13783, B1 => n7016, B2 => 
                           n13782, ZN => n9812);
   U5285 : OAI22_X1 port map( A1 => n13986, A2 => n13783, B1 => n7017, B2 => 
                           n13782, ZN => n9813);
   U5286 : OAI22_X1 port map( A1 => n13992, A2 => n13783, B1 => n7018, B2 => 
                           n13782, ZN => n9814);
   U5287 : OAI22_X1 port map( A1 => n13998, A2 => n13783, B1 => n7019, B2 => 
                           n13782, ZN => n9815);
   U5288 : OAI22_X1 port map( A1 => n14004, A2 => n13783, B1 => n7020, B2 => 
                           n13782, ZN => n9816);
   U5289 : OAI22_X1 port map( A1 => n14013, A2 => n13783, B1 => n7021, B2 => 
                           n13782, ZN => n9817);
   U5290 : OAI22_X1 port map( A1 => n13968, A2 => n13807, B1 => n6802, B2 => 
                           n13806, ZN => n9938);
   U5291 : OAI22_X1 port map( A1 => n13974, A2 => n13807, B1 => n6803, B2 => 
                           n13806, ZN => n9939);
   U5292 : OAI22_X1 port map( A1 => n13980, A2 => n13807, B1 => n6804, B2 => 
                           n13806, ZN => n9940);
   U5293 : OAI22_X1 port map( A1 => n13986, A2 => n13807, B1 => n6805, B2 => 
                           n13806, ZN => n9941);
   U5294 : OAI22_X1 port map( A1 => n13992, A2 => n13807, B1 => n6806, B2 => 
                           n13806, ZN => n9942);
   U5295 : OAI22_X1 port map( A1 => n13998, A2 => n13807, B1 => n6807, B2 => 
                           n13806, ZN => n9943);
   U5296 : OAI22_X1 port map( A1 => n14004, A2 => n13807, B1 => n6808, B2 => 
                           n13806, ZN => n9944);
   U5297 : OAI22_X1 port map( A1 => n14013, A2 => n13807, B1 => n6809, B2 => 
                           n13806, ZN => n9945);
   U5298 : OAI22_X1 port map( A1 => n13971, A2 => n13579, B1 => n5795, B2 => 
                           n13578, ZN => n8722);
   U5299 : OAI22_X1 port map( A1 => n13977, A2 => n13579, B1 => n5799, B2 => 
                           n13578, ZN => n8723);
   U5300 : OAI22_X1 port map( A1 => n13983, A2 => n13579, B1 => n5803, B2 => 
                           n13578, ZN => n8724);
   U5301 : OAI22_X1 port map( A1 => n13989, A2 => n13579, B1 => n5807, B2 => 
                           n13578, ZN => n8725);
   U5302 : OAI22_X1 port map( A1 => n13995, A2 => n13579, B1 => n5811, B2 => 
                           n13578, ZN => n8726);
   U5303 : OAI22_X1 port map( A1 => n14001, A2 => n13579, B1 => n5815, B2 => 
                           n13578, ZN => n8727);
   U5304 : OAI22_X1 port map( A1 => n14007, A2 => n13579, B1 => n5819, B2 => 
                           n13578, ZN => n8728);
   U5305 : OAI22_X1 port map( A1 => n13969, A2 => n13687, B1 => n5797, B2 => 
                           n13686, ZN => n9298);
   U5306 : OAI22_X1 port map( A1 => n13975, A2 => n13687, B1 => n5801, B2 => 
                           n13686, ZN => n9299);
   U5307 : OAI22_X1 port map( A1 => n13981, A2 => n13687, B1 => n5805, B2 => 
                           n13686, ZN => n9300);
   U5308 : OAI22_X1 port map( A1 => n13987, A2 => n13687, B1 => n5809, B2 => 
                           n13686, ZN => n9301);
   U5309 : OAI22_X1 port map( A1 => n13993, A2 => n13687, B1 => n5813, B2 => 
                           n13686, ZN => n9302);
   U5310 : OAI22_X1 port map( A1 => n13999, A2 => n13687, B1 => n5817, B2 => 
                           n13686, ZN => n9303);
   U5311 : OAI22_X1 port map( A1 => n14020, A2 => n13896, B1 => n675, B2 => 
                           n14011, ZN => n9958);
   U5312 : OAI22_X1 port map( A1 => n14020, A2 => n13902, B1 => n672, B2 => 
                           n14011, ZN => n9959);
   U5313 : OAI22_X1 port map( A1 => n14020, A2 => n13908, B1 => n669, B2 => 
                           n14011, ZN => n9960);
   U5314 : OAI22_X1 port map( A1 => n14020, A2 => n13914, B1 => n666, B2 => 
                           n14011, ZN => n9961);
   U5315 : OAI22_X1 port map( A1 => n13896, A2 => n13760, B1 => n674, B2 => 
                           n13757, ZN => n9670);
   U5316 : OAI22_X1 port map( A1 => n13902, A2 => n13760, B1 => n671, B2 => 
                           n13757, ZN => n9671);
   U5317 : OAI22_X1 port map( A1 => n13908, A2 => n13760, B1 => n668, B2 => 
                           n13757, ZN => n9672);
   U5318 : OAI22_X1 port map( A1 => n13914, A2 => n13760, B1 => n665, B2 => 
                           n13757, ZN => n9673);
   U5319 : OAI22_X1 port map( A1 => n13920, A2 => n13760, B1 => n662, B2 => 
                           n13757, ZN => n9674);
   U5320 : OAI22_X1 port map( A1 => n13926, A2 => n13760, B1 => n659, B2 => 
                           n13757, ZN => n9675);
   U5321 : OAI22_X1 port map( A1 => n13932, A2 => n13760, B1 => n656, B2 => 
                           n13757, ZN => n9676);
   U5322 : OAI22_X1 port map( A1 => n13938, A2 => n13760, B1 => n653, B2 => 
                           n13757, ZN => n9677);
   U5323 : OAI22_X1 port map( A1 => n14021, A2 => n13824, B1 => n711, B2 => 
                           n14010, ZN => n9946);
   U5324 : OAI22_X1 port map( A1 => n14021, A2 => n13830, B1 => n708, B2 => 
                           n14010, ZN => n9947);
   U5325 : OAI22_X1 port map( A1 => n14021, A2 => n13836, B1 => n705, B2 => 
                           n14010, ZN => n9948);
   U5326 : OAI22_X1 port map( A1 => n14021, A2 => n13842, B1 => n702, B2 => 
                           n14010, ZN => n9949);
   U5327 : OAI22_X1 port map( A1 => n14021, A2 => n13848, B1 => n699, B2 => 
                           n14010, ZN => n9950);
   U5328 : OAI22_X1 port map( A1 => n14021, A2 => n13854, B1 => n696, B2 => 
                           n14010, ZN => n9951);
   U5329 : OAI22_X1 port map( A1 => n14021, A2 => n13860, B1 => n693, B2 => 
                           n14010, ZN => n9952);
   U5330 : OAI22_X1 port map( A1 => n14021, A2 => n13866, B1 => n690, B2 => 
                           n14010, ZN => n9953);
   U5331 : OAI22_X1 port map( A1 => n14020, A2 => n13872, B1 => n687, B2 => 
                           n14010, ZN => n9954);
   U5332 : OAI22_X1 port map( A1 => n14020, A2 => n13878, B1 => n684, B2 => 
                           n14010, ZN => n9955);
   U5333 : OAI22_X1 port map( A1 => n14020, A2 => n13884, B1 => n681, B2 => 
                           n14010, ZN => n9956);
   U5334 : OAI22_X1 port map( A1 => n14020, A2 => n13890, B1 => n678, B2 => 
                           n14010, ZN => n9957);
   U5335 : OAI22_X1 port map( A1 => n13824, A2 => n13797, B1 => n5387, B2 => 
                           n13792, ZN => n9850);
   U5336 : OAI22_X1 port map( A1 => n13830, A2 => n13797, B1 => n5397, B2 => 
                           n13792, ZN => n9851);
   U5337 : OAI22_X1 port map( A1 => n13836, A2 => n13797, B1 => n5407, B2 => 
                           n13792, ZN => n9852);
   U5338 : OAI22_X1 port map( A1 => n13842, A2 => n13797, B1 => n5417, B2 => 
                           n13792, ZN => n9853);
   U5339 : OAI22_X1 port map( A1 => n13848, A2 => n13797, B1 => n5427, B2 => 
                           n13792, ZN => n9854);
   U5340 : OAI22_X1 port map( A1 => n13854, A2 => n13797, B1 => n5437, B2 => 
                           n13792, ZN => n9855);
   U5341 : OAI22_X1 port map( A1 => n13860, A2 => n13797, B1 => n5447, B2 => 
                           n13792, ZN => n9856);
   U5342 : OAI22_X1 port map( A1 => n13866, A2 => n13797, B1 => n5457, B2 => 
                           n13792, ZN => n9857);
   U5343 : OAI22_X1 port map( A1 => n13872, A2 => n13796, B1 => n5467, B2 => 
                           n13792, ZN => n9858);
   U5344 : OAI22_X1 port map( A1 => n13878, A2 => n13796, B1 => n5477, B2 => 
                           n13792, ZN => n9859);
   U5345 : OAI22_X1 port map( A1 => n13884, A2 => n13796, B1 => n5487, B2 => 
                           n13792, ZN => n9860);
   U5346 : OAI22_X1 port map( A1 => n13890, A2 => n13796, B1 => n5497, B2 => 
                           n13792, ZN => n9861);
   U5347 : OAI22_X1 port map( A1 => n13896, A2 => n13796, B1 => n5507, B2 => 
                           n13793, ZN => n9862);
   U5348 : OAI22_X1 port map( A1 => n13902, A2 => n13796, B1 => n5517, B2 => 
                           n13793, ZN => n9863);
   U5349 : OAI22_X1 port map( A1 => n13908, A2 => n13796, B1 => n5527, B2 => 
                           n13793, ZN => n9864);
   U5350 : OAI22_X1 port map( A1 => n13914, A2 => n13796, B1 => n5537, B2 => 
                           n13793, ZN => n9865);
   U5351 : OAI22_X1 port map( A1 => n13920, A2 => n13796, B1 => n5547, B2 => 
                           n13793, ZN => n9866);
   U5352 : OAI22_X1 port map( A1 => n13926, A2 => n13796, B1 => n5557, B2 => 
                           n13793, ZN => n9867);
   U5353 : OAI22_X1 port map( A1 => n13932, A2 => n13796, B1 => n5567, B2 => 
                           n13793, ZN => n9868);
   U5354 : OAI22_X1 port map( A1 => n13938, A2 => n13796, B1 => n5577, B2 => 
                           n13793, ZN => n9869);
   U5355 : OAI22_X1 port map( A1 => n13944, A2 => n13795, B1 => n5587, B2 => 
                           n13793, ZN => n9870);
   U5356 : OAI22_X1 port map( A1 => n13950, A2 => n13795, B1 => n5597, B2 => 
                           n13793, ZN => n9871);
   U5357 : OAI22_X1 port map( A1 => n13956, A2 => n13795, B1 => n5607, B2 => 
                           n13793, ZN => n9872);
   U5358 : OAI22_X1 port map( A1 => n13962, A2 => n13795, B1 => n5617, B2 => 
                           n13793, ZN => n9873);
   U5359 : OAI22_X1 port map( A1 => n13824, A2 => n13761, B1 => n710, B2 => 
                           n13756, ZN => n9658);
   U5360 : OAI22_X1 port map( A1 => n13830, A2 => n13761, B1 => n707, B2 => 
                           n13756, ZN => n9659);
   U5361 : OAI22_X1 port map( A1 => n13836, A2 => n13761, B1 => n704, B2 => 
                           n13756, ZN => n9660);
   U5362 : OAI22_X1 port map( A1 => n13842, A2 => n13761, B1 => n701, B2 => 
                           n13756, ZN => n9661);
   U5363 : OAI22_X1 port map( A1 => n13848, A2 => n13761, B1 => n698, B2 => 
                           n13756, ZN => n9662);
   U5364 : OAI22_X1 port map( A1 => n13854, A2 => n13761, B1 => n695, B2 => 
                           n13756, ZN => n9663);
   U5365 : OAI22_X1 port map( A1 => n13860, A2 => n13761, B1 => n692, B2 => 
                           n13756, ZN => n9664);
   U5366 : OAI22_X1 port map( A1 => n13866, A2 => n13761, B1 => n689, B2 => 
                           n13756, ZN => n9665);
   U5367 : OAI22_X1 port map( A1 => n13872, A2 => n13760, B1 => n686, B2 => 
                           n13756, ZN => n9666);
   U5368 : OAI22_X1 port map( A1 => n13878, A2 => n13760, B1 => n683, B2 => 
                           n13756, ZN => n9667);
   U5369 : OAI22_X1 port map( A1 => n13884, A2 => n13760, B1 => n680, B2 => 
                           n13756, ZN => n9668);
   U5370 : OAI22_X1 port map( A1 => n13890, A2 => n13760, B1 => n677, B2 => 
                           n13756, ZN => n9669);
   U5371 : OAI22_X1 port map( A1 => n13824, A2 => n13743, B1 => n5385, B2 => 
                           n13738, ZN => n9562);
   U5372 : OAI22_X1 port map( A1 => n13831, A2 => n13743, B1 => n5395, B2 => 
                           n13738, ZN => n9563);
   U5373 : OAI22_X1 port map( A1 => n13837, A2 => n13743, B1 => n5405, B2 => 
                           n13738, ZN => n9564);
   U5374 : OAI22_X1 port map( A1 => n13843, A2 => n13743, B1 => n5415, B2 => 
                           n13738, ZN => n9565);
   U5375 : OAI22_X1 port map( A1 => n13849, A2 => n13743, B1 => n5425, B2 => 
                           n13738, ZN => n9566);
   U5376 : OAI22_X1 port map( A1 => n13855, A2 => n13743, B1 => n5435, B2 => 
                           n13738, ZN => n9567);
   U5377 : OAI22_X1 port map( A1 => n13861, A2 => n13743, B1 => n5445, B2 => 
                           n13738, ZN => n9568);
   U5378 : OAI22_X1 port map( A1 => n13867, A2 => n13743, B1 => n5455, B2 => 
                           n13738, ZN => n9569);
   U5379 : OAI22_X1 port map( A1 => n13873, A2 => n13742, B1 => n5465, B2 => 
                           n13738, ZN => n9570);
   U5380 : OAI22_X1 port map( A1 => n13879, A2 => n13742, B1 => n5475, B2 => 
                           n13738, ZN => n9571);
   U5381 : OAI22_X1 port map( A1 => n13885, A2 => n13742, B1 => n5485, B2 => 
                           n13738, ZN => n9572);
   U5382 : OAI22_X1 port map( A1 => n13891, A2 => n13742, B1 => n5495, B2 => 
                           n13738, ZN => n9573);
   U5383 : OAI22_X1 port map( A1 => n13897, A2 => n13742, B1 => n5505, B2 => 
                           n13739, ZN => n9574);
   U5384 : OAI22_X1 port map( A1 => n13903, A2 => n13742, B1 => n5515, B2 => 
                           n13739, ZN => n9575);
   U5385 : OAI22_X1 port map( A1 => n13909, A2 => n13742, B1 => n5525, B2 => 
                           n13739, ZN => n9576);
   U5386 : OAI22_X1 port map( A1 => n13915, A2 => n13742, B1 => n5535, B2 => 
                           n13739, ZN => n9577);
   U5387 : OAI22_X1 port map( A1 => n13921, A2 => n13742, B1 => n5545, B2 => 
                           n13739, ZN => n9578);
   U5388 : OAI22_X1 port map( A1 => n13927, A2 => n13742, B1 => n5555, B2 => 
                           n13739, ZN => n9579);
   U5389 : OAI22_X1 port map( A1 => n13933, A2 => n13742, B1 => n5565, B2 => 
                           n13739, ZN => n9580);
   U5390 : OAI22_X1 port map( A1 => n13939, A2 => n13742, B1 => n5575, B2 => 
                           n13739, ZN => n9581);
   U5391 : OAI22_X1 port map( A1 => n13945, A2 => n13741, B1 => n5585, B2 => 
                           n13739, ZN => n9582);
   U5392 : OAI22_X1 port map( A1 => n13951, A2 => n13741, B1 => n5595, B2 => 
                           n13739, ZN => n9583);
   U5393 : OAI22_X1 port map( A1 => n13957, A2 => n13741, B1 => n5605, B2 => 
                           n13739, ZN => n9584);
   U5394 : OAI22_X1 port map( A1 => n13963, A2 => n13741, B1 => n5615, B2 => 
                           n13739, ZN => n9585);
   U5395 : OAI22_X1 port map( A1 => n13944, A2 => n13759, B1 => n6938, B2 => 
                           n13757, ZN => n9678);
   U5396 : OAI22_X1 port map( A1 => n13950, A2 => n13759, B1 => n6939, B2 => 
                           n13757, ZN => n9679);
   U5397 : OAI22_X1 port map( A1 => n13956, A2 => n13759, B1 => n6940, B2 => 
                           n13757, ZN => n9680);
   U5398 : OAI22_X1 port map( A1 => n13962, A2 => n13759, B1 => n6941, B2 => 
                           n13757, ZN => n9681);
   U5399 : OAI22_X1 port map( A1 => n14020, A2 => n13920, B1 => n6922, B2 => 
                           n14011, ZN => n9962);
   U5400 : OAI22_X1 port map( A1 => n14020, A2 => n13926, B1 => n6923, B2 => 
                           n14011, ZN => n9963);
   U5401 : OAI22_X1 port map( A1 => n14020, A2 => n13932, B1 => n6924, B2 => 
                           n14011, ZN => n9964);
   U5402 : OAI22_X1 port map( A1 => n14020, A2 => n13938, B1 => n6925, B2 => 
                           n14011, ZN => n9965);
   U5403 : OAI22_X1 port map( A1 => n14019, A2 => n13944, B1 => n6926, B2 => 
                           n14011, ZN => n9966);
   U5404 : OAI22_X1 port map( A1 => n14019, A2 => n13950, B1 => n6927, B2 => 
                           n14011, ZN => n9967);
   U5405 : OAI22_X1 port map( A1 => n14019, A2 => n13956, B1 => n6928, B2 => 
                           n14011, ZN => n9968);
   U5406 : OAI22_X1 port map( A1 => n14019, A2 => n13962, B1 => n6929, B2 => 
                           n14011, ZN => n9969);
   U5407 : OAI22_X1 port map( A1 => n13824, A2 => n13755, B1 => n6870, B2 => 
                           n13750, ZN => n9626);
   U5408 : OAI22_X1 port map( A1 => n13831, A2 => n13755, B1 => n6871, B2 => 
                           n13750, ZN => n9627);
   U5409 : OAI22_X1 port map( A1 => n13837, A2 => n13755, B1 => n6872, B2 => 
                           n13750, ZN => n9628);
   U5410 : OAI22_X1 port map( A1 => n13843, A2 => n13755, B1 => n6873, B2 => 
                           n13750, ZN => n9629);
   U5411 : OAI22_X1 port map( A1 => n13849, A2 => n13755, B1 => n6874, B2 => 
                           n13750, ZN => n9630);
   U5412 : OAI22_X1 port map( A1 => n13855, A2 => n13755, B1 => n6875, B2 => 
                           n13750, ZN => n9631);
   U5413 : OAI22_X1 port map( A1 => n13861, A2 => n13755, B1 => n6876, B2 => 
                           n13750, ZN => n9632);
   U5414 : OAI22_X1 port map( A1 => n13867, A2 => n13755, B1 => n6877, B2 => 
                           n13750, ZN => n9633);
   U5415 : OAI22_X1 port map( A1 => n13873, A2 => n13754, B1 => n6878, B2 => 
                           n13750, ZN => n9634);
   U5416 : OAI22_X1 port map( A1 => n13879, A2 => n13754, B1 => n6879, B2 => 
                           n13750, ZN => n9635);
   U5417 : OAI22_X1 port map( A1 => n13885, A2 => n13754, B1 => n6880, B2 => 
                           n13750, ZN => n9636);
   U5418 : OAI22_X1 port map( A1 => n13891, A2 => n13754, B1 => n6881, B2 => 
                           n13750, ZN => n9637);
   U5419 : OAI22_X1 port map( A1 => n13897, A2 => n13754, B1 => n6882, B2 => 
                           n13751, ZN => n9638);
   U5420 : OAI22_X1 port map( A1 => n13903, A2 => n13754, B1 => n6884, B2 => 
                           n13751, ZN => n9639);
   U5421 : OAI22_X1 port map( A1 => n13909, A2 => n13754, B1 => n6886, B2 => 
                           n13751, ZN => n9640);
   U5422 : OAI22_X1 port map( A1 => n13915, A2 => n13754, B1 => n6888, B2 => 
                           n13751, ZN => n9641);
   U5423 : OAI22_X1 port map( A1 => n13921, A2 => n13754, B1 => n6890, B2 => 
                           n13751, ZN => n9642);
   U5424 : OAI22_X1 port map( A1 => n13927, A2 => n13754, B1 => n6891, B2 => 
                           n13751, ZN => n9643);
   U5425 : OAI22_X1 port map( A1 => n13933, A2 => n13754, B1 => n6892, B2 => 
                           n13751, ZN => n9644);
   U5426 : OAI22_X1 port map( A1 => n13939, A2 => n13754, B1 => n6893, B2 => 
                           n13751, ZN => n9645);
   U5427 : OAI22_X1 port map( A1 => n13945, A2 => n13753, B1 => n6810, B2 => 
                           n13751, ZN => n9646);
   U5428 : OAI22_X1 port map( A1 => n13951, A2 => n13753, B1 => n6811, B2 => 
                           n13751, ZN => n9647);
   U5429 : OAI22_X1 port map( A1 => n13957, A2 => n13753, B1 => n6812, B2 => 
                           n13751, ZN => n9648);
   U5430 : OAI22_X1 port map( A1 => n13963, A2 => n13753, B1 => n6813, B2 => 
                           n13751, ZN => n9649);
   U5431 : OAI22_X1 port map( A1 => n13824, A2 => n13809, B1 => n6830, B2 => 
                           n13804, ZN => n9914);
   U5432 : OAI22_X1 port map( A1 => n13830, A2 => n13809, B1 => n6831, B2 => 
                           n13804, ZN => n9915);
   U5433 : OAI22_X1 port map( A1 => n13836, A2 => n13809, B1 => n6832, B2 => 
                           n13804, ZN => n9916);
   U5434 : OAI22_X1 port map( A1 => n13842, A2 => n13809, B1 => n6833, B2 => 
                           n13804, ZN => n9917);
   U5435 : OAI22_X1 port map( A1 => n13848, A2 => n13809, B1 => n6834, B2 => 
                           n13804, ZN => n9918);
   U5436 : OAI22_X1 port map( A1 => n13854, A2 => n13809, B1 => n6835, B2 => 
                           n13804, ZN => n9919);
   U5437 : OAI22_X1 port map( A1 => n13860, A2 => n13809, B1 => n6836, B2 => 
                           n13804, ZN => n9920);
   U5438 : OAI22_X1 port map( A1 => n13866, A2 => n13809, B1 => n6837, B2 => 
                           n13804, ZN => n9921);
   U5439 : OAI22_X1 port map( A1 => n13872, A2 => n13808, B1 => n6838, B2 => 
                           n13804, ZN => n9922);
   U5440 : OAI22_X1 port map( A1 => n13878, A2 => n13808, B1 => n6839, B2 => 
                           n13804, ZN => n9923);
   U5441 : OAI22_X1 port map( A1 => n13884, A2 => n13808, B1 => n6840, B2 => 
                           n13804, ZN => n9924);
   U5442 : OAI22_X1 port map( A1 => n13890, A2 => n13808, B1 => n6841, B2 => 
                           n13804, ZN => n9925);
   U5443 : OAI22_X1 port map( A1 => n13896, A2 => n13808, B1 => n6883, B2 => 
                           n13805, ZN => n9926);
   U5444 : OAI22_X1 port map( A1 => n13902, A2 => n13808, B1 => n6885, B2 => 
                           n13805, ZN => n9927);
   U5445 : OAI22_X1 port map( A1 => n13908, A2 => n13808, B1 => n6887, B2 => 
                           n13805, ZN => n9928);
   U5446 : OAI22_X1 port map( A1 => n13914, A2 => n13808, B1 => n6889, B2 => 
                           n13805, ZN => n9929);
   U5447 : OAI22_X1 port map( A1 => n13920, A2 => n13808, B1 => n6794, B2 => 
                           n13805, ZN => n9930);
   U5448 : OAI22_X1 port map( A1 => n13926, A2 => n13808, B1 => n6795, B2 => 
                           n13805, ZN => n9931);
   U5449 : OAI22_X1 port map( A1 => n13932, A2 => n13808, B1 => n6796, B2 => 
                           n13805, ZN => n9932);
   U5450 : OAI22_X1 port map( A1 => n13938, A2 => n13808, B1 => n6797, B2 => 
                           n13805, ZN => n9933);
   U5451 : OAI22_X1 port map( A1 => n13944, A2 => n13807, B1 => n6798, B2 => 
                           n13805, ZN => n9934);
   U5452 : OAI22_X1 port map( A1 => n13950, A2 => n13807, B1 => n6799, B2 => 
                           n13805, ZN => n9935);
   U5453 : OAI22_X1 port map( A1 => n13956, A2 => n13807, B1 => n6800, B2 => 
                           n13805, ZN => n9936);
   U5454 : OAI22_X1 port map( A1 => n13962, A2 => n13807, B1 => n6801, B2 => 
                           n13805, ZN => n9937);
   U5455 : OAI22_X1 port map( A1 => n13939, A2 => n13694, B1 => n5776, B2 => 
                           n13691, ZN => n9325);
   U5456 : OAI22_X1 port map( A1 => n13824, A2 => n13791, B1 => n840, B2 => 
                           n13786, ZN => n9818);
   U5457 : OAI22_X1 port map( A1 => n13830, A2 => n13791, B1 => n839, B2 => 
                           n13786, ZN => n9819);
   U5458 : OAI22_X1 port map( A1 => n13836, A2 => n13791, B1 => n838, B2 => 
                           n13786, ZN => n9820);
   U5459 : OAI22_X1 port map( A1 => n13842, A2 => n13791, B1 => n837, B2 => 
                           n13786, ZN => n9821);
   U5460 : OAI22_X1 port map( A1 => n13848, A2 => n13791, B1 => n836, B2 => 
                           n13786, ZN => n9822);
   U5461 : OAI22_X1 port map( A1 => n13854, A2 => n13791, B1 => n835, B2 => 
                           n13786, ZN => n9823);
   U5462 : OAI22_X1 port map( A1 => n13860, A2 => n13791, B1 => n834, B2 => 
                           n13786, ZN => n9824);
   U5463 : OAI22_X1 port map( A1 => n13866, A2 => n13791, B1 => n833, B2 => 
                           n13786, ZN => n9825);
   U5464 : OAI22_X1 port map( A1 => n13872, A2 => n13790, B1 => n832, B2 => 
                           n13786, ZN => n9826);
   U5465 : OAI22_X1 port map( A1 => n13878, A2 => n13790, B1 => n831, B2 => 
                           n13786, ZN => n9827);
   U5466 : OAI22_X1 port map( A1 => n13884, A2 => n13790, B1 => n830, B2 => 
                           n13786, ZN => n9828);
   U5467 : OAI22_X1 port map( A1 => n13890, A2 => n13790, B1 => n829, B2 => 
                           n13786, ZN => n9829);
   U5468 : OAI22_X1 port map( A1 => n13896, A2 => n13790, B1 => n828, B2 => 
                           n13787, ZN => n9830);
   U5469 : OAI22_X1 port map( A1 => n13902, A2 => n13790, B1 => n827, B2 => 
                           n13787, ZN => n9831);
   U5470 : OAI22_X1 port map( A1 => n13908, A2 => n13790, B1 => n826, B2 => 
                           n13787, ZN => n9832);
   U5471 : OAI22_X1 port map( A1 => n13914, A2 => n13790, B1 => n825, B2 => 
                           n13787, ZN => n9833);
   U5472 : OAI22_X1 port map( A1 => n13920, A2 => n13790, B1 => n824, B2 => 
                           n13787, ZN => n9834);
   U5473 : OAI22_X1 port map( A1 => n13926, A2 => n13790, B1 => n823, B2 => 
                           n13787, ZN => n9835);
   U5474 : OAI22_X1 port map( A1 => n13932, A2 => n13790, B1 => n822, B2 => 
                           n13787, ZN => n9836);
   U5475 : OAI22_X1 port map( A1 => n13938, A2 => n13790, B1 => n821, B2 => 
                           n13787, ZN => n9837);
   U5476 : OAI22_X1 port map( A1 => n13944, A2 => n13789, B1 => n820, B2 => 
                           n13787, ZN => n9838);
   U5477 : OAI22_X1 port map( A1 => n13950, A2 => n13789, B1 => n819, B2 => 
                           n13787, ZN => n9839);
   U5478 : OAI22_X1 port map( A1 => n13956, A2 => n13789, B1 => n818, B2 => 
                           n13787, ZN => n9840);
   U5479 : OAI22_X1 port map( A1 => n13962, A2 => n13789, B1 => n817, B2 => 
                           n13787, ZN => n9841);
   U5480 : OAI22_X1 port map( A1 => n13825, A2 => n13737, B1 => n872, B2 => 
                           n13732, ZN => n9530);
   U5481 : OAI22_X1 port map( A1 => n13831, A2 => n13737, B1 => n871, B2 => 
                           n13732, ZN => n9531);
   U5482 : OAI22_X1 port map( A1 => n13837, A2 => n13737, B1 => n870, B2 => 
                           n13732, ZN => n9532);
   U5483 : OAI22_X1 port map( A1 => n13843, A2 => n13737, B1 => n869, B2 => 
                           n13732, ZN => n9533);
   U5484 : OAI22_X1 port map( A1 => n13849, A2 => n13737, B1 => n868, B2 => 
                           n13732, ZN => n9534);
   U5485 : OAI22_X1 port map( A1 => n13855, A2 => n13737, B1 => n867, B2 => 
                           n13732, ZN => n9535);
   U5486 : OAI22_X1 port map( A1 => n13861, A2 => n13737, B1 => n866, B2 => 
                           n13732, ZN => n9536);
   U5487 : OAI22_X1 port map( A1 => n13867, A2 => n13737, B1 => n865, B2 => 
                           n13732, ZN => n9537);
   U5488 : OAI22_X1 port map( A1 => n13873, A2 => n13736, B1 => n864, B2 => 
                           n13732, ZN => n9538);
   U5489 : OAI22_X1 port map( A1 => n13879, A2 => n13736, B1 => n863, B2 => 
                           n13732, ZN => n9539);
   U5490 : OAI22_X1 port map( A1 => n13885, A2 => n13736, B1 => n862, B2 => 
                           n13732, ZN => n9540);
   U5491 : OAI22_X1 port map( A1 => n13891, A2 => n13736, B1 => n861, B2 => 
                           n13732, ZN => n9541);
   U5492 : OAI22_X1 port map( A1 => n13897, A2 => n13736, B1 => n860, B2 => 
                           n13733, ZN => n9542);
   U5493 : OAI22_X1 port map( A1 => n13903, A2 => n13736, B1 => n859, B2 => 
                           n13733, ZN => n9543);
   U5494 : OAI22_X1 port map( A1 => n13909, A2 => n13736, B1 => n858, B2 => 
                           n13733, ZN => n9544);
   U5495 : OAI22_X1 port map( A1 => n13915, A2 => n13736, B1 => n857, B2 => 
                           n13733, ZN => n9545);
   U5496 : OAI22_X1 port map( A1 => n13921, A2 => n13736, B1 => n856, B2 => 
                           n13733, ZN => n9546);
   U5497 : OAI22_X1 port map( A1 => n13927, A2 => n13736, B1 => n855, B2 => 
                           n13733, ZN => n9547);
   U5498 : OAI22_X1 port map( A1 => n13933, A2 => n13736, B1 => n854, B2 => 
                           n13733, ZN => n9548);
   U5499 : OAI22_X1 port map( A1 => n13939, A2 => n13736, B1 => n853, B2 => 
                           n13733, ZN => n9549);
   U5500 : OAI22_X1 port map( A1 => n13945, A2 => n13735, B1 => n852, B2 => 
                           n13733, ZN => n9550);
   U5501 : OAI22_X1 port map( A1 => n13951, A2 => n13735, B1 => n851, B2 => 
                           n13733, ZN => n9551);
   U5502 : OAI22_X1 port map( A1 => n13957, A2 => n13735, B1 => n850, B2 => 
                           n13733, ZN => n9552);
   U5503 : OAI22_X1 port map( A1 => n13963, A2 => n13735, B1 => n849, B2 => 
                           n13733, ZN => n9553);
   U5504 : OAI22_X1 port map( A1 => n13945, A2 => n13693, B1 => n5780, B2 => 
                           n13691, ZN => n9326);
   U5505 : OAI22_X1 port map( A1 => n13951, A2 => n13693, B1 => n5784, B2 => 
                           n13691, ZN => n9327);
   U5506 : OAI22_X1 port map( A1 => n13957, A2 => n13693, B1 => n5788, B2 => 
                           n13691, ZN => n9328);
   U5507 : OAI22_X1 port map( A1 => n13963, A2 => n13693, B1 => n5792, B2 => 
                           n13691, ZN => n9329);
   U5508 : OAI22_X1 port map( A1 => n13825, A2 => n13689, B1 => n5701, B2 => 
                           n13684, ZN => n9274);
   U5509 : OAI22_X1 port map( A1 => n13831, A2 => n13689, B1 => n5705, B2 => 
                           n13684, ZN => n9275);
   U5510 : OAI22_X1 port map( A1 => n13837, A2 => n13689, B1 => n5709, B2 => 
                           n13684, ZN => n9276);
   U5511 : OAI22_X1 port map( A1 => n13843, A2 => n13689, B1 => n5713, B2 => 
                           n13684, ZN => n9277);
   U5512 : OAI22_X1 port map( A1 => n13849, A2 => n13689, B1 => n5717, B2 => 
                           n13684, ZN => n9278);
   U5513 : OAI22_X1 port map( A1 => n13855, A2 => n13689, B1 => n5721, B2 => 
                           n13684, ZN => n9279);
   U5514 : OAI22_X1 port map( A1 => n13861, A2 => n13689, B1 => n5725, B2 => 
                           n13684, ZN => n9280);
   U5515 : OAI22_X1 port map( A1 => n13867, A2 => n13689, B1 => n5729, B2 => 
                           n13684, ZN => n9281);
   U5516 : OAI22_X1 port map( A1 => n13873, A2 => n13688, B1 => n5733, B2 => 
                           n13684, ZN => n9282);
   U5517 : OAI22_X1 port map( A1 => n13879, A2 => n13688, B1 => n5737, B2 => 
                           n13684, ZN => n9283);
   U5518 : OAI22_X1 port map( A1 => n13885, A2 => n13688, B1 => n5741, B2 => 
                           n13684, ZN => n9284);
   U5519 : OAI22_X1 port map( A1 => n13891, A2 => n13688, B1 => n5745, B2 => 
                           n13684, ZN => n9285);
   U5520 : OAI22_X1 port map( A1 => n13897, A2 => n13688, B1 => n5749, B2 => 
                           n13685, ZN => n9286);
   U5521 : OAI22_X1 port map( A1 => n13903, A2 => n13688, B1 => n5753, B2 => 
                           n13685, ZN => n9287);
   U5522 : OAI22_X1 port map( A1 => n13909, A2 => n13688, B1 => n5757, B2 => 
                           n13685, ZN => n9288);
   U5523 : OAI22_X1 port map( A1 => n13915, A2 => n13688, B1 => n5761, B2 => 
                           n13685, ZN => n9289);
   U5524 : OAI22_X1 port map( A1 => n13921, A2 => n13688, B1 => n5765, B2 => 
                           n13685, ZN => n9290);
   U5525 : OAI22_X1 port map( A1 => n13927, A2 => n13688, B1 => n5769, B2 => 
                           n13685, ZN => n9291);
   U5526 : OAI22_X1 port map( A1 => n13933, A2 => n13688, B1 => n5773, B2 => 
                           n13685, ZN => n9292);
   U5527 : OAI22_X1 port map( A1 => n13939, A2 => n13688, B1 => n5777, B2 => 
                           n13685, ZN => n9293);
   U5528 : OAI22_X1 port map( A1 => n13945, A2 => n13687, B1 => n5781, B2 => 
                           n13685, ZN => n9294);
   U5529 : OAI22_X1 port map( A1 => n13951, A2 => n13687, B1 => n5785, B2 => 
                           n13685, ZN => n9295);
   U5530 : OAI22_X1 port map( A1 => n13957, A2 => n13687, B1 => n5789, B2 => 
                           n13685, ZN => n9296);
   U5531 : OAI22_X1 port map( A1 => n13963, A2 => n13687, B1 => n5793, B2 => 
                           n13685, ZN => n9297);
   U5532 : OAI22_X1 port map( A1 => n13825, A2 => n13683, B1 => n904, B2 => 
                           n13678, ZN => n9242);
   U5533 : OAI22_X1 port map( A1 => n13831, A2 => n13683, B1 => n903, B2 => 
                           n13678, ZN => n9243);
   U5534 : OAI22_X1 port map( A1 => n13837, A2 => n13683, B1 => n902, B2 => 
                           n13678, ZN => n9244);
   U5535 : OAI22_X1 port map( A1 => n13843, A2 => n13683, B1 => n901, B2 => 
                           n13678, ZN => n9245);
   U5536 : OAI22_X1 port map( A1 => n13849, A2 => n13683, B1 => n900, B2 => 
                           n13678, ZN => n9246);
   U5537 : OAI22_X1 port map( A1 => n13855, A2 => n13683, B1 => n899, B2 => 
                           n13678, ZN => n9247);
   U5538 : OAI22_X1 port map( A1 => n13861, A2 => n13683, B1 => n898, B2 => 
                           n13678, ZN => n9248);
   U5539 : OAI22_X1 port map( A1 => n13867, A2 => n13683, B1 => n897, B2 => 
                           n13678, ZN => n9249);
   U5540 : OAI22_X1 port map( A1 => n13873, A2 => n13682, B1 => n896, B2 => 
                           n13678, ZN => n9250);
   U5541 : OAI22_X1 port map( A1 => n13879, A2 => n13682, B1 => n895, B2 => 
                           n13678, ZN => n9251);
   U5542 : OAI22_X1 port map( A1 => n13885, A2 => n13682, B1 => n894, B2 => 
                           n13678, ZN => n9252);
   U5543 : OAI22_X1 port map( A1 => n13891, A2 => n13682, B1 => n893, B2 => 
                           n13678, ZN => n9253);
   U5544 : OAI22_X1 port map( A1 => n13897, A2 => n13682, B1 => n892, B2 => 
                           n13679, ZN => n9254);
   U5545 : OAI22_X1 port map( A1 => n13903, A2 => n13682, B1 => n891, B2 => 
                           n13679, ZN => n9255);
   U5546 : OAI22_X1 port map( A1 => n13909, A2 => n13682, B1 => n890, B2 => 
                           n13679, ZN => n9256);
   U5547 : OAI22_X1 port map( A1 => n13915, A2 => n13682, B1 => n889, B2 => 
                           n13679, ZN => n9257);
   U5548 : OAI22_X1 port map( A1 => n13921, A2 => n13682, B1 => n888, B2 => 
                           n13679, ZN => n9258);
   U5549 : OAI22_X1 port map( A1 => n13927, A2 => n13682, B1 => n887, B2 => 
                           n13679, ZN => n9259);
   U5550 : OAI22_X1 port map( A1 => n13933, A2 => n13682, B1 => n886, B2 => 
                           n13679, ZN => n9260);
   U5551 : OAI22_X1 port map( A1 => n13939, A2 => n13682, B1 => n885, B2 => 
                           n13679, ZN => n9261);
   U5552 : OAI22_X1 port map( A1 => n13945, A2 => n13681, B1 => n884, B2 => 
                           n13679, ZN => n9262);
   U5553 : OAI22_X1 port map( A1 => n13951, A2 => n13681, B1 => n883, B2 => 
                           n13679, ZN => n9263);
   U5554 : OAI22_X1 port map( A1 => n13957, A2 => n13681, B1 => n882, B2 => 
                           n13679, ZN => n9264);
   U5555 : OAI22_X1 port map( A1 => n13963, A2 => n13681, B1 => n881, B2 => 
                           n13679, ZN => n9265);
   U5556 : OAI22_X1 port map( A1 => n13874, A2 => n13640, B1 => n5462, B2 => 
                           n13636, ZN => n9026);
   U5557 : OAI22_X1 port map( A1 => n13880, A2 => n13640, B1 => n5472, B2 => 
                           n13636, ZN => n9027);
   U5558 : OAI22_X1 port map( A1 => n13886, A2 => n13640, B1 => n5482, B2 => 
                           n13636, ZN => n9028);
   U5559 : OAI22_X1 port map( A1 => n13892, A2 => n13640, B1 => n5492, B2 => 
                           n13636, ZN => n9029);
   U5560 : OAI22_X1 port map( A1 => n13898, A2 => n13640, B1 => n5502, B2 => 
                           n13637, ZN => n9030);
   U5561 : OAI22_X1 port map( A1 => n13904, A2 => n13640, B1 => n5512, B2 => 
                           n13637, ZN => n9031);
   U5562 : OAI22_X1 port map( A1 => n13910, A2 => n13640, B1 => n5522, B2 => 
                           n13637, ZN => n9032);
   U5563 : OAI22_X1 port map( A1 => n13916, A2 => n13640, B1 => n5532, B2 => 
                           n13637, ZN => n9033);
   U5564 : OAI22_X1 port map( A1 => n13922, A2 => n13640, B1 => n5542, B2 => 
                           n13637, ZN => n9034);
   U5565 : OAI22_X1 port map( A1 => n13928, A2 => n13640, B1 => n5552, B2 => 
                           n13637, ZN => n9035);
   U5566 : OAI22_X1 port map( A1 => n13934, A2 => n13640, B1 => n5562, B2 => 
                           n13637, ZN => n9036);
   U5567 : OAI22_X1 port map( A1 => n13940, A2 => n13640, B1 => n5572, B2 => 
                           n13637, ZN => n9037);
   U5568 : OAI22_X1 port map( A1 => n13946, A2 => n13639, B1 => n5582, B2 => 
                           n13637, ZN => n9038);
   U5569 : OAI22_X1 port map( A1 => n13952, A2 => n13639, B1 => n5592, B2 => 
                           n13637, ZN => n9039);
   U5570 : OAI22_X1 port map( A1 => n13958, A2 => n13639, B1 => n5602, B2 => 
                           n13637, ZN => n9040);
   U5571 : OAI22_X1 port map( A1 => n13964, A2 => n13639, B1 => n5612, B2 => 
                           n13637, ZN => n9041);
   U5572 : OAI22_X1 port map( A1 => n13826, A2 => n13635, B1 => n5383, B2 => 
                           n13630, ZN => n8986);
   U5573 : OAI22_X1 port map( A1 => n13832, A2 => n13635, B1 => n5393, B2 => 
                           n13630, ZN => n8987);
   U5574 : OAI22_X1 port map( A1 => n13838, A2 => n13635, B1 => n5403, B2 => 
                           n13630, ZN => n8988);
   U5575 : OAI22_X1 port map( A1 => n13844, A2 => n13635, B1 => n5413, B2 => 
                           n13630, ZN => n8989);
   U5576 : OAI22_X1 port map( A1 => n13850, A2 => n13635, B1 => n5423, B2 => 
                           n13630, ZN => n8990);
   U5577 : OAI22_X1 port map( A1 => n13856, A2 => n13635, B1 => n5433, B2 => 
                           n13630, ZN => n8991);
   U5578 : OAI22_X1 port map( A1 => n13862, A2 => n13635, B1 => n5443, B2 => 
                           n13630, ZN => n8992);
   U5579 : OAI22_X1 port map( A1 => n13868, A2 => n13635, B1 => n5453, B2 => 
                           n13630, ZN => n8993);
   U5580 : OAI22_X1 port map( A1 => n13874, A2 => n13634, B1 => n5463, B2 => 
                           n13630, ZN => n8994);
   U5581 : OAI22_X1 port map( A1 => n13880, A2 => n13634, B1 => n5473, B2 => 
                           n13630, ZN => n8995);
   U5582 : OAI22_X1 port map( A1 => n13886, A2 => n13634, B1 => n5483, B2 => 
                           n13630, ZN => n8996);
   U5583 : OAI22_X1 port map( A1 => n13892, A2 => n13634, B1 => n5493, B2 => 
                           n13630, ZN => n8997);
   U5584 : OAI22_X1 port map( A1 => n13898, A2 => n13634, B1 => n5503, B2 => 
                           n13631, ZN => n8998);
   U5585 : OAI22_X1 port map( A1 => n13904, A2 => n13634, B1 => n5513, B2 => 
                           n13631, ZN => n8999);
   U5586 : OAI22_X1 port map( A1 => n13910, A2 => n13634, B1 => n5523, B2 => 
                           n13631, ZN => n9000);
   U5587 : OAI22_X1 port map( A1 => n13916, A2 => n13634, B1 => n5533, B2 => 
                           n13631, ZN => n9001);
   U5588 : OAI22_X1 port map( A1 => n13922, A2 => n13634, B1 => n5543, B2 => 
                           n13631, ZN => n9002);
   U5589 : OAI22_X1 port map( A1 => n13928, A2 => n13634, B1 => n5553, B2 => 
                           n13631, ZN => n9003);
   U5590 : OAI22_X1 port map( A1 => n13934, A2 => n13634, B1 => n5563, B2 => 
                           n13631, ZN => n9004);
   U5591 : OAI22_X1 port map( A1 => n13940, A2 => n13634, B1 => n5573, B2 => 
                           n13631, ZN => n9005);
   U5592 : OAI22_X1 port map( A1 => n13946, A2 => n13633, B1 => n5583, B2 => 
                           n13631, ZN => n9006);
   U5593 : OAI22_X1 port map( A1 => n13952, A2 => n13633, B1 => n5593, B2 => 
                           n13631, ZN => n9007);
   U5594 : OAI22_X1 port map( A1 => n13958, A2 => n13633, B1 => n5603, B2 => 
                           n13631, ZN => n9008);
   U5595 : OAI22_X1 port map( A1 => n13964, A2 => n13633, B1 => n5613, B2 => 
                           n13631, ZN => n9009);
   U5596 : OAI22_X1 port map( A1 => n13826, A2 => n13629, B1 => n936, B2 => 
                           n13624, ZN => n8954);
   U5597 : OAI22_X1 port map( A1 => n13832, A2 => n13629, B1 => n935, B2 => 
                           n13624, ZN => n8955);
   U5598 : OAI22_X1 port map( A1 => n13838, A2 => n13629, B1 => n934, B2 => 
                           n13624, ZN => n8956);
   U5599 : OAI22_X1 port map( A1 => n13844, A2 => n13629, B1 => n933, B2 => 
                           n13624, ZN => n8957);
   U5600 : OAI22_X1 port map( A1 => n13850, A2 => n13629, B1 => n932, B2 => 
                           n13624, ZN => n8958);
   U5601 : OAI22_X1 port map( A1 => n13856, A2 => n13629, B1 => n931, B2 => 
                           n13624, ZN => n8959);
   U5602 : OAI22_X1 port map( A1 => n13862, A2 => n13629, B1 => n930, B2 => 
                           n13624, ZN => n8960);
   U5603 : OAI22_X1 port map( A1 => n13868, A2 => n13629, B1 => n929, B2 => 
                           n13624, ZN => n8961);
   U5604 : OAI22_X1 port map( A1 => n13874, A2 => n13628, B1 => n928, B2 => 
                           n13624, ZN => n8962);
   U5605 : OAI22_X1 port map( A1 => n13880, A2 => n13628, B1 => n927, B2 => 
                           n13624, ZN => n8963);
   U5606 : OAI22_X1 port map( A1 => n13886, A2 => n13628, B1 => n926, B2 => 
                           n13624, ZN => n8964);
   U5607 : OAI22_X1 port map( A1 => n13892, A2 => n13628, B1 => n925, B2 => 
                           n13624, ZN => n8965);
   U5608 : OAI22_X1 port map( A1 => n13898, A2 => n13628, B1 => n924, B2 => 
                           n13625, ZN => n8966);
   U5609 : OAI22_X1 port map( A1 => n13904, A2 => n13628, B1 => n923, B2 => 
                           n13625, ZN => n8967);
   U5610 : OAI22_X1 port map( A1 => n13910, A2 => n13628, B1 => n922, B2 => 
                           n13625, ZN => n8968);
   U5611 : OAI22_X1 port map( A1 => n13916, A2 => n13628, B1 => n921, B2 => 
                           n13625, ZN => n8969);
   U5612 : OAI22_X1 port map( A1 => n13922, A2 => n13628, B1 => n920, B2 => 
                           n13625, ZN => n8970);
   U5613 : OAI22_X1 port map( A1 => n13928, A2 => n13628, B1 => n919, B2 => 
                           n13625, ZN => n8971);
   U5614 : OAI22_X1 port map( A1 => n13934, A2 => n13628, B1 => n918, B2 => 
                           n13625, ZN => n8972);
   U5615 : OAI22_X1 port map( A1 => n13940, A2 => n13628, B1 => n917, B2 => 
                           n13625, ZN => n8973);
   U5616 : OAI22_X1 port map( A1 => n13946, A2 => n13627, B1 => n916, B2 => 
                           n13625, ZN => n8974);
   U5617 : OAI22_X1 port map( A1 => n13952, A2 => n13627, B1 => n915, B2 => 
                           n13625, ZN => n8975);
   U5618 : OAI22_X1 port map( A1 => n13958, A2 => n13627, B1 => n914, B2 => 
                           n13625, ZN => n8976);
   U5619 : OAI22_X1 port map( A1 => n13964, A2 => n13627, B1 => n913, B2 => 
                           n13625, ZN => n8977);
   U5620 : OAI22_X1 port map( A1 => n13947, A2 => n13585, B1 => n5778, B2 => 
                           n13582, ZN => n8750);
   U5621 : OAI22_X1 port map( A1 => n13953, A2 => n13585, B1 => n5782, B2 => 
                           n13582, ZN => n8751);
   U5622 : OAI22_X1 port map( A1 => n13959, A2 => n13585, B1 => n5786, B2 => 
                           n13582, ZN => n8752);
   U5623 : OAI22_X1 port map( A1 => n13965, A2 => n13585, B1 => n5790, B2 => 
                           n13582, ZN => n8753);
   U5624 : OAI22_X1 port map( A1 => n13971, A2 => n13585, B1 => n5794, B2 => 
                           n13582, ZN => n8754);
   U5625 : OAI22_X1 port map( A1 => n13977, A2 => n13585, B1 => n5798, B2 => 
                           n13582, ZN => n8755);
   U5626 : OAI22_X1 port map( A1 => n13983, A2 => n13585, B1 => n5802, B2 => 
                           n13582, ZN => n8756);
   U5627 : OAI22_X1 port map( A1 => n13989, A2 => n13585, B1 => n5806, B2 => 
                           n13582, ZN => n8757);
   U5628 : OAI22_X1 port map( A1 => n13995, A2 => n13585, B1 => n5810, B2 => 
                           n13582, ZN => n8758);
   U5629 : OAI22_X1 port map( A1 => n14001, A2 => n13585, B1 => n5814, B2 => 
                           n13582, ZN => n8759);
   U5630 : OAI22_X1 port map( A1 => n14007, A2 => n13585, B1 => n5818, B2 => 
                           n13582, ZN => n8760);
   U5631 : OAI22_X1 port map( A1 => n14016, A2 => n13585, B1 => n5822, B2 => 
                           n13582, ZN => n8761);
   U5632 : OAI22_X1 port map( A1 => n13827, A2 => n13581, B1 => n5699, B2 => 
                           n13576, ZN => n8698);
   U5633 : OAI22_X1 port map( A1 => n13833, A2 => n13581, B1 => n5703, B2 => 
                           n13576, ZN => n8699);
   U5634 : OAI22_X1 port map( A1 => n13839, A2 => n13581, B1 => n5707, B2 => 
                           n13576, ZN => n8700);
   U5635 : OAI22_X1 port map( A1 => n13845, A2 => n13581, B1 => n5711, B2 => 
                           n13576, ZN => n8701);
   U5636 : OAI22_X1 port map( A1 => n13851, A2 => n13581, B1 => n5715, B2 => 
                           n13576, ZN => n8702);
   U5637 : OAI22_X1 port map( A1 => n13857, A2 => n13581, B1 => n5719, B2 => 
                           n13576, ZN => n8703);
   U5638 : OAI22_X1 port map( A1 => n13863, A2 => n13581, B1 => n5723, B2 => 
                           n13576, ZN => n8704);
   U5639 : OAI22_X1 port map( A1 => n13869, A2 => n13581, B1 => n5727, B2 => 
                           n13576, ZN => n8705);
   U5640 : OAI22_X1 port map( A1 => n13875, A2 => n13580, B1 => n5731, B2 => 
                           n13576, ZN => n8706);
   U5641 : OAI22_X1 port map( A1 => n13881, A2 => n13580, B1 => n5735, B2 => 
                           n13576, ZN => n8707);
   U5642 : OAI22_X1 port map( A1 => n13887, A2 => n13580, B1 => n5739, B2 => 
                           n13576, ZN => n8708);
   U5643 : OAI22_X1 port map( A1 => n13893, A2 => n13580, B1 => n5743, B2 => 
                           n13576, ZN => n8709);
   U5644 : OAI22_X1 port map( A1 => n13899, A2 => n13580, B1 => n5747, B2 => 
                           n13577, ZN => n8710);
   U5645 : OAI22_X1 port map( A1 => n13905, A2 => n13580, B1 => n5751, B2 => 
                           n13577, ZN => n8711);
   U5646 : OAI22_X1 port map( A1 => n13911, A2 => n13580, B1 => n5755, B2 => 
                           n13577, ZN => n8712);
   U5647 : OAI22_X1 port map( A1 => n13917, A2 => n13580, B1 => n5759, B2 => 
                           n13577, ZN => n8713);
   U5648 : OAI22_X1 port map( A1 => n13923, A2 => n13580, B1 => n5763, B2 => 
                           n13577, ZN => n8714);
   U5649 : OAI22_X1 port map( A1 => n13929, A2 => n13580, B1 => n5767, B2 => 
                           n13577, ZN => n8715);
   U5650 : OAI22_X1 port map( A1 => n13935, A2 => n13580, B1 => n5771, B2 => 
                           n13577, ZN => n8716);
   U5651 : OAI22_X1 port map( A1 => n13941, A2 => n13580, B1 => n5775, B2 => 
                           n13577, ZN => n8717);
   U5652 : OAI22_X1 port map( A1 => n13947, A2 => n13579, B1 => n5779, B2 => 
                           n13577, ZN => n8718);
   U5653 : OAI22_X1 port map( A1 => n13953, A2 => n13579, B1 => n5783, B2 => 
                           n13577, ZN => n8719);
   U5654 : OAI22_X1 port map( A1 => n13959, A2 => n13579, B1 => n5787, B2 => 
                           n13577, ZN => n8720);
   U5655 : OAI22_X1 port map( A1 => n13965, A2 => n13579, B1 => n5791, B2 => 
                           n13577, ZN => n8721);
   U5656 : OAI22_X1 port map( A1 => n13827, A2 => n13575, B1 => n968, B2 => 
                           n13570, ZN => n8666);
   U5657 : OAI22_X1 port map( A1 => n13833, A2 => n13575, B1 => n967, B2 => 
                           n13570, ZN => n8667);
   U5658 : OAI22_X1 port map( A1 => n13839, A2 => n13575, B1 => n966, B2 => 
                           n13570, ZN => n8668);
   U5659 : OAI22_X1 port map( A1 => n13845, A2 => n13575, B1 => n965, B2 => 
                           n13570, ZN => n8669);
   U5660 : OAI22_X1 port map( A1 => n13851, A2 => n13575, B1 => n964, B2 => 
                           n13570, ZN => n8670);
   U5661 : OAI22_X1 port map( A1 => n13857, A2 => n13575, B1 => n963, B2 => 
                           n13570, ZN => n8671);
   U5662 : OAI22_X1 port map( A1 => n13863, A2 => n13575, B1 => n962, B2 => 
                           n13570, ZN => n8672);
   U5663 : OAI22_X1 port map( A1 => n13869, A2 => n13575, B1 => n961, B2 => 
                           n13570, ZN => n8673);
   U5664 : OAI22_X1 port map( A1 => n13875, A2 => n13574, B1 => n960, B2 => 
                           n13570, ZN => n8674);
   U5665 : OAI22_X1 port map( A1 => n13881, A2 => n13574, B1 => n959, B2 => 
                           n13570, ZN => n8675);
   U5666 : OAI22_X1 port map( A1 => n13887, A2 => n13574, B1 => n958, B2 => 
                           n13570, ZN => n8676);
   U5667 : OAI22_X1 port map( A1 => n13893, A2 => n13574, B1 => n957, B2 => 
                           n13570, ZN => n8677);
   U5668 : OAI22_X1 port map( A1 => n13899, A2 => n13574, B1 => n956, B2 => 
                           n13571, ZN => n8678);
   U5669 : OAI22_X1 port map( A1 => n13905, A2 => n13574, B1 => n955, B2 => 
                           n13571, ZN => n8679);
   U5670 : OAI22_X1 port map( A1 => n13911, A2 => n13574, B1 => n954, B2 => 
                           n13571, ZN => n8680);
   U5671 : OAI22_X1 port map( A1 => n13917, A2 => n13574, B1 => n953, B2 => 
                           n13571, ZN => n8681);
   U5672 : OAI22_X1 port map( A1 => n13923, A2 => n13574, B1 => n952, B2 => 
                           n13571, ZN => n8682);
   U5673 : OAI22_X1 port map( A1 => n13929, A2 => n13574, B1 => n951, B2 => 
                           n13571, ZN => n8683);
   U5674 : OAI22_X1 port map( A1 => n13935, A2 => n13574, B1 => n950, B2 => 
                           n13571, ZN => n8684);
   U5675 : OAI22_X1 port map( A1 => n13941, A2 => n13574, B1 => n949, B2 => 
                           n13571, ZN => n8685);
   U5676 : OAI22_X1 port map( A1 => n13947, A2 => n13573, B1 => n948, B2 => 
                           n13571, ZN => n8686);
   U5677 : OAI22_X1 port map( A1 => n13953, A2 => n13573, B1 => n947, B2 => 
                           n13571, ZN => n8687);
   U5678 : OAI22_X1 port map( A1 => n13959, A2 => n13573, B1 => n946, B2 => 
                           n13571, ZN => n8688);
   U5679 : OAI22_X1 port map( A1 => n13965, A2 => n13573, B1 => n945, B2 => 
                           n13571, ZN => n8689);
   U5680 : OAI22_X1 port map( A1 => n13827, A2 => n13545, B1 => n712, B2 => 
                           n13540, ZN => n8506);
   U5681 : OAI22_X1 port map( A1 => n13833, A2 => n13545, B1 => n709, B2 => 
                           n13540, ZN => n8507);
   U5682 : OAI22_X1 port map( A1 => n13839, A2 => n13545, B1 => n706, B2 => 
                           n13540, ZN => n8508);
   U5683 : OAI22_X1 port map( A1 => n13845, A2 => n13545, B1 => n703, B2 => 
                           n13540, ZN => n8509);
   U5684 : OAI22_X1 port map( A1 => n13851, A2 => n13545, B1 => n700, B2 => 
                           n13540, ZN => n8510);
   U5685 : OAI22_X1 port map( A1 => n13857, A2 => n13545, B1 => n697, B2 => 
                           n13540, ZN => n8511);
   U5686 : OAI22_X1 port map( A1 => n13863, A2 => n13545, B1 => n694, B2 => 
                           n13540, ZN => n8512);
   U5687 : OAI22_X1 port map( A1 => n13869, A2 => n13545, B1 => n691, B2 => 
                           n13540, ZN => n8513);
   U5688 : OAI22_X1 port map( A1 => n13875, A2 => n13544, B1 => n688, B2 => 
                           n13540, ZN => n8514);
   U5689 : OAI22_X1 port map( A1 => n13881, A2 => n13544, B1 => n685, B2 => 
                           n13540, ZN => n8515);
   U5690 : OAI22_X1 port map( A1 => n13887, A2 => n13544, B1 => n682, B2 => 
                           n13540, ZN => n8516);
   U5691 : OAI22_X1 port map( A1 => n13893, A2 => n13544, B1 => n679, B2 => 
                           n13540, ZN => n8517);
   U5692 : OAI22_X1 port map( A1 => n13899, A2 => n13544, B1 => n676, B2 => 
                           n13541, ZN => n8518);
   U5693 : OAI22_X1 port map( A1 => n13905, A2 => n13544, B1 => n673, B2 => 
                           n13541, ZN => n8519);
   U5694 : OAI22_X1 port map( A1 => n13911, A2 => n13544, B1 => n670, B2 => 
                           n13541, ZN => n8520);
   U5695 : OAI22_X1 port map( A1 => n13917, A2 => n13544, B1 => n667, B2 => 
                           n13541, ZN => n8521);
   U5696 : OAI22_X1 port map( A1 => n13923, A2 => n13544, B1 => n664, B2 => 
                           n13541, ZN => n8522);
   U5697 : OAI22_X1 port map( A1 => n13929, A2 => n13544, B1 => n661, B2 => 
                           n13541, ZN => n8523);
   U5698 : OAI22_X1 port map( A1 => n13935, A2 => n13544, B1 => n658, B2 => 
                           n13541, ZN => n8524);
   U5699 : OAI22_X1 port map( A1 => n13941, A2 => n13544, B1 => n655, B2 => 
                           n13541, ZN => n8525);
   U5700 : OAI22_X1 port map( A1 => n13947, A2 => n13543, B1 => n652, B2 => 
                           n13541, ZN => n8526);
   U5701 : OAI22_X1 port map( A1 => n13953, A2 => n13543, B1 => n649, B2 => 
                           n13541, ZN => n8527);
   U5702 : OAI22_X1 port map( A1 => n13959, A2 => n13543, B1 => n646, B2 => 
                           n13541, ZN => n8528);
   U5703 : OAI22_X1 port map( A1 => n13965, A2 => n13543, B1 => n643, B2 => 
                           n13541, ZN => n8529);
   U5704 : OAI22_X1 port map( A1 => n13875, A2 => n13520, B1 => n992, B2 => 
                           n13516, ZN => n8386);
   U5705 : OAI22_X1 port map( A1 => n13881, A2 => n13520, B1 => n991, B2 => 
                           n13516, ZN => n8387);
   U5706 : OAI22_X1 port map( A1 => n13887, A2 => n13520, B1 => n990, B2 => 
                           n13516, ZN => n8388);
   U5707 : OAI22_X1 port map( A1 => n13893, A2 => n13520, B1 => n989, B2 => 
                           n13516, ZN => n8389);
   U5708 : OAI22_X1 port map( A1 => n13899, A2 => n13520, B1 => n988, B2 => 
                           n13517, ZN => n8390);
   U5709 : OAI22_X1 port map( A1 => n13905, A2 => n13520, B1 => n987, B2 => 
                           n13517, ZN => n8391);
   U5710 : OAI22_X1 port map( A1 => n13911, A2 => n13520, B1 => n986, B2 => 
                           n13517, ZN => n8392);
   U5711 : OAI22_X1 port map( A1 => n13917, A2 => n13520, B1 => n985, B2 => 
                           n13517, ZN => n8393);
   U5712 : OAI22_X1 port map( A1 => n13923, A2 => n13520, B1 => n984, B2 => 
                           n13517, ZN => n8394);
   U5713 : OAI22_X1 port map( A1 => n13929, A2 => n13520, B1 => n983, B2 => 
                           n13517, ZN => n8395);
   U5714 : OAI22_X1 port map( A1 => n13935, A2 => n13520, B1 => n982, B2 => 
                           n13517, ZN => n8396);
   U5715 : OAI22_X1 port map( A1 => n13941, A2 => n13520, B1 => n981, B2 => 
                           n13517, ZN => n8397);
   U5716 : OAI22_X1 port map( A1 => n13947, A2 => n13519, B1 => n980, B2 => 
                           n13517, ZN => n8398);
   U5717 : OAI22_X1 port map( A1 => n13953, A2 => n13519, B1 => n979, B2 => 
                           n13517, ZN => n8399);
   U5718 : OAI22_X1 port map( A1 => n13959, A2 => n13519, B1 => n978, B2 => 
                           n13517, ZN => n8400);
   U5719 : OAI22_X1 port map( A1 => n13965, A2 => n13519, B1 => n977, B2 => 
                           n13517, ZN => n8401);
   U5720 : OAI22_X1 port map( A1 => n13868, A2 => n13641, B1 => n5452, B2 => 
                           n13636, ZN => n9025);
   U5721 : OAI22_X1 port map( A1 => n13833, A2 => n13521, B1 => n999, B2 => 
                           n13516, ZN => n8379);
   U5722 : OAI22_X1 port map( A1 => n13839, A2 => n13521, B1 => n998, B2 => 
                           n13516, ZN => n8380);
   U5723 : OAI22_X1 port map( A1 => n13845, A2 => n13521, B1 => n997, B2 => 
                           n13516, ZN => n8381);
   U5724 : OAI22_X1 port map( A1 => n13851, A2 => n13521, B1 => n996, B2 => 
                           n13516, ZN => n8382);
   U5725 : OAI22_X1 port map( A1 => n13857, A2 => n13521, B1 => n995, B2 => 
                           n13516, ZN => n8383);
   U5726 : OAI22_X1 port map( A1 => n13863, A2 => n13521, B1 => n994, B2 => 
                           n13516, ZN => n8384);
   U5727 : OAI22_X1 port map( A1 => n13869, A2 => n13521, B1 => n993, B2 => 
                           n13516, ZN => n8385);
   U5728 : OAI22_X1 port map( A1 => n13828, A2 => n13437, B1 => n7192, B2 => 
                           n13432, ZN => n7930);
   U5729 : OAI22_X1 port map( A1 => n13828, A2 => n13467, B1 => n7224, B2 => 
                           n13462, ZN => n8090);
   U5730 : OAI22_X1 port map( A1 => n13834, A2 => n13467, B1 => n7225, B2 => 
                           n13462, ZN => n8091);
   U5731 : OAI22_X1 port map( A1 => n13840, A2 => n13467, B1 => n7226, B2 => 
                           n13462, ZN => n8092);
   U5732 : OAI22_X1 port map( A1 => n13846, A2 => n13467, B1 => n7227, B2 => 
                           n13462, ZN => n8093);
   U5733 : OAI22_X1 port map( A1 => n13852, A2 => n13467, B1 => n7228, B2 => 
                           n13462, ZN => n8094);
   U5734 : OAI22_X1 port map( A1 => n13858, A2 => n13467, B1 => n7229, B2 => 
                           n13462, ZN => n8095);
   U5735 : OAI22_X1 port map( A1 => n13864, A2 => n13467, B1 => n7230, B2 => 
                           n13462, ZN => n8096);
   U5736 : OAI22_X1 port map( A1 => n13870, A2 => n13467, B1 => n7231, B2 => 
                           n13462, ZN => n8097);
   U5737 : OAI22_X1 port map( A1 => n13876, A2 => n13466, B1 => n7232, B2 => 
                           n13462, ZN => n8098);
   U5738 : OAI22_X1 port map( A1 => n13882, A2 => n13466, B1 => n7233, B2 => 
                           n13462, ZN => n8099);
   U5739 : OAI22_X1 port map( A1 => n13888, A2 => n13466, B1 => n7234, B2 => 
                           n13462, ZN => n8100);
   U5740 : OAI22_X1 port map( A1 => n13894, A2 => n13466, B1 => n7235, B2 => 
                           n13462, ZN => n8101);
   U5741 : OAI22_X1 port map( A1 => n13900, A2 => n13466, B1 => n7236, B2 => 
                           n13463, ZN => n8102);
   U5742 : OAI22_X1 port map( A1 => n13906, A2 => n13466, B1 => n7237, B2 => 
                           n13463, ZN => n8103);
   U5743 : OAI22_X1 port map( A1 => n13912, A2 => n13466, B1 => n7238, B2 => 
                           n13463, ZN => n8104);
   U5744 : OAI22_X1 port map( A1 => n13918, A2 => n13466, B1 => n7239, B2 => 
                           n13463, ZN => n8105);
   U5745 : OAI22_X1 port map( A1 => n13924, A2 => n13466, B1 => n7240, B2 => 
                           n13463, ZN => n8106);
   U5746 : OAI22_X1 port map( A1 => n13930, A2 => n13466, B1 => n7241, B2 => 
                           n13463, ZN => n8107);
   U5747 : OAI22_X1 port map( A1 => n13936, A2 => n13466, B1 => n7242, B2 => 
                           n13463, ZN => n8108);
   U5748 : OAI22_X1 port map( A1 => n13942, A2 => n13466, B1 => n7243, B2 => 
                           n13463, ZN => n8109);
   U5749 : OAI22_X1 port map( A1 => n13948, A2 => n13465, B1 => n7244, B2 => 
                           n13463, ZN => n8110);
   U5750 : OAI22_X1 port map( A1 => n13954, A2 => n13465, B1 => n7245, B2 => 
                           n13463, ZN => n8111);
   U5751 : OAI22_X1 port map( A1 => n13960, A2 => n13465, B1 => n7246, B2 => 
                           n13463, ZN => n8112);
   U5752 : OAI22_X1 port map( A1 => n13966, A2 => n13465, B1 => n7247, B2 => 
                           n13463, ZN => n8113);
   U5753 : OAI22_X1 port map( A1 => n13827, A2 => n13515, B1 => n7022, B2 => 
                           n13510, ZN => n8346);
   U5754 : OAI22_X1 port map( A1 => n13834, A2 => n13515, B1 => n7023, B2 => 
                           n13510, ZN => n8347);
   U5755 : OAI22_X1 port map( A1 => n13840, A2 => n13515, B1 => n7024, B2 => 
                           n13510, ZN => n8348);
   U5756 : OAI22_X1 port map( A1 => n13846, A2 => n13515, B1 => n7025, B2 => 
                           n13510, ZN => n8349);
   U5757 : OAI22_X1 port map( A1 => n13852, A2 => n13515, B1 => n7026, B2 => 
                           n13510, ZN => n8350);
   U5758 : OAI22_X1 port map( A1 => n13858, A2 => n13515, B1 => n7027, B2 => 
                           n13510, ZN => n8351);
   U5759 : OAI22_X1 port map( A1 => n13864, A2 => n13515, B1 => n7028, B2 => 
                           n13510, ZN => n8352);
   U5760 : OAI22_X1 port map( A1 => n13870, A2 => n13515, B1 => n7029, B2 => 
                           n13510, ZN => n8353);
   U5761 : OAI22_X1 port map( A1 => n13876, A2 => n13514, B1 => n7030, B2 => 
                           n13510, ZN => n8354);
   U5762 : OAI22_X1 port map( A1 => n13882, A2 => n13514, B1 => n7031, B2 => 
                           n13510, ZN => n8355);
   U5763 : OAI22_X1 port map( A1 => n13888, A2 => n13514, B1 => n7032, B2 => 
                           n13510, ZN => n8356);
   U5764 : OAI22_X1 port map( A1 => n13894, A2 => n13514, B1 => n7033, B2 => 
                           n13510, ZN => n8357);
   U5765 : OAI22_X1 port map( A1 => n13900, A2 => n13514, B1 => n7034, B2 => 
                           n13511, ZN => n8358);
   U5766 : OAI22_X1 port map( A1 => n13906, A2 => n13514, B1 => n7035, B2 => 
                           n13511, ZN => n8359);
   U5767 : OAI22_X1 port map( A1 => n13912, A2 => n13514, B1 => n7036, B2 => 
                           n13511, ZN => n8360);
   U5768 : OAI22_X1 port map( A1 => n13918, A2 => n13514, B1 => n7037, B2 => 
                           n13511, ZN => n8361);
   U5769 : OAI22_X1 port map( A1 => n13924, A2 => n13514, B1 => n7038, B2 => 
                           n13511, ZN => n8362);
   U5770 : OAI22_X1 port map( A1 => n13930, A2 => n13514, B1 => n7039, B2 => 
                           n13511, ZN => n8363);
   U5771 : OAI22_X1 port map( A1 => n13936, A2 => n13514, B1 => n7040, B2 => 
                           n13511, ZN => n8364);
   U5772 : OAI22_X1 port map( A1 => n13942, A2 => n13514, B1 => n7041, B2 => 
                           n13511, ZN => n8365);
   U5773 : OAI22_X1 port map( A1 => n13948, A2 => n13513, B1 => n7042, B2 => 
                           n13511, ZN => n8366);
   U5774 : OAI22_X1 port map( A1 => n13954, A2 => n13513, B1 => n7043, B2 => 
                           n13511, ZN => n8367);
   U5775 : OAI22_X1 port map( A1 => n13960, A2 => n13513, B1 => n7044, B2 => 
                           n13511, ZN => n8368);
   U5776 : OAI22_X1 port map( A1 => n13966, A2 => n13513, B1 => n7045, B2 => 
                           n13511, ZN => n8369);
   U5777 : OAI22_X1 port map( A1 => n13827, A2 => n13521, B1 => n7256, B2 => 
                           n13516, ZN => n8378);
   U5778 : OAI22_X1 port map( A1 => n13826, A2 => n13623, B1 => n7046, B2 => 
                           n13618, ZN => n8922);
   U5779 : OAI22_X1 port map( A1 => n13832, A2 => n13623, B1 => n7047, B2 => 
                           n13618, ZN => n8923);
   U5780 : OAI22_X1 port map( A1 => n13838, A2 => n13623, B1 => n7048, B2 => 
                           n13618, ZN => n8924);
   U5781 : OAI22_X1 port map( A1 => n13844, A2 => n13623, B1 => n7049, B2 => 
                           n13618, ZN => n8925);
   U5782 : OAI22_X1 port map( A1 => n13850, A2 => n13623, B1 => n7050, B2 => 
                           n13618, ZN => n8926);
   U5783 : OAI22_X1 port map( A1 => n13856, A2 => n13623, B1 => n7051, B2 => 
                           n13618, ZN => n8927);
   U5784 : OAI22_X1 port map( A1 => n13862, A2 => n13623, B1 => n7052, B2 => 
                           n13618, ZN => n8928);
   U5785 : OAI22_X1 port map( A1 => n13868, A2 => n13623, B1 => n7053, B2 => 
                           n13618, ZN => n8929);
   U5786 : OAI22_X1 port map( A1 => n13874, A2 => n13622, B1 => n7054, B2 => 
                           n13618, ZN => n8930);
   U5787 : OAI22_X1 port map( A1 => n13880, A2 => n13622, B1 => n7055, B2 => 
                           n13618, ZN => n8931);
   U5788 : OAI22_X1 port map( A1 => n13886, A2 => n13622, B1 => n7056, B2 => 
                           n13618, ZN => n8932);
   U5789 : OAI22_X1 port map( A1 => n13892, A2 => n13622, B1 => n7057, B2 => 
                           n13618, ZN => n8933);
   U5790 : OAI22_X1 port map( A1 => n13898, A2 => n13622, B1 => n7058, B2 => 
                           n13619, ZN => n8934);
   U5791 : OAI22_X1 port map( A1 => n13904, A2 => n13622, B1 => n7059, B2 => 
                           n13619, ZN => n8935);
   U5792 : OAI22_X1 port map( A1 => n13910, A2 => n13622, B1 => n7060, B2 => 
                           n13619, ZN => n8936);
   U5793 : OAI22_X1 port map( A1 => n13916, A2 => n13622, B1 => n7061, B2 => 
                           n13619, ZN => n8937);
   U5794 : OAI22_X1 port map( A1 => n13922, A2 => n13622, B1 => n7062, B2 => 
                           n13619, ZN => n8938);
   U5795 : OAI22_X1 port map( A1 => n13928, A2 => n13622, B1 => n7063, B2 => 
                           n13619, ZN => n8939);
   U5796 : OAI22_X1 port map( A1 => n13934, A2 => n13622, B1 => n7064, B2 => 
                           n13619, ZN => n8940);
   U5797 : OAI22_X1 port map( A1 => n13940, A2 => n13622, B1 => n7065, B2 => 
                           n13619, ZN => n8941);
   U5798 : OAI22_X1 port map( A1 => n13946, A2 => n13621, B1 => n7066, B2 => 
                           n13619, ZN => n8942);
   U5799 : OAI22_X1 port map( A1 => n13952, A2 => n13621, B1 => n7067, B2 => 
                           n13619, ZN => n8943);
   U5800 : OAI22_X1 port map( A1 => n13958, A2 => n13621, B1 => n7068, B2 => 
                           n13619, ZN => n8944);
   U5801 : OAI22_X1 port map( A1 => n13964, A2 => n13621, B1 => n7069, B2 => 
                           n13619, ZN => n8945);
   U5802 : OAI22_X1 port map( A1 => n13826, A2 => n13641, B1 => n7153, B2 => 
                           n13636, ZN => n9018);
   U5803 : OAI22_X1 port map( A1 => n13832, A2 => n13641, B1 => n7154, B2 => 
                           n13636, ZN => n9019);
   U5804 : OAI22_X1 port map( A1 => n13838, A2 => n13641, B1 => n7155, B2 => 
                           n13636, ZN => n9020);
   U5805 : OAI22_X1 port map( A1 => n13844, A2 => n13641, B1 => n7156, B2 => 
                           n13636, ZN => n9021);
   U5806 : OAI22_X1 port map( A1 => n13850, A2 => n13641, B1 => n7157, B2 => 
                           n13636, ZN => n9022);
   U5807 : OAI22_X1 port map( A1 => n13856, A2 => n13641, B1 => n7158, B2 => 
                           n13636, ZN => n9023);
   U5808 : OAI22_X1 port map( A1 => n13862, A2 => n13641, B1 => n7159, B2 => 
                           n13636, ZN => n9024);
   U5809 : OAI22_X1 port map( A1 => n13825, A2 => n13677, B1 => n7070, B2 => 
                           n13672, ZN => n9210);
   U5810 : OAI22_X1 port map( A1 => n13831, A2 => n13677, B1 => n7071, B2 => 
                           n13672, ZN => n9211);
   U5811 : OAI22_X1 port map( A1 => n13837, A2 => n13677, B1 => n7072, B2 => 
                           n13672, ZN => n9212);
   U5812 : OAI22_X1 port map( A1 => n13843, A2 => n13677, B1 => n7073, B2 => 
                           n13672, ZN => n9213);
   U5813 : OAI22_X1 port map( A1 => n13849, A2 => n13677, B1 => n7074, B2 => 
                           n13672, ZN => n9214);
   U5814 : OAI22_X1 port map( A1 => n13855, A2 => n13677, B1 => n7075, B2 => 
                           n13672, ZN => n9215);
   U5815 : OAI22_X1 port map( A1 => n13861, A2 => n13677, B1 => n7076, B2 => 
                           n13672, ZN => n9216);
   U5816 : OAI22_X1 port map( A1 => n13867, A2 => n13677, B1 => n7077, B2 => 
                           n13672, ZN => n9217);
   U5817 : OAI22_X1 port map( A1 => n13873, A2 => n13676, B1 => n7078, B2 => 
                           n13672, ZN => n9218);
   U5818 : OAI22_X1 port map( A1 => n13879, A2 => n13676, B1 => n7079, B2 => 
                           n13672, ZN => n9219);
   U5819 : OAI22_X1 port map( A1 => n13885, A2 => n13676, B1 => n7080, B2 => 
                           n13672, ZN => n9220);
   U5820 : OAI22_X1 port map( A1 => n13891, A2 => n13676, B1 => n7081, B2 => 
                           n13672, ZN => n9221);
   U5821 : OAI22_X1 port map( A1 => n13897, A2 => n13676, B1 => n7082, B2 => 
                           n13673, ZN => n9222);
   U5822 : OAI22_X1 port map( A1 => n13903, A2 => n13676, B1 => n7083, B2 => 
                           n13673, ZN => n9223);
   U5823 : OAI22_X1 port map( A1 => n13909, A2 => n13676, B1 => n7084, B2 => 
                           n13673, ZN => n9224);
   U5824 : OAI22_X1 port map( A1 => n13915, A2 => n13676, B1 => n7085, B2 => 
                           n13673, ZN => n9225);
   U5825 : OAI22_X1 port map( A1 => n13921, A2 => n13676, B1 => n7086, B2 => 
                           n13673, ZN => n9226);
   U5826 : OAI22_X1 port map( A1 => n13927, A2 => n13676, B1 => n7087, B2 => 
                           n13673, ZN => n9227);
   U5827 : OAI22_X1 port map( A1 => n13933, A2 => n13676, B1 => n7088, B2 => 
                           n13673, ZN => n9228);
   U5828 : OAI22_X1 port map( A1 => n13939, A2 => n13676, B1 => n7089, B2 => 
                           n13673, ZN => n9229);
   U5829 : OAI22_X1 port map( A1 => n13945, A2 => n13675, B1 => n7090, B2 => 
                           n13673, ZN => n9230);
   U5830 : OAI22_X1 port map( A1 => n13951, A2 => n13675, B1 => n7091, B2 => 
                           n13673, ZN => n9231);
   U5831 : OAI22_X1 port map( A1 => n13957, A2 => n13675, B1 => n7092, B2 => 
                           n13673, ZN => n9232);
   U5832 : OAI22_X1 port map( A1 => n13963, A2 => n13675, B1 => n7093, B2 => 
                           n13673, ZN => n9233);
   U5833 : OAI22_X1 port map( A1 => n13825, A2 => n13695, B1 => n6998, B2 => 
                           n13690, ZN => n9306);
   U5834 : OAI22_X1 port map( A1 => n13831, A2 => n13695, B1 => n6999, B2 => 
                           n13690, ZN => n9307);
   U5835 : OAI22_X1 port map( A1 => n13837, A2 => n13695, B1 => n7000, B2 => 
                           n13690, ZN => n9308);
   U5836 : OAI22_X1 port map( A1 => n13843, A2 => n13695, B1 => n7001, B2 => 
                           n13690, ZN => n9309);
   U5837 : OAI22_X1 port map( A1 => n13849, A2 => n13695, B1 => n7002, B2 => 
                           n13690, ZN => n9310);
   U5838 : OAI22_X1 port map( A1 => n13855, A2 => n13695, B1 => n7003, B2 => 
                           n13690, ZN => n9311);
   U5839 : OAI22_X1 port map( A1 => n13861, A2 => n13695, B1 => n7004, B2 => 
                           n13690, ZN => n9312);
   U5840 : OAI22_X1 port map( A1 => n13867, A2 => n13695, B1 => n7005, B2 => 
                           n13690, ZN => n9313);
   U5841 : OAI22_X1 port map( A1 => n13873, A2 => n13694, B1 => n7094, B2 => 
                           n13690, ZN => n9314);
   U5842 : OAI22_X1 port map( A1 => n13879, A2 => n13694, B1 => n7095, B2 => 
                           n13690, ZN => n9315);
   U5843 : OAI22_X1 port map( A1 => n13885, A2 => n13694, B1 => n7096, B2 => 
                           n13690, ZN => n9316);
   U5844 : OAI22_X1 port map( A1 => n13891, A2 => n13694, B1 => n7097, B2 => 
                           n13690, ZN => n9317);
   U5845 : OAI22_X1 port map( A1 => n13897, A2 => n13694, B1 => n7098, B2 => 
                           n13691, ZN => n9318);
   U5846 : OAI22_X1 port map( A1 => n13903, A2 => n13694, B1 => n7099, B2 => 
                           n13691, ZN => n9319);
   U5847 : OAI22_X1 port map( A1 => n13909, A2 => n13694, B1 => n7100, B2 => 
                           n13691, ZN => n9320);
   U5848 : OAI22_X1 port map( A1 => n13915, A2 => n13694, B1 => n7101, B2 => 
                           n13691, ZN => n9321);
   U5849 : OAI22_X1 port map( A1 => n13921, A2 => n13694, B1 => n7102, B2 => 
                           n13691, ZN => n9322);
   U5850 : OAI22_X1 port map( A1 => n13927, A2 => n13694, B1 => n7103, B2 => 
                           n13691, ZN => n9323);
   U5851 : OAI22_X1 port map( A1 => n13933, A2 => n13694, B1 => n7104, B2 => 
                           n13691, ZN => n9324);
   U5852 : OAI22_X1 port map( A1 => n13825, A2 => n13731, B1 => n7105, B2 => 
                           n13726, ZN => n9498);
   U5853 : OAI22_X1 port map( A1 => n13831, A2 => n13731, B1 => n7106, B2 => 
                           n13726, ZN => n9499);
   U5854 : OAI22_X1 port map( A1 => n13837, A2 => n13731, B1 => n7107, B2 => 
                           n13726, ZN => n9500);
   U5855 : OAI22_X1 port map( A1 => n13843, A2 => n13731, B1 => n7108, B2 => 
                           n13726, ZN => n9501);
   U5856 : OAI22_X1 port map( A1 => n13849, A2 => n13731, B1 => n7109, B2 => 
                           n13726, ZN => n9502);
   U5857 : OAI22_X1 port map( A1 => n13855, A2 => n13731, B1 => n7110, B2 => 
                           n13726, ZN => n9503);
   U5858 : OAI22_X1 port map( A1 => n13861, A2 => n13731, B1 => n7111, B2 => 
                           n13726, ZN => n9504);
   U5859 : OAI22_X1 port map( A1 => n13867, A2 => n13731, B1 => n7112, B2 => 
                           n13726, ZN => n9505);
   U5860 : OAI22_X1 port map( A1 => n13873, A2 => n13730, B1 => n7113, B2 => 
                           n13726, ZN => n9506);
   U5861 : OAI22_X1 port map( A1 => n13879, A2 => n13730, B1 => n7114, B2 => 
                           n13726, ZN => n9507);
   U5862 : OAI22_X1 port map( A1 => n13885, A2 => n13730, B1 => n7115, B2 => 
                           n13726, ZN => n9508);
   U5863 : OAI22_X1 port map( A1 => n13891, A2 => n13730, B1 => n7116, B2 => 
                           n13726, ZN => n9509);
   U5864 : OAI22_X1 port map( A1 => n13897, A2 => n13730, B1 => n7117, B2 => 
                           n13727, ZN => n9510);
   U5865 : OAI22_X1 port map( A1 => n13903, A2 => n13730, B1 => n7118, B2 => 
                           n13727, ZN => n9511);
   U5866 : OAI22_X1 port map( A1 => n13909, A2 => n13730, B1 => n7119, B2 => 
                           n13727, ZN => n9512);
   U5867 : OAI22_X1 port map( A1 => n13915, A2 => n13730, B1 => n7120, B2 => 
                           n13727, ZN => n9513);
   U5868 : OAI22_X1 port map( A1 => n13921, A2 => n13730, B1 => n7121, B2 => 
                           n13727, ZN => n9514);
   U5869 : OAI22_X1 port map( A1 => n13927, A2 => n13730, B1 => n7122, B2 => 
                           n13727, ZN => n9515);
   U5870 : OAI22_X1 port map( A1 => n13933, A2 => n13730, B1 => n7123, B2 => 
                           n13727, ZN => n9516);
   U5871 : OAI22_X1 port map( A1 => n13939, A2 => n13730, B1 => n7124, B2 => 
                           n13727, ZN => n9517);
   U5872 : OAI22_X1 port map( A1 => n13945, A2 => n13729, B1 => n7125, B2 => 
                           n13727, ZN => n9518);
   U5873 : OAI22_X1 port map( A1 => n13951, A2 => n13729, B1 => n7126, B2 => 
                           n13727, ZN => n9519);
   U5874 : OAI22_X1 port map( A1 => n13957, A2 => n13729, B1 => n7127, B2 => 
                           n13727, ZN => n9520);
   U5875 : OAI22_X1 port map( A1 => n13963, A2 => n13729, B1 => n7128, B2 => 
                           n13727, ZN => n9521);
   U5876 : OAI22_X1 port map( A1 => n13824, A2 => n13785, B1 => n7129, B2 => 
                           n13780, ZN => n9786);
   U5877 : OAI22_X1 port map( A1 => n13830, A2 => n13785, B1 => n7130, B2 => 
                           n13780, ZN => n9787);
   U5878 : OAI22_X1 port map( A1 => n13836, A2 => n13785, B1 => n7131, B2 => 
                           n13780, ZN => n9788);
   U5879 : OAI22_X1 port map( A1 => n13842, A2 => n13785, B1 => n7132, B2 => 
                           n13780, ZN => n9789);
   U5880 : OAI22_X1 port map( A1 => n13848, A2 => n13785, B1 => n7133, B2 => 
                           n13780, ZN => n9790);
   U5881 : OAI22_X1 port map( A1 => n13854, A2 => n13785, B1 => n7134, B2 => 
                           n13780, ZN => n9791);
   U5882 : OAI22_X1 port map( A1 => n13860, A2 => n13785, B1 => n7135, B2 => 
                           n13780, ZN => n9792);
   U5883 : OAI22_X1 port map( A1 => n13866, A2 => n13785, B1 => n7136, B2 => 
                           n13780, ZN => n9793);
   U5884 : OAI22_X1 port map( A1 => n13872, A2 => n13784, B1 => n7137, B2 => 
                           n13780, ZN => n9794);
   U5885 : OAI22_X1 port map( A1 => n13878, A2 => n13784, B1 => n7138, B2 => 
                           n13780, ZN => n9795);
   U5886 : OAI22_X1 port map( A1 => n13884, A2 => n13784, B1 => n7139, B2 => 
                           n13780, ZN => n9796);
   U5887 : OAI22_X1 port map( A1 => n13890, A2 => n13784, B1 => n7140, B2 => 
                           n13780, ZN => n9797);
   U5888 : OAI22_X1 port map( A1 => n13896, A2 => n13784, B1 => n7141, B2 => 
                           n13781, ZN => n9798);
   U5889 : OAI22_X1 port map( A1 => n13902, A2 => n13784, B1 => n7142, B2 => 
                           n13781, ZN => n9799);
   U5890 : OAI22_X1 port map( A1 => n13908, A2 => n13784, B1 => n7143, B2 => 
                           n13781, ZN => n9800);
   U5891 : OAI22_X1 port map( A1 => n13914, A2 => n13784, B1 => n7144, B2 => 
                           n13781, ZN => n9801);
   U5892 : OAI22_X1 port map( A1 => n13920, A2 => n13784, B1 => n7145, B2 => 
                           n13781, ZN => n9802);
   U5893 : OAI22_X1 port map( A1 => n13926, A2 => n13784, B1 => n7146, B2 => 
                           n13781, ZN => n9803);
   U5894 : OAI22_X1 port map( A1 => n13932, A2 => n13784, B1 => n7147, B2 => 
                           n13781, ZN => n9804);
   U5895 : OAI22_X1 port map( A1 => n13938, A2 => n13784, B1 => n7148, B2 => 
                           n13781, ZN => n9805);
   U5896 : OAI22_X1 port map( A1 => n13944, A2 => n13783, B1 => n7149, B2 => 
                           n13781, ZN => n9806);
   U5897 : OAI22_X1 port map( A1 => n13950, A2 => n13783, B1 => n7150, B2 => 
                           n13781, ZN => n9807);
   U5898 : OAI22_X1 port map( A1 => n13956, A2 => n13783, B1 => n7151, B2 => 
                           n13781, ZN => n9808);
   U5899 : OAI22_X1 port map( A1 => n13962, A2 => n13783, B1 => n7152, B2 => 
                           n13781, ZN => n9809);
   U5900 : OAI22_X1 port map( A1 => n13828, A2 => n13473, B1 => n13468, B2 => 
                           n12726, ZN => n8122);
   U5901 : OAI22_X1 port map( A1 => n13834, A2 => n13473, B1 => n13468, B2 => 
                           n12727, ZN => n8123);
   U5902 : OAI22_X1 port map( A1 => n13840, A2 => n13473, B1 => n13468, B2 => 
                           n12728, ZN => n8124);
   U5903 : OAI22_X1 port map( A1 => n13846, A2 => n13473, B1 => n13468, B2 => 
                           n12729, ZN => n8125);
   U5904 : OAI22_X1 port map( A1 => n13852, A2 => n13473, B1 => n13468, B2 => 
                           n12730, ZN => n8126);
   U5905 : OAI22_X1 port map( A1 => n13858, A2 => n13473, B1 => n13468, B2 => 
                           n12731, ZN => n8127);
   U5906 : OAI22_X1 port map( A1 => n13864, A2 => n13473, B1 => n13468, B2 => 
                           n12732, ZN => n8128);
   U5907 : OAI22_X1 port map( A1 => n13870, A2 => n13473, B1 => n13468, B2 => 
                           n12733, ZN => n8129);
   U5908 : OAI22_X1 port map( A1 => n13876, A2 => n13472, B1 => n13468, B2 => 
                           n12734, ZN => n8130);
   U5909 : OAI22_X1 port map( A1 => n13882, A2 => n13472, B1 => n13468, B2 => 
                           n12735, ZN => n8131);
   U5910 : OAI22_X1 port map( A1 => n13888, A2 => n13472, B1 => n13468, B2 => 
                           n12736, ZN => n8132);
   U5911 : OAI22_X1 port map( A1 => n13894, A2 => n13472, B1 => n13468, B2 => 
                           n12737, ZN => n8133);
   U5912 : OAI22_X1 port map( A1 => n13900, A2 => n13472, B1 => n13469, B2 => 
                           n12738, ZN => n8134);
   U5913 : OAI22_X1 port map( A1 => n13906, A2 => n13472, B1 => n13469, B2 => 
                           n12739, ZN => n8135);
   U5914 : OAI22_X1 port map( A1 => n13912, A2 => n13472, B1 => n13469, B2 => 
                           n12740, ZN => n8136);
   U5915 : OAI22_X1 port map( A1 => n13918, A2 => n13472, B1 => n13469, B2 => 
                           n12741, ZN => n8137);
   U5916 : OAI22_X1 port map( A1 => n13924, A2 => n13472, B1 => n13469, B2 => 
                           n12742, ZN => n8138);
   U5917 : OAI22_X1 port map( A1 => n13930, A2 => n13472, B1 => n13469, B2 => 
                           n12743, ZN => n8139);
   U5918 : OAI22_X1 port map( A1 => n13936, A2 => n13472, B1 => n13469, B2 => 
                           n12744, ZN => n8140);
   U5919 : OAI22_X1 port map( A1 => n13942, A2 => n13472, B1 => n13469, B2 => 
                           n12745, ZN => n8141);
   U5920 : OAI22_X1 port map( A1 => n13948, A2 => n13471, B1 => n13469, B2 => 
                           n12746, ZN => n8142);
   U5921 : OAI22_X1 port map( A1 => n13954, A2 => n13471, B1 => n13469, B2 => 
                           n12747, ZN => n8143);
   U5922 : OAI22_X1 port map( A1 => n13960, A2 => n13471, B1 => n13469, B2 => 
                           n12748, ZN => n8144);
   U5923 : OAI22_X1 port map( A1 => n13966, A2 => n13471, B1 => n13469, B2 => 
                           n12749, ZN => n8145);
   U5924 : OAI22_X1 port map( A1 => n13828, A2 => n13479, B1 => n13474, B2 => 
                           n12750, ZN => n8154);
   U5925 : OAI22_X1 port map( A1 => n13834, A2 => n13479, B1 => n13474, B2 => 
                           n12751, ZN => n8155);
   U5926 : OAI22_X1 port map( A1 => n13840, A2 => n13479, B1 => n13474, B2 => 
                           n12752, ZN => n8156);
   U5927 : OAI22_X1 port map( A1 => n13846, A2 => n13479, B1 => n13474, B2 => 
                           n12753, ZN => n8157);
   U5928 : OAI22_X1 port map( A1 => n13852, A2 => n13479, B1 => n13474, B2 => 
                           n12754, ZN => n8158);
   U5929 : OAI22_X1 port map( A1 => n13858, A2 => n13479, B1 => n13474, B2 => 
                           n12755, ZN => n8159);
   U5930 : OAI22_X1 port map( A1 => n13864, A2 => n13479, B1 => n13474, B2 => 
                           n12756, ZN => n8160);
   U5931 : OAI22_X1 port map( A1 => n13870, A2 => n13479, B1 => n13474, B2 => 
                           n12757, ZN => n8161);
   U5932 : OAI22_X1 port map( A1 => n13876, A2 => n13478, B1 => n13474, B2 => 
                           n12758, ZN => n8162);
   U5933 : OAI22_X1 port map( A1 => n13882, A2 => n13478, B1 => n13474, B2 => 
                           n12759, ZN => n8163);
   U5934 : OAI22_X1 port map( A1 => n13888, A2 => n13478, B1 => n13474, B2 => 
                           n12760, ZN => n8164);
   U5935 : OAI22_X1 port map( A1 => n13894, A2 => n13478, B1 => n13474, B2 => 
                           n12761, ZN => n8165);
   U5936 : OAI22_X1 port map( A1 => n13900, A2 => n13478, B1 => n13475, B2 => 
                           n12762, ZN => n8166);
   U5937 : OAI22_X1 port map( A1 => n13906, A2 => n13478, B1 => n13475, B2 => 
                           n12763, ZN => n8167);
   U5938 : OAI22_X1 port map( A1 => n13912, A2 => n13478, B1 => n13475, B2 => 
                           n12764, ZN => n8168);
   U5939 : OAI22_X1 port map( A1 => n13918, A2 => n13478, B1 => n13475, B2 => 
                           n12765, ZN => n8169);
   U5940 : OAI22_X1 port map( A1 => n13924, A2 => n13478, B1 => n13475, B2 => 
                           n12766, ZN => n8170);
   U5941 : OAI22_X1 port map( A1 => n13930, A2 => n13478, B1 => n13475, B2 => 
                           n12767, ZN => n8171);
   U5942 : OAI22_X1 port map( A1 => n13936, A2 => n13478, B1 => n13475, B2 => 
                           n12768, ZN => n8172);
   U5943 : OAI22_X1 port map( A1 => n13942, A2 => n13478, B1 => n13475, B2 => 
                           n12769, ZN => n8173);
   U5944 : OAI22_X1 port map( A1 => n13948, A2 => n13477, B1 => n13475, B2 => 
                           n12770, ZN => n8174);
   U5945 : OAI22_X1 port map( A1 => n13954, A2 => n13477, B1 => n13475, B2 => 
                           n12771, ZN => n8175);
   U5946 : OAI22_X1 port map( A1 => n13960, A2 => n13477, B1 => n13475, B2 => 
                           n12772, ZN => n8176);
   U5947 : OAI22_X1 port map( A1 => n13966, A2 => n13477, B1 => n13475, B2 => 
                           n12773, ZN => n8177);
   U5948 : NAND4_X1 port map( A1 => n4624, A2 => n4625, A3 => n4626, A4 => 
                           n4627, ZN => n4623);
   U5949 : AOI221_X1 port map( B1 => n13101, B2 => n732, C1 => n13098, C2 => 
                           n15945, A => n4631, ZN => n4624);
   U5950 : AOI221_X1 port map( B1 => n13128, B2 => n731, C1 => n13125, C2 => 
                           n15937, A => n4629, ZN => n4626);
   U5951 : AOI221_X1 port map( B1 => n13116, B2 => n14082, C1 => n13113, C2 => 
                           n15604, A => n4630, ZN => n4625);
   U5952 : NAND4_X1 port map( A1 => n4587, A2 => n4588, A3 => n4589, A4 => 
                           n4590, ZN => n4586);
   U5953 : AOI221_X1 port map( B1 => n13101, B2 => n729, C1 => n13098, C2 => 
                           n15944, A => n4594, ZN => n4587);
   U5954 : AOI221_X1 port map( B1 => n13128, B2 => n728, C1 => n13125, C2 => 
                           n15936, A => n4592, ZN => n4589);
   U5955 : AOI221_X1 port map( B1 => n13116, B2 => n14081, C1 => n13113, C2 => 
                           n15603, A => n4593, ZN => n4588);
   U5956 : NAND4_X1 port map( A1 => n4550, A2 => n4551, A3 => n4552, A4 => 
                           n4553, ZN => n4549);
   U5957 : AOI221_X1 port map( B1 => n13101, B2 => n726, C1 => n13098, C2 => 
                           n15943, A => n4557, ZN => n4550);
   U5958 : AOI221_X1 port map( B1 => n13128, B2 => n725, C1 => n13125, C2 => 
                           n15935, A => n4555, ZN => n4552);
   U5959 : AOI221_X1 port map( B1 => n13116, B2 => n14080, C1 => n13113, C2 => 
                           n15602, A => n4556, ZN => n4551);
   U5960 : NAND4_X1 port map( A1 => n4513, A2 => n4514, A3 => n4515, A4 => 
                           n4516, ZN => n4512);
   U5961 : AOI221_X1 port map( B1 => n13101, B2 => n723, C1 => n13098, C2 => 
                           n15942, A => n4520, ZN => n4513);
   U5962 : AOI221_X1 port map( B1 => n13128, B2 => n722, C1 => n13125, C2 => 
                           n15934, A => n4518, ZN => n4515);
   U5963 : AOI221_X1 port map( B1 => n13116, B2 => n14079, C1 => n13113, C2 => 
                           n15601, A => n4519, ZN => n4514);
   U5964 : NAND4_X1 port map( A1 => n4476, A2 => n4477, A3 => n4478, A4 => 
                           n4479, ZN => n4475);
   U5965 : AOI221_X1 port map( B1 => n13101, B2 => n720, C1 => n13098, C2 => 
                           n15941, A => n4483, ZN => n4476);
   U5966 : AOI221_X1 port map( B1 => n13128, B2 => n719, C1 => n13125, C2 => 
                           n15933, A => n4481, ZN => n4478);
   U5967 : AOI221_X1 port map( B1 => n13116, B2 => n14078, C1 => n13113, C2 => 
                           n15600, A => n4482, ZN => n4477);
   U5968 : NAND4_X1 port map( A1 => n4439, A2 => n4440, A3 => n4441, A4 => 
                           n4442, ZN => n4438);
   U5969 : AOI221_X1 port map( B1 => n13101, B2 => n717, C1 => n13098, C2 => 
                           n15940, A => n4446, ZN => n4439);
   U5970 : AOI221_X1 port map( B1 => n13128, B2 => n716, C1 => n13125, C2 => 
                           n15932, A => n4444, ZN => n4441);
   U5971 : AOI221_X1 port map( B1 => n13116, B2 => n14077, C1 => n13113, C2 => 
                           n15599, A => n4445, ZN => n4440);
   U5972 : NAND4_X1 port map( A1 => n4330, A2 => n4331, A3 => n4332, A4 => 
                           n4333, ZN => n4329);
   U5973 : AOI221_X1 port map( B1 => n13101, B2 => n714, C1 => n13098, C2 => 
                           n15939, A => n4353, ZN => n4330);
   U5974 : AOI221_X1 port map( B1 => n13128, B2 => n713, C1 => n13125, C2 => 
                           n15931, A => n4342, ZN => n4332);
   U5975 : AOI221_X1 port map( B1 => n13116, B2 => n14076, C1 => n13113, C2 => 
                           n15598, A => n4347, ZN => n4331);
   U5976 : NAND4_X1 port map( A1 => n5650, A2 => n5651, A3 => n5654, A4 => 
                           n5656, ZN => n5649);
   U5977 : AOI221_X1 port map( B1 => n13099, B2 => n807, C1 => n13096, C2 => 
                           n16030, A => n5680, ZN => n5650);
   U5978 : AOI221_X1 port map( B1 => n13126, B2 => n806, C1 => n13123, C2 => 
                           n15994, A => n5670, ZN => n5654);
   U5979 : AOI221_X1 port map( B1 => n13114, B2 => n14107, C1 => n13111, C2 => 
                           n15921, A => n5678, ZN => n5651);
   U5980 : NAND4_X1 port map( A1 => n5589, A2 => n5590, A3 => n5591, A4 => 
                           n5594, ZN => n5588);
   U5981 : AOI221_X1 port map( B1 => n13099, B2 => n804, C1 => n13096, C2 => 
                           n16029, A => n5600, ZN => n5589);
   U5982 : AOI221_X1 port map( B1 => n13126, B2 => n803, C1 => n13123, C2 => 
                           n15993, A => n5598, ZN => n5591);
   U5983 : AOI221_X1 port map( B1 => n13114, B2 => n14106, C1 => n13111, C2 => 
                           n15920, A => n5599, ZN => n5590);
   U5984 : NAND4_X1 port map( A1 => n5528, A2 => n5529, A3 => n5530, A4 => 
                           n5531, ZN => n5526);
   U5985 : AOI221_X1 port map( B1 => n13099, B2 => n801, C1 => n13096, C2 => 
                           n16028, A => n5539, ZN => n5528);
   U5986 : AOI221_X1 port map( B1 => n13126, B2 => n800, C1 => n13123, C2 => 
                           n15992, A => n5536, ZN => n5530);
   U5987 : AOI221_X1 port map( B1 => n13114, B2 => n14105, C1 => n13111, C2 => 
                           n15919, A => n5538, ZN => n5529);
   U5988 : NAND4_X1 port map( A1 => n5466, A2 => n5468, A3 => n5469, A4 => 
                           n5470, ZN => n5464);
   U5989 : AOI221_X1 port map( B1 => n13099, B2 => n798, C1 => n13096, C2 => 
                           n16027, A => n5478, ZN => n5466);
   U5990 : AOI221_X1 port map( B1 => n13126, B2 => n797, C1 => n13123, C2 => 
                           n15991, A => n5474, ZN => n5469);
   U5991 : AOI221_X1 port map( B1 => n13114, B2 => n14104, C1 => n13111, C2 => 
                           n15918, A => n5476, ZN => n5468);
   U5992 : NAND4_X1 port map( A1 => n5410, A2 => n5411, A3 => n5412, A4 => 
                           n5414, ZN => n5409);
   U5993 : AOI221_X1 port map( B1 => n13099, B2 => n795, C1 => n13096, C2 => 
                           n16026, A => n5420, ZN => n5410);
   U5994 : AOI221_X1 port map( B1 => n13126, B2 => n794, C1 => n13123, C2 => 
                           n15990, A => n5418, ZN => n5412);
   U5995 : AOI221_X1 port map( B1 => n13114, B2 => n14103, C1 => n13111, C2 => 
                           n15917, A => n5419, ZN => n5411);
   U5996 : NAND4_X1 port map( A1 => n5364, A2 => n5365, A3 => n5366, A4 => 
                           n5367, ZN => n5363);
   U5997 : AOI221_X1 port map( B1 => n13099, B2 => n792, C1 => n13096, C2 => 
                           n16025, A => n5371, ZN => n5364);
   U5998 : AOI221_X1 port map( B1 => n13126, B2 => n791, C1 => n13123, C2 => 
                           n15989, A => n5369, ZN => n5366);
   U5999 : AOI221_X1 port map( B1 => n13114, B2 => n14102, C1 => n13111, C2 => 
                           n15916, A => n5370, ZN => n5365);
   U6000 : NAND4_X1 port map( A1 => n5327, A2 => n5328, A3 => n5329, A4 => 
                           n5330, ZN => n5326);
   U6001 : AOI221_X1 port map( B1 => n13099, B2 => n789, C1 => n13096, C2 => 
                           n16024, A => n5334, ZN => n5327);
   U6002 : AOI221_X1 port map( B1 => n13126, B2 => n788, C1 => n13123, C2 => 
                           n15988, A => n5332, ZN => n5329);
   U6003 : AOI221_X1 port map( B1 => n13114, B2 => n14101, C1 => n13111, C2 => 
                           n15915, A => n5333, ZN => n5328);
   U6004 : NAND4_X1 port map( A1 => n5290, A2 => n5291, A3 => n5292, A4 => 
                           n5293, ZN => n5289);
   U6005 : AOI221_X1 port map( B1 => n13099, B2 => n786, C1 => n13096, C2 => 
                           n16023, A => n5297, ZN => n5290);
   U6006 : AOI221_X1 port map( B1 => n13126, B2 => n785, C1 => n13123, C2 => 
                           n15987, A => n5295, ZN => n5292);
   U6007 : AOI221_X1 port map( B1 => n13114, B2 => n14100, C1 => n13111, C2 => 
                           n15914, A => n5296, ZN => n5291);
   U6008 : NAND4_X1 port map( A1 => n5253, A2 => n5254, A3 => n5255, A4 => 
                           n5256, ZN => n5252);
   U6009 : AOI221_X1 port map( B1 => n13099, B2 => n783, C1 => n13096, C2 => 
                           n16022, A => n5260, ZN => n5253);
   U6010 : AOI221_X1 port map( B1 => n13126, B2 => n782, C1 => n13123, C2 => 
                           n15986, A => n5258, ZN => n5255);
   U6011 : AOI221_X1 port map( B1 => n13114, B2 => n14099, C1 => n13111, C2 => 
                           n15913, A => n5259, ZN => n5254);
   U6012 : NAND4_X1 port map( A1 => n5216, A2 => n5217, A3 => n5218, A4 => 
                           n5219, ZN => n5215);
   U6013 : AOI221_X1 port map( B1 => n13099, B2 => n780, C1 => n13096, C2 => 
                           n16021, A => n5223, ZN => n5216);
   U6014 : AOI221_X1 port map( B1 => n13126, B2 => n779, C1 => n13123, C2 => 
                           n15985, A => n5221, ZN => n5218);
   U6015 : AOI221_X1 port map( B1 => n13114, B2 => n14098, C1 => n13111, C2 => 
                           n15912, A => n5222, ZN => n5217);
   U6016 : NAND4_X1 port map( A1 => n5179, A2 => n5180, A3 => n5181, A4 => 
                           n5182, ZN => n5178);
   U6017 : AOI221_X1 port map( B1 => n13099, B2 => n777, C1 => n13096, C2 => 
                           n16020, A => n5186, ZN => n5179);
   U6018 : AOI221_X1 port map( B1 => n13126, B2 => n776, C1 => n13123, C2 => 
                           n15984, A => n5184, ZN => n5181);
   U6019 : AOI221_X1 port map( B1 => n13114, B2 => n14097, C1 => n13111, C2 => 
                           n15911, A => n5185, ZN => n5180);
   U6020 : NAND4_X1 port map( A1 => n5142, A2 => n5143, A3 => n5144, A4 => 
                           n5145, ZN => n5141);
   U6021 : AOI221_X1 port map( B1 => n13099, B2 => n774, C1 => n13096, C2 => 
                           n16019, A => n5149, ZN => n5142);
   U6022 : AOI221_X1 port map( B1 => n13126, B2 => n773, C1 => n13123, C2 => 
                           n15983, A => n5147, ZN => n5144);
   U6023 : AOI221_X1 port map( B1 => n13114, B2 => n14096, C1 => n13111, C2 => 
                           n15910, A => n5148, ZN => n5143);
   U6024 : NAND4_X1 port map( A1 => n5105, A2 => n5106, A3 => n5107, A4 => 
                           n5108, ZN => n5104);
   U6025 : AOI221_X1 port map( B1 => n13100, B2 => n771, C1 => n13097, C2 => 
                           n16018, A => n5112, ZN => n5105);
   U6026 : AOI221_X1 port map( B1 => n13127, B2 => n770, C1 => n13124, C2 => 
                           n15982, A => n5110, ZN => n5107);
   U6027 : AOI221_X1 port map( B1 => n13115, B2 => n14095, C1 => n13112, C2 => 
                           n15909, A => n5111, ZN => n5106);
   U6028 : NAND4_X1 port map( A1 => n5068, A2 => n5069, A3 => n5070, A4 => 
                           n5071, ZN => n5067);
   U6029 : AOI221_X1 port map( B1 => n13100, B2 => n768, C1 => n13097, C2 => 
                           n16017, A => n5075, ZN => n5068);
   U6030 : AOI221_X1 port map( B1 => n13127, B2 => n767, C1 => n13124, C2 => 
                           n15981, A => n5073, ZN => n5070);
   U6031 : AOI221_X1 port map( B1 => n13115, B2 => n14094, C1 => n13112, C2 => 
                           n15908, A => n5074, ZN => n5069);
   U6032 : NAND4_X1 port map( A1 => n5031, A2 => n5032, A3 => n5033, A4 => 
                           n5034, ZN => n5030);
   U6033 : AOI221_X1 port map( B1 => n13100, B2 => n765, C1 => n13097, C2 => 
                           n16016, A => n5038, ZN => n5031);
   U6034 : AOI221_X1 port map( B1 => n13127, B2 => n764, C1 => n13124, C2 => 
                           n15980, A => n5036, ZN => n5033);
   U6035 : AOI221_X1 port map( B1 => n13115, B2 => n14093, C1 => n13112, C2 => 
                           n15907, A => n5037, ZN => n5032);
   U6036 : NAND4_X1 port map( A1 => n4994, A2 => n4995, A3 => n4996, A4 => 
                           n4997, ZN => n4993);
   U6037 : AOI221_X1 port map( B1 => n13100, B2 => n762, C1 => n13097, C2 => 
                           n16015, A => n5001, ZN => n4994);
   U6038 : AOI221_X1 port map( B1 => n13127, B2 => n761, C1 => n13124, C2 => 
                           n15979, A => n4999, ZN => n4996);
   U6039 : AOI221_X1 port map( B1 => n13115, B2 => n14092, C1 => n13112, C2 => 
                           n15906, A => n5000, ZN => n4995);
   U6040 : NAND4_X1 port map( A1 => n4957, A2 => n4958, A3 => n4959, A4 => 
                           n4960, ZN => n4956);
   U6041 : AOI221_X1 port map( B1 => n13100, B2 => n759, C1 => n13097, C2 => 
                           n16014, A => n4964, ZN => n4957);
   U6042 : AOI221_X1 port map( B1 => n13127, B2 => n758, C1 => n13124, C2 => 
                           n15978, A => n4962, ZN => n4959);
   U6043 : AOI221_X1 port map( B1 => n13115, B2 => n14091, C1 => n13112, C2 => 
                           n15905, A => n4963, ZN => n4958);
   U6044 : NAND4_X1 port map( A1 => n4920, A2 => n4921, A3 => n4922, A4 => 
                           n4923, ZN => n4919);
   U6045 : AOI221_X1 port map( B1 => n13100, B2 => n756, C1 => n13097, C2 => 
                           n16013, A => n4927, ZN => n4920);
   U6046 : AOI221_X1 port map( B1 => n13127, B2 => n755, C1 => n13124, C2 => 
                           n15977, A => n4925, ZN => n4922);
   U6047 : AOI221_X1 port map( B1 => n13115, B2 => n14090, C1 => n13112, C2 => 
                           n15904, A => n4926, ZN => n4921);
   U6048 : NAND4_X1 port map( A1 => n4883, A2 => n4884, A3 => n4885, A4 => 
                           n4886, ZN => n4882);
   U6049 : AOI221_X1 port map( B1 => n13100, B2 => n753, C1 => n13097, C2 => 
                           n16012, A => n4890, ZN => n4883);
   U6050 : AOI221_X1 port map( B1 => n13127, B2 => n752, C1 => n13124, C2 => 
                           n15976, A => n4888, ZN => n4885);
   U6051 : AOI221_X1 port map( B1 => n13115, B2 => n14089, C1 => n13112, C2 => 
                           n15903, A => n4889, ZN => n4884);
   U6052 : NAND4_X1 port map( A1 => n4846, A2 => n4847, A3 => n4848, A4 => 
                           n4849, ZN => n4845);
   U6053 : AOI221_X1 port map( B1 => n13100, B2 => n750, C1 => n13097, C2 => 
                           n16011, A => n4853, ZN => n4846);
   U6054 : AOI221_X1 port map( B1 => n13127, B2 => n749, C1 => n13124, C2 => 
                           n15975, A => n4851, ZN => n4848);
   U6055 : AOI221_X1 port map( B1 => n13115, B2 => n14088, C1 => n13112, C2 => 
                           n15902, A => n4852, ZN => n4847);
   U6056 : NAND4_X1 port map( A1 => n4809, A2 => n4810, A3 => n4811, A4 => 
                           n4812, ZN => n4808);
   U6057 : AOI221_X1 port map( B1 => n13100, B2 => n747, C1 => n13097, C2 => 
                           n16010, A => n4816, ZN => n4809);
   U6058 : AOI221_X1 port map( B1 => n13127, B2 => n746, C1 => n13124, C2 => 
                           n15974, A => n4814, ZN => n4811);
   U6059 : AOI221_X1 port map( B1 => n13115, B2 => n14087, C1 => n13112, C2 => 
                           n15901, A => n4815, ZN => n4810);
   U6060 : NAND4_X1 port map( A1 => n4772, A2 => n4773, A3 => n4774, A4 => 
                           n4775, ZN => n4771);
   U6061 : AOI221_X1 port map( B1 => n13100, B2 => n744, C1 => n13097, C2 => 
                           n16009, A => n4779, ZN => n4772);
   U6062 : AOI221_X1 port map( B1 => n13127, B2 => n743, C1 => n13124, C2 => 
                           n15973, A => n4777, ZN => n4774);
   U6063 : AOI221_X1 port map( B1 => n13115, B2 => n14086, C1 => n13112, C2 => 
                           n15900, A => n4778, ZN => n4773);
   U6064 : NAND4_X1 port map( A1 => n4735, A2 => n4736, A3 => n4737, A4 => 
                           n4738, ZN => n4734);
   U6065 : AOI221_X1 port map( B1 => n13100, B2 => n741, C1 => n13097, C2 => 
                           n16008, A => n4742, ZN => n4735);
   U6066 : AOI221_X1 port map( B1 => n13127, B2 => n740, C1 => n13124, C2 => 
                           n15972, A => n4740, ZN => n4737);
   U6067 : AOI221_X1 port map( B1 => n13115, B2 => n14085, C1 => n13112, C2 => 
                           n15899, A => n4741, ZN => n4736);
   U6068 : NAND4_X1 port map( A1 => n4698, A2 => n4699, A3 => n4700, A4 => 
                           n4701, ZN => n4697);
   U6069 : AOI221_X1 port map( B1 => n13100, B2 => n738, C1 => n13097, C2 => 
                           n16007, A => n4705, ZN => n4698);
   U6070 : AOI221_X1 port map( B1 => n13127, B2 => n737, C1 => n13124, C2 => 
                           n15971, A => n4703, ZN => n4700);
   U6071 : AOI221_X1 port map( B1 => n13115, B2 => n14084, C1 => n13112, C2 => 
                           n15898, A => n4704, ZN => n4699);
   U6072 : NAND4_X1 port map( A1 => n4661, A2 => n4662, A3 => n4663, A4 => 
                           n4664, ZN => n4660);
   U6073 : AOI221_X1 port map( B1 => n13101, B2 => n735, C1 => n13098, C2 => 
                           n15946, A => n4668, ZN => n4661);
   U6074 : AOI221_X1 port map( B1 => n13128, B2 => n734, C1 => n13125, C2 => 
                           n15938, A => n4666, ZN => n4663);
   U6075 : AOI221_X1 port map( B1 => n13116, B2 => n14083, C1 => n13113, C2 => 
                           n15605, A => n4667, ZN => n4662);
   U6076 : NAND4_X1 port map( A1 => n3163, A2 => n3164, A3 => n3165, A4 => 
                           n3166, ZN => n3153);
   U6077 : AOI221_X1 port map( B1 => n13275, B2 => n15863, C1 => n13272, C2 => 
                           n99, A => n3170, ZN => n3163);
   U6078 : AOI221_X1 port map( B1 => n13302, B2 => n15575, C1 => n13299, C2 => 
                           n15791, A => n3168, ZN => n3165);
   U6079 : AOI221_X1 port map( B1 => n13290, B2 => n14462, C1 => n13287, C2 => 
                           n15583, A => n3169, ZN => n3164);
   U6080 : NAND4_X1 port map( A1 => n3072, A2 => n3073, A3 => n3074, A4 => 
                           n3075, ZN => n3044);
   U6081 : AOI221_X1 port map( B1 => n13275, B2 => n15862, C1 => n13272, C2 => 
                           n97, A => n3095, ZN => n3072);
   U6082 : AOI221_X1 port map( B1 => n13302, B2 => n15574, C1 => n13299, C2 => 
                           n15790, A => n3084, ZN => n3074);
   U6083 : AOI221_X1 port map( B1 => n13290, B2 => n14461, C1 => n13287, C2 => 
                           n15582, A => n3089, ZN => n3073);
   U6084 : NAND4_X1 port map( A1 => n4447, A2 => n4448, A3 => n4449, A4 => 
                           n4450, ZN => n4437);
   U6085 : AOI221_X1 port map( B1 => n13047, B2 => n15863, C1 => n13044, C2 => 
                           n99, A => n4454, ZN => n4447);
   U6086 : AOI221_X1 port map( B1 => n13074, B2 => n15791, C1 => n13071, C2 => 
                           n15575, A => n4452, ZN => n4449);
   U6087 : AOI221_X1 port map( B1 => n13062, B2 => n14462, C1 => n13059, C2 => 
                           n15583, A => n4453, ZN => n4448);
   U6088 : NAND4_X1 port map( A1 => n4356, A2 => n4357, A3 => n4358, A4 => 
                           n4359, ZN => n4328);
   U6089 : AOI221_X1 port map( B1 => n13047, B2 => n15862, C1 => n13044, C2 => 
                           n97, A => n4379, ZN => n4356);
   U6090 : AOI221_X1 port map( B1 => n13074, B2 => n15790, C1 => n13071, C2 => 
                           n15574, A => n4368, ZN => n4358);
   U6091 : AOI221_X1 port map( B1 => n13062, B2 => n14461, C1 => n13059, C2 => 
                           n15582, A => n4373, ZN => n4357);
   U6092 : OAI21_X1 port map( B1 => n13149, B2 => n1576, A => n14026, ZN => 
                           n7546);
   U6093 : OAI21_X1 port map( B1 => n13149, B2 => n1545, A => n14024, ZN => 
                           n7608);
   U6094 : OAI21_X1 port map( B1 => n13377, B2 => n1544, A => n14024, ZN => 
                           n7610);
   U6095 : OAI21_X1 port map( B1 => n13377, B2 => n1513, A => n14022, ZN => 
                           n7672);
   U6096 : OAI21_X1 port map( B1 => n13148, B2 => n1575, A => n14026, ZN => 
                           n7548);
   U6097 : OAI21_X1 port map( B1 => n13148, B2 => n1574, A => n14026, ZN => 
                           n7550);
   U6098 : OAI21_X1 port map( B1 => n13148, B2 => n1573, A => n14026, ZN => 
                           n7552);
   U6099 : OAI21_X1 port map( B1 => n13148, B2 => n1572, A => n14026, ZN => 
                           n7554);
   U6100 : OAI21_X1 port map( B1 => n13147, B2 => n1571, A => n14026, ZN => 
                           n7556);
   U6101 : OAI21_X1 port map( B1 => n13147, B2 => n1570, A => n14026, ZN => 
                           n7558);
   U6102 : OAI21_X1 port map( B1 => n13147, B2 => n1569, A => n14026, ZN => 
                           n7560);
   U6103 : OAI21_X1 port map( B1 => n13147, B2 => n1568, A => n14026, ZN => 
                           n7562);
   U6104 : OAI21_X1 port map( B1 => n13147, B2 => n1566, A => n14026, ZN => 
                           n7566);
   U6105 : OAI21_X1 port map( B1 => n13147, B2 => n1564, A => n14026, ZN => 
                           n7570);
   U6106 : OAI21_X1 port map( B1 => n13147, B2 => n1561, A => n14025, ZN => 
                           n7576);
   U6107 : OAI21_X1 port map( B1 => n13147, B2 => n1560, A => n14025, ZN => 
                           n7578);
   U6108 : OAI21_X1 port map( B1 => n13147, B2 => n1559, A => n14025, ZN => 
                           n7580);
   U6109 : OAI21_X1 port map( B1 => n13147, B2 => n1558, A => n14025, ZN => 
                           n7582);
   U6110 : OAI21_X1 port map( B1 => n13147, B2 => n1557, A => n14025, ZN => 
                           n7584);
   U6111 : OAI21_X1 port map( B1 => n13147, B2 => n1556, A => n14025, ZN => 
                           n7586);
   U6112 : OAI21_X1 port map( B1 => n13148, B2 => n1555, A => n14025, ZN => 
                           n7588);
   U6113 : OAI21_X1 port map( B1 => n13147, B2 => n1554, A => n14025, ZN => 
                           n7590);
   U6114 : OAI21_X1 port map( B1 => n13148, B2 => n1553, A => n14025, ZN => 
                           n7592);
   U6115 : OAI21_X1 port map( B1 => n13148, B2 => n1552, A => n14025, ZN => 
                           n7594);
   U6116 : OAI21_X1 port map( B1 => n13148, B2 => n1551, A => n14025, ZN => 
                           n7596);
   U6117 : OAI21_X1 port map( B1 => n13148, B2 => n1550, A => n14024, ZN => 
                           n7598);
   U6118 : OAI21_X1 port map( B1 => n13148, B2 => n1549, A => n14024, ZN => 
                           n7600);
   U6119 : OAI21_X1 port map( B1 => n13148, B2 => n1548, A => n14024, ZN => 
                           n7602);
   U6120 : OAI21_X1 port map( B1 => n13148, B2 => n1547, A => n14024, ZN => 
                           n7604);
   U6121 : OAI21_X1 port map( B1 => n13148, B2 => n1546, A => n14024, ZN => 
                           n7606);
   U6122 : OAI21_X1 port map( B1 => n13376, B2 => n1543, A => n14024, ZN => 
                           n7612);
   U6123 : OAI21_X1 port map( B1 => n13376, B2 => n1542, A => n14024, ZN => 
                           n7614);
   U6124 : OAI21_X1 port map( B1 => n13376, B2 => n1541, A => n14024, ZN => 
                           n7616);
   U6125 : OAI21_X1 port map( B1 => n13376, B2 => n1540, A => n14024, ZN => 
                           n7618);
   U6126 : OAI21_X1 port map( B1 => n13375, B2 => n1539, A => n14024, ZN => 
                           n7620);
   U6127 : OAI21_X1 port map( B1 => n13375, B2 => n1538, A => n14023, ZN => 
                           n7622);
   U6128 : OAI21_X1 port map( B1 => n13375, B2 => n1537, A => n14023, ZN => 
                           n7624);
   U6129 : OAI21_X1 port map( B1 => n13375, B2 => n1536, A => n14023, ZN => 
                           n7626);
   U6130 : OAI21_X1 port map( B1 => n13375, B2 => n1534, A => n14023, ZN => 
                           n7630);
   U6131 : OAI21_X1 port map( B1 => n13375, B2 => n1532, A => n14023, ZN => 
                           n7634);
   U6132 : OAI21_X1 port map( B1 => n13375, B2 => n1529, A => n14023, ZN => 
                           n7640);
   U6133 : OAI21_X1 port map( B1 => n13375, B2 => n1528, A => n14024, ZN => 
                           n7642);
   U6134 : OAI21_X1 port map( B1 => n13375, B2 => n1527, A => n14023, ZN => 
                           n7644);
   U6135 : OAI21_X1 port map( B1 => n13375, B2 => n1526, A => n14023, ZN => 
                           n7646);
   U6136 : OAI21_X1 port map( B1 => n13375, B2 => n1525, A => n14022, ZN => 
                           n7648);
   U6137 : OAI21_X1 port map( B1 => n13375, B2 => n1524, A => n14023, ZN => 
                           n7650);
   U6138 : OAI21_X1 port map( B1 => n13376, B2 => n1523, A => n14022, ZN => 
                           n7652);
   U6139 : OAI21_X1 port map( B1 => n13375, B2 => n1522, A => n14022, ZN => 
                           n7654);
   U6140 : OAI21_X1 port map( B1 => n13376, B2 => n1521, A => n14022, ZN => 
                           n7656);
   U6141 : OAI21_X1 port map( B1 => n13376, B2 => n1520, A => n14022, ZN => 
                           n7658);
   U6142 : OAI21_X1 port map( B1 => n13376, B2 => n1519, A => n14022, ZN => 
                           n7660);
   U6143 : OAI21_X1 port map( B1 => n13376, B2 => n1518, A => n14022, ZN => 
                           n7662);
   U6144 : OAI21_X1 port map( B1 => n13376, B2 => n1517, A => n14022, ZN => 
                           n7664);
   U6145 : OAI21_X1 port map( B1 => n13376, B2 => n1516, A => n14022, ZN => 
                           n7666);
   U6146 : OAI21_X1 port map( B1 => n13376, B2 => n1515, A => n14022, ZN => 
                           n7668);
   U6147 : OAI21_X1 port map( B1 => n13376, B2 => n1514, A => n14022, ZN => 
                           n7670);
   U6148 : OAI21_X1 port map( B1 => n13146, B2 => n1567, A => n14026, ZN => 
                           n7564);
   U6149 : OAI21_X1 port map( B1 => n13146, B2 => n1565, A => n14026, ZN => 
                           n7568);
   U6150 : OAI21_X1 port map( B1 => n13146, B2 => n1563, A => n14025, ZN => 
                           n7572);
   U6151 : OAI21_X1 port map( B1 => n13146, B2 => n1562, A => n14025, ZN => 
                           n7574);
   U6152 : OAI21_X1 port map( B1 => n13374, B2 => n1535, A => n14023, ZN => 
                           n7628);
   U6153 : OAI21_X1 port map( B1 => n13374, B2 => n1533, A => n14023, ZN => 
                           n7632);
   U6154 : OAI21_X1 port map( B1 => n13374, B2 => n1531, A => n14023, ZN => 
                           n7636);
   U6155 : OAI21_X1 port map( B1 => n13374, B2 => n1530, A => n14023, ZN => 
                           n7638);
   U6156 : OAI22_X1 port map( A1 => n13828, A2 => n13431, B1 => n13426, B2 => 
                           n12774, ZN => n7898);
   U6157 : OAI22_X1 port map( A1 => n13835, A2 => n13431, B1 => n13426, B2 => 
                           n12775, ZN => n7899);
   U6158 : OAI22_X1 port map( A1 => n13841, A2 => n13431, B1 => n13426, B2 => 
                           n12776, ZN => n7900);
   U6159 : OAI22_X1 port map( A1 => n13847, A2 => n13431, B1 => n13426, B2 => 
                           n12777, ZN => n7901);
   U6160 : OAI22_X1 port map( A1 => n13853, A2 => n13431, B1 => n13426, B2 => 
                           n12778, ZN => n7902);
   U6161 : OAI22_X1 port map( A1 => n13859, A2 => n13431, B1 => n13426, B2 => 
                           n12779, ZN => n7903);
   U6162 : OAI22_X1 port map( A1 => n13865, A2 => n13431, B1 => n13426, B2 => 
                           n12780, ZN => n7904);
   U6163 : OAI22_X1 port map( A1 => n13871, A2 => n13431, B1 => n13426, B2 => 
                           n12781, ZN => n7905);
   U6164 : OAI22_X1 port map( A1 => n13877, A2 => n13430, B1 => n13426, B2 => 
                           n12782, ZN => n7906);
   U6165 : OAI22_X1 port map( A1 => n13883, A2 => n13430, B1 => n13426, B2 => 
                           n12783, ZN => n7907);
   U6166 : OAI22_X1 port map( A1 => n13889, A2 => n13430, B1 => n13426, B2 => 
                           n12784, ZN => n7908);
   U6167 : OAI22_X1 port map( A1 => n13895, A2 => n13430, B1 => n13426, B2 => 
                           n12785, ZN => n7909);
   U6168 : OAI22_X1 port map( A1 => n13901, A2 => n13430, B1 => n13427, B2 => 
                           n12786, ZN => n7910);
   U6169 : OAI22_X1 port map( A1 => n13907, A2 => n13430, B1 => n13427, B2 => 
                           n12787, ZN => n7911);
   U6170 : OAI22_X1 port map( A1 => n13913, A2 => n13430, B1 => n13427, B2 => 
                           n12788, ZN => n7912);
   U6171 : OAI22_X1 port map( A1 => n13919, A2 => n13430, B1 => n13427, B2 => 
                           n12789, ZN => n7913);
   U6172 : OAI22_X1 port map( A1 => n13925, A2 => n13430, B1 => n13427, B2 => 
                           n12790, ZN => n7914);
   U6173 : OAI22_X1 port map( A1 => n13931, A2 => n13430, B1 => n13427, B2 => 
                           n12791, ZN => n7915);
   U6174 : OAI22_X1 port map( A1 => n13937, A2 => n13430, B1 => n13427, B2 => 
                           n12792, ZN => n7916);
   U6175 : OAI22_X1 port map( A1 => n13943, A2 => n13430, B1 => n13427, B2 => 
                           n12793, ZN => n7917);
   U6176 : OAI22_X1 port map( A1 => n13949, A2 => n13429, B1 => n13427, B2 => 
                           n12794, ZN => n7918);
   U6177 : OAI22_X1 port map( A1 => n13955, A2 => n13429, B1 => n13427, B2 => 
                           n12795, ZN => n7919);
   U6178 : OAI22_X1 port map( A1 => n13961, A2 => n13429, B1 => n13427, B2 => 
                           n12796, ZN => n7920);
   U6179 : OAI22_X1 port map( A1 => n13967, A2 => n13429, B1 => n13427, B2 => 
                           n12797, ZN => n7921);
   U6180 : OAI22_X1 port map( A1 => n13973, A2 => n13429, B1 => n13428, B2 => 
                           n12798, ZN => n7922);
   U6181 : OAI22_X1 port map( A1 => n13979, A2 => n13429, B1 => n13428, B2 => 
                           n12799, ZN => n7923);
   U6182 : OAI22_X1 port map( A1 => n13985, A2 => n13429, B1 => n13428, B2 => 
                           n12800, ZN => n7924);
   U6183 : OAI22_X1 port map( A1 => n13991, A2 => n13429, B1 => n13428, B2 => 
                           n12801, ZN => n7925);
   U6184 : OAI22_X1 port map( A1 => n13997, A2 => n13429, B1 => n13428, B2 => 
                           n12802, ZN => n7926);
   U6185 : OAI22_X1 port map( A1 => n14003, A2 => n13429, B1 => n13428, B2 => 
                           n12803, ZN => n7927);
   U6186 : OAI22_X1 port map( A1 => n14009, A2 => n13429, B1 => n13428, B2 => 
                           n12804, ZN => n7928);
   U6187 : OAI22_X1 port map( A1 => n14018, A2 => n13429, B1 => n13428, B2 => 
                           n12805, ZN => n7929);
   U6188 : OAI22_X1 port map( A1 => n13828, A2 => n13461, B1 => n13456, B2 => 
                           n12806, ZN => n8058);
   U6189 : OAI22_X1 port map( A1 => n13834, A2 => n13461, B1 => n13456, B2 => 
                           n12807, ZN => n8059);
   U6190 : OAI22_X1 port map( A1 => n13840, A2 => n13461, B1 => n13456, B2 => 
                           n12808, ZN => n8060);
   U6191 : OAI22_X1 port map( A1 => n13846, A2 => n13461, B1 => n13456, B2 => 
                           n12809, ZN => n8061);
   U6192 : OAI22_X1 port map( A1 => n13852, A2 => n13461, B1 => n13456, B2 => 
                           n12810, ZN => n8062);
   U6193 : OAI22_X1 port map( A1 => n13858, A2 => n13461, B1 => n13456, B2 => 
                           n12811, ZN => n8063);
   U6194 : OAI22_X1 port map( A1 => n13864, A2 => n13461, B1 => n13456, B2 => 
                           n12812, ZN => n8064);
   U6195 : OAI22_X1 port map( A1 => n13870, A2 => n13461, B1 => n13456, B2 => 
                           n12813, ZN => n8065);
   U6196 : OAI22_X1 port map( A1 => n13876, A2 => n13460, B1 => n13456, B2 => 
                           n12814, ZN => n8066);
   U6197 : OAI22_X1 port map( A1 => n13882, A2 => n13460, B1 => n13456, B2 => 
                           n12815, ZN => n8067);
   U6198 : OAI22_X1 port map( A1 => n13888, A2 => n13460, B1 => n13456, B2 => 
                           n12816, ZN => n8068);
   U6199 : OAI22_X1 port map( A1 => n13894, A2 => n13460, B1 => n13456, B2 => 
                           n12817, ZN => n8069);
   U6200 : OAI22_X1 port map( A1 => n13900, A2 => n13460, B1 => n13457, B2 => 
                           n12818, ZN => n8070);
   U6201 : OAI22_X1 port map( A1 => n13906, A2 => n13460, B1 => n13457, B2 => 
                           n12819, ZN => n8071);
   U6202 : OAI22_X1 port map( A1 => n13912, A2 => n13460, B1 => n13457, B2 => 
                           n12820, ZN => n8072);
   U6203 : OAI22_X1 port map( A1 => n13918, A2 => n13460, B1 => n13457, B2 => 
                           n12821, ZN => n8073);
   U6204 : OAI22_X1 port map( A1 => n13924, A2 => n13460, B1 => n13457, B2 => 
                           n12822, ZN => n8074);
   U6205 : OAI22_X1 port map( A1 => n13930, A2 => n13460, B1 => n13457, B2 => 
                           n12823, ZN => n8075);
   U6206 : OAI22_X1 port map( A1 => n13936, A2 => n13460, B1 => n13457, B2 => 
                           n12824, ZN => n8076);
   U6207 : OAI22_X1 port map( A1 => n13942, A2 => n13460, B1 => n13457, B2 => 
                           n12825, ZN => n8077);
   U6208 : OAI22_X1 port map( A1 => n13948, A2 => n13459, B1 => n13457, B2 => 
                           n12826, ZN => n8078);
   U6209 : OAI22_X1 port map( A1 => n13954, A2 => n13459, B1 => n13457, B2 => 
                           n12827, ZN => n8079);
   U6210 : OAI22_X1 port map( A1 => n13960, A2 => n13459, B1 => n13457, B2 => 
                           n12828, ZN => n8080);
   U6211 : OAI22_X1 port map( A1 => n13966, A2 => n13459, B1 => n13457, B2 => 
                           n12829, ZN => n8081);
   U6212 : OAI22_X1 port map( A1 => n13972, A2 => n13459, B1 => n13458, B2 => 
                           n12830, ZN => n8082);
   U6213 : OAI22_X1 port map( A1 => n13978, A2 => n13459, B1 => n13458, B2 => 
                           n12831, ZN => n8083);
   U6214 : OAI22_X1 port map( A1 => n13984, A2 => n13459, B1 => n13458, B2 => 
                           n12832, ZN => n8084);
   U6215 : OAI22_X1 port map( A1 => n13990, A2 => n13459, B1 => n13458, B2 => 
                           n12833, ZN => n8085);
   U6216 : OAI22_X1 port map( A1 => n13996, A2 => n13459, B1 => n13458, B2 => 
                           n12834, ZN => n8086);
   U6217 : OAI22_X1 port map( A1 => n14002, A2 => n13459, B1 => n13458, B2 => 
                           n12835, ZN => n8087);
   U6218 : OAI22_X1 port map( A1 => n14008, A2 => n13459, B1 => n13458, B2 => 
                           n12836, ZN => n8088);
   U6219 : OAI22_X1 port map( A1 => n14017, A2 => n13459, B1 => n13458, B2 => 
                           n12837, ZN => n8089);
   U6220 : OAI22_X1 port map( A1 => n13827, A2 => n13539, B1 => n13534, B2 => 
                           n12838, ZN => n8474);
   U6221 : OAI22_X1 port map( A1 => n13833, A2 => n13539, B1 => n13534, B2 => 
                           n12839, ZN => n8475);
   U6222 : OAI22_X1 port map( A1 => n13839, A2 => n13539, B1 => n13534, B2 => 
                           n12840, ZN => n8476);
   U6223 : OAI22_X1 port map( A1 => n13845, A2 => n13539, B1 => n13534, B2 => 
                           n12841, ZN => n8477);
   U6224 : OAI22_X1 port map( A1 => n13851, A2 => n13539, B1 => n13534, B2 => 
                           n12842, ZN => n8478);
   U6225 : OAI22_X1 port map( A1 => n13857, A2 => n13539, B1 => n13534, B2 => 
                           n12843, ZN => n8479);
   U6226 : OAI22_X1 port map( A1 => n13863, A2 => n13539, B1 => n13534, B2 => 
                           n12844, ZN => n8480);
   U6227 : OAI22_X1 port map( A1 => n13869, A2 => n13539, B1 => n13534, B2 => 
                           n12845, ZN => n8481);
   U6228 : OAI22_X1 port map( A1 => n13875, A2 => n13538, B1 => n13534, B2 => 
                           n12846, ZN => n8482);
   U6229 : OAI22_X1 port map( A1 => n13881, A2 => n13538, B1 => n13534, B2 => 
                           n12847, ZN => n8483);
   U6230 : OAI22_X1 port map( A1 => n13887, A2 => n13538, B1 => n13534, B2 => 
                           n12848, ZN => n8484);
   U6231 : OAI22_X1 port map( A1 => n13893, A2 => n13538, B1 => n13534, B2 => 
                           n12849, ZN => n8485);
   U6232 : OAI22_X1 port map( A1 => n13899, A2 => n13538, B1 => n13535, B2 => 
                           n12850, ZN => n8486);
   U6233 : OAI22_X1 port map( A1 => n13905, A2 => n13538, B1 => n13535, B2 => 
                           n12851, ZN => n8487);
   U6234 : OAI22_X1 port map( A1 => n13911, A2 => n13538, B1 => n13535, B2 => 
                           n12852, ZN => n8488);
   U6235 : OAI22_X1 port map( A1 => n13917, A2 => n13538, B1 => n13535, B2 => 
                           n12853, ZN => n8489);
   U6236 : OAI22_X1 port map( A1 => n13923, A2 => n13538, B1 => n13535, B2 => 
                           n12854, ZN => n8490);
   U6237 : OAI22_X1 port map( A1 => n13929, A2 => n13538, B1 => n13535, B2 => 
                           n12855, ZN => n8491);
   U6238 : OAI22_X1 port map( A1 => n13935, A2 => n13538, B1 => n13535, B2 => 
                           n12856, ZN => n8492);
   U6239 : OAI22_X1 port map( A1 => n13941, A2 => n13538, B1 => n13535, B2 => 
                           n12857, ZN => n8493);
   U6240 : OAI22_X1 port map( A1 => n13947, A2 => n13537, B1 => n13535, B2 => 
                           n12858, ZN => n8494);
   U6241 : OAI22_X1 port map( A1 => n13953, A2 => n13537, B1 => n13535, B2 => 
                           n12859, ZN => n8495);
   U6242 : OAI22_X1 port map( A1 => n13959, A2 => n13537, B1 => n13535, B2 => 
                           n12860, ZN => n8496);
   U6243 : OAI22_X1 port map( A1 => n13965, A2 => n13537, B1 => n13535, B2 => 
                           n12861, ZN => n8497);
   U6244 : OAI22_X1 port map( A1 => n13971, A2 => n13537, B1 => n13536, B2 => 
                           n12862, ZN => n8498);
   U6245 : OAI22_X1 port map( A1 => n13977, A2 => n13537, B1 => n13536, B2 => 
                           n12863, ZN => n8499);
   U6246 : OAI22_X1 port map( A1 => n13983, A2 => n13537, B1 => n13536, B2 => 
                           n12864, ZN => n8500);
   U6247 : OAI22_X1 port map( A1 => n13989, A2 => n13537, B1 => n13536, B2 => 
                           n12865, ZN => n8501);
   U6248 : OAI22_X1 port map( A1 => n13995, A2 => n13537, B1 => n13536, B2 => 
                           n12866, ZN => n8502);
   U6249 : OAI22_X1 port map( A1 => n14001, A2 => n13537, B1 => n13536, B2 => 
                           n12867, ZN => n8503);
   U6250 : OAI22_X1 port map( A1 => n14007, A2 => n13537, B1 => n13536, B2 => 
                           n12868, ZN => n8504);
   U6251 : OAI22_X1 port map( A1 => n14016, A2 => n13537, B1 => n13536, B2 => 
                           n12869, ZN => n8505);
   U6252 : OAI22_X1 port map( A1 => n13827, A2 => n13569, B1 => n13564, B2 => 
                           n12870, ZN => n8634);
   U6253 : OAI22_X1 port map( A1 => n13833, A2 => n13569, B1 => n13564, B2 => 
                           n12871, ZN => n8635);
   U6254 : OAI22_X1 port map( A1 => n13839, A2 => n13569, B1 => n13564, B2 => 
                           n12872, ZN => n8636);
   U6255 : OAI22_X1 port map( A1 => n13845, A2 => n13569, B1 => n13564, B2 => 
                           n12873, ZN => n8637);
   U6256 : OAI22_X1 port map( A1 => n13851, A2 => n13569, B1 => n13564, B2 => 
                           n12874, ZN => n8638);
   U6257 : OAI22_X1 port map( A1 => n13857, A2 => n13569, B1 => n13564, B2 => 
                           n12875, ZN => n8639);
   U6258 : OAI22_X1 port map( A1 => n13863, A2 => n13569, B1 => n13564, B2 => 
                           n12876, ZN => n8640);
   U6259 : OAI22_X1 port map( A1 => n13869, A2 => n13569, B1 => n13564, B2 => 
                           n12877, ZN => n8641);
   U6260 : OAI22_X1 port map( A1 => n13875, A2 => n13568, B1 => n13564, B2 => 
                           n12878, ZN => n8642);
   U6261 : OAI22_X1 port map( A1 => n13881, A2 => n13568, B1 => n13564, B2 => 
                           n12879, ZN => n8643);
   U6262 : OAI22_X1 port map( A1 => n13887, A2 => n13568, B1 => n13564, B2 => 
                           n12880, ZN => n8644);
   U6263 : OAI22_X1 port map( A1 => n13893, A2 => n13568, B1 => n13564, B2 => 
                           n12881, ZN => n8645);
   U6264 : OAI22_X1 port map( A1 => n13899, A2 => n13568, B1 => n13565, B2 => 
                           n12882, ZN => n8646);
   U6265 : OAI22_X1 port map( A1 => n13905, A2 => n13568, B1 => n13565, B2 => 
                           n12883, ZN => n8647);
   U6266 : OAI22_X1 port map( A1 => n13911, A2 => n13568, B1 => n13565, B2 => 
                           n12884, ZN => n8648);
   U6267 : OAI22_X1 port map( A1 => n13917, A2 => n13568, B1 => n13565, B2 => 
                           n12885, ZN => n8649);
   U6268 : OAI22_X1 port map( A1 => n13923, A2 => n13568, B1 => n13565, B2 => 
                           n12886, ZN => n8650);
   U6269 : OAI22_X1 port map( A1 => n13929, A2 => n13568, B1 => n13565, B2 => 
                           n12887, ZN => n8651);
   U6270 : OAI22_X1 port map( A1 => n13935, A2 => n13568, B1 => n13565, B2 => 
                           n12888, ZN => n8652);
   U6271 : OAI22_X1 port map( A1 => n13941, A2 => n13568, B1 => n13565, B2 => 
                           n12889, ZN => n8653);
   U6272 : OAI22_X1 port map( A1 => n13947, A2 => n13567, B1 => n13565, B2 => 
                           n12890, ZN => n8654);
   U6273 : OAI22_X1 port map( A1 => n13953, A2 => n13567, B1 => n13565, B2 => 
                           n12891, ZN => n8655);
   U6274 : OAI22_X1 port map( A1 => n13959, A2 => n13567, B1 => n13565, B2 => 
                           n12892, ZN => n8656);
   U6275 : OAI22_X1 port map( A1 => n13965, A2 => n13567, B1 => n13565, B2 => 
                           n12893, ZN => n8657);
   U6276 : OAI22_X1 port map( A1 => n13971, A2 => n13567, B1 => n13566, B2 => 
                           n12894, ZN => n8658);
   U6277 : OAI22_X1 port map( A1 => n13977, A2 => n13567, B1 => n13566, B2 => 
                           n12895, ZN => n8659);
   U6278 : OAI22_X1 port map( A1 => n13983, A2 => n13567, B1 => n13566, B2 => 
                           n12896, ZN => n8660);
   U6279 : OAI22_X1 port map( A1 => n13989, A2 => n13567, B1 => n13566, B2 => 
                           n12897, ZN => n8661);
   U6280 : OAI22_X1 port map( A1 => n13995, A2 => n13567, B1 => n13566, B2 => 
                           n12898, ZN => n8662);
   U6281 : OAI22_X1 port map( A1 => n14001, A2 => n13567, B1 => n13566, B2 => 
                           n12899, ZN => n8663);
   U6282 : OAI22_X1 port map( A1 => n14007, A2 => n13567, B1 => n13566, B2 => 
                           n12900, ZN => n8664);
   U6283 : OAI22_X1 port map( A1 => n14016, A2 => n13567, B1 => n13566, B2 => 
                           n12901, ZN => n8665);
   U6284 : OAI22_X1 port map( A1 => n13826, A2 => n13587, B1 => n13584, B2 => 
                           n12902, ZN => n8730);
   U6285 : OAI22_X1 port map( A1 => n13833, A2 => n13587, B1 => n13584, B2 => 
                           n12903, ZN => n8731);
   U6286 : OAI22_X1 port map( A1 => n13839, A2 => n13587, B1 => n13584, B2 => 
                           n12904, ZN => n8732);
   U6287 : OAI22_X1 port map( A1 => n13845, A2 => n13587, B1 => n13584, B2 => 
                           n12905, ZN => n8733);
   U6288 : OAI22_X1 port map( A1 => n13851, A2 => n13587, B1 => n13584, B2 => 
                           n12906, ZN => n8734);
   U6289 : OAI22_X1 port map( A1 => n13857, A2 => n13587, B1 => n13584, B2 => 
                           n12907, ZN => n8735);
   U6290 : OAI22_X1 port map( A1 => n13863, A2 => n13587, B1 => n13584, B2 => 
                           n12908, ZN => n8736);
   U6291 : OAI22_X1 port map( A1 => n13869, A2 => n13587, B1 => n13583, B2 => 
                           n12909, ZN => n8737);
   U6292 : OAI22_X1 port map( A1 => n13875, A2 => n13586, B1 => n13583, B2 => 
                           n12910, ZN => n8738);
   U6293 : OAI22_X1 port map( A1 => n13881, A2 => n13586, B1 => n13583, B2 => 
                           n12911, ZN => n8739);
   U6294 : OAI22_X1 port map( A1 => n13887, A2 => n13586, B1 => n13583, B2 => 
                           n12912, ZN => n8740);
   U6295 : OAI22_X1 port map( A1 => n13893, A2 => n13586, B1 => n13583, B2 => 
                           n12913, ZN => n8741);
   U6296 : OAI22_X1 port map( A1 => n13899, A2 => n13586, B1 => n13583, B2 => 
                           n12914, ZN => n8742);
   U6297 : OAI22_X1 port map( A1 => n13905, A2 => n13586, B1 => n13583, B2 => 
                           n12915, ZN => n8743);
   U6298 : OAI22_X1 port map( A1 => n13911, A2 => n13586, B1 => n13583, B2 => 
                           n12916, ZN => n8744);
   U6299 : OAI22_X1 port map( A1 => n13917, A2 => n13586, B1 => n13583, B2 => 
                           n12917, ZN => n8745);
   U6300 : OAI22_X1 port map( A1 => n13923, A2 => n13586, B1 => n13583, B2 => 
                           n12918, ZN => n8746);
   U6301 : OAI22_X1 port map( A1 => n13929, A2 => n13586, B1 => n13583, B2 => 
                           n12919, ZN => n8747);
   U6302 : OAI22_X1 port map( A1 => n13935, A2 => n13586, B1 => n13583, B2 => 
                           n12920, ZN => n8748);
   U6303 : OAI22_X1 port map( A1 => n13941, A2 => n13586, B1 => n13583, B2 => 
                           n12921, ZN => n8749);
   U6304 : BUF_X1 port map( A => ENABLE, Z => n14022);
   U6305 : BUF_X1 port map( A => ENABLE, Z => n14026);
   U6306 : BUF_X1 port map( A => ENABLE, Z => n14025);
   U6307 : BUF_X1 port map( A => ENABLE, Z => n14024);
   U6308 : BUF_X1 port map( A => ENABLE, Z => n14023);
   U6309 : NAND2_X1 port map( A1 => DATAIN(0), A2 => n13821, ZN => n2865);
   U6310 : NAND2_X1 port map( A1 => DATAIN(1), A2 => n13821, ZN => n2864);
   U6311 : NAND2_X1 port map( A1 => DATAIN(2), A2 => n13821, ZN => n2863);
   U6312 : NAND2_X1 port map( A1 => DATAIN(3), A2 => n13821, ZN => n2862);
   U6313 : NAND2_X1 port map( A1 => DATAIN(4), A2 => n13820, ZN => n2861);
   U6314 : NAND2_X1 port map( A1 => DATAIN(5), A2 => n13820, ZN => n2860);
   U6315 : NAND2_X1 port map( A1 => DATAIN(6), A2 => n13820, ZN => n2859);
   U6316 : NAND2_X1 port map( A1 => DATAIN(7), A2 => n13820, ZN => n2858);
   U6317 : NAND2_X1 port map( A1 => DATAIN(8), A2 => n13819, ZN => n2857);
   U6318 : NAND2_X1 port map( A1 => DATAIN(9), A2 => n13819, ZN => n2856);
   U6319 : NAND2_X1 port map( A1 => DATAIN(10), A2 => n13819, ZN => n2855);
   U6320 : NAND2_X1 port map( A1 => DATAIN(11), A2 => n13819, ZN => n2854);
   U6321 : NAND2_X1 port map( A1 => DATAIN(12), A2 => n13818, ZN => n2853);
   U6322 : NAND2_X1 port map( A1 => DATAIN(13), A2 => n13818, ZN => n2852);
   U6323 : NAND2_X1 port map( A1 => DATAIN(14), A2 => n13818, ZN => n2851);
   U6324 : NAND2_X1 port map( A1 => DATAIN(15), A2 => n13818, ZN => n2850);
   U6325 : NAND2_X1 port map( A1 => DATAIN(16), A2 => n13817, ZN => n2849);
   U6326 : NAND2_X1 port map( A1 => DATAIN(17), A2 => n13817, ZN => n2848);
   U6327 : NAND2_X1 port map( A1 => DATAIN(18), A2 => n13817, ZN => n2847);
   U6328 : NAND2_X1 port map( A1 => DATAIN(19), A2 => n13817, ZN => n2846);
   U6329 : NAND2_X1 port map( A1 => DATAIN(20), A2 => n13816, ZN => n2845);
   U6330 : NAND2_X1 port map( A1 => DATAIN(21), A2 => n13816, ZN => n2844);
   U6331 : NAND2_X1 port map( A1 => DATAIN(22), A2 => n13816, ZN => n2843);
   U6332 : NAND2_X1 port map( A1 => DATAIN(23), A2 => n13816, ZN => n2842);
   U6333 : NAND2_X1 port map( A1 => DATAIN(24), A2 => n13815, ZN => n2841);
   U6334 : NAND2_X1 port map( A1 => DATAIN(25), A2 => n13815, ZN => n2840);
   U6335 : NAND2_X1 port map( A1 => DATAIN(26), A2 => n13815, ZN => n2839);
   U6336 : NAND2_X1 port map( A1 => DATAIN(27), A2 => n13815, ZN => n2838);
   U6337 : NAND2_X1 port map( A1 => DATAIN(28), A2 => n13814, ZN => n2837);
   U6338 : NAND2_X1 port map( A1 => DATAIN(29), A2 => n13814, ZN => n2836);
   U6339 : NAND2_X1 port map( A1 => DATAIN(30), A2 => n13814, ZN => n2835);
   U6340 : NAND2_X1 port map( A1 => DATAIN(31), A2 => n13814, ZN => n2833);
   U6341 : INV_X1 port map( A => RESET, ZN => n16063);
   U6342 : BUF_X1 port map( A => n2866, Z => n13810);
   U6343 : NAND2_X1 port map( A1 => WR, A2 => n14022, ZN => n2866);
   U6344 : INV_X1 port map( A => RD2, ZN => n16074);
   U6345 : INV_X1 port map( A => RD1, ZN => n16073);
   U6346 : INV_X1 port map( A => WR, ZN => n16075);
   U6347 : INV_X1 port map( A => DATAIN(28), ZN => n16079);
   U6348 : INV_X1 port map( A => DATAIN(29), ZN => n16078);
   U6349 : INV_X1 port map( A => DATAIN(30), ZN => n16077);
   U6350 : INV_X1 port map( A => DATAIN(31), ZN => n16076);
   U6351 : INV_X1 port map( A => DATAIN(0), ZN => n16107);
   U6352 : INV_X1 port map( A => DATAIN(1), ZN => n16106);
   U6353 : INV_X1 port map( A => DATAIN(2), ZN => n16105);
   U6354 : INV_X1 port map( A => DATAIN(3), ZN => n16104);
   U6355 : INV_X1 port map( A => DATAIN(4), ZN => n16103);
   U6356 : INV_X1 port map( A => DATAIN(5), ZN => n16102);
   U6357 : INV_X1 port map( A => DATAIN(6), ZN => n16101);
   U6358 : INV_X1 port map( A => DATAIN(7), ZN => n16100);
   U6359 : INV_X1 port map( A => DATAIN(8), ZN => n16099);
   U6360 : INV_X1 port map( A => DATAIN(9), ZN => n16098);
   U6361 : INV_X1 port map( A => DATAIN(10), ZN => n16097);
   U6362 : INV_X1 port map( A => DATAIN(11), ZN => n16096);
   U6363 : INV_X1 port map( A => DATAIN(12), ZN => n16095);
   U6364 : INV_X1 port map( A => DATAIN(13), ZN => n16094);
   U6365 : INV_X1 port map( A => DATAIN(14), ZN => n16093);
   U6366 : INV_X1 port map( A => DATAIN(15), ZN => n16092);
   U6367 : INV_X1 port map( A => DATAIN(16), ZN => n16091);
   U6368 : INV_X1 port map( A => DATAIN(17), ZN => n16090);
   U6369 : INV_X1 port map( A => DATAIN(18), ZN => n16089);
   U6370 : INV_X1 port map( A => DATAIN(19), ZN => n16088);
   U6371 : INV_X1 port map( A => DATAIN(20), ZN => n16087);
   U6372 : INV_X1 port map( A => DATAIN(21), ZN => n16086);
   U6373 : INV_X1 port map( A => DATAIN(22), ZN => n16085);
   U6374 : INV_X1 port map( A => DATAIN(23), ZN => n16084);
   U6375 : INV_X1 port map( A => DATAIN(24), ZN => n16083);
   U6376 : INV_X1 port map( A => DATAIN(25), ZN => n16082);
   U6377 : INV_X1 port map( A => DATAIN(26), ZN => n16081);
   U6378 : INV_X1 port map( A => DATAIN(27), ZN => n16080);
   U6379 : NOR3_X4 port map( A1 => n16060, A2 => ADD_WR(6), A3 => n16059, ZN =>
                           n2982);
   U6380 : NOR3_X4 port map( A1 => ADD_WR(4), A2 => ADD_WR(6), A3 => n16059, ZN
                           => n2949);
   U6381 : NOR3_X4 port map( A1 => ADD_WR(5), A2 => ADD_WR(6), A3 => n16060, ZN
                           => n2916);
   U6382 : NOR3_X4 port map( A1 => ADD_WR(5), A2 => ADD_WR(6), A3 => ADD_WR(4),
                           ZN => n2868);
   U6383 : CLKBUF_X1 port map( A => n4325, Z => n13149);
   U6384 : CLKBUF_X1 port map( A => n3041, Z => n13377);
   U6385 : CLKBUF_X1 port map( A => n2865, Z => n13829);
   U6386 : CLKBUF_X1 port map( A => n2864, Z => n13835);
   U6387 : CLKBUF_X1 port map( A => n2863, Z => n13841);
   U6388 : CLKBUF_X1 port map( A => n2862, Z => n13847);
   U6389 : CLKBUF_X1 port map( A => n2861, Z => n13853);
   U6390 : CLKBUF_X1 port map( A => n2860, Z => n13859);
   U6391 : CLKBUF_X1 port map( A => n2859, Z => n13865);
   U6392 : CLKBUF_X1 port map( A => n2858, Z => n13871);
   U6393 : CLKBUF_X1 port map( A => n2857, Z => n13877);
   U6394 : CLKBUF_X1 port map( A => n2856, Z => n13883);
   U6395 : CLKBUF_X1 port map( A => n2855, Z => n13889);
   U6396 : CLKBUF_X1 port map( A => n2854, Z => n13895);
   U6397 : CLKBUF_X1 port map( A => n2853, Z => n13901);
   U6398 : CLKBUF_X1 port map( A => n2852, Z => n13907);
   U6399 : CLKBUF_X1 port map( A => n2851, Z => n13913);
   U6400 : CLKBUF_X1 port map( A => n2850, Z => n13919);
   U6401 : CLKBUF_X1 port map( A => n2849, Z => n13925);
   U6402 : CLKBUF_X1 port map( A => n2848, Z => n13931);
   U6403 : CLKBUF_X1 port map( A => n2847, Z => n13937);
   U6404 : CLKBUF_X1 port map( A => n2846, Z => n13943);
   U6405 : CLKBUF_X1 port map( A => n2845, Z => n13949);
   U6406 : CLKBUF_X1 port map( A => n2844, Z => n13955);
   U6407 : CLKBUF_X1 port map( A => n2843, Z => n13961);
   U6408 : CLKBUF_X1 port map( A => n2842, Z => n13967);
   U6409 : CLKBUF_X1 port map( A => n2841, Z => n13973);
   U6410 : CLKBUF_X1 port map( A => n2840, Z => n13979);
   U6411 : CLKBUF_X1 port map( A => n2839, Z => n13985);
   U6412 : CLKBUF_X1 port map( A => n2838, Z => n13991);
   U6413 : CLKBUF_X1 port map( A => n2837, Z => n13997);
   U6414 : CLKBUF_X1 port map( A => n2836, Z => n14003);
   U6415 : CLKBUF_X1 port map( A => n2835, Z => n14009);
   U6416 : CLKBUF_X1 port map( A => n2833, Z => n14018);
   U6417 : CLKBUF_X1 port map( A => ENABLE, Z => n14027);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_registerFile_TLE.all;

entity 
   translationUnit_RF_N8_M8_windowBlocks3_F4_NAddr_Windowed5_NAddr_Physical7 is

   port( clk, reset, enable, rd1, rd2, wr : in std_logic;  add_wr, add_rd1, 
         add_rd2 : in std_logic_vector (4 downto 0);  cwp : in std_logic_vector
         (3 downto 0);  add_wr_out, add_rd1_out, add_rd2_out : out 
         std_logic_vector (6 downto 0));

end translationUnit_RF_N8_M8_windowBlocks3_F4_NAddr_Windowed5_NAddr_Physical7;

architecture SYN_beh of 
   translationUnit_RF_N8_M8_windowBlocks3_F4_NAddr_Windowed5_NAddr_Physical7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal N49, N50, N97, N98, N127, N128, r31_B_AS_3_port, r31_B_AS_4_port, 
      r31_carry_4_port, r31_carry_5_port, r186_B_AS_3_port, r186_B_AS_4_port, 
      r186_carry_4_port, r186_carry_5_port, r32_B_AS_4_port, r32_carry_4_port, 
      r32_carry_5_port, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, 
      n25, n26, n27, n28, n29, n30, n33, n34, n35, n36, n37, n38, n39, n40, n41
      , n42, n43, n44, n45 : std_logic;

begin
   
   r31_U1_3 : FA_X1 port map( A => add_rd2(3), B => r31_B_AS_3_port, CI => n38,
                           CO => r31_carry_4_port, S => N127);
   r31_U1_4 : FA_X1 port map( A => add_rd2(4), B => r31_B_AS_4_port, CI => 
                           r31_carry_4_port, CO => r31_carry_5_port, S => N128)
                           ;
   r186_U1_3 : FA_X1 port map( A => add_wr(3), B => r186_B_AS_3_port, CI => n39
                           , CO => r186_carry_4_port, S => N49);
   r186_U1_4 : FA_X1 port map( A => add_wr(4), B => r186_B_AS_4_port, CI => 
                           r186_carry_4_port, CO => r186_carry_5_port, S => N50
                           );
   r32_U1_3 : FA_X1 port map( A => add_rd1(3), B => n37, CI => n30, CO => 
                           r32_carry_4_port, S => N97);
   r32_U1_4 : FA_X1 port map( A => add_rd1(4), B => r32_B_AS_4_port, CI => 
                           r32_carry_4_port, CO => r32_carry_5_port, S => N98);
   U9 : NOR2_X2 port map( A1 => n17, A2 => n33, ZN => add_wr_out(6));
   U56 : NAND3_X1 port map( A1 => n20, A2 => n42, A3 => add_wr(4), ZN => n16);
   U57 : NAND3_X1 port map( A1 => n20, A2 => n45, A3 => add_rd2(4), ZN => n15);
   U58 : XOR2_X1 port map( A => n27, B => n30, Z => n26);
   U3 : NOR2_X1 port map( A1 => n22, A2 => n33, ZN => add_rd2_out(6));
   U4 : NOR2_X1 port map( A1 => n26, A2 => n33, ZN => add_rd1_out(6));
   U5 : XNOR2_X1 port map( A => n39, B => n18, ZN => n17);
   U6 : NOR2_X1 port map( A1 => n19, A2 => n35, ZN => n18);
   U7 : XNOR2_X1 port map( A => n38, B => n23, ZN => n22);
   U8 : NOR2_X1 port map( A1 => n24, A2 => n34, ZN => n23);
   U10 : NAND2_X1 port map( A1 => r32_carry_5_port, A2 => n40, ZN => n27);
   U11 : NOR2_X1 port map( A1 => n33, A2 => n21, ZN => add_wr_out(5));
   U12 : XNOR2_X1 port map( A => n35, B => n19, ZN => n21);
   U13 : NOR2_X1 port map( A1 => n33, A2 => n25, ZN => add_rd2_out(5));
   U14 : XNOR2_X1 port map( A => n34, B => n24, ZN => n25);
   U15 : NOR2_X1 port map( A1 => n33, A2 => n28, ZN => add_rd1_out(5));
   U16 : XNOR2_X1 port map( A => r32_carry_5_port, B => n40, ZN => n28);
   U17 : AND2_X1 port map( A1 => N50, A2 => enable, ZN => add_wr_out(4));
   U18 : AND2_X1 port map( A1 => N128, A2 => enable, ZN => add_rd2_out(4));
   U19 : AND2_X1 port map( A1 => N98, A2 => enable, ZN => add_rd1_out(4));
   U20 : AND2_X1 port map( A1 => N127, A2 => enable, ZN => add_rd2_out(3));
   U21 : AND2_X1 port map( A1 => N97, A2 => enable, ZN => add_rd1_out(3));
   U22 : AND2_X1 port map( A1 => N49, A2 => enable, ZN => add_wr_out(3));
   U23 : INV_X1 port map( A => n15, ZN => n38);
   U24 : INV_X1 port map( A => n16, ZN => n39);
   U25 : INV_X1 port map( A => r31_carry_5_port, ZN => n34);
   U26 : INV_X1 port map( A => r186_carry_5_port, ZN => n35);
   U27 : AND2_X1 port map( A1 => add_rd1(0), A2 => enable, ZN => add_rd1_out(0)
                           );
   U28 : AND2_X1 port map( A1 => add_rd2(1), A2 => enable, ZN => add_rd2_out(1)
                           );
   U29 : AND2_X1 port map( A1 => add_rd1(1), A2 => enable, ZN => add_rd1_out(1)
                           );
   U30 : AND2_X1 port map( A1 => add_rd2(2), A2 => enable, ZN => add_rd2_out(2)
                           );
   U31 : AND2_X1 port map( A1 => add_rd1(2), A2 => enable, ZN => add_rd1_out(2)
                           );
   U32 : AND2_X1 port map( A1 => add_rd2(0), A2 => enable, ZN => add_rd2_out(0)
                           );
   U33 : AOI21_X1 port map( B1 => add_rd2(4), B2 => add_rd2(3), A => cwp(1), ZN
                           => n24);
   U34 : AOI21_X1 port map( B1 => add_wr(3), B2 => add_wr(4), A => cwp(1), ZN 
                           => n19);
   U35 : OAI21_X1 port map( B1 => n44, B2 => n45, A => n15, ZN => 
                           r31_B_AS_3_port);
   U36 : INV_X1 port map( A => add_rd2(4), ZN => n44);
   U37 : OAI21_X1 port map( B1 => n42, B2 => n41, A => n16, ZN => 
                           r186_B_AS_3_port);
   U38 : INV_X1 port map( A => add_wr(4), ZN => n41);
   U39 : NOR2_X1 port map( A1 => n37, A2 => n36, ZN => r32_B_AS_4_port);
   U40 : AND2_X1 port map( A1 => add_wr(0), A2 => enable, ZN => add_wr_out(0));
   U41 : AND2_X1 port map( A1 => add_wr(1), A2 => enable, ZN => add_wr_out(1));
   U42 : AND3_X1 port map( A1 => add_rd1(4), A2 => n43, A3 => n20, ZN => n30);
   U43 : INV_X1 port map( A => add_rd1(3), ZN => n43);
   U44 : INV_X1 port map( A => cwp(0), ZN => n36);
   U45 : NOR2_X1 port map( A1 => r31_B_AS_3_port, A2 => n36, ZN => 
                           r31_B_AS_4_port);
   U46 : NOR2_X1 port map( A1 => r186_B_AS_3_port, A2 => n36, ZN => 
                           r186_B_AS_4_port);
   U47 : AND2_X1 port map( A1 => add_wr(2), A2 => enable, ZN => add_wr_out(2));
   U48 : INV_X1 port map( A => n29, ZN => n40);
   U49 : AOI21_X1 port map( B1 => add_rd1(3), B2 => add_rd1(4), A => cwp(1), ZN
                           => n29);
   U50 : AND2_X1 port map( A1 => cwp(1), A2 => cwp(0), ZN => n20);
   U51 : INV_X1 port map( A => n14, ZN => n37);
   U52 : AOI21_X1 port map( B1 => add_rd1(3), B2 => add_rd1(4), A => n30, ZN =>
                           n14);
   U53 : INV_X1 port map( A => add_rd2(3), ZN => n45);
   U54 : INV_X1 port map( A => add_wr(3), ZN => n42);
   U55 : INV_X1 port map( A => enable, ZN => n33);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_registerFile_TLE.all;

entity controlUnit_RF_N8_M8_F4_windowBlocks3_NData32_NAddr_Windowed5 is

   port( clk, reset, enable : in std_logic;  cwpOut, swpOut : out 
         std_logic_vector (3 downto 0);  call, ret : in std_logic;  fill, spill
         : out std_logic;  MMUStrobe : in std_logic;  dataACK : out std_logic);

end controlUnit_RF_N8_M8_F4_windowBlocks3_NData32_NAddr_Windowed5;

architecture SYN_beh of 
   controlUnit_RF_N8_M8_F4_windowBlocks3_NData32_NAddr_Windowed5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component 
      controlUnit_RF_N8_M8_F4_windowBlocks3_NData32_NAddr_Windowed5_DW01_incdec_0
      port( A : in std_logic_vector (31 downto 0);  INC_DEC : in std_logic;  
            SUM : out std_logic_vector (31 downto 0));
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal cwpOut_3_port, cwpOut_2_port, cwpOut_1_port, cwpOut_0_port, 
      swpOut_3_port, swpOut_2_port, swpOut_1_port, swpOut_0_port, 
      need_to_fill_0_port, need_to_spill_0_port, nextState_2_port, 
      nextState_1_port, nextState_0_port, cansaveNext_3_port, 
      cansaveNext_2_port, cansaveNext_1_port, cansaveNext_0_port, 
      canrestoreNext_3_port, canrestoreNext_2_port, canrestoreNext_1_port, 
      canrestoreNext_0_port, actual_round_31_port, actual_round_30_port, 
      actual_round_29_port, actual_round_28_port, actual_round_27_port, 
      actual_round_26_port, actual_round_25_port, actual_round_24_port, 
      actual_round_23_port, actual_round_22_port, actual_round_21_port, 
      actual_round_20_port, actual_round_19_port, actual_round_18_port, 
      actual_round_17_port, actual_round_16_port, actual_round_15_port, 
      actual_round_14_port, actual_round_13_port, actual_round_12_port, 
      actual_round_11_port, actual_round_10_port, actual_round_9_port, 
      actual_round_8_port, actual_round_7_port, actual_round_6_port, 
      actual_round_5_port, actual_round_4_port, actual_round_3_port, 
      actual_round_2_port, actual_round_1_port, actual_round_0_port, N436, N437
      , N438, N440, N441, N442, N443, N444, N445, N446, N447, N448, N449, N450,
      N451, N452, N453, N454, N455, N456, N457, N458, N459, N460, N461, N462, 
      N463, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473, N474, 
      N475, N476, N477, N478, N479, N480, N481, N482, N483, N484, N485, N486, 
      N487, N488, N489, N490, N491, N492, N493, N494, N495, N496, N497, n65, 
      n66, n73, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, 
      n230, n4, n6, n8, n9, n192, n205, n214, n43, n44, n45, n46, n47, n48, n49
      , n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, 
      n64, n67, n68, n69, n70, n71, n72, n74, n75, n76, n77, n78, n79, n80, n81
      , n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, 
      n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n219, n231, n232, n233, n234, n235, n236, n237, n238, 
      n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, 
      n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, 
      n263, n264, n265, n266, n267, n268, n269, n270, n271, n_2218, n_2219 : 
      std_logic;

begin
   cwpOut <= ( cwpOut_3_port, cwpOut_2_port, cwpOut_1_port, cwpOut_0_port );
   swpOut <= ( swpOut_3_port, swpOut_2_port, swpOut_1_port, swpOut_0_port );
   
   cansaveNext_reg_2_inst : DLH_X1 port map( G => N442, D => N445, Q => 
                           cansaveNext_2_port);
   cansaveNext_reg_3_inst : DLH_X1 port map( G => N442, D => N446, Q => 
                           cansaveNext_3_port);
   cansave_reg_3_inst : DFF_X1 port map( D => n227, CK => clk, Q => n8, QN => 
                           n244);
   nextState_reg_1_inst : DLH_X1 port map( G => N447, D => N449, Q => 
                           nextState_1_port);
   nextState_reg_0_inst : DLH_X1 port map( G => N447, D => N448, Q => 
                           nextState_0_port);
   nextState_reg_2_inst : DLH_X1 port map( G => N447, D => N450, Q => 
                           nextState_2_port);
   swp_reg_0_inst : DLH_X1 port map( G => N460, D => N461, Q => swpOut_0_port);
   swp_reg_1_inst : DLH_X1 port map( G => N460, D => N462, Q => swpOut_1_port);
   actual_round_reg_31_inst : DLH_X1 port map( G => n233, D => N497, Q => 
                           actual_round_31_port);
   actual_round_reg_0_inst : DLH_X1 port map( G => n234, D => N466, Q => 
                           actual_round_0_port);
   actual_round_reg_1_inst : DLH_X1 port map( G => n233, D => N467, Q => 
                           actual_round_1_port);
   actual_round_reg_2_inst : DLH_X1 port map( G => n233, D => N468, Q => 
                           actual_round_2_port);
   actual_round_reg_3_inst : DLH_X1 port map( G => n233, D => N469, Q => 
                           actual_round_3_port);
   actual_round_reg_4_inst : DLH_X1 port map( G => n233, D => N470, Q => 
                           actual_round_4_port);
   actual_round_reg_5_inst : DLH_X1 port map( G => n233, D => N471, Q => 
                           actual_round_5_port);
   actual_round_reg_6_inst : DLH_X1 port map( G => n233, D => N472, Q => 
                           actual_round_6_port);
   actual_round_reg_7_inst : DLH_X1 port map( G => n233, D => N473, Q => 
                           actual_round_7_port);
   actual_round_reg_8_inst : DLH_X1 port map( G => n233, D => N474, Q => 
                           actual_round_8_port);
   actual_round_reg_9_inst : DLH_X1 port map( G => n233, D => N475, Q => 
                           actual_round_9_port);
   actual_round_reg_10_inst : DLH_X1 port map( G => n233, D => N476, Q => 
                           actual_round_10_port);
   actual_round_reg_11_inst : DLH_X1 port map( G => n232, D => N477, Q => 
                           actual_round_11_port);
   actual_round_reg_12_inst : DLH_X1 port map( G => n232, D => N478, Q => 
                           actual_round_12_port);
   actual_round_reg_13_inst : DLH_X1 port map( G => n232, D => N479, Q => 
                           actual_round_13_port);
   actual_round_reg_14_inst : DLH_X1 port map( G => n232, D => N480, Q => 
                           actual_round_14_port);
   actual_round_reg_15_inst : DLH_X1 port map( G => n232, D => N481, Q => 
                           actual_round_15_port);
   actual_round_reg_16_inst : DLH_X1 port map( G => n232, D => N482, Q => 
                           actual_round_16_port);
   actual_round_reg_17_inst : DLH_X1 port map( G => n232, D => N483, Q => 
                           actual_round_17_port);
   actual_round_reg_18_inst : DLH_X1 port map( G => n232, D => N484, Q => 
                           actual_round_18_port);
   actual_round_reg_19_inst : DLH_X1 port map( G => n232, D => N485, Q => 
                           actual_round_19_port);
   actual_round_reg_20_inst : DLH_X1 port map( G => n232, D => N486, Q => 
                           actual_round_20_port);
   actual_round_reg_21_inst : DLH_X1 port map( G => n232, D => N487, Q => 
                           actual_round_21_port);
   actual_round_reg_22_inst : DLH_X1 port map( G => n234, D => N488, Q => 
                           actual_round_22_port);
   actual_round_reg_23_inst : DLH_X1 port map( G => n234, D => N489, Q => 
                           actual_round_23_port);
   actual_round_reg_24_inst : DLH_X1 port map( G => n234, D => N490, Q => 
                           actual_round_24_port);
   actual_round_reg_25_inst : DLH_X1 port map( G => n234, D => N491, Q => 
                           actual_round_25_port);
   actual_round_reg_26_inst : DLH_X1 port map( G => n234, D => N492, Q => 
                           actual_round_26_port);
   actual_round_reg_27_inst : DLH_X1 port map( G => n234, D => N493, Q => 
                           actual_round_27_port);
   actual_round_reg_28_inst : DLH_X1 port map( G => n234, D => N494, Q => 
                           actual_round_28_port);
   actual_round_reg_29_inst : DLH_X1 port map( G => n234, D => N495, Q => 
                           actual_round_29_port);
   actual_round_reg_30_inst : DLH_X1 port map( G => n234, D => N496, Q => 
                           actual_round_30_port);
   swp_reg_2_inst : DLH_X1 port map( G => N460, D => N463, Q => swpOut_2_port);
   swp_reg_3_inst : DLH_X1 port map( G => N460, D => N464, Q => swpOut_3_port);
   need_to_spill_reg_0_inst : DLH_X1 port map( G => N438, D => n157, Q => 
                           need_to_spill_0_port);
   canrestoreNext_reg_0_inst : DLH_X1 port map( G => N442, D => N451, Q => 
                           canrestoreNext_0_port);
   canrestore_reg_0_inst : DFF_X1 port map( D => n223, CK => clk, Q => n9, QN 
                           => n259);
   canrestoreNext_reg_2_inst : DLH_X1 port map( G => N442, D => N453, Q => 
                           canrestoreNext_2_port);
   canrestoreNext_reg_3_inst : DLH_X1 port map( G => N442, D => N454, Q => 
                           canrestoreNext_3_port);
   canrestore_reg_3_inst : DFF_X1 port map( D => n220, CK => clk, Q => n6, QN 
                           => n260);
   need_to_fill_reg_0_inst : DLH_X1 port map( G => N436, D => N437, Q => 
                           need_to_fill_0_port);
   canrestoreNext_reg_1_inst : DLH_X1 port map( G => N442, D => N452, Q => 
                           canrestoreNext_1_port);
   spill_reg : DLH_X1 port map( G => N440, D => n158, Q => spill);
   fill_reg : DLH_X1 port map( G => N440, D => n159, Q => fill);
   dataACK_reg : DLH_X1 port map( G => N440, D => N441, Q => dataACK);
   cwp_reg_3_inst : DLH_X1 port map( G => N455, D => N459, Q => cwpOut_3_port);
   cwp_reg_0_inst : DLH_X1 port map( G => N455, D => N456, Q => cwpOut_0_port);
   cwp_reg_1_inst : DLH_X1 port map( G => N455, D => N457, Q => cwpOut_1_port);
   cansaveNext_reg_1_inst : DLH_X1 port map( G => N442, D => N444, Q => 
                           cansaveNext_1_port);
   cansaveNext_reg_0_inst : DLH_X1 port map( G => N442, D => N443, Q => 
                           cansaveNext_0_port);
   cwp_reg_2_inst : DLH_X1 port map( G => N455, D => N458, Q => cwpOut_2_port);
   cansave_reg_1_inst : DFF_X1 port map( D => n229, CK => clk, Q => n156, QN =>
                           n264);
   U183 : XOR2_X1 port map( A => n88, B => n89, Z => n85);
   U184 : XOR2_X1 port map( A => n119, B => n120, Z => n118);
   U185 : XOR2_X1 port map( A => n124, B => n125, Z => n75);
   U186 : XOR2_X1 port map( A => n127, B => n134, Z => n76);
   U187 : XOR2_X1 port map( A => n140, B => n137, Z => n77);
   U188 : NAND3_X1 port map( A1 => n142, A2 => n253, A3 => n145, ZN => n79);
   U189 : NAND3_X1 port map( A1 => n245, A2 => n111, A3 => n109, ZN => N442);
   U190 : NAND3_X1 port map( A1 => n150, A2 => n107, A3 => call, ZN => n145);
   U191 : NAND3_X1 port map( A1 => n151, A2 => n248, A3 => n152, ZN => n89);
   U192 : NAND3_X1 port map( A1 => n110, A2 => ret, A3 => n100, ZN => n152);
   U193 : NAND3_X1 port map( A1 => n249, A2 => n245, A3 => n74, ZN => N440);
   U194 : NAND3_X1 port map( A1 => n133, A2 => n244, A3 => n192, ZN => n107);
   r243 : 
                           controlUnit_RF_N8_M8_F4_windowBlocks3_NData32_NAddr_Windowed5_DW01_incdec_0 
                           port map( A(31) => actual_round_31_port, A(30) => 
                           actual_round_30_port, A(29) => actual_round_29_port,
                           A(28) => actual_round_28_port, A(27) => 
                           actual_round_27_port, A(26) => actual_round_26_port,
                           A(25) => actual_round_25_port, A(24) => 
                           actual_round_24_port, A(23) => actual_round_23_port,
                           A(22) => actual_round_22_port, A(21) => 
                           actual_round_21_port, A(20) => actual_round_20_port,
                           A(19) => actual_round_19_port, A(18) => 
                           actual_round_18_port, A(17) => actual_round_17_port,
                           A(16) => actual_round_16_port, A(15) => 
                           actual_round_15_port, A(14) => actual_round_14_port,
                           A(13) => actual_round_13_port, A(12) => 
                           actual_round_12_port, A(11) => actual_round_11_port,
                           A(10) => actual_round_10_port, A(9) => 
                           actual_round_9_port, A(8) => actual_round_8_port, 
                           A(7) => actual_round_7_port, A(6) => 
                           actual_round_6_port, A(5) => actual_round_5_port, 
                           A(4) => actual_round_4_port, A(3) => 
                           actual_round_3_port, A(2) => actual_round_2_port, 
                           A(1) => actual_round_1_port, A(0) => 
                           actual_round_0_port, INC_DEC => n231, SUM(31) => 
                           N497, SUM(30) => N496, SUM(29) => N495, SUM(28) => 
                           N494, SUM(27) => N493, SUM(26) => N492, SUM(25) => 
                           N491, SUM(24) => N490, SUM(23) => N489, SUM(22) => 
                           N488, SUM(21) => N487, SUM(20) => N486, SUM(19) => 
                           N485, SUM(18) => N484, SUM(17) => N483, SUM(16) => 
                           N482, SUM(15) => N481, SUM(14) => N480, SUM(13) => 
                           N479, SUM(12) => N478, SUM(11) => N477, SUM(10) => 
                           N476, SUM(9) => N475, SUM(8) => N474, SUM(7) => N473
                           , SUM(6) => N472, SUM(5) => N471, SUM(4) => N470, 
                           SUM(3) => N469, SUM(2) => N468, SUM(1) => N467, 
                           SUM(0) => N466);
   canrestore_reg_1_inst : DFF_X1 port map( D => n222, CK => clk, Q => n_2218, 
                           QN => n214);
   currentState_reg_1_inst : DFF_X1 port map( D => n225, CK => clk, Q => n265, 
                           QN => n65);
   canrestore_reg_2_inst : DFF_X1 port map( D => n221, CK => clk, Q => n262, QN
                           => n4);
   cansave_reg_2_inst : DFF_X1 port map( D => n228, CK => clk, Q => n_2219, QN 
                           => n192);
   currentState_reg_2_inst : DFF_X1 port map( D => n224, CK => clk, Q => n251, 
                           QN => n205);
   cansave_reg_0_inst : DFF_X1 port map( D => n230, CK => clk, Q => n263, QN =>
                           n73);
   currentState_reg_0_inst : DFF_X1 port map( D => n226, CK => clk, Q => n261, 
                           QN => n66);
   U3 : NOR3_X1 port map( A1 => n205, A2 => n66, A3 => n265, ZN => n159);
   U4 : NOR3_X1 port map( A1 => n261, A2 => n205, A3 => n265, ZN => n158);
   U5 : INV_X1 port map( A => n130, ZN => n248);
   U6 : INV_X1 port map( A => n103, ZN => n249);
   U7 : NAND2_X1 port map( A1 => n99, A2 => n248, ZN => n83);
   U8 : XNOR2_X1 port map( A => n238, B => n91, ZN => n94);
   U9 : AND2_X1 port map( A1 => n72, A2 => n99, ZN => n74);
   U10 : INV_X1 port map( A => n122, ZN => n243);
   U11 : AND2_X1 port map( A1 => n99, A2 => n247, ZN => n117);
   U12 : NOR2_X1 port map( A1 => n258, A2 => n250, ZN => N437);
   U13 : INV_X1 port map( A => n136, ZN => n240);
   U14 : BUF_X1 port map( A => N465, Z => n232);
   U15 : BUF_X1 port map( A => N465, Z => n233);
   U16 : BUF_X1 port map( A => N465, Z => n234);
   U17 : NAND2_X1 port map( A1 => n253, A2 => n245, ZN => N460);
   U18 : INV_X1 port map( A => n95, ZN => n247);
   U19 : NOR2_X1 port map( A1 => n74, A2 => n76, ZN => N458);
   U20 : NOR2_X1 port map( A1 => n74, A2 => n77, ZN => N457);
   U21 : INV_X1 port map( A => N441, ZN => n253);
   U22 : OR2_X1 port map( A1 => n235, A2 => n127, ZN => n126);
   U23 : NOR3_X1 port map( A1 => n261, A2 => n251, A3 => n265, ZN => n103);
   U24 : XNOR2_X1 port map( A => n240, B => n128, ZN => n134);
   U25 : XNOR2_X1 port map( A => n78, B => n136, ZN => n140);
   U26 : AOI21_X1 port map( B1 => n258, B2 => n146, A => n249, ZN => n95);
   U27 : OAI21_X1 port map( B1 => n252, B2 => n271, A => n142, ZN => n136);
   U28 : AOI21_X1 port map( B1 => n96, B2 => n89, A => n87, ZN => n91);
   U29 : NOR3_X1 port map( A1 => n249, A2 => n148, A3 => n269, ZN => n130);
   U30 : INV_X1 port map( A => n50, ZN => n266);
   U31 : INV_X1 port map( A => n80, ZN => n245);
   U32 : NAND2_X1 port map( A1 => n267, A2 => n50, ZN => n43);
   U33 : AOI22_X1 port map( A1 => n136, A2 => n137, B1 => n78, B2 => n138, ZN 
                           => n127);
   U34 : OR2_X1 port map( A1 => n137, A2 => n136, ZN => n138);
   U35 : NOR2_X1 port map( A1 => n110, A2 => n150, ZN => n99);
   U36 : NOR2_X1 port map( A1 => n246, A2 => n107, ZN => n157);
   U37 : OAI221_X1 port map( B1 => n248, B2 => n78, C1 => n117, C2 => n263, A 
                           => n245, ZN => N443);
   U38 : NOR2_X1 port map( A1 => n159, A2 => n158, ZN => n72);
   U39 : NAND2_X1 port map( A1 => n111, A2 => n145, ZN => n122);
   U40 : INV_X1 port map( A => n159, ZN => n252);
   U41 : AOI21_X1 port map( B1 => n219, B2 => n57, A => n271, ZN => N465);
   U42 : NAND2_X1 port map( A1 => n158, A2 => n255, ZN => n57);
   U43 : INV_X1 port map( A => n89, ZN => n238);
   U44 : INV_X1 port map( A => n110, ZN => n250);
   U45 : OAI22_X1 port map( A1 => n238, A2 => n256, B1 => n97, B2 => n98, ZN =>
                           N452);
   U46 : INV_X1 port map( A => n98, ZN => n256);
   U47 : NAND2_X1 port map( A1 => n257, A2 => n96, ZN => n98);
   U48 : AOI21_X1 port map( B1 => n238, B2 => n83, A => n95, ZN => n97);
   U49 : XNOR2_X1 port map( A => N467, B => n67, ZN => n64);
   U50 : NOR2_X1 port map( A1 => n271, A2 => n72, ZN => N441);
   U51 : INV_X1 port map( A => n158, ZN => n254);
   U52 : NAND2_X1 port map( A1 => n43, A2 => n50, ZN => n44);
   U53 : NAND2_X1 port map( A1 => n231, A2 => n68, ZN => n60);
   U54 : INV_X1 port map( A => n148, ZN => n258);
   U55 : INV_X1 port map( A => n150, ZN => n246);
   U56 : OAI211_X1 port map( C1 => n250, C2 => n149, A => n249, B => n155, ZN 
                           => N436);
   U57 : NOR2_X1 port map( A1 => N437, A2 => n159, ZN => n155);
   U58 : OAI211_X1 port map( C1 => n231, C2 => n68, A => n60, B => n245, ZN => 
                           N463);
   U59 : OAI211_X1 port map( C1 => n246, C2 => n268, A => n249, B => n154, ZN 
                           => N438);
   U60 : NOR2_X1 port map( A1 => n157, A2 => n158, ZN => n154);
   U61 : INV_X1 port map( A => n63, ZN => n255);
   U62 : INV_X1 port map( A => n87, ZN => n257);
   U63 : OAI21_X1 port map( B1 => n108, B2 => n268, A => n109, ZN => N449);
   U64 : AOI21_X1 port map( B1 => n100, B2 => n110, A => n241, ZN => n108);
   U65 : INV_X1 port map( A => n111, ZN => n241);
   U66 : NOR2_X1 port map( A1 => n74, A2 => n78, ZN => N456);
   U67 : OR3_X1 port map( A1 => n250, A2 => n148, A3 => n149, ZN => n142);
   U68 : NOR2_X1 port map( A1 => n74, A2 => n75, ZN => N459);
   U69 : INV_X1 port map( A => n85, ZN => n236);
   U70 : INV_X1 port map( A => n146, ZN => n269);
   U71 : AND2_X1 port map( A1 => n238, A2 => n145, ZN => n109);
   U72 : OR2_X1 port map( A1 => n79, A2 => n80, ZN => N455);
   U73 : INV_X1 port map( A => n128, ZN => n235);
   U74 : OAI211_X1 port map( C1 => n73, C2 => n43, A => n44, B => n45, ZN => 
                           n230);
   U75 : NAND2_X1 port map( A1 => cansaveNext_0_port, A2 => n43, ZN => n45);
   U76 : OAI211_X1 port map( C1 => n66, C2 => n43, A => n44, B => n49, ZN => 
                           n226);
   U77 : NAND2_X1 port map( A1 => nextState_0_port, A2 => n43, ZN => n49);
   U78 : OAI211_X1 port map( C1 => n43, C2 => n264, A => n44, B => n46, ZN => 
                           n229);
   U79 : NAND2_X1 port map( A1 => cansaveNext_1_port, A2 => n43, ZN => n46);
   U80 : OAI21_X1 port map( B1 => n205, B2 => n43, A => n52, ZN => n224);
   U81 : NAND2_X1 port map( A1 => nextState_2_port, A2 => n266, ZN => n52);
   U82 : OAI21_X1 port map( B1 => n43, B2 => n260, A => n56, ZN => n220);
   U83 : NAND2_X1 port map( A1 => canrestoreNext_3_port, A2 => n266, ZN => n56)
                           ;
   U84 : OAI21_X1 port map( B1 => n43, B2 => n259, A => n53, ZN => n223);
   U85 : NAND2_X1 port map( A1 => canrestoreNext_0_port, A2 => n266, ZN => n53)
                           ;
   U86 : OAI21_X1 port map( B1 => n43, B2 => n244, A => n48, ZN => n227);
   U87 : NAND2_X1 port map( A1 => cansaveNext_3_port, A2 => n266, ZN => n48);
   U88 : OAI21_X1 port map( B1 => n4, B2 => n43, A => n55, ZN => n221);
   U89 : NAND2_X1 port map( A1 => canrestoreNext_2_port, A2 => n266, ZN => n55)
                           ;
   U90 : OAI21_X1 port map( B1 => n192, B2 => n43, A => n47, ZN => n228);
   U91 : NAND2_X1 port map( A1 => cansaveNext_2_port, A2 => n266, ZN => n47);
   U92 : OAI21_X1 port map( B1 => n65, B2 => n43, A => n51, ZN => n225);
   U93 : NAND2_X1 port map( A1 => nextState_1_port, A2 => n266, ZN => n51);
   U94 : OAI21_X1 port map( B1 => n214, B2 => n43, A => n54, ZN => n222);
   U95 : NAND2_X1 port map( A1 => canrestoreNext_1_port, A2 => n266, ZN => n54)
                           ;
   U96 : NOR3_X1 port map( A1 => n65, A2 => n66, A3 => n251, ZN => n110);
   U97 : NOR3_X1 port map( A1 => n251, A2 => n66, A3 => n265, ZN => n80);
   U98 : NOR3_X1 port map( A1 => n251, A2 => n65, A3 => n261, ZN => n150);
   U99 : OAI22_X1 port map( A1 => actual_round_0_port, A2 => n255, B1 => N466, 
                           B2 => n63, ZN => n67);
   U100 : NOR3_X1 port map( A1 => n96, A2 => n6, A3 => n262, ZN => n148);
   U101 : OAI22_X1 port map( A1 => n73, A2 => n264, B1 => n133, B2 => n243, ZN 
                           => n121);
   U102 : XNOR2_X1 port map( A => n240, B => n129, ZN => n124);
   U103 : AOI22_X1 port map( A1 => n240, A2 => n126, B1 => n235, B2 => n127, ZN
                           => n125);
   U104 : AOI22_X1 port map( A1 => cwpOut_3_port, A2 => n79, B1 => n130, B2 => 
                           n8, ZN => n129);
   U105 : OAI21_X1 port map( B1 => n89, B2 => n239, A => n90, ZN => n88);
   U106 : INV_X1 port map( A => n91, ZN => n239);
   U107 : OAI21_X1 port map( B1 => n91, B2 => n238, A => n4, ZN => n90);
   U108 : OAI21_X1 port map( B1 => n73, B2 => n248, A => n147, ZN => n78);
   U109 : NAND2_X1 port map( A1 => cwpOut_0_port, A2 => n79, ZN => n147);
   U110 : NAND4_X1 port map( A1 => n146, A2 => n150, A3 => n101, A4 => n107, ZN
                           => n151);
   U111 : NOR2_X1 port map( A1 => n259, A2 => n214, ZN => n87);
   U112 : AOI22_X1 port map( A1 => n159, A2 => swpOut_2_port, B1 => n67, B2 => 
                           n158, ZN => n68);
   U113 : NOR2_X1 port map( A1 => n270, A2 => call, ZN => n146);
   U114 : OAI21_X1 port map( B1 => n192, B2 => n248, A => n135, ZN => n128);
   U115 : NAND2_X1 port map( A1 => cwpOut_2_port, A2 => n79, ZN => n135);
   U116 : NAND4_X1 port map( A1 => n103, A2 => call, A3 => n107, A4 => n270, ZN
                           => n111);
   U117 : OAI221_X1 port map( B1 => n100, B2 => n250, C1 => n246, C2 => n101, A
                           => n102, ZN => N450);
   U118 : AOI211_X1 port map( C1 => n103, C2 => n104, A => n157, B => n105, ZN 
                           => n102);
   U119 : OAI21_X1 port map( B1 => n269, B2 => n258, A => n106, ZN => n104);
   U120 : NOR3_X1 port map( A1 => n265, A2 => n205, A3 => MMUStrobe, ZN => n105
                           );
   U121 : OAI21_X1 port map( B1 => n264, B2 => n248, A => n141, ZN => n137);
   U122 : NAND2_X1 port map( A1 => cwpOut_1_port, A2 => n79, ZN => n141);
   U123 : OAI221_X1 port map( B1 => n112, B2 => n270, C1 => n100, C2 => n250, A
                           => n113, ZN => N448);
   U124 : NOR2_X1 port map( A1 => n114, A2 => n110, ZN => n112);
   U125 : AOI22_X1 port map( A1 => reset, A2 => n80, B1 => n159, B2 => n271, ZN
                           => n113);
   U126 : AOI21_X1 port map( B1 => n249, B2 => n115, A => call, ZN => n114);
   U127 : OAI221_X1 port map( B1 => n117, B2 => n139, C1 => n248, C2 => n77, A 
                           => n245, ZN => N444);
   U128 : AOI221_X1 port map( B1 => n133, B2 => n122, C1 => n143, C2 => n156, A
                           => n144, ZN => n139);
   U129 : XNOR2_X1 port map( A => n243, B => n73, ZN => n143);
   U130 : NOR3_X1 port map( A1 => n122, A2 => n156, A3 => n73, ZN => n144);
   U131 : NAND2_X1 port map( A1 => ret, A2 => n107, ZN => n149);
   U132 : NOR2_X1 port map( A1 => n263, A2 => n156, ZN => n133);
   U133 : NOR3_X1 port map( A1 => n247, A2 => n4, A3 => n257, ZN => n84);
   U134 : NAND4_X1 port map( A1 => n66, A2 => n205, A3 => n101, A4 => n107, ZN 
                           => n115);
   U135 : OAI22_X1 port map( A1 => n92, A2 => n262, B1 => n4, B2 => n93, ZN => 
                           N453);
   U136 : AOI22_X1 port map( A1 => n237, A2 => n83, B1 => n95, B2 => n87, ZN =>
                           n92);
   U137 : AOI22_X1 port map( A1 => n94, A2 => n83, B1 => n95, B2 => n257, ZN =>
                           n93);
   U138 : INV_X1 port map( A => n94, ZN => n237);
   U139 : OAI22_X1 port map( A1 => n81, A2 => n260, B1 => n6, B2 => n82, ZN => 
                           N454);
   U140 : AOI21_X1 port map( B1 => n85, B2 => n83, A => n86, ZN => n81);
   U141 : AOI21_X1 port map( B1 => n236, B2 => n83, A => n84, ZN => n82);
   U142 : AOI21_X1 port map( B1 => n87, B2 => n262, A => n247, ZN => n86);
   U143 : OAI22_X1 port map( A1 => n75, A2 => n248, B1 => n117, B2 => n118, ZN 
                           => N446);
   U144 : XNOR2_X1 port map( A => n243, B => n8, ZN => n120);
   U145 : OAI21_X1 port map( B1 => n121, B2 => n122, A => n123, ZN => n119);
   U146 : OAI22_X1 port map( A1 => n248, A2 => n76, B1 => n117, B2 => n131, ZN 
                           => N445);
   U147 : XNOR2_X1 port map( A => n121, B => n132, ZN => n131);
   U148 : XNOR2_X1 port map( A => n192, B => n122, ZN => n132);
   U149 : NAND2_X1 port map( A1 => enable, A2 => n267, ZN => n50);
   U150 : NAND2_X1 port map( A1 => swpOut_1_port, A2 => swpOut_0_port, ZN => 
                           n63);
   U151 : INV_X1 port map( A => call, ZN => n268);
   U152 : INV_X1 port map( A => MMUStrobe, ZN => n271);
   U153 : NAND4_X1 port map( A1 => n74, A2 => call, A3 => n116, A4 => ret, ZN 
                           => N447);
   U154 : NOR2_X1 port map( A1 => n80, A2 => n265, ZN => n116);
   U155 : XNOR2_X1 port map( A => actual_round_1_port, B => n67, ZN => n62);
   U156 : OAI21_X1 port map( B1 => n242, B2 => n243, A => n192, ZN => n123);
   U157 : INV_X1 port map( A => n121, ZN => n242);
   U158 : AND2_X1 port map( A1 => n153, A2 => n258, ZN => n100);
   U159 : NAND2_X1 port map( A1 => need_to_fill_0_port, A2 => n149, ZN => n153)
                           ;
   U160 : NAND2_X1 port map( A1 => need_to_spill_0_port, A2 => n268, ZN => n101
                           );
   U161 : NAND2_X1 port map( A1 => n214, A2 => n259, ZN => n96);
   U162 : AOI21_X1 port map( B1 => n99, B2 => n249, A => n9, ZN => N451);
   U163 : OAI21_X1 port map( B1 => swpOut_0_port, B2 => n72, A => n245, ZN => 
                           N461);
   U164 : INV_X1 port map( A => ret, ZN => n270);
   U165 : OR3_X1 port map( A1 => swpOut_0_port, A2 => swpOut_1_port, A3 => n252
                           , ZN => n219);
   U166 : INV_X1 port map( A => reset, ZN => n267);
   U167 : OR3_X1 port map( A1 => n107, A2 => ret, A3 => n268, ZN => n106);
   U168 : NAND2_X1 port map( A1 => n58, A2 => n245, ZN => N464);
   U169 : XNOR2_X1 port map( A => n59, B => n60, ZN => n58);
   U170 : AOI22_X1 port map( A1 => n61, A2 => n158, B1 => swpOut_3_port, B2 => 
                           n159, ZN => n59);
   U171 : AOI22_X1 port map( A1 => n62, A2 => n63, B1 => n255, B2 => n64, ZN =>
                           n61);
   U172 : NAND2_X1 port map( A1 => n245, A2 => n69, ZN => N462);
   U173 : OAI21_X1 port map( B1 => n70, B2 => n252, A => n71, ZN => n69);
   U174 : OAI21_X1 port map( B1 => n70, B2 => n254, A => n252, ZN => n71);
   U175 : XNOR2_X1 port map( A => swpOut_1_port, B => swpOut_0_port, ZN => n70)
                           ;
   U176 : INV_X1 port map( A => n219, ZN => n231);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_registerFile_TLE.all;

entity registerFile_TLE is

   port( clk, reset, enable, rd1, rd2, wr1 : in std_logic;  add_wr, add_rd1, 
         add_rd2 : in std_logic_vector (4 downto 0);  dataIn : in 
         std_logic_vector (31 downto 0);  dataOut1, dataOut2 : out 
         std_logic_vector (31 downto 0);  fill, spill : out std_logic;  call, 
         ret : in std_logic;  dataACK : out std_logic;  MMUStrobe : in 
         std_logic);

end registerFile_TLE;

architecture SYN_struct of registerFile_TLE is

   component physical_RF_NData32_NRegs72_NAddr7
      port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
            ADD_RD2 : in std_logic_vector (6 downto 0);  DATAIN : in 
            std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component 
      translationUnit_RF_N8_M8_windowBlocks3_F4_NAddr_Windowed5_NAddr_Physical7
      port( clk, reset, enable, rd1, rd2, wr : in std_logic;  add_wr, add_rd1, 
            add_rd2 : in std_logic_vector (4 downto 0);  cwp : in 
            std_logic_vector (3 downto 0);  add_wr_out, add_rd1_out, 
            add_rd2_out : out std_logic_vector (6 downto 0));
   end component;
   
   component controlUnit_RF_N8_M8_F4_windowBlocks3_NData32_NAddr_Windowed5
      port( clk, reset, enable : in std_logic;  cwpOut, swpOut : out 
            std_logic_vector (3 downto 0);  call, ret : in std_logic;  fill, 
            spill : out std_logic;  MMUStrobe : in std_logic;  dataACK : out 
            std_logic);
   end component;
   
   signal cwp_s_3_port, cwp_s_2_port, cwp_s_1_port, cwp_s_0_port, 
      add_wr_out_s_6_port, add_wr_out_s_5_port, add_wr_out_s_4_port, 
      add_wr_out_s_3_port, add_wr_out_s_2_port, add_wr_out_s_1_port, 
      add_wr_out_s_0_port, add_rd1_out_s_6_port, add_rd1_out_s_5_port, 
      add_rd1_out_s_4_port, add_rd1_out_s_3_port, add_rd1_out_s_2_port, 
      add_rd1_out_s_1_port, add_rd1_out_s_0_port, add_rd2_out_s_6_port, 
      add_rd2_out_s_5_port, add_rd2_out_s_4_port, add_rd2_out_s_3_port, 
      add_rd2_out_s_2_port, add_rd2_out_s_1_port, add_rd2_out_s_0_port, n_2220,
      n_2221, n_2222, n_2223 : std_logic;

begin
   
   contrU : controlUnit_RF_N8_M8_F4_windowBlocks3_NData32_NAddr_Windowed5 port 
                           map( clk => clk, reset => reset, enable => enable, 
                           cwpOut(3) => cwp_s_3_port, cwpOut(2) => cwp_s_2_port
                           , cwpOut(1) => cwp_s_1_port, cwpOut(0) => 
                           cwp_s_0_port, swpOut(3) => n_2220, swpOut(2) => 
                           n_2221, swpOut(1) => n_2222, swpOut(0) => n_2223, 
                           call => call, ret => ret, fill => fill, spill => 
                           spill, MMUStrobe => MMUStrobe, dataACK => dataACK);
   translU : 
                           translationUnit_RF_N8_M8_windowBlocks3_F4_NAddr_Windowed5_NAddr_Physical7 
                           port map( clk => clk, reset => reset, enable => 
                           enable, rd1 => rd1, rd2 => rd2, wr => wr1, add_wr(4)
                           => add_wr(4), add_wr(3) => add_wr(3), add_wr(2) => 
                           add_wr(2), add_wr(1) => add_wr(1), add_wr(0) => 
                           add_wr(0), add_rd1(4) => add_rd1(4), add_rd1(3) => 
                           add_rd1(3), add_rd1(2) => add_rd1(2), add_rd1(1) => 
                           add_rd1(1), add_rd1(0) => add_rd1(0), add_rd2(4) => 
                           add_rd2(4), add_rd2(3) => add_rd2(3), add_rd2(2) => 
                           add_rd2(2), add_rd2(1) => add_rd2(1), add_rd2(0) => 
                           add_rd2(0), cwp(3) => cwp_s_3_port, cwp(2) => 
                           cwp_s_2_port, cwp(1) => cwp_s_1_port, cwp(0) => 
                           cwp_s_0_port, add_wr_out(6) => add_wr_out_s_6_port, 
                           add_wr_out(5) => add_wr_out_s_5_port, add_wr_out(4) 
                           => add_wr_out_s_4_port, add_wr_out(3) => 
                           add_wr_out_s_3_port, add_wr_out(2) => 
                           add_wr_out_s_2_port, add_wr_out(1) => 
                           add_wr_out_s_1_port, add_wr_out(0) => 
                           add_wr_out_s_0_port, add_rd1_out(6) => 
                           add_rd1_out_s_6_port, add_rd1_out(5) => 
                           add_rd1_out_s_5_port, add_rd1_out(4) => 
                           add_rd1_out_s_4_port, add_rd1_out(3) => 
                           add_rd1_out_s_3_port, add_rd1_out(2) => 
                           add_rd1_out_s_2_port, add_rd1_out(1) => 
                           add_rd1_out_s_1_port, add_rd1_out(0) => 
                           add_rd1_out_s_0_port, add_rd2_out(6) => 
                           add_rd2_out_s_6_port, add_rd2_out(5) => 
                           add_rd2_out_s_5_port, add_rd2_out(4) => 
                           add_rd2_out_s_4_port, add_rd2_out(3) => 
                           add_rd2_out_s_3_port, add_rd2_out(2) => 
                           add_rd2_out_s_2_port, add_rd2_out(1) => 
                           add_rd2_out_s_1_port, add_rd2_out(0) => 
                           add_rd2_out_s_0_port);
   physRF : physical_RF_NData32_NRegs72_NAddr7 port map( CLK => clk, RESET => 
                           reset, ENABLE => enable, RD1 => rd1, RD2 => rd2, WR 
                           => wr1, ADD_WR(6) => add_wr_out_s_6_port, ADD_WR(5) 
                           => add_wr_out_s_5_port, ADD_WR(4) => 
                           add_wr_out_s_4_port, ADD_WR(3) => 
                           add_wr_out_s_3_port, ADD_WR(2) => 
                           add_wr_out_s_2_port, ADD_WR(1) => 
                           add_wr_out_s_1_port, ADD_WR(0) => 
                           add_wr_out_s_0_port, ADD_RD1(6) => 
                           add_rd1_out_s_6_port, ADD_RD1(5) => 
                           add_rd1_out_s_5_port, ADD_RD1(4) => 
                           add_rd1_out_s_4_port, ADD_RD1(3) => 
                           add_rd1_out_s_3_port, ADD_RD1(2) => 
                           add_rd1_out_s_2_port, ADD_RD1(1) => 
                           add_rd1_out_s_1_port, ADD_RD1(0) => 
                           add_rd1_out_s_0_port, ADD_RD2(6) => 
                           add_rd2_out_s_6_port, ADD_RD2(5) => 
                           add_rd2_out_s_5_port, ADD_RD2(4) => 
                           add_rd2_out_s_4_port, ADD_RD2(3) => 
                           add_rd2_out_s_3_port, ADD_RD2(2) => 
                           add_rd2_out_s_2_port, ADD_RD2(1) => 
                           add_rd2_out_s_1_port, ADD_RD2(0) => 
                           add_rd2_out_s_0_port, DATAIN(31) => dataIn(31), 
                           DATAIN(30) => dataIn(30), DATAIN(29) => dataIn(29), 
                           DATAIN(28) => dataIn(28), DATAIN(27) => dataIn(27), 
                           DATAIN(26) => dataIn(26), DATAIN(25) => dataIn(25), 
                           DATAIN(24) => dataIn(24), DATAIN(23) => dataIn(23), 
                           DATAIN(22) => dataIn(22), DATAIN(21) => dataIn(21), 
                           DATAIN(20) => dataIn(20), DATAIN(19) => dataIn(19), 
                           DATAIN(18) => dataIn(18), DATAIN(17) => dataIn(17), 
                           DATAIN(16) => dataIn(16), DATAIN(15) => dataIn(15), 
                           DATAIN(14) => dataIn(14), DATAIN(13) => dataIn(13), 
                           DATAIN(12) => dataIn(12), DATAIN(11) => dataIn(11), 
                           DATAIN(10) => dataIn(10), DATAIN(9) => dataIn(9), 
                           DATAIN(8) => dataIn(8), DATAIN(7) => dataIn(7), 
                           DATAIN(6) => dataIn(6), DATAIN(5) => dataIn(5), 
                           DATAIN(4) => dataIn(4), DATAIN(3) => dataIn(3), 
                           DATAIN(2) => dataIn(2), DATAIN(1) => dataIn(1), 
                           DATAIN(0) => dataIn(0), OUT1(31) => dataOut1(31), 
                           OUT1(30) => dataOut1(30), OUT1(29) => dataOut1(29), 
                           OUT1(28) => dataOut1(28), OUT1(27) => dataOut1(27), 
                           OUT1(26) => dataOut1(26), OUT1(25) => dataOut1(25), 
                           OUT1(24) => dataOut1(24), OUT1(23) => dataOut1(23), 
                           OUT1(22) => dataOut1(22), OUT1(21) => dataOut1(21), 
                           OUT1(20) => dataOut1(20), OUT1(19) => dataOut1(19), 
                           OUT1(18) => dataOut1(18), OUT1(17) => dataOut1(17), 
                           OUT1(16) => dataOut1(16), OUT1(15) => dataOut1(15), 
                           OUT1(14) => dataOut1(14), OUT1(13) => dataOut1(13), 
                           OUT1(12) => dataOut1(12), OUT1(11) => dataOut1(11), 
                           OUT1(10) => dataOut1(10), OUT1(9) => dataOut1(9), 
                           OUT1(8) => dataOut1(8), OUT1(7) => dataOut1(7), 
                           OUT1(6) => dataOut1(6), OUT1(5) => dataOut1(5), 
                           OUT1(4) => dataOut1(4), OUT1(3) => dataOut1(3), 
                           OUT1(2) => dataOut1(2), OUT1(1) => dataOut1(1), 
                           OUT1(0) => dataOut1(0), OUT2(31) => dataOut2(31), 
                           OUT2(30) => dataOut2(30), OUT2(29) => dataOut2(29), 
                           OUT2(28) => dataOut2(28), OUT2(27) => dataOut2(27), 
                           OUT2(26) => dataOut2(26), OUT2(25) => dataOut2(25), 
                           OUT2(24) => dataOut2(24), OUT2(23) => dataOut2(23), 
                           OUT2(22) => dataOut2(22), OUT2(21) => dataOut2(21), 
                           OUT2(20) => dataOut2(20), OUT2(19) => dataOut2(19), 
                           OUT2(18) => dataOut2(18), OUT2(17) => dataOut2(17), 
                           OUT2(16) => dataOut2(16), OUT2(15) => dataOut2(15), 
                           OUT2(14) => dataOut2(14), OUT2(13) => dataOut2(13), 
                           OUT2(12) => dataOut2(12), OUT2(11) => dataOut2(11), 
                           OUT2(10) => dataOut2(10), OUT2(9) => dataOut2(9), 
                           OUT2(8) => dataOut2(8), OUT2(7) => dataOut2(7), 
                           OUT2(6) => dataOut2(6), OUT2(5) => dataOut2(5), 
                           OUT2(4) => dataOut2(4), OUT2(3) => dataOut2(3), 
                           OUT2(2) => dataOut2(2), OUT2(1) => dataOut2(1), 
                           OUT2(0) => dataOut2(0));

end SYN_struct;
