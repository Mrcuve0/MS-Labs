package constants is

  constant numBit : integer := 4;
  constant radixN : integer := 3;

end package constants;
