package constants is
  
  constant numBit : integer := 4;
  constant CSSG_NBIT : integer := 32;

end package constants;
