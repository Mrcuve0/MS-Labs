library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.constants.all;


entity translationUnit_RF is
  
end entity translationUnit_RF;


architecture beh of translationUnit_RF is

begin  -- architecture beh

  

end architecture beh;
