package constants is

  constant numBit : integer := 8;
  constant radixN : integer := 3;

end package constants;
