
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_register_file is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_register_file;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_register_file.all;

entity register_file is

   port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
         std_logic_vector (63 downto 0);  OUT1, OUT2 : out std_logic_vector (63
         downto 0));

end register_file;

architecture SYN_beh of register_file is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component TBUF_X1
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107,
      n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, 
      n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, 
      n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, 
      n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, 
      n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, 
      n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, 
      n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, 
      n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, 
      n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, 
      n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, 
      n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, 
      n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, 
      n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, 
      n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, 
      n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, 
      n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, 
      n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, 
      n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, 
      n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, 
      n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, 
      n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, 
      n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, 
      n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, 
      n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, 
      n4348, n4349, n4350, n4351, n4352, n4353, n5763, n5765, n5767, n5769, 
      n5771, n5773, n5775, n5777, n5779, n5781, n5783, n5785, n5787, n5789, 
      n5791, n5793, n5795, n5797, n5799, n5801, n5803, n5805, n5807, n5809, 
      n5811, n5813, n5815, n5817, n5819, n5821, n5823, n5825, n5827, n5829, 
      n5831, n5833, n5835, n5837, n5839, n5841, n5843, n5845, n5847, n5849, 
      n5851, n5853, n5855, n5857, n5859, n5861, n5863, n5865, n5867, n5869, 
      n5871, n5873, n5875, n5877, n5879, n5881, n5883, n5885, n5887, n5889, 
      n5891, n5893, n5895, n5897, n5899, n5901, n5903, n5905, n5907, n5909, 
      n5911, n5913, n5915, n5917, n5919, n5921, n5923, n5925, n5927, n5929, 
      n5931, n5933, n5935, n5937, n5939, n5941, n5943, n5945, n5947, n5949, 
      n5951, n5953, n5955, n5957, n5959, n5961, n5963, n5965, n5967, n5969, 
      n5971, n5973, n5975, n5977, n5979, n5981, n5983, n5985, n5987, n5989, 
      n5991, n5993, n5995, n5997, n5999, n6001, n6003, n6005, n6007, n6009, 
      n6011, n6013, n6015, n6017, n6018, n6019, n6020, n6021, n6022, n6023, 
      n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, 
      n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, 
      n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, 
      n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, 
      n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, 
      n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, 
      n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, 
      n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, 
      n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, 
      n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, 
      n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, 
      n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, 
      n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, 
      n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, 
      n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, 
      n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, 
      n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, 
      n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, 
      n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, 
      n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, 
      n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, 
      n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, 
      n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, 
      n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, 
      n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, 
      n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, 
      n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, 
      n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, 
      n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, 
      n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, 
      n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, 
      n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, 
      n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, 
      n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, 
      n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, 
      n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, 
      n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, 
      n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, 
      n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, 
      n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, 
      n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, 
      n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, 
      n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, 
      n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, 
      n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, 
      n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, 
      n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, 
      n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, 
      n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, 
      n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, 
      n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, 
      n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, 
      n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, 
      n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, 
      n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, 
      n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, 
      n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, 
      n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, 
      n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, 
      n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, 
      n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, 
      n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, 
      n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, 
      n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, 
      n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, 
      n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, 
      n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, 
      n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, 
      n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, 
      n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, 
      n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, 
      n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, 
      n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, 
      n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, 
      n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, 
      n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, 
      n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, 
      n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, 
      n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, 
      n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, 
      n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, 
      n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, 
      n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, 
      n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, 
      n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, 
      n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, 
      n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, 
      n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, 
      n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, 
      n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, 
      n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, 
      n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, 
      n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, 
      n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, 
      n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, 
      n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, 
      n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, 
      n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, 
      n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, 
      n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, 
      n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, 
      n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, 
      n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, 
      n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, 
      n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, 
      n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, 
      n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, 
      n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, 
      n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, 
      n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, 
      n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, 
      n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, 
      n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, 
      n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, 
      n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, 
      n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, 
      n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, 
      n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, 
      n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, 
      n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, 
      n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, 
      n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, 
      n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, 
      n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, 
      n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, 
      n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, 
      n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, 
      n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, 
      n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, 
      n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, 
      n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, 
      n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, 
      n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, 
      n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, 
      n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, 
      n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, 
      n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, 
      n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, 
      n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, 
      n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, 
      n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, 
      n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, 
      n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, 
      n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, 
      n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, 
      n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, 
      n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, 
      n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, 
      n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, 
      n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, 
      n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, 
      n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, 
      n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, 
      n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, 
      n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, 
      n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, 
      n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, 
      n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, 
      n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, 
      n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, 
      n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, 
      n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, 
      n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, 
      n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, 
      n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, 
      n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, 
      n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, 
      n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, 
      n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, 
      n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, 
      n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, 
      n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, 
      n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, 
      n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, 
      n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, 
      n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, 
      n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, 
      n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, 
      n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, 
      n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, 
      n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, 
      n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, 
      n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, 
      n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, 
      n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, 
      n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, 
      n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, 
      n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, 
      n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, 
      n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, 
      n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, 
      n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, 
      n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, 
      n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, 
      n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, 
      n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, 
      n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, 
      n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, 
      n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, 
      n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, 
      n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, 
      n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, 
      n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, 
      n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, 
      n8064, n8065, n8450, n8453, n8456, n8459, n8462, n8465, n8468, n8471, 
      n8474, n8477, n8480, n8483, n8486, n8489, n8492, n8495, n8498, n8501, 
      n8504, n8507, n8510, n8513, n8516, n8519, n8522, n8525, n8528, n8531, 
      n8534, n8537, n8540, n8543, n8546, n8549, n8552, n8555, n8558, n8561, 
      n8564, n8567, n8570, n8573, n8576, n8579, n8582, n8585, n8588, n8591, 
      n8594, n8597, n8600, n8603, n8606, n8609, n8612, n8615, n8618, n8621, 
      n8624, n8627, n8630, n8633, n8636, n8639, n9249, n9252, n9255, n9258, 
      n9261, n9264, n9267, n9270, n9273, n9276, n9279, n9282, n9285, n9288, 
      n9291, n9294, n9297, n9300, n9303, n9306, n9309, n9312, n9315, n9318, 
      n9321, n9324, n9327, n9330, n9333, n9336, n9339, n9342, n9345, n9348, 
      n9351, n9354, n9357, n9360, n9363, n9366, n9369, n9372, n9375, n9378, 
      n9381, n9384, n9387, n9390, n9393, n9396, n9399, n9402, n9405, n9408, 
      n9411, n9414, n9417, n9420, n9423, n9426, n9429, n9432, n9435, n9438, 
      n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, 
      n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, 
      n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, 
      n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, 
      n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, 
      n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, 
      n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, 
      n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, 
      n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, 
      n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, 
      n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, 
      n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, 
      n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, 
      n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, 
      n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, 
      n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, 
      n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, 
      n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, 
      n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, 
      n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, 
      n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, 
      n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, 
      n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, 
      n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, 
      n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, 
      n9755, n9756, n9757, n9758, n9759, n9760, n18303, n18304, n18305, n18306,
      n18307, n18308, n18309, n18310, n18311, n18312, n18313, n18314, n18315, 
      n18316, n18317, n18318, n18319, n18320, n18321, n18322, n18323, n18324, 
      n18325, n18326, n18327, n18328, n18329, n18330, n18331, n18332, n18333, 
      n18334, n18335, n18336, n18337, n18338, n18339, n18340, n18341, n18342, 
      n18343, n18344, n18345, n18346, n18347, n18348, n18349, n18350, n18351, 
      n18352, n18353, n18354, n18355, n18356, n18357, n18358, n18359, n18360, 
      n18361, n18362, n18363, n18364, n18365, n18366, n18367, n18382, n18383, 
      n18384, n18399, n18400, n18401, n18416, n18417, n18418, n18433, n18434, 
      n18435, n18450, n18451, n18452, n18467, n18468, n18469, n18484, n18485, 
      n18486, n18501, n18502, n18503, n18518, n18519, n18520, n18535, n18536, 
      n18537, n18552, n18553, n18554, n18569, n18570, n18571, n18586, n18587, 
      n18588, n18603, n18604, n18605, n18620, n18621, n18622, n18637, n18638, 
      n18639, n18654, n18655, n18656, n18671, n18672, n18673, n18688, n18689, 
      n18690, n18705, n18706, n18707, n18722, n18723, n18724, n18739, n18740, 
      n18741, n18756, n18757, n18758, n18773, n18774, n18775, n18790, n18791, 
      n18792, n18807, n18808, n18809, n18824, n18825, n18826, n18841, n18842, 
      n18843, n18858, n18859, n18860, n18875, n18876, n18877, n18892, n18893, 
      n18894, n18909, n18910, n18911, n18926, n18927, n18928, n18943, n18944, 
      n18945, n18960, n18961, n18962, n18977, n18978, n18979, n18994, n18995, 
      n18996, n19011, n19012, n19013, n19028, n19029, n19030, n19045, n19046, 
      n19047, n19062, n19063, n19064, n19079, n19080, n19081, n19096, n19097, 
      n19098, n19113, n19114, n19115, n19130, n19131, n19132, n19147, n19148, 
      n19149, n19164, n19165, n19166, n19181, n19182, n19183, n19198, n19199, 
      n19200, n19215, n19216, n19217, n19232, n19233, n19234, n19249, n19250, 
      n19251, n19266, n19267, n19268, n19283, n19284, n19285, n19300, n19301, 
      n19302, n19317, n19318, n19319, n19334, n19335, n19336, n19351, n19352, 
      n19353, n19368, n19369, n19370, n19385, n19386, n19387, n19402, n19403, 
      n19404, n19419, n19420, n19421, n19436, n19437, n19438, n19453, n19454, 
      n19455, n19456, n19457, n19458, n19459, n19460, n19461, n19462, n19463, 
      n19464, n19465, n19466, n19467, n19468, n19469, n19470, n19471, n19472, 
      n19473, n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481, 
      n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489, n19490, 
      n19491, n19492, n19493, n19494, n19495, n19496, n19497, n19498, n19499, 
      n19500, n19501, n19502, n19503, n19504, n19505, n19506, n19507, n19508, 
      n19509, n19510, n19511, n19512, n19513, n19514, n19515, n19516, n19517, 
      n19518, n19519, n19520, n19521, n19522, n19523, n19524, n19525, n19526, 
      n19527, n19528, n19529, n19530, n19531, n19532, n19533, n19534, n19535, 
      n19536, n19537, n19538, n19539, n19540, n19541, n19542, n19543, n19544, 
      n19545, n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553, 
      n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561, n19562, 
      n19563, n19564, n19565, n19566, n19567, n19568, n19569, n19570, n19571, 
      n19572, n19573, n19574, n19575, n19576, n19577, n19578, n19579, n19580, 
      n19581, n19582, n20626, n20630, n20631, n20632, n20633, n20634, n20635, 
      n20636, n20637, n20638, n20639, n20640, n20641, n20642, n20643, n20644, 
      n20645, n20646, n20647, n20648, n20649, n20650, n20651, n20652, n20653, 
      n20654, n20655, n20656, n20657, n20658, n20659, n20660, n20661, n20662, 
      n20663, n20664, n20665, n20666, n20667, n20668, n20669, n20670, n20671, 
      n20672, n20673, n20674, n20675, n20676, n20677, n20678, n20679, n20680, 
      n20681, n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689, 
      n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697, n20698, 
      n20699, n20700, n20701, n20702, n20703, n20704, n20705, n20706, n20707, 
      n20708, n20709, n20710, n20711, n20712, n20713, n20714, n20715, n20716, 
      n20717, n20718, n20719, n20720, n20721, n20722, n20723, n20724, n20725, 
      n20726, n20727, n20728, n20729, n20730, n20731, n20732, n20733, n20734, 
      n20735, n20736, n20737, n20738, n20739, n20740, n20741, n20742, n20743, 
      n20744, n20745, n20746, n20747, n20748, n20749, n20750, n20751, n20752, 
      n20753, n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761, 
      n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769, n20770, 
      n20771, n20772, n20773, n20774, n20775, n20776, n20777, n20778, n20779, 
      n20780, n20781, n20782, n20783, n20784, n20785, n20786, n20787, n20788, 
      n20789, n20790, n20791, n20792, n20793, n20794, n20795, n20796, n20797, 
      n20798, n20799, n20800, n20801, n20802, n20803, n20804, n20805, n20806, 
      n20807, n20808, n20809, n20810, n20811, n20812, n20813, n20814, n20815, 
      n20816, n20817, n20818, n20819, n20820, n20821, n20822, n20823, n20824, 
      n20825, n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833, 
      n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841, n20842, 
      n20843, n20844, n20845, n20846, n20847, n20848, n20849, n20850, n20851, 
      n20852, n20853, n20854, n20855, n20856, n20857, n20858, n20859, n20860, 
      n20861, n20862, n20863, n20864, n20865, n20866, n20867, n20868, n20869, 
      n20870, n20871, n20872, n20873, n20874, n20875, n20876, n20877, n20878, 
      n20879, n20880, n20881, n20882, n20883, n20884, n20885, n20886, n20887, 
      n20888, n20889, n20890, n20891, n20892, n20893, n20894, n20895, n20896, 
      n20897, n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905, 
      n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913, n20914, 
      n20915, n20916, n20917, n20918, n20919, n20920, n20921, n20922, n20923, 
      n20924, n20925, n20926, n20927, n20928, n20929, n20930, n20931, n20932, 
      n20933, n20934, n20935, n20936, n20937, n20938, n20939, n20940, n20941, 
      n20942, n20943, n20944, n20945, n20946, n20947, n20948, n20949, n20950, 
      n20951, n20952, n20953, n20954, n20955, n20956, n20957, n20958, n20959, 
      n20960, n20961, n20962, n20963, n20964, n20965, n20966, n20967, n20968, 
      n20969, n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977, 
      n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985, n20986, 
      n20987, n20988, n20989, n20990, n20991, n20992, n20993, n20994, n20995, 
      n20996, n20997, n20998, n20999, n21000, n21001, n21002, n21003, n21004, 
      n21005, n21006, n21007, n21008, n21009, n21010, n21011, n21012, n21013, 
      n21014, n21015, n21016, n21017, n21018, n21019, n21020, n21021, n21022, 
      n21023, n21024, n21025, n21026, n21027, n21028, n21029, n21030, n21031, 
      n21032, n21033, n21034, n21035, n21036, n21037, n21038, n21039, n21040, 
      n21041, n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049, 
      n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057, n21058, 
      n21059, n21060, n21061, n21062, n21063, n21064, n21065, n21066, n21067, 
      n21068, n21069, n21070, n21071, n21072, n21073, n21074, n21075, n21076, 
      n21077, n21078, n21079, n21080, n21081, n21082, n21083, n21084, n21085, 
      n21086, n21087, n21088, n21089, n21090, n21091, n21092, n21093, n21094, 
      n21095, n21096, n21097, n21098, n21099, n21100, n21101, n21102, n21103, 
      n21104, n21105, n21106, n21107, n21108, n21109, n21110, n21111, n21112, 
      n21113, n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121, 
      n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129, n21130, 
      n21131, n21132, n21133, n21134, n21135, n21136, n21137, n21138, n21139, 
      n21140, n21141, n21142, n21143, n21144, n21145, n21146, n21147, n21148, 
      n21149, n21150, n21151, n21152, n21153, n21154, n21155, n21156, n21157, 
      n21158, n21159, n21160, n21161, n21162, n21163, n21164, n21165, n21166, 
      n21167, n21168, n21169, n21170, n21171, n21172, n21173, n21174, n21175, 
      n21176, n21177, n21178, n21179, n21180, n21181, n21182, n21183, n21184, 
      n21185, n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193, 
      n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201, n21202, 
      n21203, n21204, n21205, n21206, n21207, n21208, n21209, n21210, n21211, 
      n21212, n21213, n21214, n21215, n21216, n21217, n21218, n21219, n21220, 
      n21221, n21222, n21223, n21224, n21225, n21226, n21227, n21228, n21229, 
      n21230, n21231, n21232, n21233, n21234, n21235, n21236, n21237, n21238, 
      n21239, n21240, n21241, n21242, n21243, n21244, n21245, n21246, n21247, 
      n21248, n21249, n21250, n21251, n21252, n21253, n21254, n21255, n21256, 
      n21257, n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265, 
      n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273, n21274, 
      n21275, n21276, n21277, n21278, n21279, n21280, n21281, n21282, n21283, 
      n21284, n21285, n21286, n21287, n21288, n21289, n21290, n21291, n21292, 
      n21293, n21294, n21295, n21296, n21297, n21298, n21299, n21300, n21301, 
      n21302, n21303, n21304, n21305, n21306, n21307, n21308, n21309, n21310, 
      n21311, n21312, n21313, n21314, n21315, n21316, n21317, n21318, n21319, 
      n21320, n21321, n21322, n21323, n21324, n21325, n21326, n21327, n21328, 
      n21329, n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337, 
      n21338, n21339, n21340, n21341, n21342, n21343, n21344, n21345, n21346, 
      n21347, n21348, n21349, n21350, n21351, n21352, n21353, n21354, n21355, 
      n21356, n21357, n21358, n21359, n21360, n21361, n21362, n21363, n21364, 
      n21365, n21366, n21367, n21368, n21369, n21370, n21371, n21372, n21373, 
      n21374, n21375, n21376, n21377, n21378, n21379, n21380, n21381, n21382, 
      n21383, n21384, n21385, n21386, n21387, n21388, n21389, n21390, n21391, 
      n21392, n21393, n21394, n21395, n21396, n21397, n21398, n21399, n21400, 
      n21401, n21402, n21403, n21404, n21405, n21406, n21407, n21408, n21409, 
      n21410, n21411, n21412, n21413, n21414, n21415, n21416, n21417, n21418, 
      n21419, n21420, n21421, n21422, n21423, n21424, n21425, n21426, n21427, 
      n21428, n21429, n21430, n21431, n21432, n21433, n21434, n21435, n21436, 
      n21437, n21438, n21439, n21440, n21441, n21442, n21443, n21444, n21445, 
      n21446, n21447, n21448, n21449, n21450, n21451, n21452, n21453, n21454, 
      n21455, n21456, n21457, n21458, n21459, n21460, n21461, n21462, n21463, 
      n21464, n21465, n21466, n21467, n21468, n21469, n21470, n21471, n21472, 
      n21473, n21474, n21475, n21476, n21477, n21478, n21479, n21480, n21481, 
      n21482, n21483, n21484, n21485, n21486, n21487, n21488, n21489, n21490, 
      n21491, n21492, n21493, n21494, n21495, n21496, n21497, n21498, n21499, 
      n21500, n21501, n21502, n21503, n21504, n21505, n21506, n21507, n21508, 
      n21509, n21510, n21511, n21512, n21513, n21514, n21515, n21516, n21517, 
      n21518, n21519, n21520, n21521, n21522, n21523, n21524, n21525, n21526, 
      n21527, n21528, n21529, n21530, n21531, n21532, n21533, n21534, n21535, 
      n21536, n21537, n21538, n21539, n21540, n21541, n21542, n21543, n21544, 
      n21545, n21546, n21547, n21548, n21549, n21550, n21551, n21552, n21553, 
      n21554, n21555, n21556, n21557, n21558, n21559, n21560, n21561, n21562, 
      n21563, n21564, n21565, n21566, n21567, n21568, n21569, n21570, n21571, 
      n21572, n21573, n21574, n21575, n21576, n21577, n21578, n21579, n21580, 
      n21581, n21582, n21583, n21584, n21585, n21586, n21587, n21588, n21589, 
      n21590, n21591, n21592, n21593, n21594, n21595, n21596, n21597, n21598, 
      n21599, n21600, n21601, n21602, n21603, n21604, n21605, n21606, n21607, 
      n21608, n21609, n21610, n21611, n21612, n21613, n21614, n21615, n21616, 
      n21617, n21618, n21619, n21620, n21621, n21622, n21623, n21624, n21625, 
      n21626, n21627, n21628, n21629, n21630, n21631, n21632, n21633, n21634, 
      n21635, n21636, n21637, n21638, n21639, n21640, n21641, n21642, n21643, 
      n21644, n21645, n21646, n21647, n21648, n21649, n21650, n21651, n21652, 
      n21653, n21654, n21655, n21656, n21657, n21658, n21659, n21660, n21661, 
      n21662, n21663, n21664, n21665, n21666, n21667, n21668, n21669, n21670, 
      n21671, n21672, n21673, n21674, n21675, n21676, n21677, n21678, n21679, 
      n21680, n21681, n21682, n21683, n21684, n21685, n21686, n21687, n21688, 
      n21689, n21690, n21691, n21692, n21693, n21694, n21695, n21696, n21697, 
      n21698, n21699, n21700, n21701, n21702, n21703, n21704, n21705, n21706, 
      n21707, n21708, n21709, n21710, n21711, n21712, n21713, n21714, n21715, 
      n21716, n21717, n21718, n21719, n21720, n21721, n21722, n21723, n21724, 
      n21725, n21726, n21727, n21728, n21729, n21730, n21731, n21732, n21733, 
      n21734, n21735, n21736, n21737, n21738, n21739, n21740, n21741, n21742, 
      n21743, n21744, n21745, n21746, n21747, n21748, n21749, n21750, n21751, 
      n21752, n21753, n21754, n21755, n21756, n21757, n21758, n21759, n21760, 
      n21761, n21762, n21763, n21764, n21765, n21766, n21767, n21768, n21769, 
      n21770, n21771, n21772, n21773, n21774, n21775, n21776, n21777, n21778, 
      n21779, n21780, n21781, n21782, n21783, n21784, n21785, n21786, n21787, 
      n21788, n21789, n21790, n21791, n21792, n21793, n21794, n21795, n21796, 
      n21797, n21798, n21799, n21800, n21801, n21802, n21803, n21804, n21805, 
      n21806, n21807, n21808, n21809, n21810, n21811, n21812, n21813, n21814, 
      n21815, n21816, n21817, n21818, n21819, n21820, n21821, n21822, n21823, 
      n21824, n21825, n21826, n21827, n21828, n21829, n21830, n21831, n21832, 
      n21833, n21834, n21835, n21836, n21837, n21838, n21839, n21840, n21841, 
      n21842, n21843, n21844, n21845, n21846, n21847, n21848, n21849, n21850, 
      n21851, n21852, n21853, n21854, n21855, n21856, n21857, n21858, n21859, 
      n21860, n21861, n21862, n21863, n21864, n21865, n21866, n21867, n21868, 
      n21869, n21870, n21871, n21872, n21873, n21874, n21875, n21876, n21877, 
      n21878, n21879, n21880, n21881, n21882, n21883, n21884, n21885, n21886, 
      n21887, n21888, n21889, n21890, n21891, n21892, n21893, n21894, n21895, 
      n21896, n21897, n21898, n21899, n21900, n21901, n21902, n21903, n21904, 
      n21905, n21906, n21907, n21908, n21909, n21910, n21911, n21912, n21913, 
      n21914, n21915, n21916, n21917, n21918, n21919, n21920, n21921, n21922, 
      n21923, n21924, n21925, n21926, n21927, n21928, n21929, n21930, n21931, 
      n21932, n21933, n21934, n21935, n21936, n21937, n21938, n21939, n21940, 
      n21941, n21942, n21943, n21944, n21945, n21946, n21947, n21948, n21949, 
      n21950, n21951, n21952, n21953, n21954, n21955, n21956, n21957, n21958, 
      n21959, n21960, n21961, n21962, n21963, n21964, n21965, n21966, n21967, 
      n21968, n21969, n21970, n21971, n21972, n21973, n21974, n21975, n21976, 
      n21977, n21978, n21979, n21980, n21981, n21982, n21983, n21984, n21985, 
      n21986, n21987, n21988, n21989, n21990, n21991, n21992, n21993, n21994, 
      n21995, n21996, n21997, n21998, n21999, n22000, n22001, n22002, n22003, 
      n22004, n22005, n22006, n22007, n22008, n22009, n22010, n22011, n22012, 
      n22013, n22014, n22015, n22016, n22017, n22018, n22019, n22020, n22021, 
      n22022, n22023, n22024, n22025, n22026, n22027, n22028, n22029, n22030, 
      n22031, n22032, n22033, n22034, n22035, n22036, n22037, n22038, n22039, 
      n22040, n22041, n22042, n22043, n22044, n22045, n22046, n22047, n22048, 
      n22049, n22050, n22051, n22052, n22053, n22054, n22055, n22056, n22057, 
      n22058, n22059, n22060, n22061, n22062, n22063, n22064, n22065, n22066, 
      n22067, n22068, n22069, n22070, n22071, n22072, n22073, n22074, n22075, 
      n22076, n22077, n22078, n22079, n22080, n22081, n22082, n22083, n22084, 
      n22085, n22086, n22087, n22088, n22089, n22090, n22091, n22092, n22093, 
      n22094, n22095, n22096, n22097, n22098, n22099, n22100, n22101, n22102, 
      n22103, n22104, n22105, n22106, n22107, n22108, n22109, n22110, n22111, 
      n22112, n22113, n22114, n22115, n22116, n22117, n22118, n22119, n22120, 
      n22121, n22122, n22123, n22124, n22125, n22126, n22127, n22128, n22129, 
      n22130, n22131, n22132, n22133, n22134, n22135, n22136, n22137, n22138, 
      n22139, n22140, n22141, n22142, n22143, n22144, n22145, n22146, n22147, 
      n22148, n22149, n22150, n22151, n22152, n22153, n22154, n22155, n22156, 
      n22157, n22158, n22159, n22160, n22161, n22162, n22163, n22164, n22165, 
      n22166, n22167, n22168, n22169, n22170, n22171, n22172, n22173, n22174, 
      n22175, n22176, n22177, n22178, n22179, n22180, n22181, n22182, n22183, 
      n22184, n22185, n22186, n22187, n22188, n22189, n22190, n22191, n22192, 
      n22193, n22194, n22195, n22196, n22197, n22198, n22199, n22200, n22201, 
      n22202, n22203, n22204, n22205, n22206, n22207, n22208, n22209, n22210, 
      n22211, n22212, n22213, n22214, n22215, n22216, n22217, n22218, n22219, 
      n22220, n22221, n22222, n22223, n22224, n22225, n22226, n22227, n22228, 
      n22229, n22230, n22231, n22232, n22233, n22234, n22235, n22236, n22237, 
      n22238, n22239, n22240, n22241, n22242, n22243, n22244, n22245, n22246, 
      n22247, n22248, n22249, n22250, n22251, n22252, n22253, n22254, n22255, 
      n22256, n22257, n22258, n22259, n22260, n22261, n22262, n22263, n22264, 
      n22265, n22266, n22267, n22268, n22269, n22270, n22271, n22272, n22273, 
      n22274, n22275, n22276, n22277, n22278, n22279, n22280, n22281, n22282, 
      n22283, n22284, n22285, n22286, n22287, n22288, n22289, n22290, n22291, 
      n22292, n22293, n22294, n22295, n22296, n22297, n22298, n22299, n22300, 
      n22301, n22302, n22303, n22304, n22305, n22306, n22307, n22308, n22309, 
      n22310, n22311, n22312, n22313, n22314, n22315, n22316, n22317, n22318, 
      n22319, n22320, n22321, n22322, n22323, n22324, n22325, n22326, n22327, 
      n22328, n22329, n22330, n22331, n22332, n22333, n22334, n22335, n22336, 
      n22337, n22338, n22339, n22340, n22341, n22342, n22343, n22344, n22345, 
      n22346, n22347, n22348, n22349, n22350, n22351, n22352, n22353, n22354, 
      n22355, n22356, n22357, n22358, n22359, n22360, n22361, n22362, n22363, 
      n22364, n22365, n22366, n22367, n22368, n22369, n22370, n22371, n22372, 
      n22373, n22374, n22375, n22376, n22377, n22378, n22379, n22380, n22381, 
      n22382, n22383, n22384, n22385, n22386, n22387, n22388, n22389, n22390, 
      n22391, n22392, n22393, n22394, n22395, n22396, n22397, n22398, n22399, 
      n22400, n22401, n22402, n22403, n22404, n22405, n22406, n22407, n22408, 
      n22409, n22410, n22411, n22412, n22413, n22414, n22415, n22416, n22417, 
      n22418, n22419, n22420, n22421, n22422, n22423, n22424, n22425, n22426, 
      n22427, n22428, n22429, n22430, n22431, n22432, n22433, n22434, n22435, 
      n22436, n22437, n22438, n22439, n22440, n22441, n22442, n22443, n22444, 
      n22445, n22446, n22447, n22448, n22449, n22450, n22451, n22452, n22453, 
      n22454, n22455, n22456, n22457, n22458, n22459, n22460, n22461, n22462, 
      n22463, n22464, n22465, n22466, n22467, n22468, n22469, n22470, n22471, 
      n22472, n22473, n22474, n22475, n22476, n22477, n22478, n22479, n22480, 
      n22481, n22482, n22483, n22484, n22485, n22486, n22487, n22488, n22489, 
      n22490, n22491, n22492, n22493, n22494, n22495, n22496, n22497, n22498, 
      n22499, n22500, n22501, n22502, n22503, n22504, n22505, n22506, n22507, 
      n22508, n22509, n22510, n22511, n22512, n22513, n22514, n22515, n22516, 
      n22517, n22518, n22519, n22520, n22521, n22522, n22523, n22524, n22525, 
      n22526, n22527, n22528, n22529, n22530, n22531, n22532, n22533, n22534, 
      n22535, n22536, n22537, n22538, n22539, n22540, n22541, n22542, n22543, 
      n22544, n22545, n22546, n22547, n22548, n22549, n22550, n22551, n22552, 
      n22553, n22554, n22555, n22556, n22557, n22558, n22559, n22560, n22561, 
      n22562, n22563, n22564, n22565, n22566, n22567, n22568, n22569, n22570, 
      n22571, n22572, n22573, n22574, n22575, n22576, n22577, n22578, n22579, 
      n22580, n22581, n22582, n22583, n22584, n22585, n22586, n22587, n22588, 
      n22589, n22590, n22591, n22592, n22593, n22594, n22595, n22596, n22597, 
      n22598, n22599, n22600, n22601, n22602, n22603, n22604, n22605, n22606, 
      n22607, n22608, n22609, n22610, n22611, n22612, n22613, n22614, n22615, 
      n22616, n22617, n22618, n22619, n22620, n22621, n22622, n22623, n22624, 
      n22625, n22626, n22627, n22628, n22629, n22630, n22631, n22632, n22633, 
      n22634, n22635, n22636, n22637, n22638, n22639, n22640, n22641, n22642, 
      n22643, n22644, n22645, n22646, n22647, n22648, n22649, n22650, n22651, 
      n22652, n22653, n22654, n22655, n22656, n22657, n22658, n22659, n22660, 
      n22661, n22662, n22663, n22664, n22665, n22666, n22667, n22668, n22669, 
      n22670, n22671, n22672, n22673, n22674, n22675, n22676, n22677, n22678, 
      n22679, n22680, n22681, n22682, n22683, n22684, n22685, n22686, n22687, 
      n22688, n22689, n22690, n22691, n22692, n22693, n22694, n22695, n22696, 
      n22697, n22698, n22699, n22700, n22701, n22702, n22703, n22704, n22705, 
      n22706, n22707, n22708, n22709, n22710, n22711, n22712, n22713, n22714, 
      n22715, n22716, n22717, n22718, n22719, n22720, n22721, n22722, n22723, 
      n22724, n22725, n22726, n22727, n22728, n22729, n22730, n22731, n22732, 
      n22733, n22734, n22735, n22736, n22737, n22738, n22739, n22740, n22741, 
      n22742, n22743, n22744, n22745, n22746, n22747, n22748, n22749, n22750, 
      n22751, n22752, n22753, n22754, n22755, n22756, n22757, n22758, n22759, 
      n22760, n22761, n22762, n22763, n22764, n22765, n22766, n22767, n22768, 
      n22769, n22770, n22771, n22772, n22773, n22774, n22775, n22776, n22777, 
      n22778, n22779, n22780, n22781, n22782, n22783, n22784, n22785, n22786, 
      n22787, n22788, n22789, n22790, n22791, n22792, n22793, n22794, n22795, 
      n22796, n22797, n22798, n22799, n22800, n22801, n22802, n22803, n22804, 
      n22805, n22806, n22807, n22808, n22809, n22810, n22811, n22812, n22813, 
      n22814, n22815, n22816, n22817, n22818, n22819, n22820, n22821, n22822, 
      n22823, n22824, n22825, n22826, n22827, n22828, n22829, n22830, n22831, 
      n22832, n22833, n22834, n22835, n22836, n22837, n22838, n22839, n22840, 
      n22841, n22842, n22843, n22844, n22845, n22846, n22847, n22848, n22849, 
      n22850, n22851, n22852, n22853, n22854, n22855, n22856, n22857, n22858, 
      n22859, n22860, n22861, n22862, n22863, n22864, n22865, n22866, n22867, 
      n22868, n22869, n22870, n22871, n22872, n22873, n22874, n22875, n22876, 
      n22877, n22878, n22879, n22880, n22881, n22882, n22883, n22884, n22885, 
      n22886, n22887, n22888, n22889, n22890, n22891, n22892, n22893, n22894, 
      n22895, n22896, n22897, n22898, n22899, n22900, n22901, n22902, n22903, 
      n22904, n22905, n22906, n22907, n22908, n22909, n22910, n22911, n22912, 
      n22913, n22914, n22915, n22916, n22917, n22918, n22919, n22920, n22921, 
      n22922, n22923, n22924, n22925, n22926, n22927, n22928, n22929, n22930, 
      n22931, n22932, n22933, n22934, n22935, n22936, n22937, n22938, n22939, 
      n22940, n22941, n22942, n22943, n22944, n22945, n22946, n22947, n22948, 
      n22949, n22950, n22951, n22952, n22953, n22954, n22955, n22956, n22957, 
      n22958, n22959, n22960, n22961, n22962, n22963, n22964, n22965, n22966, 
      n22967, n22968, n22969, n22970, n22971, n22972, n22973, n22974, n22975, 
      n22976, n22977, n22978, n22979, n22980, n22981, n22982, n22983, n22984, 
      n22985, n22986, n22987, n22988, n22989, n22990, n22991, n22992, n22993, 
      n22994, n22995, n22996, n22997, n22998, n22999, n23000, n23001, n23002, 
      n23003, n23004, n23005, n23006, n23007, n23008, n23009, n23010, n23011, 
      n23012, n23013, n23014, n23015, n23016, n23017, n23018, n23019, n23020, 
      n23021, n23022, n23023, n23024, n23025, n23026, n23027, n23028, n23029, 
      n23030, n23031, n23032, n23033, n23034, n23035, n23036, n23037, n23038, 
      n23039, n23040, n23041, n23042, n23043, n23044, n23045, n23046, n23047, 
      n23048, n23049, n23050, n23051, n23052, n23053, n23054, n23055, n23056, 
      n23057, n23058, n23059, n23060, n23061, n23062, n23063, n23064, n23065, 
      n23066, n23067, n23068, n23069, n23070, n23071, n23072, n23073, n23074, 
      n23075, n23076, n23077, n23078, n23079, n23080, n23081, n23082, n23083, 
      n23084, n23085, n23086, n23087, n23088, n23089, n23090, n23091, n23092, 
      n23093, n23094, n23095, n23096, n23097, n23098, n23099, n23100, n23101, 
      n23102, n23103, n23104, n23105, n23106, n23107, n23108, n23109, n23110, 
      n23111, n23112, n23113, n23114, n23115, n23116, n23117, n23118, n23119, 
      n23120, n23121, n23122, n23123, n23124, n23125, n23126, n23127, n23128, 
      n23129, n23130, n23131, n23132, n23133, n23134, n23135, n23136, n23137, 
      n23138, n23139, n23140, n23141, n23142, n23143, n23144, n23145, n23146, 
      n23147, n23148, n23149, n23150, n23151, n23152, n23153, n23154, n23155, 
      n23156, n23157, n23158, n23159, n23160, n23161, n23162, n23163, n23164, 
      n23165, n23166, n23167, n23168, n23169, n23170, n23171, n23172, n23173, 
      n23174, n23175, n23176, n23177, n23178, n23179, n23180, n23181, n23182, 
      n23183, n23184, n23185, n23186, n23187, n23188, n23189, n23190, n23191, 
      n23192, n23193, n23194, n23195, n23196, n23197, n23198, n23199, n23200, 
      n23201, n23202, n23203, n23204, n23205, n23206, n23207, n23208, n23209, 
      n23210, n23211, n23212, n23213, n23214, n23215, n23216, n23217, n23218, 
      n23219, n23220, n23221, n23222, n23223, n23224, n23225, n23226, n23227, 
      n23228, n23229, n23230, n23231, n23232, n23233, n23234, n23235, n23236, 
      n23237, n23238, n23239, n23240, n23241, n23242, n23243, n23244, n23245, 
      n23246, n23247, n23248, n23249, n23250, n23251, n23252, n23253, n23254, 
      n23255, n23256, n23257, n23258, n23259, n23260, n23261, n23262, n23263, 
      n23264, n23265, n23266, n23267, n23268, n23269, n23270, n23271, n23272, 
      n23273, n23274, n23275, n23276, n23277, n23278, n23279, n23280, n23281, 
      n23282, n23283, n23284, n23285, n23286, n23287, n23288, n23289, n23290, 
      n23291, n23292, n23293, n23294, n23295, n23296, n23297, n23298, n23299, 
      n23300, n23301, n23302, n23303, n23304, n23305, n23306, n23307, n23308, 
      n23309, n23310, n23311, n23312, n23313, n23314, n23315, n23316, n23317, 
      n23318, n23319, n23320, n23321, n23322, n23323, n23324, n23325, n23326, 
      n23327, n23328, n23329, n23330, n23331, n23332, n23333, n23334, n23335, 
      n23336, n23337, n23338, n23339, n23340, n23341, n23342, n23343, n23344, 
      n23345, n23346, n23347, n23348, n23349, n23350, n23351, n23352, n23353, 
      n23354, n23355, n23356, n23357, n23358, n23359, n23360, n23361, n23362, 
      n23363, n23364, n23365, n23366, n23367, n23368, n23369, n23370, n23371, 
      n23372, n23373, n23374, n23375, n23376, n23377, n23378, n23379, n23380, 
      n23381, n23382, n23383, n23384, n23385, n23386, n23387, n23388, n23389, 
      n23390, n23391, n23392, n23393, n23394, n23395, n23396, n23397, n23398, 
      n23399, n23400, n23401, n23402, n23403, n23404, n23405, n23406, n23407, 
      n23408, n23409, n23410, n23411, n23412, n23413, n23414, n23415, n23416, 
      n23417, n23418, n23419, n23420, n23421, n23422, n23423, n23424, n23425, 
      n23426, n23427, n23428, n23429, n23430, n23431, n23432, n23433, n23434, 
      n23435, n23436, n23437, n23438, n23439, n23440, n23441, n23442, n23443, 
      n23444, n23445, n23446, n23447, n23448, n23449, n23450, n23451, n23452, 
      n23453, n23454, n23455, n23456, n23457, n23458, n23459, n23460, n23461, 
      n23462, n23463, n23464, n23465, n23466, n23467, n23468, n23469, n23470, 
      n23471, n23472, n23473, n23474, n23475, n23476, n23477, n23478, n23479, 
      n23480, n23481, n23482, n23483, n23484, n23485, n23486, n23487, n23488, 
      n23489, n23490, n23491, n23492, n23493, n23494, n23495, n23496, n23497, 
      n23498, n23499, n23500, n23501, n23502, n23503, n23504, n23505, n23506, 
      n23507, n23508, n23509, n23510, n23511, n23512, n23513, n23514, n23515, 
      n23516, n23517, n23518, n23519, n23520, n23521, n23522, n23523, n23524, 
      n23525, n23526, n23527, n23528, n23529, n23530, n23531, n23532, n23533, 
      n23534, n23535, n23536, n23537, n23538, n23539, n23540, n23541, n23542, 
      n23543, n23544, n23545, n23546, n23547, n23548, n23549, n23550, n23551, 
      n23552, n23553, n23554, n23555, n23556, n23557, n23558, n23559, n23560, 
      n23561, n23562, n23563, n23564, n23565, n23566, n23567, n23568, n23569, 
      n23570, n23571, n23572, n23573, n23574, n23575, n23576, n23577, n23578, 
      n23579, n23580, n23581, n23582, n23583, n23584, n23585, n23586, n23587, 
      n23588, n23589, n23590, n23591, n23592, n23593, n23594, n23595, n23596, 
      n23597, n23598, n23599, n23600, n23601, n23602, n23603, n23604, n23605, 
      n23606, n23607, n23608, n23609, n23610, n23611, n23612, n23613, n23614, 
      n23615, n23616, n23617, n23618, n23619, n23620, n23621, n23622, n23623, 
      n23624, n23625, n23626, n23627, n23628, n23629, n23630, n23631, n23632, 
      n23633, n23634, n23635, n23636, n23637, n23638, n23639, n23640, n23641, 
      n23642, n23643, n23644, n23645, n23646, n23647, n23648, n23649, n23650, 
      n23651, n23652, n23653, n23654, n23655, n23656, n23657, n23658, n23659, 
      n23660, n23661, n23662, n23663, n23664, n23665, n23666, n23667, n23668, 
      n23669, n23670, n23671, n23672, n23673, n23674, n23675, n23676, n23677, 
      n23678, n23679, n23680, n23681, n23682, n23683, n23684, n23685, n23686, 
      n23687, n23688, n23689, n23690, n23691, n23692, n23693, n23694, n23695, 
      n23696, n23697, n23698, n23699, n23700, n23701, n23702, n23703, n23704, 
      n23705, n23706, n23707, n23708, n23709, n23710, n23711, n23712, n23713, 
      n23714, n23715, n23716, n23717, n23718, n23719, n23720, n23721, n23722, 
      n23723, n23724, n23725, n23726, n23727, n23728, n23729, n23730, n23731, 
      n23732, n23733, n23734, n23735, n23736, n23737, n23738, n23739, n23740, 
      n23741, n23742, n23743, n23744, n23745, n23746, n23747, n23748, n23749, 
      n23750, n23751, n23752, n23753, n23754, n23755, n23756, n23757, n23758, 
      n23759, n23760, n23761, n23762, n23763, n23764, n23765, n23766, n23767, 
      n23768, n23769, n23770, n23771, n23772, n23773, n23774, n23775, n23776, 
      n23777, n23778, n23779, n23780, n23781, n23782, n23783, n23784, n23785, 
      n23786, n23787, n23788, n23789, n23790, n23791, n23792, n23793, n23794, 
      n23795, n23796, n23797, n23798, n23799, n23800, n23801, n23802, n23803, 
      n23804, n23805, n23806, n23807, n23808, n23809, n23810, n23811, n23812, 
      n23813, n23814, n23815, n23816, n23817, n23818, n23819, n23820, n23821, 
      n23822, n23823, n23824, n23825, n23826, n23827, n23828, n23829, n23830, 
      n23831, n23832, n23833, n23834, n23835, n23836, n23837, n23838, n23839, 
      n23840, n23841, n23842, n23843, n23844, n23845, n23846, n23847, n23848, 
      n23849, n23850, n23851, n23852, n23853, n23854, n23855, n23856, n23857, 
      n23858, n23859, n23860, n23861, n23862, n23863, n23864, n23865, n23866, 
      n23867, n23868, n23869, n23870, n23871, n23872, n23873, n23874, n23875, 
      n23876, n23877, n23878, n23879, n23880, n23881, n23882, n23883, n23884, 
      n23885, n23886, n23887, n23888, n23889, n23890, n23891, n23892, n23893, 
      n23894, n23895, n23896, n23897, n23898, n23899, n23900, n23901, n23902, 
      n23903, n23904, n23905, n23906, n23907, n23908, n23909, n23910, n23911, 
      n23912, n23913, n23914, n23915, n23916, n23917, n23918, n23919, n23920, 
      n23921, n23922, n23923, n23924, n23925, n23926, n23927, n23928, n23929, 
      n23930, n23931, n23932, n23933, n23934, n23935, n23936, n23937, n23938, 
      n23939, n23940, n23941, n23942, n23943, n23944, n23945, n23946, n23947, 
      n23948, n23949, n23950, n23951, n23952, n23953, n23954, n23955, n23956, 
      n23957, n23958, n23959, n23960, n23961, n23962, n23963, n23964, n23965, 
      n23966, n23967, n23968, n23969, n23970, n23971, n23972, n23973, n23974, 
      n23975, n23976, n23977, n23978, n23979, n23980, n23981, n23982, n23983, 
      n23984, n23985, n23986, n23987, n23988, n23989, n23990, n23991, n23992, 
      n23993, n23994, n23995, n23996, n23997, n23998, n23999, n24000, n24001, 
      n24002, n24003, n24004, n24005, n24006, n24007, n24008, n24009, n24010, 
      n24011, n24012, n24013, n24014, n24015, n24016, n24017, n24018, n24019, 
      n24020, n24021, n24022, n24023, n24024, n24025, n24026, n24027, n24028, 
      n24029, n24030, n24031, n24032, n24033, n24034, n24035, n24036, n24037, 
      n24038, n24039, n24040, n24041, n24042, n24043, n24044, n24045, n24046, 
      n24047, n24048, n24049, n24050, n24051, n24052, n24053, n24054, n24055, 
      n24056, n24057, n24058, n24059, n24060, n24061, n24062, n24063, n24064, 
      n24065, n24066, n24067, n24068, n24069, n24070, n24071, n24072, n24073, 
      n24074, n24075, n24076, n24077, n24078, n24079, n24080, n24081, n24082, 
      n24083, n24084, n24085, n24086, n24087, n24088, n24089, n24090, n24091, 
      n24092, n24093, n24094, n24095, n24096, n24097, n24098, n24099, n24100, 
      n24101, n24102, n24103, n24104, n24105, n24106, n24107, n24108, n24109, 
      n24110, n24111, n24112, n24113, n24114, n24115, n24116, n24117, n24118, 
      n24119, n24120, n24121, n24122, n24123, n24124, n24125, n24126, n24127, 
      n24128, n24129, n24130, n24131, n24132, n24133, n24134, n24135, n24136, 
      n24137, n24138, n24139, n24140, n24141, n24142, n24143, n24144, n24145, 
      n24146, n24147, n24148, n24149, n24150, n24151, n24152, n24153, n24154, 
      n24155, n24156, n24157, n24158, n24159, n24160, n24161, n24162, n24163, 
      n24164, n24165, n24166, n24167, n24168, n24169, n24170, n24171, n24172, 
      n24173, n24174, n24175, n24176, n24177, n24178, n24179, n24180, n24181, 
      n24182, n24183, n24184, n24185, n24186, n24187, n24188, n24189, n24190, 
      n24191, n24192, n24193, n24194, n24195, n24196, n24197, n24198, n24199, 
      n24200, n24201, n24202, n24203, n24204, n24205, n24206, n24207, n24208, 
      n24209, n24210, n24211, n24212, n24213, n24214, n24215, n24216, n24217, 
      n24218, n24219, n24220, n24221, n24222, n24223, n24224, n24225, n24226, 
      n24227, n24228, n24229, n24230, n24231, n24232, n24233, n24234, n24235, 
      n24236, n24237, n24238, n24239, n24240, n24241, n24242, n24243, n24244, 
      n24245, n24246, n24247, n24248, n24249, n24250, n24251, n24252, n24253, 
      n24254, n24255, n24256, n24257, n24258, n24259, n24260, n24261, n24262, 
      n24263, n24264, n24265, n24266, n24267, n24268, n24269, n24270, n24271, 
      n24272, n24273, n24274, n24275, n24276, n24277, n24278, n24279, n24280, 
      n24281, n24282, n24283, n24284, n24285, n24286, n24287, n24288, n24289, 
      n24290, n24291, n24292, n24293, n24294, n24295, n24296, n24297, n24298, 
      n24299, n24300, n24301, n24302, n24303, n24304, n24305, n24306, n24307, 
      n24308, n24309, n24310, n24311, n24312, n24313, n24314, n24315, n24316, 
      n24317, n24318, n24319, n24320, n24321, n24322, n24323, n24324, n24325, 
      n24326, n24327, n24328, n24329, n24330, n24331, n24332, n24333, n24334, 
      n24335, n24336, n24337, n24338, n24339, n24340, n24341, n24342, n24343, 
      n24344, n24345, n24346, n24347, n24348, n24349, n24350, n24351, n24352, 
      n24353, n24354, n24355, n24356, n24357, n24358, n24359, n24360, n24361, 
      n24362, n24363, n24364, n24365, n24366, n24367, n24368, n24369, n24370, 
      n24371, n24372, n24373, n24374, n24375, n24376, n24377, n24378, n24379, 
      n24380, n24381, n24382, n24383, n24384, n24385, n24386, n24387, n24388, 
      n24389, n24390, n24391, n24392, n24393, n24394, n24395, n24396, n24397, 
      n24398, n24399, n24400, n24401, n24402, n24403, n24404, n24405, n24406, 
      n24407, n24408, n24409, n24410, n24411, n24412, n24413, n24414, n24415, 
      n24416, n24417, n24418, n24419, n24420, n24421, n24422, n24423, n24424, 
      n24425, n24426, n24427, n24428, n24429, n24430, n24431, n24432, n24433, 
      n24434, n24435, n24436, n24437, n24438, n24439, n24440, n24441, n24442, 
      n24443, n24444, n24445, n24446, n24447, n24448, n24449, n24450, n24451, 
      n24452, n24453, n24454, n24455, n24456, n24457, n24458, n24459, n24460, 
      n24461, n24462, n24463, n24464, n24465, n24466, n24467, n24468, n24469, 
      n24470, n24471, n24472, n24473, n24474, n24475, n24476, n24477, n24478, 
      n24479, n24480, n24481, n24482, n24483, n24484, n24485, n24486, n24487, 
      n24488, n24489, n24490, n24491, n24492, n24493, n24494, n24495, n24496, 
      n24497, n24498, n24499, n24500, n24501, n24502, n24503, n24504, n24505, 
      n24506, n24507, n24508, n24509, n24510, n24511, n24512, n24513, n24514, 
      n24515, n24516, n24517, n24518, n24519, n24520, n24521, n24522, n24523, 
      n24524, n24525, n24526, n24527, n24528, n24529, n24530, n24531, n24532, 
      n24533, n24534, n24535, n24536, n24537, n24538, n24539, n24540, n24541, 
      n24542, n24543, n24544, n24545, n24546, n24547, n24548, n24549, n24550, 
      n24551, n24552, n24553, n24554, n24555, n24556, n24557, n24558, n24559, 
      n24560, n24561, n24562, n24563, n24564, n24565, n24566, n24567, n24568, 
      n24569, n24570, n24571, n24572, n24573, n24574, n24575, n24576, n24577, 
      n24578, n24579, n24580, n24581, n24582, n24583, n24584, n24585, n24586, 
      n24587, n24588, n24589, n24590, n24591, n24592, n24593, n24594, n24595, 
      n24596, n24597, n24598, n24599, n24600, n24601, n24602, n24603, n24604, 
      n24605, n24606, n24607, n24608, n24609, n24610, n24611, n24612, n24613, 
      n24614, n24615, n24616, n24617, n24618, n24619, n24620, n24621, n24622, 
      n24623, n24624, n24625, n24626, n24627, n24628, n24629, n24630, n24631, 
      n24632, n24633, n24634, n24635, n24636, n24637, n24638, n24639, n24640, 
      n24641, n24642, n24643, n24644, n24645, n24646, n24647, n24648, n24649, 
      n24650, n24651, n24652, n24653, n24654, n24655, n24656, n24657, n24658, 
      n24659, n24660, n24661, n24662, n24663, n24664, n24665, n24666, n24667, 
      n24668, n24669, n24670, n24671, n24672, n24673, n24674, n24675, n24676, 
      n24677, n24678, n24679, n24680, n24681, n24682, n24683, n24684, n24685, 
      n24686, n24687, n24688, n24689, n24690, n24691, n24692, n24693, n24694, 
      n24695, n24696, n24697, n24698, n24699, n24700, n24701, n24702, n24703, 
      n24704, n24705, n24706, n24707, n24708, n24709, n24710, n24711, n24712, 
      n24713, n24714, n24715, n24716, n24717, n24718, n24719, n24720, n24721, 
      n24722, n24723, n24724, n24725, n24726, n24727, n24728, n24729, n24730, 
      n24731, n24732, n24733, n24734, n24735, n24736, n24737, n24738, n24739, 
      n24740, n24741, n24742, n24743, n24744, n24745, n24746, n24747, n24748, 
      n24749, n24750, n24751, n24752, n24753, n24754, n24755, n24756, n24757, 
      n24758, n24759, n24760, n24761, n24762, n24763, n24764, n24765, n24766, 
      n24767, n24768, n24769, n24770, n24771, n24772, n24773, n24774, n24775, 
      n24776, n24777, n24778, n24779, n24780, n24781, n24782, n24783, n24784, 
      n24785, n24786, n24787, n24788, n24789, n24790, n24791, n24792, n24793, 
      n24794, n24795, n24796, n24797, n24798, n24799, n24800, n24801, n24802, 
      n24803, n24804, n24805, n24806, n24807, n24808, n24809, n24810, n24811, 
      n24812, n24813, n24814, n24815, n24816, n24817, n24818, n24819, n24820, 
      n24821, n24822, n24823, n24824, n24825, n24826, n24827, n24828, n24829, 
      n24830, n24831, n24832, n24833, n24834, n24835, n24836, n24837, n24838, 
      n24839, n24840, n24841, n24842, n24843, n24844, n24845, n24846, n24847, 
      n24848, n24849, n24850, n24851, n24852, n24853, n24854, n24855, n24856, 
      n24857, n24858, n24859, n24860, n24861, n24862, n24863, n24864, n24865, 
      n24866, n24867, n24868, n24869, n24870, n24871, n24872, n24873, n24874, 
      n24875, n24876, n24877, n24878, n24879, n24880, n24881, n24882, n24883, 
      n24884, n24885, n24886, n24887, n24888, n24889, n24890, n24891, n24892, 
      n24893, n24894, n24895, n24896, n24897, n24898, n24899, n24900, n24901, 
      n24902, n24903, n24904, n24905, n24906, n24907, n24908, n24909, n24910, 
      n24911, n24912, n24913, n24914, n24915, n24916, n24917, n24918, n24919, 
      n24920, n24921, n24922, n24923, n24924, n24925, n24926, n24927, n24928, 
      n24929, n24930, n24931, n24932, n24933, n24934, n24935, n24936, n24937, 
      n24938, n24939, n24940, n24941, n24942, n24943, n24944, n24945, n24946, 
      n24947, n24948, n24949, n24950, n24951, n24952, n24953, n24954, n24955, 
      n24956, n24957, n24958, n24959, n24960, n24961, n24962, n24963, n24964, 
      n24965, n24966, n24967, n24968, n24969, n24970, n24971, n24972, n24973, 
      n24974, n24975, n24976, n24977, n24978, n24979, n24980, n24981, n24982, 
      n24983, n24984, n24985, n24986, n24987, n24988, n24989, n24990, n24991, 
      n24992, n24993, n24994, n24995, n24996, n24997, n24998, n24999, n25000, 
      n25001, n25002, n25003, n25004, n25005, n25006, n25007, n25008, n25009, 
      n25010, n25011, n25012, n25013, n25014, n25015, n25016, n25017, n25018, 
      n25019, n25020, n25021, n25022, n25023, n25024, n25025, n25026, n25027, 
      n25028, n25029, n25030, n25031, n25032, n25033, n25034, n25035, n25036, 
      n25037, n25038, n25039, n25040, n25041, n25042, n25043, n25044, n25045, 
      n25046, n25047, n25048, n25049, n25050, n25051, n25052, n25053, n25054, 
      n25055, n25056, n25057, n25058, n25059, n25060, n25061, n25062, n25063, 
      n25064, n25065, n25066, n25067, n25068, n25069, n25070, n25071, n25072, 
      n25073, n25074, n25075, n25076, n25077, n25078, n25079, n25080, n25081, 
      n25082, n25083, n25084, n25085, n25086, n25087, n25088, n25089, n25090, 
      n25091, n25092, n25093, n25094, n25095, n25096, n25097, n25098, n25099, 
      n25100, n25101, n25102, n25103, n25104, n25105, n25106, n25107, n25108, 
      n25109, n25110, n25111, n25112, n25113, n25114, n25115, n25116, n25117, 
      n25118, n25119, n25120, n25121, n25122, n25123, n25124, n25125, n25126, 
      n25127, n25128, n25129, n25130, n25131, n25132, n25133, n25134, n25135, 
      n25136, n25137, n25138, n25139, n25140, n25141, n25142, n25143, n25144, 
      n25145, n25146, n25147, n25148, n25149, n25150, n25151, n25152, n25153, 
      n25154, n25155, n25156, n25157, n25158, n25159, n25160, n25161, n25162, 
      n25163, n25164, n25165, n25166, n25215, n25216, n25217, n25218, n25219, 
      n25220, n25221, n25222, n25223, n25224, n25225, n25226, n25227, n25228, 
      n25229, n25230, n25231, n25232, n25233, n25234, n25235, n25236, n25237, 
      n25238, n25239, n25240, n25241, n25242, n25243, n25244, n25245, n25246, 
      n25247, n25248, n25249, n25250, n25251, n25252, n25253, n25254, n25255, 
      n25256, n25257, n25258, n25259, n25260, n25261, n25262, n25311, n25312, 
      n25313, n25314, n25315, n25316, n25317, n25318, n25319, n25320, n25321, 
      n25322, n25323, n25324, n25325, n25326, n25327, n25328, n25329, n25330, 
      n25331, n25332, n25333, n25334, n25335, n25336, n25337, n25338, n25339, 
      n25340, n25341, n25342, n25343, n25344, n25345, n25346, n25347, n25348, 
      n25349, n25350, n25351, n25352, n25353, n25354, n25355, n25356, n25357, 
      n25358, n25407, n25408, n25409, n25410, n25411, n25412, n25413, n25414, 
      n25415, n25416, n25417, n25418, n25419, n25420, n25421, n25422, n25423, 
      n25424, n25425, n25426, n25427, n25428, n25429, n25430, n25431, n25432, 
      n25433, n25434, n25435, n25436, n25437, n25438, n25439, n25440, n25441, 
      n25442, n25443, n25444, n25445, n25446, n25447, n25448, n25449, n25450, 
      n25451, n25452, n25453, n25454, n25455, n25456, n25457, n25458, n25459, 
      n25460, n25461, n25462, n25463, n25464, n25465, n25466, n25467, n25468, 
      n25469, n25470, n25471, n25472, n25473, n25474, n25475, n25476, n25477, 
      n25478, n25479, n25480, n25481, n25482, n25483, n25484, n25485, n25486, 
      n25487, n25488, n25489, n25490, n25491, n25492, n25493, n25494, n25495, 
      n25496, n25497, n25498, n25499, n25500, n25501, n25502, n25503, n25504, 
      n25505, n25506, n25507, n25508, n25509, n25510, n25511, n25512, n25513, 
      n25514, n25515, n25516, n25517, n25518, n25519, n25520, n25521, n25522, 
      n25523, n25524, n25525, n25526, n25527, n25528, n25529, n25530, n25531, 
      n25532, n25533, n25534, n25535, n25536, n25537, n25538, n25539, n25540, 
      n25541, n25542, n25543, n25544, n25545, n25546, n25547, n25548, n25549, 
      n25550, n25555, n25556, n25557, n25558, n25563, n25564, n25565, n25566, 
      n25571, n25572, n25573, n25574, n25575, n25576, n25577, n25578, n25579, 
      n25580, n25581, n25582, n25595, n25596, n25597, n25598, n25599, n25600, 
      n25601, n25602, n25603, n25604, n25605, n25606, n25619, n25620, n25621, 
      n25622, n25623, n25624, n25625, n25626, n25627, n25628, n25629, n25630, 
      n25643, n25644, n25645, n25646, n25647, n25648, n25649, n25650, n25651, 
      n25652, n25653, n25654, n25655, n25656, n25657, n25658, n25659, n25660, 
      n25661, n25662, n25663, n25664, n25665, n25666, n25667, n25668, n25669, 
      n25670, n25671, n25672, n25673, n25674, n25675, n25676, n25677, n25678, 
      n25680, n25681, n25682, n25685, n25686, n25687, n25690, n25691, n25692, 
      n25695, n25696, n25697, n25700, n25701, n25702, n25705, n25706, n25707, 
      n25710, n25711, n25712, n25715, n25716, n25717, n25720, n25721, n25722, 
      n25725, n25726, n25727, n25730, n25731, n25732, n25735, n25736, n25737, 
      n25740, n25741, n25742, n25745, n25746, n25747, n25750, n25751, n25752, 
      n25755, n25756, n25757, n25760, n25761, n25762, n25765, n25766, n25767, 
      n25770, n25771, n25772, n25775, n25776, n25777, n25780, n25781, n25782, 
      n25785, n25786, n25787, n25790, n25791, n25792, n25795, n25796, n25797, 
      n25800, n25801, n25802, n25805, n25806, n25807, n25810, n25811, n25812, 
      n25815, n25816, n25817, n25820, n25821, n25822, n25825, n25826, n25827, 
      n25830, n25831, n25832, n25835, n25836, n25837, n25840, n25841, n25842, 
      n25845, n25846, n25847, n25850, n25851, n25852, n25855, n25856, n25857, 
      n25860, n25861, n25862, n25865, n25866, n25867, n25870, n25871, n25872, 
      n25875, n25876, n25877, n25880, n25881, n25882, n25885, n25886, n25887, 
      n25890, n25891, n25892, n25895, n25896, n25897, n25900, n25901, n25902, 
      n25905, n25906, n25907, n25910, n25911, n25912, n25915, n25916, n25917, 
      n25920, n25921, n25922, n25925, n25926, n25927, n25930, n25931, n25932, 
      n25935, n25936, n25937, n25940, n25941, n25942, n25945, n25946, n25947, 
      n25950, n25951, n25952, n25955, n25956, n25957, n25960, n25961, n25962, 
      n25965, n25966, n25967, n25970, n25971, n25972, n25975, n25976, n25977, 
      n25980, n25981, n25982, n25985, n25986, n25987, n25990, n25991, n25992, 
      n25995, n25996, n25997, n26191, n26192, n26193, n26194, n26195, n26196, 
      n26197, n26198, n26207, n26208, n26209, n26210, n26211, n26212, n26213, 
      n26214, n26215, n26216, n26217, n26218, n26219, n26220, n26221, n26222, 
      n26223, n26224, n26225, n26226, n26227, n26228, n26229, n26230, n26231, 
      n26232, n26233, n26234, n26235, n26236, n26237, n26238, n26239, n26240, 
      n26241, n26242, n26243, n26244, n26245, n26246, n26247, n26248, n26249, 
      n26250, n26251, n26252, n26253, n26254, n26255, n26256, n26257, n26258, 
      n26259, n26260, n26261, n26262, n26263, n26264, n26265, n26266, n26327, 
      n26328, n26329, n26330, n26331, n26332, n26333, n26334, n26335, n26336, 
      n26337, n26338, n26339, n26340, n26341, n26342, n26343, n26344, n26345, 
      n26346, n26347, n26348, n26349, n26350, n26351, n26352, n26353, n26354, 
      n26355, n26356, n26357, n26358, n26359, n26360, n26361, n26362, n26363, 
      n26364, n26365, n26366, n26367, n26368, n26369, n26370, n26371, n26372, 
      n26373, n26374, n26375, n26376, n26377, n26378, n26379, n26380, n26381, 
      n26382, n26383, n26384, n26385, n26386, n26447, n26448, n26449, n26450, 
      n26451, n26452, n26453, n26454, n26455, n26456, n26457, n26458, n26459, 
      n26460, n26461, n26462, n26463, n26464, n26465, n26466, n26467, n26468, 
      n26469, n26470, n26471, n26472, n26473, n26474, n26475, n26476, n26477, 
      n26478, n26479, n26480, n26481, n26482, n26483, n26484, n26485, n26486, 
      n26487, n26488, n26489, n26490, n26491, n26492, n26493, n26494, n26495, 
      n26496, n26497, n26498, n26499, n26500, n26501, n26502, n26503, n26504, 
      n26505, n26506, n26507, n26508, n26509, n26510, n26511, n26512, n26513, 
      n26514, n26515, n26516, n26517, n26518, n26519, n26520, n26521, n26522, 
      n26523, n26524, n26525, n26526, n26527, n26528, n26529, n26530, n26531, 
      n26532, n26533, n26534, n26535, n26536, n26537, n26538, n26539, n26540, 
      n26541, n26542, n26543, n26544, n26545, n26546, n26547, n26548, n26549, 
      n26550, n26551, n26552, n26553, n26554, n26555, n26556, n26557, n26558, 
      n26559, n26560, n26561, n26562, n26563, n26564, n26565, n26566, n26567, 
      n26568, n26569, n26570, n26571, n26572, n26573, n26574, n26575, n26576, 
      n26577, n26578, n26579, n26580, n26581, n26582, n26583, n26584, n26585, 
      n26586, n26587, n26588, n26589, n26590, n26591, n26592, n26593, n26594, 
      n26595, n26596, n26597, n26598, n26599, n26600, n26601, n26602, n26603, 
      n26604, n26605, n26606, n26607, n26608, n26609, n26610, n26611, n26612, 
      n26613, n26614, n26615, n26616, n26617, n26618, n26619, n26620, n26621, 
      n26622, n26623, n26624, n26625, n26626, n26627, n26628, n26629, n26630, 
      n26631, n26632, n26633, n26634, n26635, n26636, n26637, n26638, n26639, 
      n26640, n26641, n26642, n26643, n26644, n26645, n26646, n26647, n26648, 
      n26649, n26650, n26651, n26652, n26653, n26654, n26655, n26656, n26657, 
      n26658, n26659, n26660, n26661, n26662, n26663, n26664, n26665, n26666, 
      n26667, n26668, n26669, n26670, n26671, n26672, n26673, n26674, n26675, 
      n26676, n26677, n26678, n26679, n26680, n26681, n26682, n26683, n26684, 
      n26685, n26686, n26687, n26688, n26689, n26690, n26691, n26692, n26693, 
      n26694, n26695, n26696, n26697, n26698, n26699, n26700, n26701, n26702, 
      n26703, n26704, n26705, n26706, n26707, n26708, n26709, n26710, n26711, 
      n26712, n26713, n26714, n26715, n26716, n26717, n26718, n26719, n26720, 
      n26721, n26722, n26723, n26724, n26725, n26726, n26727, n26728, n26729, 
      n26730, n26731, n26732, n26733, n26734, n26735, n26736, n26737, n26738, 
      n26739, n26740, n26741, n26742, n26743, n26744, n26745, n26746, n26747, 
      n26748, n26749, n26750, n26751, n26752, n26753, n26754, n26755, n26756, 
      n26757, n26758, n26759, n26760, n26761, n26762, n26763, n26764, n26765, 
      n26766, n26767, n26768, n26769, n26770, n26771, n26772, n26773, n26774, 
      n26775, n26776, n26777, n26778, n26779, n26780, n26781, n26782, n26783, 
      n26784, n26785, n26786, n26787, n26788, n26789, n26790, n26791, n26792, 
      n26793, n26794, n26795, n26796, n26797, n26798, n26799, n26800, n26801, 
      n26802, n26803, n26804, n26805, n26806, n26807, n26808, n26809, n26810, 
      n26811, n26812, n26813, n26814, n26815, n26816, n26817, n26818, n26819, 
      n26820, n26821, n26822, n26823, n26824, n26825, n26826, n26827, n26828, 
      n26829, n26830, n26831, n26832, n26833, n26834, n26835, n26836, n26837, 
      n26838, n26839, n26840, n26841, n26842, n26843, n26844, n26845, n26846, 
      n26847, n26848, n26849, n26850, n26851, n26852, n26853, n26854, n26855, 
      n26856, n26857, n26858, n26859, n26860, n26861, n26862, n26863, n26864, 
      n26865, n26866, n26867, n26868, n26869, n26870, n26871, n26872, n26873, 
      n26874, n26875, n26876, n26877, n26878, n26879, n26880, n26881, n26882, 
      n26883, n26884, n26885, n26886, n26887, n26888, n26889, n26890, n26891, 
      n26892, n26893, n26894, n26895, n26896, n26897, n26898, n26899, n26900, 
      n26901, n26902, n26903, n26904, n26905, n26906, n26907, n26908, n26909, 
      n26910, n26911, n26912, n26913, n26914, n26915, n26916, n26917, n26918, 
      n26919, n26920, n26921, n26922, n26923, n26924, n26925, n26926, n26927, 
      n26928, n26929, n26930, n26931, n26932, n26933, n26934, n26935, n26936, 
      n26937, n26938, n26939, n26940, n26941, n26942, n26943, n26944, n26945, 
      n26946, n26947, n26948, n26949, n26950, n26951, n26952, n26953, n26954, 
      n26955, n26956, n26957, n26958, n26959, n26960, n26961, n26962, n26963, 
      n26964, n26965, n26966, n26967, n26968, n26969, n26970, n26971, n26972, 
      n26973, n26974, n26975, n26976, n26977, n26978, n26979, n26980, n26981, 
      n26982, n26983, n26984, n26985, n26986, n26987, n26988, n26989, n26990, 
      n26991, n26992, n26993, n26994, n26995, n26996, n26997, n26998, n26999, 
      n27000, n27001, n27002, n27003, n27004, n27005, n27006, n27007, n27008, 
      n27009, n27010, n27011, n27012, n27013, n27014, n27015, n27016, n27017, 
      n27018, n27019, n27020, n27021, n27022, n27023, n27024, n27025, n27026, 
      n27027, n27028, n27029, n27030, n27031, n27032, n27033, n27034, n27035, 
      n27036, n27037, n27038, n27039, n27040, n27041, n27042, n27043, n27044, 
      n27045, n27046, n27047, n27048, n27049, n27050, n27051, n27052, n27053, 
      n27054, n27055, n27056, n27057, n27058, n27059, n27060, n27061, n27062, 
      n27063, n27064, n27065, n27066, n27067, n27068, n27069, n27070, n27071, 
      n27072, n27073, n27074, n27075, n27076, n27077, n27078, n27079, n27080, 
      n27081, n27082, n27083, n27084, n27085, n27086, n27087, n27088, n27089, 
      n27090, n27091, n27092, n27093, n27094, n27095, n27096, n27097, n27098, 
      n27099, n27100, n27101, n27102, n27103, n27104, n27105, n27106, n27107, 
      n27108, n27109, n27110, n27111, n27112, n27113, n27114, n27115, n27116, 
      n27117, n27118, n27119, n27120, n27121, n27122, n27123, n27124, n27125, 
      n27126, n27127, n27128, n27129, n27130, n27131, n27132, n27133, n27134, 
      n27135, n27136, n27137, n27138, n27139, n27140, n27141, n27142, n27143, 
      n27144, n27145, n27146, n27147, n27148, n27149, n27150, n27151, n27152, 
      n27153, n27154, n27155, n27156, n27157, n27158, n27159, n27160, n27161, 
      n27162, n27163, n27164, n27165, n27166, n27167, n27168, n27169, n27170, 
      n27171, n27172, n27173, n27174, n27175, n27176, n27177, n27178, n27179, 
      n27180, n27181, n27182, n27183, n27184, n27185, n27186, n27187, n27188, 
      n27189, n27190, n27191, n27192, n27193, n27194, n27195, n27196, n27197, 
      n27198, n27199, n27200, n27201, n27202, n27203, n27204, n27205, n27206, 
      n27207, n27208, n27209, n27210, n27211, n27212, n27213, n27214, n27215, 
      n27216, n27217, n27218, n27219, n27220, n27221, n27222, n27223, n27224, 
      n27225, n27226, n27227, n27228, n27229, n27230, n27231, n27232, n27233, 
      n27234, n27235, n27236, n27237, n27238, n27239, n27240, n27241, n27242, 
      n27243, n27244, n27245, n27246, n27247, n27248, n27249, n27250, n27251, 
      n27252, n27253, n27254, n27255, n27256, n27257, n27258, n27259, n27260, 
      n27261, n27262, n27263, n27264, n27265, n27266, n27267, n27268, n27269, 
      n27270, n27271, n27272, n27273, n27274, n27275, n27276, n27277, n27278, 
      n27279, n27280, n27281, n27282, n27283, n27284, n27285, n27286, n27287, 
      n27288, n27289, n27290, n27291, n27292, n27293, n27294, n27295, n27296, 
      n27297, n27298, n27299, n27300, n27301, n27302, n27303, n27304, n27305, 
      n27306, n27307, n27308, n27309, n27310, n27311, n27312, n27313, n27314, 
      n27315, n27316, n27317, n27318, n27319, n27320, n27321, n27322, n27323, 
      n27324, n27325, n27326, n27327, n27328, n27329, n27330, n27331, n27332, 
      n27333, n27334, n27335, n27336, n27337, n27338, n27339, n27340, n27341, 
      n27342, n27343, n27344, n27345, n27346, n27347, n27348, n27349, n27350, 
      n27351, n27352, n27353, n27354, n27355, n27356, n27357, n27358, n27359, 
      n27360, n27361, n27362, n27363, n27364, n27365, n27366, n27367, n27368, 
      n27369, n27370, n27371, n27372, n27373, n27374, n27375, n27376, n27377, 
      n27378, n27379, n27380, n27381, n27382, n27383, n27384, n27385, n27386, 
      n27387, n27388, n27389, n27390, n27391, n27392, n27393, n27394, n27395, 
      n27396, n27397, n27398, n27399, n27400, n27401, n27402, n27403, n27404, 
      n27405, n27406, n27407, n27408, n27409, n27410, n27411, n27412, n27413, 
      n27414, n27415, n27416, n27417, n27418, n27419, n27420, n27421, n27422, 
      n27423, n27424, n27425, n27426, n27427, n27428, n27429, n27430, n27431, 
      n27432, n27433, n27434, n27435, n27436, n27437, n27438, n27439, n27440, 
      n27441, n27442, n27443, n27444, n27445, n27446, n27447, n27448, n27449, 
      n27450, n27451, n27452, n27453, n27454, n27455, n27456, n27457, n27458, 
      n27459, n27460, n27461, n27462, n27463, n27464, n27465, n27466, n27467, 
      n27468, n27469, n27470, n27471, n27472, n27473, n27474, n27475, n27476, 
      n27477, n27478, n27479, n27480, n27481, n27482, n27483, n27484, n27485, 
      n27486, n27487, n_1000, n_1001, n_1002, n_1003, n_1004, n_1005, n_1006, 
      n_1007, n_1008, n_1009, n_1010, n_1011, n_1012, n_1013, n_1014, n_1015, 
      n_1016, n_1017, n_1018, n_1019, n_1020, n_1021, n_1022, n_1023, n_1024, 
      n_1025, n_1026, n_1027, n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, 
      n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, 
      n_1043, n_1044, n_1045, n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, 
      n_1052, n_1053, n_1054, n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, 
      n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, n_1068, n_1069, 
      n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, 
      n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, 
      n_1088, n_1089, n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, 
      n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, 
      n_1106, n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, 
      n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, 
      n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, 
      n_1133, n_1134, n_1135, n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, 
      n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, 
      n_1151, n_1152, n_1153, n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, 
      n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, 
      n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, 
      n_1178, n_1179, n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, 
      n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, 
      n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, 
      n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, 
      n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, 
      n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, 
      n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, 
      n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, 
      n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, 
      n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, 
      n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, 
      n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, 
      n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, 
      n_1295, n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, 
      n_1304, n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, 
      n_1313, n_1314, n_1315, n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, 
      n_1322, n_1323, n_1324, n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, 
      n_1331, n_1332, n_1333, n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, 
      n_1340, n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, 
      n_1349, n_1350, n_1351, n_1352, n_1353, n_1354, n_1355, n_1356, n_1357, 
      n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, n_1364, n_1365, n_1366, 
      n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, n_1373, n_1374, n_1375, 
      n_1376, n_1377, n_1378, n_1379, n_1380, n_1381, n_1382, n_1383, n_1384, 
      n_1385, n_1386, n_1387, n_1388, n_1389, n_1390, n_1391, n_1392, n_1393, 
      n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, n_1400, n_1401, n_1402, 
      n_1403, n_1404, n_1405, n_1406, n_1407, n_1408, n_1409, n_1410, n_1411, 
      n_1412, n_1413, n_1414, n_1415, n_1416, n_1417, n_1418, n_1419, n_1420, 
      n_1421, n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, n_1428, n_1429, 
      n_1430, n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, n_1437, n_1438, 
      n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, n_1445, n_1446, n_1447, 
      n_1448, n_1449, n_1450, n_1451, n_1452, n_1453, n_1454, n_1455, n_1456, 
      n_1457, n_1458, n_1459, n_1460, n_1461, n_1462, n_1463, n_1464, n_1465, 
      n_1466, n_1467, n_1468, n_1469, n_1470, n_1471, n_1472, n_1473, n_1474, 
      n_1475, n_1476, n_1477, n_1478, n_1479, n_1480, n_1481, n_1482, n_1483, 
      n_1484, n_1485, n_1486, n_1487, n_1488, n_1489, n_1490, n_1491, n_1492, 
      n_1493, n_1494, n_1495, n_1496, n_1497, n_1498, n_1499, n_1500, n_1501, 
      n_1502, n_1503, n_1504, n_1505, n_1506, n_1507, n_1508, n_1509, n_1510, 
      n_1511, n_1512, n_1513, n_1514, n_1515, n_1516, n_1517, n_1518, n_1519, 
      n_1520, n_1521, n_1522, n_1523, n_1524, n_1525, n_1526, n_1527, n_1528, 
      n_1529, n_1530, n_1531, n_1532, n_1533, n_1534, n_1535, n_1536, n_1537, 
      n_1538, n_1539, n_1540, n_1541, n_1542, n_1543, n_1544, n_1545, n_1546, 
      n_1547, n_1548, n_1549, n_1550, n_1551, n_1552, n_1553, n_1554, n_1555, 
      n_1556, n_1557, n_1558, n_1559, n_1560, n_1561, n_1562, n_1563, n_1564, 
      n_1565, n_1566, n_1567, n_1568, n_1569, n_1570, n_1571, n_1572, n_1573, 
      n_1574, n_1575, n_1576, n_1577, n_1578, n_1579, n_1580, n_1581, n_1582, 
      n_1583, n_1584, n_1585, n_1586, n_1587, n_1588, n_1589, n_1590, n_1591, 
      n_1592, n_1593, n_1594, n_1595, n_1596, n_1597, n_1598, n_1599, n_1600, 
      n_1601, n_1602, n_1603, n_1604, n_1605, n_1606, n_1607, n_1608, n_1609, 
      n_1610, n_1611, n_1612, n_1613, n_1614, n_1615, n_1616, n_1617, n_1618, 
      n_1619, n_1620, n_1621, n_1622, n_1623, n_1624, n_1625, n_1626, n_1627, 
      n_1628, n_1629, n_1630, n_1631, n_1632, n_1633, n_1634, n_1635, n_1636, 
      n_1637, n_1638, n_1639, n_1640, n_1641, n_1642, n_1643, n_1644, n_1645, 
      n_1646, n_1647, n_1648, n_1649, n_1650, n_1651, n_1652, n_1653, n_1654, 
      n_1655, n_1656, n_1657, n_1658, n_1659, n_1660, n_1661, n_1662, n_1663, 
      n_1664, n_1665, n_1666, n_1667, n_1668, n_1669, n_1670, n_1671, n_1672, 
      n_1673, n_1674, n_1675, n_1676, n_1677, n_1678, n_1679, n_1680, n_1681, 
      n_1682, n_1683, n_1684, n_1685, n_1686, n_1687, n_1688, n_1689, n_1690, 
      n_1691, n_1692, n_1693, n_1694, n_1695, n_1696, n_1697, n_1698, n_1699, 
      n_1700, n_1701, n_1702, n_1703, n_1704, n_1705, n_1706, n_1707, n_1708, 
      n_1709, n_1710, n_1711, n_1712, n_1713, n_1714, n_1715, n_1716, n_1717, 
      n_1718, n_1719, n_1720, n_1721, n_1722, n_1723, n_1724, n_1725, n_1726, 
      n_1727, n_1728, n_1729, n_1730, n_1731, n_1732, n_1733, n_1734, n_1735, 
      n_1736, n_1737, n_1738, n_1739, n_1740, n_1741, n_1742, n_1743, n_1744, 
      n_1745, n_1746, n_1747, n_1748, n_1749, n_1750, n_1751, n_1752, n_1753, 
      n_1754, n_1755, n_1756, n_1757, n_1758, n_1759, n_1760, n_1761, n_1762, 
      n_1763, n_1764, n_1765, n_1766, n_1767, n_1768, n_1769, n_1770, n_1771, 
      n_1772, n_1773, n_1774, n_1775, n_1776, n_1777, n_1778, n_1779, n_1780, 
      n_1781, n_1782, n_1783, n_1784, n_1785, n_1786, n_1787, n_1788, n_1789, 
      n_1790, n_1791, n_1792, n_1793, n_1794, n_1795, n_1796, n_1797, n_1798, 
      n_1799, n_1800, n_1801, n_1802, n_1803, n_1804, n_1805, n_1806, n_1807, 
      n_1808, n_1809, n_1810, n_1811, n_1812, n_1813, n_1814, n_1815, n_1816, 
      n_1817, n_1818, n_1819, n_1820, n_1821, n_1822, n_1823, n_1824, n_1825, 
      n_1826, n_1827, n_1828, n_1829, n_1830, n_1831, n_1832, n_1833, n_1834, 
      n_1835, n_1836, n_1837, n_1838, n_1839, n_1840, n_1841, n_1842, n_1843, 
      n_1844, n_1845, n_1846, n_1847, n_1848, n_1849, n_1850, n_1851, n_1852, 
      n_1853, n_1854, n_1855, n_1856, n_1857, n_1858, n_1859, n_1860, n_1861, 
      n_1862, n_1863, n_1864, n_1865, n_1866, n_1867, n_1868, n_1869, n_1870, 
      n_1871, n_1872, n_1873, n_1874, n_1875, n_1876, n_1877, n_1878, n_1879, 
      n_1880, n_1881, n_1882, n_1883, n_1884, n_1885, n_1886, n_1887, n_1888, 
      n_1889, n_1890, n_1891, n_1892, n_1893, n_1894, n_1895, n_1896, n_1897, 
      n_1898, n_1899, n_1900, n_1901, n_1902, n_1903, n_1904, n_1905, n_1906, 
      n_1907, n_1908, n_1909, n_1910, n_1911, n_1912, n_1913, n_1914, n_1915, 
      n_1916, n_1917, n_1918, n_1919, n_1920, n_1921, n_1922, n_1923, n_1924, 
      n_1925, n_1926, n_1927, n_1928, n_1929, n_1930, n_1931, n_1932, n_1933, 
      n_1934, n_1935, n_1936, n_1937, n_1938, n_1939, n_1940, n_1941, n_1942, 
      n_1943, n_1944, n_1945, n_1946, n_1947, n_1948, n_1949, n_1950, n_1951, 
      n_1952, n_1953, n_1954, n_1955, n_1956, n_1957, n_1958, n_1959, n_1960, 
      n_1961, n_1962, n_1963, n_1964, n_1965, n_1966, n_1967, n_1968, n_1969, 
      n_1970, n_1971, n_1972, n_1973, n_1974, n_1975, n_1976, n_1977, n_1978, 
      n_1979, n_1980, n_1981, n_1982, n_1983, n_1984, n_1985, n_1986, n_1987, 
      n_1988, n_1989, n_1990, n_1991, n_1992, n_1993, n_1994, n_1995, n_1996, 
      n_1997, n_1998, n_1999, n_2000, n_2001, n_2002, n_2003, n_2004, n_2005, 
      n_2006, n_2007, n_2008, n_2009, n_2010, n_2011, n_2012, n_2013, n_2014, 
      n_2015, n_2016, n_2017, n_2018, n_2019, n_2020, n_2021, n_2022, n_2023, 
      n_2024, n_2025, n_2026, n_2027, n_2028, n_2029, n_2030, n_2031, n_2032, 
      n_2033, n_2034, n_2035, n_2036, n_2037, n_2038, n_2039, n_2040, n_2041, 
      n_2042, n_2043, n_2044, n_2045, n_2046, n_2047, n_2048, n_2049, n_2050, 
      n_2051, n_2052, n_2053, n_2054, n_2055, n_2056, n_2057, n_2058, n_2059, 
      n_2060, n_2061, n_2062, n_2063, n_2064, n_2065, n_2066, n_2067, n_2068, 
      n_2069, n_2070, n_2071, n_2072, n_2073, n_2074, n_2075, n_2076, n_2077, 
      n_2078, n_2079, n_2080, n_2081, n_2082, n_2083, n_2084, n_2085, n_2086, 
      n_2087 : std_logic;

begin
   
   OUT1_reg_63_inst : DFF_X1 port map( D => n6017, CK => CLK, Q => n4098, QN =>
                           n_1000);
   OUT1_tri_enable_reg_63_inst : DFF_X1 port map( D => n19582, CK => CLK, Q => 
                           n4099, QN => n18303);
   OUT1_reg_62_inst : DFF_X1 port map( D => n6015, CK => CLK, Q => n4100, QN =>
                           n_1001);
   OUT1_tri_enable_reg_62_inst : DFF_X1 port map( D => n19578, CK => CLK, Q => 
                           n4101, QN => n18304);
   OUT1_reg_61_inst : DFF_X1 port map( D => n6013, CK => CLK, Q => n4102, QN =>
                           n_1002);
   OUT1_tri_enable_reg_61_inst : DFF_X1 port map( D => n19581, CK => CLK, Q => 
                           n4103, QN => n18305);
   OUT1_reg_60_inst : DFF_X1 port map( D => n6011, CK => CLK, Q => n4104, QN =>
                           n_1003);
   OUT1_tri_enable_reg_60_inst : DFF_X1 port map( D => n19576, CK => CLK, Q => 
                           n4105, QN => n18306);
   OUT1_reg_59_inst : DFF_X1 port map( D => n6009, CK => CLK, Q => n4106, QN =>
                           n_1004);
   OUT1_tri_enable_reg_59_inst : DFF_X1 port map( D => n19579, CK => CLK, Q => 
                           n4107, QN => n18307);
   OUT1_reg_58_inst : DFF_X1 port map( D => n6007, CK => CLK, Q => n4108, QN =>
                           n_1005);
   OUT1_tri_enable_reg_58_inst : DFF_X1 port map( D => n19549, CK => CLK, Q => 
                           n4109, QN => n18308);
   OUT1_reg_57_inst : DFF_X1 port map( D => n6005, CK => CLK, Q => n4110, QN =>
                           n_1006);
   OUT1_tri_enable_reg_57_inst : DFF_X1 port map( D => n19577, CK => CLK, Q => 
                           n4111, QN => n18309);
   OUT1_reg_56_inst : DFF_X1 port map( D => n6003, CK => CLK, Q => n4112, QN =>
                           n_1007);
   OUT1_tri_enable_reg_56_inst : DFF_X1 port map( D => n19574, CK => CLK, Q => 
                           n4113, QN => n18310);
   OUT1_reg_55_inst : DFF_X1 port map( D => n6001, CK => CLK, Q => n4114, QN =>
                           n_1008);
   OUT1_tri_enable_reg_55_inst : DFF_X1 port map( D => n19575, CK => CLK, Q => 
                           n4115, QN => n18311);
   OUT1_reg_54_inst : DFF_X1 port map( D => n5999, CK => CLK, Q => n4116, QN =>
                           n_1009);
   OUT1_tri_enable_reg_54_inst : DFF_X1 port map( D => n19572, CK => CLK, Q => 
                           n4117, QN => n18312);
   OUT1_reg_53_inst : DFF_X1 port map( D => n5997, CK => CLK, Q => n4118, QN =>
                           n_1010);
   OUT1_tri_enable_reg_53_inst : DFF_X1 port map( D => n19573, CK => CLK, Q => 
                           n4119, QN => n18313);
   OUT1_reg_52_inst : DFF_X1 port map( D => n5995, CK => CLK, Q => n4120, QN =>
                           n_1011);
   OUT1_tri_enable_reg_52_inst : DFF_X1 port map( D => n19570, CK => CLK, Q => 
                           n4121, QN => n18314);
   OUT1_reg_51_inst : DFF_X1 port map( D => n5993, CK => CLK, Q => n4122, QN =>
                           n_1012);
   OUT1_tri_enable_reg_51_inst : DFF_X1 port map( D => n19571, CK => CLK, Q => 
                           n4123, QN => n18315);
   OUT1_reg_50_inst : DFF_X1 port map( D => n5991, CK => CLK, Q => n4124, QN =>
                           n_1013);
   OUT1_tri_enable_reg_50_inst : DFF_X1 port map( D => n19568, CK => CLK, Q => 
                           n4125, QN => n18316);
   OUT1_reg_49_inst : DFF_X1 port map( D => n5989, CK => CLK, Q => n4126, QN =>
                           n_1014);
   OUT1_tri_enable_reg_49_inst : DFF_X1 port map( D => n19569, CK => CLK, Q => 
                           n4127, QN => n18317);
   OUT1_reg_48_inst : DFF_X1 port map( D => n5987, CK => CLK, Q => n4128, QN =>
                           n_1015);
   OUT1_tri_enable_reg_48_inst : DFF_X1 port map( D => n19566, CK => CLK, Q => 
                           n4129, QN => n18318);
   OUT1_reg_47_inst : DFF_X1 port map( D => n5985, CK => CLK, Q => n4130, QN =>
                           n_1016);
   OUT1_tri_enable_reg_47_inst : DFF_X1 port map( D => n19567, CK => CLK, Q => 
                           n4131, QN => n18319);
   OUT1_reg_46_inst : DFF_X1 port map( D => n5983, CK => CLK, Q => n4132, QN =>
                           n_1017);
   OUT1_tri_enable_reg_46_inst : DFF_X1 port map( D => n19564, CK => CLK, Q => 
                           n4133, QN => n18320);
   OUT1_reg_45_inst : DFF_X1 port map( D => n5981, CK => CLK, Q => n4134, QN =>
                           n_1018);
   OUT1_tri_enable_reg_45_inst : DFF_X1 port map( D => n19565, CK => CLK, Q => 
                           n4135, QN => n18321);
   OUT1_reg_44_inst : DFF_X1 port map( D => n5979, CK => CLK, Q => n4136, QN =>
                           n_1019);
   OUT1_tri_enable_reg_44_inst : DFF_X1 port map( D => n19562, CK => CLK, Q => 
                           n4137, QN => n18322);
   OUT1_reg_43_inst : DFF_X1 port map( D => n5977, CK => CLK, Q => n4138, QN =>
                           n_1020);
   OUT1_tri_enable_reg_43_inst : DFF_X1 port map( D => n19563, CK => CLK, Q => 
                           n4139, QN => n18323);
   OUT1_reg_42_inst : DFF_X1 port map( D => n5975, CK => CLK, Q => n4140, QN =>
                           n_1021);
   OUT1_tri_enable_reg_42_inst : DFF_X1 port map( D => n19560, CK => CLK, Q => 
                           n4141, QN => n18324);
   OUT1_reg_41_inst : DFF_X1 port map( D => n5973, CK => CLK, Q => n4142, QN =>
                           n_1022);
   OUT1_tri_enable_reg_41_inst : DFF_X1 port map( D => n19561, CK => CLK, Q => 
                           n4143, QN => n18325);
   OUT1_reg_40_inst : DFF_X1 port map( D => n5971, CK => CLK, Q => n4144, QN =>
                           n_1023);
   OUT1_tri_enable_reg_40_inst : DFF_X1 port map( D => n19558, CK => CLK, Q => 
                           n4145, QN => n18326);
   OUT1_reg_39_inst : DFF_X1 port map( D => n5969, CK => CLK, Q => n4146, QN =>
                           n_1024);
   OUT1_tri_enable_reg_39_inst : DFF_X1 port map( D => n19559, CK => CLK, Q => 
                           n4147, QN => n18327);
   OUT1_reg_38_inst : DFF_X1 port map( D => n5967, CK => CLK, Q => n4148, QN =>
                           n_1025);
   OUT1_tri_enable_reg_38_inst : DFF_X1 port map( D => n19556, CK => CLK, Q => 
                           n4149, QN => n18328);
   OUT1_reg_37_inst : DFF_X1 port map( D => n5965, CK => CLK, Q => n4150, QN =>
                           n_1026);
   OUT1_tri_enable_reg_37_inst : DFF_X1 port map( D => n19557, CK => CLK, Q => 
                           n4151, QN => n18329);
   OUT1_reg_36_inst : DFF_X1 port map( D => n5963, CK => CLK, Q => n4152, QN =>
                           n_1027);
   OUT1_tri_enable_reg_36_inst : DFF_X1 port map( D => n19554, CK => CLK, Q => 
                           n4153, QN => n18330);
   OUT1_reg_35_inst : DFF_X1 port map( D => n5961, CK => CLK, Q => n4154, QN =>
                           n_1028);
   OUT1_tri_enable_reg_35_inst : DFF_X1 port map( D => n19555, CK => CLK, Q => 
                           n4155, QN => n18331);
   OUT1_reg_34_inst : DFF_X1 port map( D => n5959, CK => CLK, Q => n4156, QN =>
                           n_1029);
   OUT1_tri_enable_reg_34_inst : DFF_X1 port map( D => n19552, CK => CLK, Q => 
                           n4157, QN => n18332);
   OUT1_reg_33_inst : DFF_X1 port map( D => n5957, CK => CLK, Q => n4158, QN =>
                           n_1030);
   OUT1_tri_enable_reg_33_inst : DFF_X1 port map( D => n19553, CK => CLK, Q => 
                           n4159, QN => n18333);
   OUT1_reg_32_inst : DFF_X1 port map( D => n5955, CK => CLK, Q => n4160, QN =>
                           n_1031);
   OUT1_tri_enable_reg_32_inst : DFF_X1 port map( D => n19519, CK => CLK, Q => 
                           n4161, QN => n18334);
   OUT1_reg_31_inst : DFF_X1 port map( D => n5953, CK => CLK, Q => n4162, QN =>
                           n_1032);
   OUT1_tri_enable_reg_31_inst : DFF_X1 port map( D => n19551, CK => CLK, Q => 
                           n4163, QN => n18335);
   OUT1_reg_30_inst : DFF_X1 port map( D => n5951, CK => CLK, Q => n4164, QN =>
                           n_1033);
   OUT1_tri_enable_reg_30_inst : DFF_X1 port map( D => n19550, CK => CLK, Q => 
                           n4165, QN => n18336);
   OUT1_reg_29_inst : DFF_X1 port map( D => n5949, CK => CLK, Q => n4166, QN =>
                           n_1034);
   OUT1_tri_enable_reg_29_inst : DFF_X1 port map( D => n19520, CK => CLK, Q => 
                           n4167, QN => n18337);
   OUT1_reg_28_inst : DFF_X1 port map( D => n5947, CK => CLK, Q => n4168, QN =>
                           n_1035);
   OUT1_tri_enable_reg_28_inst : DFF_X1 port map( D => n19548, CK => CLK, Q => 
                           n4169, QN => n18338);
   OUT1_reg_27_inst : DFF_X1 port map( D => n5945, CK => CLK, Q => n4170, QN =>
                           n_1036);
   OUT1_tri_enable_reg_27_inst : DFF_X1 port map( D => n19547, CK => CLK, Q => 
                           n4171, QN => n18339);
   OUT1_reg_26_inst : DFF_X1 port map( D => n5943, CK => CLK, Q => n4172, QN =>
                           n_1037);
   OUT1_tri_enable_reg_26_inst : DFF_X1 port map( D => n19546, CK => CLK, Q => 
                           n4173, QN => n18340);
   OUT1_reg_25_inst : DFF_X1 port map( D => n5941, CK => CLK, Q => n4174, QN =>
                           n_1038);
   OUT1_tri_enable_reg_25_inst : DFF_X1 port map( D => n19545, CK => CLK, Q => 
                           n4175, QN => n18341);
   OUT1_reg_24_inst : DFF_X1 port map( D => n5939, CK => CLK, Q => n4176, QN =>
                           n_1039);
   OUT1_tri_enable_reg_24_inst : DFF_X1 port map( D => n19544, CK => CLK, Q => 
                           n4177, QN => n18342);
   OUT1_reg_23_inst : DFF_X1 port map( D => n5937, CK => CLK, Q => n4178, QN =>
                           n_1040);
   OUT1_tri_enable_reg_23_inst : DFF_X1 port map( D => n19543, CK => CLK, Q => 
                           n4179, QN => n18343);
   OUT1_reg_22_inst : DFF_X1 port map( D => n5935, CK => CLK, Q => n4180, QN =>
                           n_1041);
   OUT1_tri_enable_reg_22_inst : DFF_X1 port map( D => n19542, CK => CLK, Q => 
                           n4181, QN => n18344);
   OUT1_reg_21_inst : DFF_X1 port map( D => n5933, CK => CLK, Q => n4182, QN =>
                           n_1042);
   OUT1_tri_enable_reg_21_inst : DFF_X1 port map( D => n19541, CK => CLK, Q => 
                           n4183, QN => n18345);
   OUT1_reg_20_inst : DFF_X1 port map( D => n5931, CK => CLK, Q => n4184, QN =>
                           n_1043);
   OUT1_tri_enable_reg_20_inst : DFF_X1 port map( D => n19540, CK => CLK, Q => 
                           n4185, QN => n18346);
   OUT1_reg_19_inst : DFF_X1 port map( D => n5929, CK => CLK, Q => n4186, QN =>
                           n_1044);
   OUT1_tri_enable_reg_19_inst : DFF_X1 port map( D => n19539, CK => CLK, Q => 
                           n4187, QN => n18347);
   OUT1_reg_18_inst : DFF_X1 port map( D => n5927, CK => CLK, Q => n4188, QN =>
                           n_1045);
   OUT1_tri_enable_reg_18_inst : DFF_X1 port map( D => n19538, CK => CLK, Q => 
                           n4189, QN => n18348);
   OUT1_reg_17_inst : DFF_X1 port map( D => n5925, CK => CLK, Q => n4190, QN =>
                           n_1046);
   OUT1_tri_enable_reg_17_inst : DFF_X1 port map( D => n19537, CK => CLK, Q => 
                           n4191, QN => n18349);
   OUT1_reg_16_inst : DFF_X1 port map( D => n5923, CK => CLK, Q => n4192, QN =>
                           n_1047);
   OUT1_tri_enable_reg_16_inst : DFF_X1 port map( D => n19536, CK => CLK, Q => 
                           n4193, QN => n18350);
   OUT1_reg_15_inst : DFF_X1 port map( D => n5921, CK => CLK, Q => n4194, QN =>
                           n_1048);
   OUT1_tri_enable_reg_15_inst : DFF_X1 port map( D => n19535, CK => CLK, Q => 
                           n4195, QN => n18351);
   OUT1_reg_14_inst : DFF_X1 port map( D => n5919, CK => CLK, Q => n4196, QN =>
                           n_1049);
   OUT1_tri_enable_reg_14_inst : DFF_X1 port map( D => n19534, CK => CLK, Q => 
                           n4197, QN => n18352);
   OUT1_reg_13_inst : DFF_X1 port map( D => n5917, CK => CLK, Q => n4198, QN =>
                           n_1050);
   OUT1_tri_enable_reg_13_inst : DFF_X1 port map( D => n19533, CK => CLK, Q => 
                           n4199, QN => n18353);
   OUT1_reg_12_inst : DFF_X1 port map( D => n5915, CK => CLK, Q => n4200, QN =>
                           n_1051);
   OUT1_tri_enable_reg_12_inst : DFF_X1 port map( D => n19532, CK => CLK, Q => 
                           n4201, QN => n18354);
   OUT1_reg_11_inst : DFF_X1 port map( D => n5913, CK => CLK, Q => n4202, QN =>
                           n_1052);
   OUT1_tri_enable_reg_11_inst : DFF_X1 port map( D => n19531, CK => CLK, Q => 
                           n4203, QN => n18355);
   OUT1_reg_10_inst : DFF_X1 port map( D => n5911, CK => CLK, Q => n4204, QN =>
                           n_1053);
   OUT1_tri_enable_reg_10_inst : DFF_X1 port map( D => n19530, CK => CLK, Q => 
                           n4205, QN => n18356);
   OUT1_reg_9_inst : DFF_X1 port map( D => n5909, CK => CLK, Q => n4206, QN => 
                           n_1054);
   OUT1_tri_enable_reg_9_inst : DFF_X1 port map( D => n19529, CK => CLK, Q => 
                           n4207, QN => n18357);
   OUT1_reg_8_inst : DFF_X1 port map( D => n5907, CK => CLK, Q => n4208, QN => 
                           n_1055);
   OUT1_tri_enable_reg_8_inst : DFF_X1 port map( D => n19528, CK => CLK, Q => 
                           n4209, QN => n18358);
   OUT1_reg_7_inst : DFF_X1 port map( D => n5905, CK => CLK, Q => n4210, QN => 
                           n_1056);
   OUT1_tri_enable_reg_7_inst : DFF_X1 port map( D => n19527, CK => CLK, Q => 
                           n4211, QN => n18359);
   OUT1_reg_6_inst : DFF_X1 port map( D => n5903, CK => CLK, Q => n4212, QN => 
                           n_1057);
   OUT1_tri_enable_reg_6_inst : DFF_X1 port map( D => n19526, CK => CLK, Q => 
                           n4213, QN => n18360);
   OUT1_reg_5_inst : DFF_X1 port map( D => n5901, CK => CLK, Q => n4214, QN => 
                           n_1058);
   OUT1_tri_enable_reg_5_inst : DFF_X1 port map( D => n19525, CK => CLK, Q => 
                           n4215, QN => n18361);
   OUT1_reg_4_inst : DFF_X1 port map( D => n5899, CK => CLK, Q => n4216, QN => 
                           n_1059);
   OUT1_tri_enable_reg_4_inst : DFF_X1 port map( D => n19524, CK => CLK, Q => 
                           n4217, QN => n18362);
   OUT1_reg_3_inst : DFF_X1 port map( D => n5897, CK => CLK, Q => n4218, QN => 
                           n_1060);
   OUT1_tri_enable_reg_3_inst : DFF_X1 port map( D => n19523, CK => CLK, Q => 
                           n4219, QN => n18363);
   OUT1_reg_2_inst : DFF_X1 port map( D => n5895, CK => CLK, Q => n4220, QN => 
                           n_1061);
   OUT1_tri_enable_reg_2_inst : DFF_X1 port map( D => n19522, CK => CLK, Q => 
                           n4221, QN => n18364);
   OUT1_reg_1_inst : DFF_X1 port map( D => n5893, CK => CLK, Q => n4222, QN => 
                           n_1062);
   OUT1_tri_enable_reg_1_inst : DFF_X1 port map( D => n19521, CK => CLK, Q => 
                           n4223, QN => n18365);
   OUT1_reg_0_inst : DFF_X1 port map( D => n5891, CK => CLK, Q => n4224, QN => 
                           n_1063);
   OUT1_tri_enable_reg_0_inst : DFF_X1 port map( D => n19518, CK => CLK, Q => 
                           n4225, QN => n18366);
   OUT2_tri_enable_reg_63_inst : DFF_X1 port map( D => n19517, CK => CLK, Q => 
                           n4227, QN => n18383);
   OUT2_reg_62_inst : DFF_X1 port map( D => n5887, CK => CLK, Q => n4228, QN =>
                           n_1064);
   OUT2_tri_enable_reg_62_inst : DFF_X1 port map( D => n19516, CK => CLK, Q => 
                           n4229, QN => n18400);
   OUT2_reg_61_inst : DFF_X1 port map( D => n5885, CK => CLK, Q => n4230, QN =>
                           n_1065);
   OUT2_tri_enable_reg_61_inst : DFF_X1 port map( D => n19515, CK => CLK, Q => 
                           n4231, QN => n18417);
   OUT2_reg_60_inst : DFF_X1 port map( D => n5883, CK => CLK, Q => n4232, QN =>
                           n_1066);
   OUT2_tri_enable_reg_60_inst : DFF_X1 port map( D => n19514, CK => CLK, Q => 
                           n4233, QN => n18434);
   OUT2_reg_59_inst : DFF_X1 port map( D => n5881, CK => CLK, Q => n4234, QN =>
                           n_1067);
   OUT2_tri_enable_reg_59_inst : DFF_X1 port map( D => n19513, CK => CLK, Q => 
                           n4235, QN => n18451);
   OUT2_reg_58_inst : DFF_X1 port map( D => n5879, CK => CLK, Q => n4236, QN =>
                           n_1068);
   OUT2_tri_enable_reg_58_inst : DFF_X1 port map( D => n19512, CK => CLK, Q => 
                           n4237, QN => n18468);
   OUT2_reg_57_inst : DFF_X1 port map( D => n5877, CK => CLK, Q => n4238, QN =>
                           n_1069);
   OUT2_tri_enable_reg_57_inst : DFF_X1 port map( D => n19511, CK => CLK, Q => 
                           n4239, QN => n18485);
   OUT2_reg_56_inst : DFF_X1 port map( D => n5875, CK => CLK, Q => n4240, QN =>
                           n_1070);
   OUT2_tri_enable_reg_56_inst : DFF_X1 port map( D => n19510, CK => CLK, Q => 
                           n4241, QN => n18502);
   OUT2_reg_55_inst : DFF_X1 port map( D => n5873, CK => CLK, Q => n4242, QN =>
                           n_1071);
   OUT2_tri_enable_reg_55_inst : DFF_X1 port map( D => n19509, CK => CLK, Q => 
                           n4243, QN => n18519);
   OUT2_reg_54_inst : DFF_X1 port map( D => n5871, CK => CLK, Q => n4244, QN =>
                           n_1072);
   OUT2_tri_enable_reg_54_inst : DFF_X1 port map( D => n19508, CK => CLK, Q => 
                           n4245, QN => n18536);
   OUT2_reg_53_inst : DFF_X1 port map( D => n5869, CK => CLK, Q => n4246, QN =>
                           n_1073);
   OUT2_tri_enable_reg_53_inst : DFF_X1 port map( D => n19507, CK => CLK, Q => 
                           n4247, QN => n18553);
   OUT2_reg_52_inst : DFF_X1 port map( D => n5867, CK => CLK, Q => n4248, QN =>
                           n_1074);
   OUT2_tri_enable_reg_52_inst : DFF_X1 port map( D => n19506, CK => CLK, Q => 
                           n4249, QN => n18570);
   OUT2_reg_51_inst : DFF_X1 port map( D => n5865, CK => CLK, Q => n4250, QN =>
                           n_1075);
   OUT2_tri_enable_reg_51_inst : DFF_X1 port map( D => n19505, CK => CLK, Q => 
                           n4251, QN => n18587);
   OUT2_reg_50_inst : DFF_X1 port map( D => n5863, CK => CLK, Q => n4252, QN =>
                           n_1076);
   OUT2_tri_enable_reg_50_inst : DFF_X1 port map( D => n19504, CK => CLK, Q => 
                           n4253, QN => n18604);
   OUT2_reg_49_inst : DFF_X1 port map( D => n5861, CK => CLK, Q => n4254, QN =>
                           n_1077);
   OUT2_tri_enable_reg_49_inst : DFF_X1 port map( D => n19503, CK => CLK, Q => 
                           n4255, QN => n18621);
   OUT2_reg_48_inst : DFF_X1 port map( D => n5859, CK => CLK, Q => n4256, QN =>
                           n_1078);
   OUT2_tri_enable_reg_48_inst : DFF_X1 port map( D => n19502, CK => CLK, Q => 
                           n4257, QN => n18638);
   OUT2_reg_47_inst : DFF_X1 port map( D => n5857, CK => CLK, Q => n4258, QN =>
                           n_1079);
   OUT2_tri_enable_reg_47_inst : DFF_X1 port map( D => n19501, CK => CLK, Q => 
                           n4259, QN => n18655);
   OUT2_reg_46_inst : DFF_X1 port map( D => n5855, CK => CLK, Q => n4260, QN =>
                           n_1080);
   OUT2_tri_enable_reg_46_inst : DFF_X1 port map( D => n19500, CK => CLK, Q => 
                           n4261, QN => n18672);
   OUT2_reg_45_inst : DFF_X1 port map( D => n5853, CK => CLK, Q => n4262, QN =>
                           n_1081);
   OUT2_tri_enable_reg_45_inst : DFF_X1 port map( D => n19499, CK => CLK, Q => 
                           n4263, QN => n18689);
   OUT2_reg_44_inst : DFF_X1 port map( D => n5851, CK => CLK, Q => n4264, QN =>
                           n_1082);
   OUT2_tri_enable_reg_44_inst : DFF_X1 port map( D => n19498, CK => CLK, Q => 
                           n4265, QN => n18706);
   OUT2_reg_43_inst : DFF_X1 port map( D => n5849, CK => CLK, Q => n4266, QN =>
                           n_1083);
   OUT2_tri_enable_reg_43_inst : DFF_X1 port map( D => n19497, CK => CLK, Q => 
                           n4267, QN => n18723);
   OUT2_reg_42_inst : DFF_X1 port map( D => n5847, CK => CLK, Q => n4268, QN =>
                           n_1084);
   OUT2_tri_enable_reg_42_inst : DFF_X1 port map( D => n19496, CK => CLK, Q => 
                           n4269, QN => n18740);
   OUT2_reg_41_inst : DFF_X1 port map( D => n5845, CK => CLK, Q => n4270, QN =>
                           n_1085);
   OUT2_tri_enable_reg_41_inst : DFF_X1 port map( D => n19495, CK => CLK, Q => 
                           n4271, QN => n18757);
   OUT2_reg_40_inst : DFF_X1 port map( D => n5843, CK => CLK, Q => n4272, QN =>
                           n_1086);
   OUT2_tri_enable_reg_40_inst : DFF_X1 port map( D => n19494, CK => CLK, Q => 
                           n4273, QN => n18774);
   OUT2_reg_39_inst : DFF_X1 port map( D => n5841, CK => CLK, Q => n4274, QN =>
                           n_1087);
   OUT2_tri_enable_reg_39_inst : DFF_X1 port map( D => n19493, CK => CLK, Q => 
                           n4275, QN => n18791);
   OUT2_reg_38_inst : DFF_X1 port map( D => n5839, CK => CLK, Q => n4276, QN =>
                           n_1088);
   OUT2_tri_enable_reg_38_inst : DFF_X1 port map( D => n19492, CK => CLK, Q => 
                           n4277, QN => n18808);
   OUT2_reg_37_inst : DFF_X1 port map( D => n5837, CK => CLK, Q => n4278, QN =>
                           n_1089);
   OUT2_tri_enable_reg_37_inst : DFF_X1 port map( D => n19491, CK => CLK, Q => 
                           n4279, QN => n18825);
   OUT2_reg_36_inst : DFF_X1 port map( D => n5835, CK => CLK, Q => n4280, QN =>
                           n_1090);
   OUT2_tri_enable_reg_36_inst : DFF_X1 port map( D => n19490, CK => CLK, Q => 
                           n4281, QN => n18842);
   OUT2_reg_35_inst : DFF_X1 port map( D => n5833, CK => CLK, Q => n4282, QN =>
                           n_1091);
   OUT2_tri_enable_reg_35_inst : DFF_X1 port map( D => n19489, CK => CLK, Q => 
                           n4283, QN => n18859);
   OUT2_reg_34_inst : DFF_X1 port map( D => n5831, CK => CLK, Q => n4284, QN =>
                           n_1092);
   OUT2_tri_enable_reg_34_inst : DFF_X1 port map( D => n19488, CK => CLK, Q => 
                           n4285, QN => n18876);
   OUT2_reg_33_inst : DFF_X1 port map( D => n5829, CK => CLK, Q => n4286, QN =>
                           n_1093);
   OUT2_tri_enable_reg_33_inst : DFF_X1 port map( D => n19487, CK => CLK, Q => 
                           n4287, QN => n18893);
   OUT2_reg_32_inst : DFF_X1 port map( D => n5827, CK => CLK, Q => n4288, QN =>
                           n_1094);
   OUT2_tri_enable_reg_32_inst : DFF_X1 port map( D => n19486, CK => CLK, Q => 
                           n4289, QN => n18910);
   OUT2_reg_31_inst : DFF_X1 port map( D => n5825, CK => CLK, Q => n4290, QN =>
                           n_1095);
   OUT2_tri_enable_reg_31_inst : DFF_X1 port map( D => n19485, CK => CLK, Q => 
                           n4291, QN => n18927);
   OUT2_reg_30_inst : DFF_X1 port map( D => n5823, CK => CLK, Q => n4292, QN =>
                           n_1096);
   OUT2_tri_enable_reg_30_inst : DFF_X1 port map( D => n19484, CK => CLK, Q => 
                           n4293, QN => n18944);
   OUT2_reg_29_inst : DFF_X1 port map( D => n5821, CK => CLK, Q => n4294, QN =>
                           n_1097);
   OUT2_tri_enable_reg_29_inst : DFF_X1 port map( D => n19483, CK => CLK, Q => 
                           n4295, QN => n18961);
   OUT2_reg_28_inst : DFF_X1 port map( D => n5819, CK => CLK, Q => n4296, QN =>
                           n_1098);
   OUT2_tri_enable_reg_28_inst : DFF_X1 port map( D => n19482, CK => CLK, Q => 
                           n4297, QN => n18978);
   OUT2_reg_27_inst : DFF_X1 port map( D => n5817, CK => CLK, Q => n4298, QN =>
                           n_1099);
   OUT2_tri_enable_reg_27_inst : DFF_X1 port map( D => n19481, CK => CLK, Q => 
                           n4299, QN => n18995);
   OUT2_reg_26_inst : DFF_X1 port map( D => n5815, CK => CLK, Q => n4300, QN =>
                           n_1100);
   OUT2_tri_enable_reg_26_inst : DFF_X1 port map( D => n19480, CK => CLK, Q => 
                           n4301, QN => n19012);
   OUT2_reg_25_inst : DFF_X1 port map( D => n5813, CK => CLK, Q => n4302, QN =>
                           n_1101);
   OUT2_tri_enable_reg_25_inst : DFF_X1 port map( D => n19479, CK => CLK, Q => 
                           n4303, QN => n19029);
   OUT2_reg_24_inst : DFF_X1 port map( D => n5811, CK => CLK, Q => n4304, QN =>
                           n_1102);
   OUT2_tri_enable_reg_24_inst : DFF_X1 port map( D => n19478, CK => CLK, Q => 
                           n4305, QN => n19046);
   OUT2_reg_23_inst : DFF_X1 port map( D => n5809, CK => CLK, Q => n4306, QN =>
                           n_1103);
   OUT2_tri_enable_reg_23_inst : DFF_X1 port map( D => n19477, CK => CLK, Q => 
                           n4307, QN => n19063);
   OUT2_reg_22_inst : DFF_X1 port map( D => n5807, CK => CLK, Q => n4308, QN =>
                           n_1104);
   OUT2_tri_enable_reg_22_inst : DFF_X1 port map( D => n19476, CK => CLK, Q => 
                           n4309, QN => n19080);
   OUT2_reg_21_inst : DFF_X1 port map( D => n5805, CK => CLK, Q => n4310, QN =>
                           n_1105);
   OUT2_tri_enable_reg_21_inst : DFF_X1 port map( D => n19475, CK => CLK, Q => 
                           n4311, QN => n19097);
   OUT2_reg_20_inst : DFF_X1 port map( D => n5803, CK => CLK, Q => n4312, QN =>
                           n_1106);
   OUT2_tri_enable_reg_20_inst : DFF_X1 port map( D => n19474, CK => CLK, Q => 
                           n4313, QN => n19114);
   OUT2_reg_19_inst : DFF_X1 port map( D => n5801, CK => CLK, Q => n4314, QN =>
                           n_1107);
   OUT2_tri_enable_reg_19_inst : DFF_X1 port map( D => n19473, CK => CLK, Q => 
                           n4315, QN => n19131);
   OUT2_reg_18_inst : DFF_X1 port map( D => n5799, CK => CLK, Q => n4316, QN =>
                           n_1108);
   OUT2_tri_enable_reg_18_inst : DFF_X1 port map( D => n19472, CK => CLK, Q => 
                           n4317, QN => n19148);
   OUT2_reg_17_inst : DFF_X1 port map( D => n5797, CK => CLK, Q => n4318, QN =>
                           n_1109);
   OUT2_tri_enable_reg_17_inst : DFF_X1 port map( D => n19471, CK => CLK, Q => 
                           n4319, QN => n19165);
   OUT2_reg_16_inst : DFF_X1 port map( D => n5795, CK => CLK, Q => n4320, QN =>
                           n_1110);
   OUT2_tri_enable_reg_16_inst : DFF_X1 port map( D => n19470, CK => CLK, Q => 
                           n4321, QN => n19182);
   OUT2_reg_15_inst : DFF_X1 port map( D => n5793, CK => CLK, Q => n4322, QN =>
                           n_1111);
   OUT2_tri_enable_reg_15_inst : DFF_X1 port map( D => n19469, CK => CLK, Q => 
                           n4323, QN => n19199);
   OUT2_reg_14_inst : DFF_X1 port map( D => n5791, CK => CLK, Q => n4324, QN =>
                           n_1112);
   OUT2_tri_enable_reg_14_inst : DFF_X1 port map( D => n19468, CK => CLK, Q => 
                           n4325, QN => n19216);
   OUT2_reg_13_inst : DFF_X1 port map( D => n5789, CK => CLK, Q => n4326, QN =>
                           n_1113);
   OUT2_tri_enable_reg_13_inst : DFF_X1 port map( D => n19467, CK => CLK, Q => 
                           n4327, QN => n19233);
   OUT2_reg_12_inst : DFF_X1 port map( D => n5787, CK => CLK, Q => n4328, QN =>
                           n_1114);
   OUT2_tri_enable_reg_12_inst : DFF_X1 port map( D => n19466, CK => CLK, Q => 
                           n4329, QN => n19250);
   OUT2_reg_11_inst : DFF_X1 port map( D => n5785, CK => CLK, Q => n4330, QN =>
                           n_1115);
   OUT2_tri_enable_reg_11_inst : DFF_X1 port map( D => n19465, CK => CLK, Q => 
                           n4331, QN => n19267);
   OUT2_reg_10_inst : DFF_X1 port map( D => n5783, CK => CLK, Q => n4332, QN =>
                           n_1116);
   OUT2_tri_enable_reg_10_inst : DFF_X1 port map( D => n19464, CK => CLK, Q => 
                           n4333, QN => n19284);
   OUT2_reg_9_inst : DFF_X1 port map( D => n5781, CK => CLK, Q => n4334, QN => 
                           n_1117);
   OUT2_tri_enable_reg_9_inst : DFF_X1 port map( D => n19463, CK => CLK, Q => 
                           n4335, QN => n19301);
   OUT2_reg_8_inst : DFF_X1 port map( D => n5779, CK => CLK, Q => n4336, QN => 
                           n_1118);
   OUT2_tri_enable_reg_8_inst : DFF_X1 port map( D => n19462, CK => CLK, Q => 
                           n4337, QN => n19318);
   OUT2_reg_7_inst : DFF_X1 port map( D => n5777, CK => CLK, Q => n4338, QN => 
                           n_1119);
   OUT2_tri_enable_reg_7_inst : DFF_X1 port map( D => n19461, CK => CLK, Q => 
                           n4339, QN => n19335);
   OUT2_reg_6_inst : DFF_X1 port map( D => n5775, CK => CLK, Q => n4340, QN => 
                           n_1120);
   OUT2_tri_enable_reg_6_inst : DFF_X1 port map( D => n19460, CK => CLK, Q => 
                           n4341, QN => n19352);
   OUT2_reg_5_inst : DFF_X1 port map( D => n5773, CK => CLK, Q => n4342, QN => 
                           n_1121);
   OUT2_tri_enable_reg_5_inst : DFF_X1 port map( D => n19459, CK => CLK, Q => 
                           n4343, QN => n19369);
   OUT2_reg_4_inst : DFF_X1 port map( D => n5771, CK => CLK, Q => n4344, QN => 
                           n_1122);
   OUT2_tri_enable_reg_4_inst : DFF_X1 port map( D => n19458, CK => CLK, Q => 
                           n4345, QN => n19386);
   OUT2_reg_3_inst : DFF_X1 port map( D => n5769, CK => CLK, Q => n4346, QN => 
                           n_1123);
   OUT2_tri_enable_reg_3_inst : DFF_X1 port map( D => n19457, CK => CLK, Q => 
                           n4347, QN => n19403);
   OUT2_reg_2_inst : DFF_X1 port map( D => n5767, CK => CLK, Q => n4348, QN => 
                           n_1124);
   OUT2_tri_enable_reg_2_inst : DFF_X1 port map( D => n19456, CK => CLK, Q => 
                           n4349, QN => n19420);
   OUT2_reg_1_inst : DFF_X1 port map( D => n5765, CK => CLK, Q => n4350, QN => 
                           n_1125);
   OUT2_tri_enable_reg_1_inst : DFF_X1 port map( D => n19455, CK => CLK, Q => 
                           n4351, QN => n19437);
   OUT2_reg_0_inst : DFF_X1 port map( D => n5763, CK => CLK, Q => n4352, QN => 
                           n_1126);
   OUT2_tri_enable_reg_0_inst : DFF_X1 port map( D => n19580, CK => CLK, Q => 
                           n4353, QN => n19454);
   REGISTERS_reg_20_62_inst : DFF_X1 port map( D => n6784, CK => CLK, Q => 
                           n_1127, QN => n9570);
   REGISTERS_reg_20_61_inst : DFF_X1 port map( D => n6783, CK => CLK, Q => 
                           n_1128, QN => n9571);
   REGISTERS_reg_20_60_inst : DFF_X1 port map( D => n6782, CK => CLK, Q => 
                           n_1129, QN => n9572);
   REGISTERS_reg_20_59_inst : DFF_X1 port map( D => n6781, CK => CLK, Q => 
                           n_1130, QN => n9573);
   REGISTERS_reg_20_58_inst : DFF_X1 port map( D => n6780, CK => CLK, Q => 
                           n_1131, QN => n9574);
   REGISTERS_reg_20_57_inst : DFF_X1 port map( D => n6779, CK => CLK, Q => 
                           n_1132, QN => n9575);
   REGISTERS_reg_20_56_inst : DFF_X1 port map( D => n6778, CK => CLK, Q => 
                           n_1133, QN => n9576);
   REGISTERS_reg_20_55_inst : DFF_X1 port map( D => n6777, CK => CLK, Q => 
                           n_1134, QN => n9577);
   REGISTERS_reg_20_54_inst : DFF_X1 port map( D => n6776, CK => CLK, Q => 
                           n_1135, QN => n9578);
   REGISTERS_reg_20_53_inst : DFF_X1 port map( D => n6775, CK => CLK, Q => 
                           n_1136, QN => n9579);
   REGISTERS_reg_20_52_inst : DFF_X1 port map( D => n6774, CK => CLK, Q => 
                           n_1137, QN => n9580);
   REGISTERS_reg_20_51_inst : DFF_X1 port map( D => n6773, CK => CLK, Q => 
                           n_1138, QN => n9581);
   REGISTERS_reg_20_50_inst : DFF_X1 port map( D => n6772, CK => CLK, Q => 
                           n_1139, QN => n9582);
   REGISTERS_reg_20_49_inst : DFF_X1 port map( D => n6771, CK => CLK, Q => 
                           n_1140, QN => n9583);
   REGISTERS_reg_20_48_inst : DFF_X1 port map( D => n6770, CK => CLK, Q => 
                           n_1141, QN => n9584);
   REGISTERS_reg_20_47_inst : DFF_X1 port map( D => n6769, CK => CLK, Q => 
                           n_1142, QN => n9585);
   REGISTERS_reg_20_46_inst : DFF_X1 port map( D => n6768, CK => CLK, Q => 
                           n_1143, QN => n9586);
   REGISTERS_reg_20_45_inst : DFF_X1 port map( D => n6767, CK => CLK, Q => 
                           n_1144, QN => n9587);
   REGISTERS_reg_20_44_inst : DFF_X1 port map( D => n6766, CK => CLK, Q => 
                           n_1145, QN => n9588);
   REGISTERS_reg_20_43_inst : DFF_X1 port map( D => n6765, CK => CLK, Q => 
                           n_1146, QN => n9589);
   REGISTERS_reg_20_42_inst : DFF_X1 port map( D => n6764, CK => CLK, Q => 
                           n_1147, QN => n9590);
   REGISTERS_reg_20_41_inst : DFF_X1 port map( D => n6763, CK => CLK, Q => 
                           n_1148, QN => n9591);
   REGISTERS_reg_20_40_inst : DFF_X1 port map( D => n6762, CK => CLK, Q => 
                           n_1149, QN => n9592);
   REGISTERS_reg_20_39_inst : DFF_X1 port map( D => n6761, CK => CLK, Q => 
                           n_1150, QN => n9593);
   REGISTERS_reg_20_38_inst : DFF_X1 port map( D => n6760, CK => CLK, Q => 
                           n_1151, QN => n9594);
   REGISTERS_reg_20_37_inst : DFF_X1 port map( D => n6759, CK => CLK, Q => 
                           n_1152, QN => n9595);
   REGISTERS_reg_20_36_inst : DFF_X1 port map( D => n6758, CK => CLK, Q => 
                           n_1153, QN => n9596);
   REGISTERS_reg_20_35_inst : DFF_X1 port map( D => n6757, CK => CLK, Q => 
                           n_1154, QN => n9597);
   REGISTERS_reg_20_34_inst : DFF_X1 port map( D => n6756, CK => CLK, Q => 
                           n_1155, QN => n9598);
   REGISTERS_reg_20_33_inst : DFF_X1 port map( D => n6755, CK => CLK, Q => 
                           n_1156, QN => n9599);
   REGISTERS_reg_20_32_inst : DFF_X1 port map( D => n6754, CK => CLK, Q => 
                           n_1157, QN => n9600);
   REGISTERS_reg_20_31_inst : DFF_X1 port map( D => n6753, CK => CLK, Q => 
                           n_1158, QN => n9601);
   REGISTERS_reg_20_30_inst : DFF_X1 port map( D => n6752, CK => CLK, Q => 
                           n_1159, QN => n9602);
   REGISTERS_reg_20_29_inst : DFF_X1 port map( D => n6751, CK => CLK, Q => 
                           n_1160, QN => n9603);
   REGISTERS_reg_20_28_inst : DFF_X1 port map( D => n6750, CK => CLK, Q => 
                           n_1161, QN => n9604);
   REGISTERS_reg_20_27_inst : DFF_X1 port map( D => n6749, CK => CLK, Q => 
                           n_1162, QN => n9605);
   REGISTERS_reg_20_26_inst : DFF_X1 port map( D => n6748, CK => CLK, Q => 
                           n_1163, QN => n9606);
   REGISTERS_reg_20_25_inst : DFF_X1 port map( D => n6747, CK => CLK, Q => 
                           n_1164, QN => n9607);
   REGISTERS_reg_20_24_inst : DFF_X1 port map( D => n6746, CK => CLK, Q => 
                           n_1165, QN => n9608);
   REGISTERS_reg_20_23_inst : DFF_X1 port map( D => n6745, CK => CLK, Q => 
                           n_1166, QN => n9609);
   REGISTERS_reg_20_22_inst : DFF_X1 port map( D => n6744, CK => CLK, Q => 
                           n_1167, QN => n9610);
   REGISTERS_reg_20_21_inst : DFF_X1 port map( D => n6743, CK => CLK, Q => 
                           n_1168, QN => n9611);
   REGISTERS_reg_20_20_inst : DFF_X1 port map( D => n6742, CK => CLK, Q => 
                           n_1169, QN => n9612);
   REGISTERS_reg_20_19_inst : DFF_X1 port map( D => n6741, CK => CLK, Q => 
                           n_1170, QN => n9613);
   REGISTERS_reg_20_18_inst : DFF_X1 port map( D => n6740, CK => CLK, Q => 
                           n_1171, QN => n9614);
   REGISTERS_reg_20_17_inst : DFF_X1 port map( D => n6739, CK => CLK, Q => 
                           n_1172, QN => n9615);
   REGISTERS_reg_20_16_inst : DFF_X1 port map( D => n6738, CK => CLK, Q => 
                           n_1173, QN => n9616);
   REGISTERS_reg_20_15_inst : DFF_X1 port map( D => n6737, CK => CLK, Q => 
                           n_1174, QN => n9617);
   REGISTERS_reg_20_14_inst : DFF_X1 port map( D => n6736, CK => CLK, Q => 
                           n_1175, QN => n9618);
   REGISTERS_reg_20_13_inst : DFF_X1 port map( D => n6735, CK => CLK, Q => 
                           n_1176, QN => n9619);
   REGISTERS_reg_20_12_inst : DFF_X1 port map( D => n6734, CK => CLK, Q => 
                           n_1177, QN => n9620);
   REGISTERS_reg_20_11_inst : DFF_X1 port map( D => n6733, CK => CLK, Q => 
                           n_1178, QN => n9621);
   REGISTERS_reg_20_10_inst : DFF_X1 port map( D => n6732, CK => CLK, Q => 
                           n_1179, QN => n9622);
   REGISTERS_reg_20_9_inst : DFF_X1 port map( D => n6731, CK => CLK, Q => 
                           n_1180, QN => n9623);
   REGISTERS_reg_20_8_inst : DFF_X1 port map( D => n6730, CK => CLK, Q => 
                           n_1181, QN => n9624);
   REGISTERS_reg_20_7_inst : DFF_X1 port map( D => n6729, CK => CLK, Q => 
                           n_1182, QN => n9625);
   REGISTERS_reg_20_6_inst : DFF_X1 port map( D => n6728, CK => CLK, Q => 
                           n_1183, QN => n9626);
   REGISTERS_reg_20_5_inst : DFF_X1 port map( D => n6727, CK => CLK, Q => 
                           n_1184, QN => n9627);
   REGISTERS_reg_20_4_inst : DFF_X1 port map( D => n6726, CK => CLK, Q => 
                           n_1185, QN => n9628);
   REGISTERS_reg_20_3_inst : DFF_X1 port map( D => n6725, CK => CLK, Q => 
                           n_1186, QN => n9629);
   REGISTERS_reg_20_2_inst : DFF_X1 port map( D => n6724, CK => CLK, Q => 
                           n_1187, QN => n9630);
   REGISTERS_reg_20_1_inst : DFF_X1 port map( D => n6723, CK => CLK, Q => 
                           n_1188, QN => n9631);
   REGISTERS_reg_20_0_inst : DFF_X1 port map( D => n6722, CK => CLK, Q => 
                           n_1189, QN => n9632);
   U19260 : NAND3_X1 port map( A1 => ADD_RD1(1), A2 => n20636, A3 => n23966, ZN
                           => n22811);
   U19261 : NAND3_X1 port map( A1 => ADD_RD1(2), A2 => n20637, A3 => n23966, ZN
                           => n22810);
   U19262 : NAND3_X1 port map( A1 => ADD_RD1(2), A2 => ADD_RD1(1), A3 => n23966
                           , ZN => n22815);
   U19263 : NAND3_X1 port map( A1 => ADD_RD2(1), A2 => n20641, A3 => n25165, ZN
                           => n24010);
   U19264 : NAND3_X1 port map( A1 => ADD_RD2(2), A2 => n20642, A3 => n25165, ZN
                           => n24009);
   U19265 : NAND3_X1 port map( A1 => ADD_RD2(2), A2 => ADD_RD2(1), A3 => n25165
                           , ZN => n24014);
   OUT2_tri_0_inst : TBUF_X1 port map( A => n4352, EN => n4353, Z => OUT2(0));
   OUT2_tri_1_inst : TBUF_X1 port map( A => n4350, EN => n4351, Z => OUT2(1));
   OUT2_tri_2_inst : TBUF_X1 port map( A => n4348, EN => n4349, Z => OUT2(2));
   OUT2_tri_3_inst : TBUF_X1 port map( A => n4346, EN => n4347, Z => OUT2(3));
   OUT2_tri_4_inst : TBUF_X1 port map( A => n4344, EN => n4345, Z => OUT2(4));
   OUT2_tri_5_inst : TBUF_X1 port map( A => n4342, EN => n4343, Z => OUT2(5));
   OUT2_tri_6_inst : TBUF_X1 port map( A => n4340, EN => n4341, Z => OUT2(6));
   OUT2_tri_7_inst : TBUF_X1 port map( A => n4338, EN => n4339, Z => OUT2(7));
   OUT2_tri_8_inst : TBUF_X1 port map( A => n4336, EN => n4337, Z => OUT2(8));
   OUT2_tri_9_inst : TBUF_X1 port map( A => n4334, EN => n4335, Z => OUT2(9));
   OUT2_tri_10_inst : TBUF_X1 port map( A => n4332, EN => n4333, Z => OUT2(10))
                           ;
   OUT2_tri_11_inst : TBUF_X1 port map( A => n4330, EN => n4331, Z => OUT2(11))
                           ;
   OUT2_tri_12_inst : TBUF_X1 port map( A => n4328, EN => n4329, Z => OUT2(12))
                           ;
   OUT2_tri_13_inst : TBUF_X1 port map( A => n4326, EN => n4327, Z => OUT2(13))
                           ;
   OUT2_tri_14_inst : TBUF_X1 port map( A => n4324, EN => n4325, Z => OUT2(14))
                           ;
   OUT2_tri_15_inst : TBUF_X1 port map( A => n4322, EN => n4323, Z => OUT2(15))
                           ;
   OUT2_tri_16_inst : TBUF_X1 port map( A => n4320, EN => n4321, Z => OUT2(16))
                           ;
   OUT2_tri_17_inst : TBUF_X1 port map( A => n4318, EN => n4319, Z => OUT2(17))
                           ;
   OUT2_tri_18_inst : TBUF_X1 port map( A => n4316, EN => n4317, Z => OUT2(18))
                           ;
   OUT2_tri_19_inst : TBUF_X1 port map( A => n4314, EN => n4315, Z => OUT2(19))
                           ;
   OUT2_tri_20_inst : TBUF_X1 port map( A => n4312, EN => n4313, Z => OUT2(20))
                           ;
   OUT2_tri_21_inst : TBUF_X1 port map( A => n4310, EN => n4311, Z => OUT2(21))
                           ;
   OUT2_tri_22_inst : TBUF_X1 port map( A => n4308, EN => n4309, Z => OUT2(22))
                           ;
   OUT2_tri_23_inst : TBUF_X1 port map( A => n4306, EN => n4307, Z => OUT2(23))
                           ;
   OUT2_tri_24_inst : TBUF_X1 port map( A => n4304, EN => n4305, Z => OUT2(24))
                           ;
   OUT2_tri_25_inst : TBUF_X1 port map( A => n4302, EN => n4303, Z => OUT2(25))
                           ;
   OUT2_tri_26_inst : TBUF_X1 port map( A => n4300, EN => n4301, Z => OUT2(26))
                           ;
   OUT2_tri_27_inst : TBUF_X1 port map( A => n4298, EN => n4299, Z => OUT2(27))
                           ;
   OUT2_tri_28_inst : TBUF_X1 port map( A => n4296, EN => n4297, Z => OUT2(28))
                           ;
   OUT2_tri_29_inst : TBUF_X1 port map( A => n4294, EN => n4295, Z => OUT2(29))
                           ;
   OUT2_tri_30_inst : TBUF_X1 port map( A => n4292, EN => n4293, Z => OUT2(30))
                           ;
   OUT2_tri_31_inst : TBUF_X1 port map( A => n4290, EN => n4291, Z => OUT2(31))
                           ;
   OUT2_tri_32_inst : TBUF_X1 port map( A => n4288, EN => n4289, Z => OUT2(32))
                           ;
   OUT2_tri_33_inst : TBUF_X1 port map( A => n4286, EN => n4287, Z => OUT2(33))
                           ;
   OUT2_tri_34_inst : TBUF_X1 port map( A => n4284, EN => n4285, Z => OUT2(34))
                           ;
   OUT2_tri_35_inst : TBUF_X1 port map( A => n4282, EN => n4283, Z => OUT2(35))
                           ;
   OUT2_tri_36_inst : TBUF_X1 port map( A => n4280, EN => n4281, Z => OUT2(36))
                           ;
   OUT2_tri_37_inst : TBUF_X1 port map( A => n4278, EN => n4279, Z => OUT2(37))
                           ;
   OUT2_tri_38_inst : TBUF_X1 port map( A => n4276, EN => n4277, Z => OUT2(38))
                           ;
   OUT2_tri_39_inst : TBUF_X1 port map( A => n4274, EN => n4275, Z => OUT2(39))
                           ;
   OUT2_tri_40_inst : TBUF_X1 port map( A => n4272, EN => n4273, Z => OUT2(40))
                           ;
   OUT2_tri_41_inst : TBUF_X1 port map( A => n4270, EN => n4271, Z => OUT2(41))
                           ;
   OUT2_tri_42_inst : TBUF_X1 port map( A => n4268, EN => n4269, Z => OUT2(42))
                           ;
   OUT2_tri_43_inst : TBUF_X1 port map( A => n4266, EN => n4267, Z => OUT2(43))
                           ;
   OUT2_tri_44_inst : TBUF_X1 port map( A => n4264, EN => n4265, Z => OUT2(44))
                           ;
   OUT2_tri_45_inst : TBUF_X1 port map( A => n4262, EN => n4263, Z => OUT2(45))
                           ;
   OUT2_tri_46_inst : TBUF_X1 port map( A => n4260, EN => n4261, Z => OUT2(46))
                           ;
   OUT2_tri_47_inst : TBUF_X1 port map( A => n4258, EN => n4259, Z => OUT2(47))
                           ;
   OUT2_tri_48_inst : TBUF_X1 port map( A => n4256, EN => n4257, Z => OUT2(48))
                           ;
   OUT2_tri_49_inst : TBUF_X1 port map( A => n4254, EN => n4255, Z => OUT2(49))
                           ;
   OUT2_tri_50_inst : TBUF_X1 port map( A => n4252, EN => n4253, Z => OUT2(50))
                           ;
   OUT2_tri_51_inst : TBUF_X1 port map( A => n4250, EN => n4251, Z => OUT2(51))
                           ;
   OUT2_tri_52_inst : TBUF_X1 port map( A => n4248, EN => n4249, Z => OUT2(52))
                           ;
   OUT2_tri_53_inst : TBUF_X1 port map( A => n4246, EN => n4247, Z => OUT2(53))
                           ;
   OUT2_tri_54_inst : TBUF_X1 port map( A => n4244, EN => n4245, Z => OUT2(54))
                           ;
   OUT2_tri_55_inst : TBUF_X1 port map( A => n4242, EN => n4243, Z => OUT2(55))
                           ;
   OUT2_tri_56_inst : TBUF_X1 port map( A => n4240, EN => n4241, Z => OUT2(56))
                           ;
   OUT2_tri_57_inst : TBUF_X1 port map( A => n4238, EN => n4239, Z => OUT2(57))
                           ;
   OUT2_tri_58_inst : TBUF_X1 port map( A => n4236, EN => n4237, Z => OUT2(58))
                           ;
   OUT2_tri_59_inst : TBUF_X1 port map( A => n4234, EN => n4235, Z => OUT2(59))
                           ;
   OUT2_tri_60_inst : TBUF_X1 port map( A => n4232, EN => n4233, Z => OUT2(60))
                           ;
   OUT2_tri_61_inst : TBUF_X1 port map( A => n4230, EN => n4231, Z => OUT2(61))
                           ;
   OUT2_tri_62_inst : TBUF_X1 port map( A => n4228, EN => n4229, Z => OUT2(62))
                           ;
   OUT2_tri_63_inst : TBUF_X1 port map( A => n4226, EN => n4227, Z => OUT2(63))
                           ;
   OUT1_tri_0_inst : TBUF_X1 port map( A => n4224, EN => n4225, Z => OUT1(0));
   OUT1_tri_1_inst : TBUF_X1 port map( A => n4222, EN => n4223, Z => OUT1(1));
   OUT1_tri_2_inst : TBUF_X1 port map( A => n4220, EN => n4221, Z => OUT1(2));
   OUT1_tri_3_inst : TBUF_X1 port map( A => n4218, EN => n4219, Z => OUT1(3));
   OUT1_tri_4_inst : TBUF_X1 port map( A => n4216, EN => n4217, Z => OUT1(4));
   OUT1_tri_5_inst : TBUF_X1 port map( A => n4214, EN => n4215, Z => OUT1(5));
   OUT1_tri_6_inst : TBUF_X1 port map( A => n4212, EN => n4213, Z => OUT1(6));
   OUT1_tri_7_inst : TBUF_X1 port map( A => n4210, EN => n4211, Z => OUT1(7));
   OUT1_tri_8_inst : TBUF_X1 port map( A => n4208, EN => n4209, Z => OUT1(8));
   OUT1_tri_9_inst : TBUF_X1 port map( A => n4206, EN => n4207, Z => OUT1(9));
   OUT1_tri_10_inst : TBUF_X1 port map( A => n4204, EN => n4205, Z => OUT1(10))
                           ;
   OUT1_tri_11_inst : TBUF_X1 port map( A => n4202, EN => n4203, Z => OUT1(11))
                           ;
   OUT1_tri_12_inst : TBUF_X1 port map( A => n4200, EN => n4201, Z => OUT1(12))
                           ;
   OUT1_tri_13_inst : TBUF_X1 port map( A => n4198, EN => n4199, Z => OUT1(13))
                           ;
   OUT1_tri_14_inst : TBUF_X1 port map( A => n4196, EN => n4197, Z => OUT1(14))
                           ;
   OUT1_tri_15_inst : TBUF_X1 port map( A => n4194, EN => n4195, Z => OUT1(15))
                           ;
   OUT1_tri_16_inst : TBUF_X1 port map( A => n4192, EN => n4193, Z => OUT1(16))
                           ;
   OUT1_tri_17_inst : TBUF_X1 port map( A => n4190, EN => n4191, Z => OUT1(17))
                           ;
   OUT1_tri_18_inst : TBUF_X1 port map( A => n4188, EN => n4189, Z => OUT1(18))
                           ;
   OUT1_tri_19_inst : TBUF_X1 port map( A => n4186, EN => n4187, Z => OUT1(19))
                           ;
   OUT1_tri_20_inst : TBUF_X1 port map( A => n4184, EN => n4185, Z => OUT1(20))
                           ;
   OUT1_tri_21_inst : TBUF_X1 port map( A => n4182, EN => n4183, Z => OUT1(21))
                           ;
   OUT1_tri_22_inst : TBUF_X1 port map( A => n4180, EN => n4181, Z => OUT1(22))
                           ;
   OUT1_tri_23_inst : TBUF_X1 port map( A => n4178, EN => n4179, Z => OUT1(23))
                           ;
   OUT1_tri_24_inst : TBUF_X1 port map( A => n4176, EN => n4177, Z => OUT1(24))
                           ;
   OUT1_tri_25_inst : TBUF_X1 port map( A => n4174, EN => n4175, Z => OUT1(25))
                           ;
   OUT1_tri_26_inst : TBUF_X1 port map( A => n4172, EN => n4173, Z => OUT1(26))
                           ;
   OUT1_tri_27_inst : TBUF_X1 port map( A => n4170, EN => n4171, Z => OUT1(27))
                           ;
   OUT1_tri_28_inst : TBUF_X1 port map( A => n4168, EN => n4169, Z => OUT1(28))
                           ;
   OUT1_tri_29_inst : TBUF_X1 port map( A => n4166, EN => n4167, Z => OUT1(29))
                           ;
   OUT1_tri_30_inst : TBUF_X1 port map( A => n4164, EN => n4165, Z => OUT1(30))
                           ;
   OUT1_tri_31_inst : TBUF_X1 port map( A => n4162, EN => n4163, Z => OUT1(31))
                           ;
   OUT1_tri_32_inst : TBUF_X1 port map( A => n4160, EN => n4161, Z => OUT1(32))
                           ;
   OUT1_tri_33_inst : TBUF_X1 port map( A => n4158, EN => n4159, Z => OUT1(33))
                           ;
   OUT1_tri_34_inst : TBUF_X1 port map( A => n4156, EN => n4157, Z => OUT1(34))
                           ;
   OUT1_tri_35_inst : TBUF_X1 port map( A => n4154, EN => n4155, Z => OUT1(35))
                           ;
   OUT1_tri_36_inst : TBUF_X1 port map( A => n4152, EN => n4153, Z => OUT1(36))
                           ;
   OUT1_tri_37_inst : TBUF_X1 port map( A => n4150, EN => n4151, Z => OUT1(37))
                           ;
   OUT1_tri_38_inst : TBUF_X1 port map( A => n4148, EN => n4149, Z => OUT1(38))
                           ;
   OUT1_tri_39_inst : TBUF_X1 port map( A => n4146, EN => n4147, Z => OUT1(39))
                           ;
   OUT1_tri_40_inst : TBUF_X1 port map( A => n4144, EN => n4145, Z => OUT1(40))
                           ;
   OUT1_tri_41_inst : TBUF_X1 port map( A => n4142, EN => n4143, Z => OUT1(41))
                           ;
   OUT1_tri_42_inst : TBUF_X1 port map( A => n4140, EN => n4141, Z => OUT1(42))
                           ;
   OUT1_tri_43_inst : TBUF_X1 port map( A => n4138, EN => n4139, Z => OUT1(43))
                           ;
   OUT1_tri_44_inst : TBUF_X1 port map( A => n4136, EN => n4137, Z => OUT1(44))
                           ;
   OUT1_tri_45_inst : TBUF_X1 port map( A => n4134, EN => n4135, Z => OUT1(45))
                           ;
   OUT1_tri_46_inst : TBUF_X1 port map( A => n4132, EN => n4133, Z => OUT1(46))
                           ;
   OUT1_tri_47_inst : TBUF_X1 port map( A => n4130, EN => n4131, Z => OUT1(47))
                           ;
   OUT1_tri_48_inst : TBUF_X1 port map( A => n4128, EN => n4129, Z => OUT1(48))
                           ;
   OUT1_tri_49_inst : TBUF_X1 port map( A => n4126, EN => n4127, Z => OUT1(49))
                           ;
   OUT1_tri_50_inst : TBUF_X1 port map( A => n4124, EN => n4125, Z => OUT1(50))
                           ;
   OUT1_tri_51_inst : TBUF_X1 port map( A => n4122, EN => n4123, Z => OUT1(51))
                           ;
   OUT1_tri_52_inst : TBUF_X1 port map( A => n4120, EN => n4121, Z => OUT1(52))
                           ;
   OUT1_tri_53_inst : TBUF_X1 port map( A => n4118, EN => n4119, Z => OUT1(53))
                           ;
   OUT1_tri_54_inst : TBUF_X1 port map( A => n4116, EN => n4117, Z => OUT1(54))
                           ;
   OUT1_tri_55_inst : TBUF_X1 port map( A => n4114, EN => n4115, Z => OUT1(55))
                           ;
   OUT1_tri_56_inst : TBUF_X1 port map( A => n4112, EN => n4113, Z => OUT1(56))
                           ;
   OUT1_tri_57_inst : TBUF_X1 port map( A => n4110, EN => n4111, Z => OUT1(57))
                           ;
   OUT1_tri_58_inst : TBUF_X1 port map( A => n4108, EN => n4109, Z => OUT1(58))
                           ;
   OUT1_tri_59_inst : TBUF_X1 port map( A => n4106, EN => n4107, Z => OUT1(59))
                           ;
   OUT1_tri_60_inst : TBUF_X1 port map( A => n4104, EN => n4105, Z => OUT1(60))
                           ;
   OUT1_tri_61_inst : TBUF_X1 port map( A => n4102, EN => n4103, Z => OUT1(61))
                           ;
   OUT1_tri_62_inst : TBUF_X1 port map( A => n4100, EN => n4101, Z => OUT1(62))
                           ;
   OUT1_tri_63_inst : TBUF_X1 port map( A => n4098, EN => n4099, Z => OUT1(63))
                           ;
   REGISTERS_reg_21_63_inst : DFF_X1 port map( D => n6721, CK => CLK, Q => 
                           n20963, QN => n9633);
   REGISTERS_reg_21_62_inst : DFF_X1 port map( D => n6720, CK => CLK, Q => 
                           n20964, QN => n9634);
   REGISTERS_reg_21_61_inst : DFF_X1 port map( D => n6719, CK => CLK, Q => 
                           n20965, QN => n9635);
   REGISTERS_reg_21_60_inst : DFF_X1 port map( D => n6718, CK => CLK, Q => 
                           n20966, QN => n9636);
   REGISTERS_reg_15_63_inst : DFF_X1 port map( D => n7105, CK => CLK, Q => 
                           n20967, QN => n9505);
   REGISTERS_reg_15_62_inst : DFF_X1 port map( D => n7104, CK => CLK, Q => 
                           n20968, QN => n9506);
   REGISTERS_reg_15_61_inst : DFF_X1 port map( D => n7103, CK => CLK, Q => 
                           n20969, QN => n9507);
   REGISTERS_reg_15_60_inst : DFF_X1 port map( D => n7102, CK => CLK, Q => 
                           n20970, QN => n9508);
   REGISTERS_reg_13_63_inst : DFF_X1 port map( D => n7233, CK => CLK, Q => 
                           n20971, QN => n9697);
   REGISTERS_reg_13_62_inst : DFF_X1 port map( D => n7232, CK => CLK, Q => 
                           n20972, QN => n9698);
   REGISTERS_reg_13_61_inst : DFF_X1 port map( D => n7231, CK => CLK, Q => 
                           n20973, QN => n9699);
   REGISTERS_reg_13_60_inst : DFF_X1 port map( D => n7230, CK => CLK, Q => 
                           n20974, QN => n9700);
   REGISTERS_reg_21_59_inst : DFF_X1 port map( D => n6717, CK => CLK, Q => 
                           n20975, QN => n9637);
   REGISTERS_reg_21_58_inst : DFF_X1 port map( D => n6716, CK => CLK, Q => 
                           n20976, QN => n9638);
   REGISTERS_reg_21_57_inst : DFF_X1 port map( D => n6715, CK => CLK, Q => 
                           n20977, QN => n9639);
   REGISTERS_reg_21_56_inst : DFF_X1 port map( D => n6714, CK => CLK, Q => 
                           n20978, QN => n9640);
   REGISTERS_reg_21_55_inst : DFF_X1 port map( D => n6713, CK => CLK, Q => 
                           n20979, QN => n9641);
   REGISTERS_reg_21_54_inst : DFF_X1 port map( D => n6712, CK => CLK, Q => 
                           n20980, QN => n9642);
   REGISTERS_reg_21_53_inst : DFF_X1 port map( D => n6711, CK => CLK, Q => 
                           n20981, QN => n9643);
   REGISTERS_reg_21_52_inst : DFF_X1 port map( D => n6710, CK => CLK, Q => 
                           n20982, QN => n9644);
   REGISTERS_reg_21_51_inst : DFF_X1 port map( D => n6709, CK => CLK, Q => 
                           n20983, QN => n9645);
   REGISTERS_reg_21_50_inst : DFF_X1 port map( D => n6708, CK => CLK, Q => 
                           n20984, QN => n9646);
   REGISTERS_reg_21_49_inst : DFF_X1 port map( D => n6707, CK => CLK, Q => 
                           n20985, QN => n9647);
   REGISTERS_reg_21_48_inst : DFF_X1 port map( D => n6706, CK => CLK, Q => 
                           n20986, QN => n9648);
   REGISTERS_reg_21_47_inst : DFF_X1 port map( D => n6705, CK => CLK, Q => 
                           n20987, QN => n9649);
   REGISTERS_reg_21_46_inst : DFF_X1 port map( D => n6704, CK => CLK, Q => 
                           n20988, QN => n9650);
   REGISTERS_reg_21_45_inst : DFF_X1 port map( D => n6703, CK => CLK, Q => 
                           n20989, QN => n9651);
   REGISTERS_reg_21_44_inst : DFF_X1 port map( D => n6702, CK => CLK, Q => 
                           n20990, QN => n9652);
   REGISTERS_reg_21_43_inst : DFF_X1 port map( D => n6701, CK => CLK, Q => 
                           n20991, QN => n9653);
   REGISTERS_reg_21_42_inst : DFF_X1 port map( D => n6700, CK => CLK, Q => 
                           n20992, QN => n9654);
   REGISTERS_reg_21_41_inst : DFF_X1 port map( D => n6699, CK => CLK, Q => 
                           n20993, QN => n9655);
   REGISTERS_reg_21_40_inst : DFF_X1 port map( D => n6698, CK => CLK, Q => 
                           n20994, QN => n9656);
   REGISTERS_reg_21_39_inst : DFF_X1 port map( D => n6697, CK => CLK, Q => 
                           n20995, QN => n9657);
   REGISTERS_reg_21_38_inst : DFF_X1 port map( D => n6696, CK => CLK, Q => 
                           n20996, QN => n9658);
   REGISTERS_reg_21_37_inst : DFF_X1 port map( D => n6695, CK => CLK, Q => 
                           n20997, QN => n9659);
   REGISTERS_reg_21_36_inst : DFF_X1 port map( D => n6694, CK => CLK, Q => 
                           n20998, QN => n9660);
   REGISTERS_reg_21_35_inst : DFF_X1 port map( D => n6693, CK => CLK, Q => 
                           n20999, QN => n9661);
   REGISTERS_reg_21_34_inst : DFF_X1 port map( D => n6692, CK => CLK, Q => 
                           n21000, QN => n9662);
   REGISTERS_reg_21_33_inst : DFF_X1 port map( D => n6691, CK => CLK, Q => 
                           n21001, QN => n9663);
   REGISTERS_reg_21_32_inst : DFF_X1 port map( D => n6690, CK => CLK, Q => 
                           n21002, QN => n9664);
   REGISTERS_reg_21_31_inst : DFF_X1 port map( D => n6689, CK => CLK, Q => 
                           n21003, QN => n9665);
   REGISTERS_reg_21_30_inst : DFF_X1 port map( D => n6688, CK => CLK, Q => 
                           n21004, QN => n9666);
   REGISTERS_reg_21_29_inst : DFF_X1 port map( D => n6687, CK => CLK, Q => 
                           n21005, QN => n9667);
   REGISTERS_reg_21_28_inst : DFF_X1 port map( D => n6686, CK => CLK, Q => 
                           n21006, QN => n9668);
   REGISTERS_reg_21_27_inst : DFF_X1 port map( D => n6685, CK => CLK, Q => 
                           n21007, QN => n9669);
   REGISTERS_reg_21_26_inst : DFF_X1 port map( D => n6684, CK => CLK, Q => 
                           n21008, QN => n9670);
   REGISTERS_reg_21_25_inst : DFF_X1 port map( D => n6683, CK => CLK, Q => 
                           n21009, QN => n9671);
   REGISTERS_reg_21_24_inst : DFF_X1 port map( D => n6682, CK => CLK, Q => 
                           n21010, QN => n9672);
   REGISTERS_reg_21_23_inst : DFF_X1 port map( D => n6681, CK => CLK, Q => 
                           n21011, QN => n9673);
   REGISTERS_reg_21_22_inst : DFF_X1 port map( D => n6680, CK => CLK, Q => 
                           n21012, QN => n9674);
   REGISTERS_reg_21_21_inst : DFF_X1 port map( D => n6679, CK => CLK, Q => 
                           n21013, QN => n9675);
   REGISTERS_reg_21_20_inst : DFF_X1 port map( D => n6678, CK => CLK, Q => 
                           n21014, QN => n9676);
   REGISTERS_reg_21_19_inst : DFF_X1 port map( D => n6677, CK => CLK, Q => 
                           n21015, QN => n9677);
   REGISTERS_reg_21_18_inst : DFF_X1 port map( D => n6676, CK => CLK, Q => 
                           n21016, QN => n9678);
   REGISTERS_reg_21_17_inst : DFF_X1 port map( D => n6675, CK => CLK, Q => 
                           n21017, QN => n9679);
   REGISTERS_reg_21_16_inst : DFF_X1 port map( D => n6674, CK => CLK, Q => 
                           n21018, QN => n9680);
   REGISTERS_reg_21_15_inst : DFF_X1 port map( D => n6673, CK => CLK, Q => 
                           n21019, QN => n9681);
   REGISTERS_reg_21_14_inst : DFF_X1 port map( D => n6672, CK => CLK, Q => 
                           n21020, QN => n9682);
   REGISTERS_reg_21_13_inst : DFF_X1 port map( D => n6671, CK => CLK, Q => 
                           n21021, QN => n9683);
   REGISTERS_reg_21_12_inst : DFF_X1 port map( D => n6670, CK => CLK, Q => 
                           n21022, QN => n9684);
   REGISTERS_reg_21_11_inst : DFF_X1 port map( D => n6669, CK => CLK, Q => 
                           n21023, QN => n9685);
   REGISTERS_reg_21_10_inst : DFF_X1 port map( D => n6668, CK => CLK, Q => 
                           n21024, QN => n9686);
   REGISTERS_reg_21_9_inst : DFF_X1 port map( D => n6667, CK => CLK, Q => 
                           n21025, QN => n9687);
   REGISTERS_reg_21_8_inst : DFF_X1 port map( D => n6666, CK => CLK, Q => 
                           n21026, QN => n9688);
   REGISTERS_reg_21_7_inst : DFF_X1 port map( D => n6665, CK => CLK, Q => 
                           n21027, QN => n9689);
   REGISTERS_reg_21_6_inst : DFF_X1 port map( D => n6664, CK => CLK, Q => 
                           n21028, QN => n9690);
   REGISTERS_reg_21_5_inst : DFF_X1 port map( D => n6663, CK => CLK, Q => 
                           n21029, QN => n9691);
   REGISTERS_reg_21_4_inst : DFF_X1 port map( D => n6662, CK => CLK, Q => 
                           n21030, QN => n9692);
   REGISTERS_reg_21_3_inst : DFF_X1 port map( D => n6661, CK => CLK, Q => 
                           n21031, QN => n9693);
   REGISTERS_reg_21_2_inst : DFF_X1 port map( D => n6660, CK => CLK, Q => 
                           n21032, QN => n9694);
   REGISTERS_reg_21_1_inst : DFF_X1 port map( D => n6659, CK => CLK, Q => 
                           n21033, QN => n9695);
   REGISTERS_reg_21_0_inst : DFF_X1 port map( D => n6658, CK => CLK, Q => 
                           n21034, QN => n9696);
   REGISTERS_reg_15_59_inst : DFF_X1 port map( D => n7101, CK => CLK, Q => 
                           n21035, QN => n9509);
   REGISTERS_reg_15_58_inst : DFF_X1 port map( D => n7100, CK => CLK, Q => 
                           n21036, QN => n9510);
   REGISTERS_reg_15_57_inst : DFF_X1 port map( D => n7099, CK => CLK, Q => 
                           n21037, QN => n9511);
   REGISTERS_reg_15_56_inst : DFF_X1 port map( D => n7098, CK => CLK, Q => 
                           n21038, QN => n9512);
   REGISTERS_reg_15_55_inst : DFF_X1 port map( D => n7097, CK => CLK, Q => 
                           n21039, QN => n9513);
   REGISTERS_reg_15_54_inst : DFF_X1 port map( D => n7096, CK => CLK, Q => 
                           n21040, QN => n9514);
   REGISTERS_reg_15_53_inst : DFF_X1 port map( D => n7095, CK => CLK, Q => 
                           n21041, QN => n9515);
   REGISTERS_reg_15_52_inst : DFF_X1 port map( D => n7094, CK => CLK, Q => 
                           n21042, QN => n9516);
   REGISTERS_reg_15_51_inst : DFF_X1 port map( D => n7093, CK => CLK, Q => 
                           n21043, QN => n9517);
   REGISTERS_reg_15_50_inst : DFF_X1 port map( D => n7092, CK => CLK, Q => 
                           n21044, QN => n9518);
   REGISTERS_reg_15_49_inst : DFF_X1 port map( D => n7091, CK => CLK, Q => 
                           n21045, QN => n9519);
   REGISTERS_reg_15_48_inst : DFF_X1 port map( D => n7090, CK => CLK, Q => 
                           n21046, QN => n9520);
   REGISTERS_reg_15_47_inst : DFF_X1 port map( D => n7089, CK => CLK, Q => 
                           n21047, QN => n9521);
   REGISTERS_reg_15_46_inst : DFF_X1 port map( D => n7088, CK => CLK, Q => 
                           n21048, QN => n9522);
   REGISTERS_reg_15_45_inst : DFF_X1 port map( D => n7087, CK => CLK, Q => 
                           n21049, QN => n9523);
   REGISTERS_reg_15_44_inst : DFF_X1 port map( D => n7086, CK => CLK, Q => 
                           n21050, QN => n9524);
   REGISTERS_reg_15_43_inst : DFF_X1 port map( D => n7085, CK => CLK, Q => 
                           n21051, QN => n9525);
   REGISTERS_reg_15_42_inst : DFF_X1 port map( D => n7084, CK => CLK, Q => 
                           n21052, QN => n9526);
   REGISTERS_reg_15_41_inst : DFF_X1 port map( D => n7083, CK => CLK, Q => 
                           n21053, QN => n9527);
   REGISTERS_reg_15_40_inst : DFF_X1 port map( D => n7082, CK => CLK, Q => 
                           n21054, QN => n9528);
   REGISTERS_reg_15_39_inst : DFF_X1 port map( D => n7081, CK => CLK, Q => 
                           n21055, QN => n9529);
   REGISTERS_reg_15_38_inst : DFF_X1 port map( D => n7080, CK => CLK, Q => 
                           n21056, QN => n9530);
   REGISTERS_reg_15_37_inst : DFF_X1 port map( D => n7079, CK => CLK, Q => 
                           n21057, QN => n9531);
   REGISTERS_reg_15_36_inst : DFF_X1 port map( D => n7078, CK => CLK, Q => 
                           n21058, QN => n9532);
   REGISTERS_reg_15_35_inst : DFF_X1 port map( D => n7077, CK => CLK, Q => 
                           n21059, QN => n9533);
   REGISTERS_reg_15_34_inst : DFF_X1 port map( D => n7076, CK => CLK, Q => 
                           n21060, QN => n9534);
   REGISTERS_reg_15_33_inst : DFF_X1 port map( D => n7075, CK => CLK, Q => 
                           n21061, QN => n9535);
   REGISTERS_reg_15_32_inst : DFF_X1 port map( D => n7074, CK => CLK, Q => 
                           n21062, QN => n9536);
   REGISTERS_reg_15_31_inst : DFF_X1 port map( D => n7073, CK => CLK, Q => 
                           n21063, QN => n9537);
   REGISTERS_reg_15_30_inst : DFF_X1 port map( D => n7072, CK => CLK, Q => 
                           n21064, QN => n9538);
   REGISTERS_reg_15_29_inst : DFF_X1 port map( D => n7071, CK => CLK, Q => 
                           n21065, QN => n9539);
   REGISTERS_reg_15_28_inst : DFF_X1 port map( D => n7070, CK => CLK, Q => 
                           n21066, QN => n9540);
   REGISTERS_reg_15_27_inst : DFF_X1 port map( D => n7069, CK => CLK, Q => 
                           n21067, QN => n9541);
   REGISTERS_reg_15_26_inst : DFF_X1 port map( D => n7068, CK => CLK, Q => 
                           n21068, QN => n9542);
   REGISTERS_reg_15_25_inst : DFF_X1 port map( D => n7067, CK => CLK, Q => 
                           n21069, QN => n9543);
   REGISTERS_reg_15_24_inst : DFF_X1 port map( D => n7066, CK => CLK, Q => 
                           n21070, QN => n9544);
   REGISTERS_reg_15_23_inst : DFF_X1 port map( D => n7065, CK => CLK, Q => 
                           n21071, QN => n9545);
   REGISTERS_reg_15_22_inst : DFF_X1 port map( D => n7064, CK => CLK, Q => 
                           n21072, QN => n9546);
   REGISTERS_reg_15_21_inst : DFF_X1 port map( D => n7063, CK => CLK, Q => 
                           n21073, QN => n9547);
   REGISTERS_reg_15_20_inst : DFF_X1 port map( D => n7062, CK => CLK, Q => 
                           n21074, QN => n9548);
   REGISTERS_reg_15_19_inst : DFF_X1 port map( D => n7061, CK => CLK, Q => 
                           n21075, QN => n9549);
   REGISTERS_reg_15_18_inst : DFF_X1 port map( D => n7060, CK => CLK, Q => 
                           n21076, QN => n9550);
   REGISTERS_reg_15_17_inst : DFF_X1 port map( D => n7059, CK => CLK, Q => 
                           n21077, QN => n9551);
   REGISTERS_reg_15_16_inst : DFF_X1 port map( D => n7058, CK => CLK, Q => 
                           n21078, QN => n9552);
   REGISTERS_reg_15_15_inst : DFF_X1 port map( D => n7057, CK => CLK, Q => 
                           n21079, QN => n9553);
   REGISTERS_reg_15_14_inst : DFF_X1 port map( D => n7056, CK => CLK, Q => 
                           n21080, QN => n9554);
   REGISTERS_reg_15_13_inst : DFF_X1 port map( D => n7055, CK => CLK, Q => 
                           n21081, QN => n9555);
   REGISTERS_reg_15_12_inst : DFF_X1 port map( D => n7054, CK => CLK, Q => 
                           n21082, QN => n9556);
   REGISTERS_reg_15_11_inst : DFF_X1 port map( D => n7053, CK => CLK, Q => 
                           n21083, QN => n9557);
   REGISTERS_reg_15_10_inst : DFF_X1 port map( D => n7052, CK => CLK, Q => 
                           n21084, QN => n9558);
   REGISTERS_reg_15_9_inst : DFF_X1 port map( D => n7051, CK => CLK, Q => 
                           n21085, QN => n9559);
   REGISTERS_reg_15_8_inst : DFF_X1 port map( D => n7050, CK => CLK, Q => 
                           n21086, QN => n9560);
   REGISTERS_reg_15_7_inst : DFF_X1 port map( D => n7049, CK => CLK, Q => 
                           n21087, QN => n9561);
   REGISTERS_reg_15_6_inst : DFF_X1 port map( D => n7048, CK => CLK, Q => 
                           n21088, QN => n9562);
   REGISTERS_reg_15_5_inst : DFF_X1 port map( D => n7047, CK => CLK, Q => 
                           n21089, QN => n9563);
   REGISTERS_reg_15_4_inst : DFF_X1 port map( D => n7046, CK => CLK, Q => 
                           n21090, QN => n9564);
   REGISTERS_reg_15_3_inst : DFF_X1 port map( D => n7045, CK => CLK, Q => 
                           n21091, QN => n9565);
   REGISTERS_reg_15_2_inst : DFF_X1 port map( D => n7044, CK => CLK, Q => 
                           n21092, QN => n9566);
   REGISTERS_reg_15_1_inst : DFF_X1 port map( D => n7043, CK => CLK, Q => 
                           n21093, QN => n9567);
   REGISTERS_reg_15_0_inst : DFF_X1 port map( D => n7042, CK => CLK, Q => 
                           n21094, QN => n9568);
   REGISTERS_reg_13_59_inst : DFF_X1 port map( D => n7229, CK => CLK, Q => 
                           n21095, QN => n9701);
   REGISTERS_reg_13_58_inst : DFF_X1 port map( D => n7228, CK => CLK, Q => 
                           n21096, QN => n9702);
   REGISTERS_reg_13_57_inst : DFF_X1 port map( D => n7227, CK => CLK, Q => 
                           n21097, QN => n9703);
   REGISTERS_reg_13_56_inst : DFF_X1 port map( D => n7226, CK => CLK, Q => 
                           n21098, QN => n9704);
   REGISTERS_reg_13_55_inst : DFF_X1 port map( D => n7225, CK => CLK, Q => 
                           n21099, QN => n9705);
   REGISTERS_reg_13_54_inst : DFF_X1 port map( D => n7224, CK => CLK, Q => 
                           n21100, QN => n9706);
   REGISTERS_reg_13_53_inst : DFF_X1 port map( D => n7223, CK => CLK, Q => 
                           n21101, QN => n9707);
   REGISTERS_reg_13_52_inst : DFF_X1 port map( D => n7222, CK => CLK, Q => 
                           n21102, QN => n9708);
   REGISTERS_reg_13_51_inst : DFF_X1 port map( D => n7221, CK => CLK, Q => 
                           n21103, QN => n9709);
   REGISTERS_reg_13_50_inst : DFF_X1 port map( D => n7220, CK => CLK, Q => 
                           n21104, QN => n9710);
   REGISTERS_reg_13_49_inst : DFF_X1 port map( D => n7219, CK => CLK, Q => 
                           n21105, QN => n9711);
   REGISTERS_reg_13_48_inst : DFF_X1 port map( D => n7218, CK => CLK, Q => 
                           n21106, QN => n9712);
   REGISTERS_reg_13_47_inst : DFF_X1 port map( D => n7217, CK => CLK, Q => 
                           n21107, QN => n9713);
   REGISTERS_reg_13_46_inst : DFF_X1 port map( D => n7216, CK => CLK, Q => 
                           n21108, QN => n9714);
   REGISTERS_reg_13_45_inst : DFF_X1 port map( D => n7215, CK => CLK, Q => 
                           n21109, QN => n9715);
   REGISTERS_reg_13_44_inst : DFF_X1 port map( D => n7214, CK => CLK, Q => 
                           n21110, QN => n9716);
   REGISTERS_reg_13_43_inst : DFF_X1 port map( D => n7213, CK => CLK, Q => 
                           n21111, QN => n9717);
   REGISTERS_reg_13_42_inst : DFF_X1 port map( D => n7212, CK => CLK, Q => 
                           n21112, QN => n9718);
   REGISTERS_reg_13_41_inst : DFF_X1 port map( D => n7211, CK => CLK, Q => 
                           n21113, QN => n9719);
   REGISTERS_reg_13_40_inst : DFF_X1 port map( D => n7210, CK => CLK, Q => 
                           n21114, QN => n9720);
   REGISTERS_reg_13_39_inst : DFF_X1 port map( D => n7209, CK => CLK, Q => 
                           n21115, QN => n9721);
   REGISTERS_reg_13_38_inst : DFF_X1 port map( D => n7208, CK => CLK, Q => 
                           n21116, QN => n9722);
   REGISTERS_reg_13_37_inst : DFF_X1 port map( D => n7207, CK => CLK, Q => 
                           n21117, QN => n9723);
   REGISTERS_reg_13_36_inst : DFF_X1 port map( D => n7206, CK => CLK, Q => 
                           n21118, QN => n9724);
   REGISTERS_reg_13_35_inst : DFF_X1 port map( D => n7205, CK => CLK, Q => 
                           n21119, QN => n9725);
   REGISTERS_reg_13_34_inst : DFF_X1 port map( D => n7204, CK => CLK, Q => 
                           n21120, QN => n9726);
   REGISTERS_reg_13_33_inst : DFF_X1 port map( D => n7203, CK => CLK, Q => 
                           n21121, QN => n9727);
   REGISTERS_reg_13_32_inst : DFF_X1 port map( D => n7202, CK => CLK, Q => 
                           n21122, QN => n9728);
   REGISTERS_reg_13_31_inst : DFF_X1 port map( D => n7201, CK => CLK, Q => 
                           n21123, QN => n9729);
   REGISTERS_reg_13_30_inst : DFF_X1 port map( D => n7200, CK => CLK, Q => 
                           n21124, QN => n9730);
   REGISTERS_reg_13_29_inst : DFF_X1 port map( D => n7199, CK => CLK, Q => 
                           n21125, QN => n9731);
   REGISTERS_reg_13_28_inst : DFF_X1 port map( D => n7198, CK => CLK, Q => 
                           n21126, QN => n9732);
   REGISTERS_reg_13_27_inst : DFF_X1 port map( D => n7197, CK => CLK, Q => 
                           n21127, QN => n9733);
   REGISTERS_reg_13_26_inst : DFF_X1 port map( D => n7196, CK => CLK, Q => 
                           n21128, QN => n9734);
   REGISTERS_reg_13_25_inst : DFF_X1 port map( D => n7195, CK => CLK, Q => 
                           n21129, QN => n9735);
   REGISTERS_reg_13_24_inst : DFF_X1 port map( D => n7194, CK => CLK, Q => 
                           n21130, QN => n9736);
   REGISTERS_reg_13_23_inst : DFF_X1 port map( D => n7193, CK => CLK, Q => 
                           n21131, QN => n9737);
   REGISTERS_reg_13_22_inst : DFF_X1 port map( D => n7192, CK => CLK, Q => 
                           n21132, QN => n9738);
   REGISTERS_reg_13_21_inst : DFF_X1 port map( D => n7191, CK => CLK, Q => 
                           n21133, QN => n9739);
   REGISTERS_reg_13_20_inst : DFF_X1 port map( D => n7190, CK => CLK, Q => 
                           n21134, QN => n9740);
   REGISTERS_reg_13_19_inst : DFF_X1 port map( D => n7189, CK => CLK, Q => 
                           n21135, QN => n9741);
   REGISTERS_reg_13_18_inst : DFF_X1 port map( D => n7188, CK => CLK, Q => 
                           n21136, QN => n9742);
   REGISTERS_reg_13_17_inst : DFF_X1 port map( D => n7187, CK => CLK, Q => 
                           n21137, QN => n9743);
   REGISTERS_reg_13_16_inst : DFF_X1 port map( D => n7186, CK => CLK, Q => 
                           n21138, QN => n9744);
   REGISTERS_reg_13_15_inst : DFF_X1 port map( D => n7185, CK => CLK, Q => 
                           n21139, QN => n9745);
   REGISTERS_reg_13_14_inst : DFF_X1 port map( D => n7184, CK => CLK, Q => 
                           n21140, QN => n9746);
   REGISTERS_reg_13_13_inst : DFF_X1 port map( D => n7183, CK => CLK, Q => 
                           n21141, QN => n9747);
   REGISTERS_reg_13_12_inst : DFF_X1 port map( D => n7182, CK => CLK, Q => 
                           n21142, QN => n9748);
   REGISTERS_reg_13_11_inst : DFF_X1 port map( D => n7181, CK => CLK, Q => 
                           n21143, QN => n9749);
   REGISTERS_reg_13_10_inst : DFF_X1 port map( D => n7180, CK => CLK, Q => 
                           n21144, QN => n9750);
   REGISTERS_reg_13_9_inst : DFF_X1 port map( D => n7179, CK => CLK, Q => 
                           n21145, QN => n9751);
   REGISTERS_reg_13_8_inst : DFF_X1 port map( D => n7178, CK => CLK, Q => 
                           n21146, QN => n9752);
   REGISTERS_reg_13_7_inst : DFF_X1 port map( D => n7177, CK => CLK, Q => 
                           n21147, QN => n9753);
   REGISTERS_reg_13_6_inst : DFF_X1 port map( D => n7176, CK => CLK, Q => 
                           n21148, QN => n9754);
   REGISTERS_reg_13_5_inst : DFF_X1 port map( D => n7175, CK => CLK, Q => 
                           n21149, QN => n9755);
   REGISTERS_reg_13_4_inst : DFF_X1 port map( D => n7174, CK => CLK, Q => 
                           n21150, QN => n9756);
   REGISTERS_reg_13_3_inst : DFF_X1 port map( D => n7173, CK => CLK, Q => 
                           n21151, QN => n9757);
   REGISTERS_reg_13_2_inst : DFF_X1 port map( D => n7172, CK => CLK, Q => 
                           n21152, QN => n9758);
   REGISTERS_reg_13_1_inst : DFF_X1 port map( D => n7171, CK => CLK, Q => 
                           n21153, QN => n9759);
   REGISTERS_reg_13_0_inst : DFF_X1 port map( D => n7170, CK => CLK, Q => 
                           n21154, QN => n9760);
   REGISTERS_reg_20_63_inst : DFF_X1 port map( D => n6785, CK => CLK, Q => 
                           n_1190, QN => n9569);
   REGISTERS_reg_26_63_inst : DFF_X1 port map( D => n6401, CK => CLK, Q => 
                           n_1191, QN => n21480);
   REGISTERS_reg_26_62_inst : DFF_X1 port map( D => n6400, CK => CLK, Q => 
                           n_1192, QN => n21481);
   REGISTERS_reg_26_61_inst : DFF_X1 port map( D => n6399, CK => CLK, Q => 
                           n_1193, QN => n21482);
   REGISTERS_reg_26_60_inst : DFF_X1 port map( D => n6398, CK => CLK, Q => 
                           n_1194, QN => n21483);
   REGISTERS_reg_25_63_inst : DFF_X1 port map( D => n6465, CK => CLK, Q => 
                           n_1195, QN => n21156);
   REGISTERS_reg_25_62_inst : DFF_X1 port map( D => n6464, CK => CLK, Q => 
                           n_1196, QN => n21157);
   REGISTERS_reg_25_61_inst : DFF_X1 port map( D => n6463, CK => CLK, Q => 
                           n_1197, QN => n21158);
   REGISTERS_reg_25_60_inst : DFF_X1 port map( D => n6462, CK => CLK, Q => 
                           n_1198, QN => n21159);
   REGISTERS_reg_19_63_inst : DFF_X1 port map( D => n6849, CK => CLK, Q => 
                           n_1199, QN => n22248);
   REGISTERS_reg_19_62_inst : DFF_X1 port map( D => n6848, CK => CLK, Q => 
                           n_1200, QN => n22249);
   REGISTERS_reg_19_61_inst : DFF_X1 port map( D => n6847, CK => CLK, Q => 
                           n_1201, QN => n22250);
   REGISTERS_reg_19_60_inst : DFF_X1 port map( D => n6846, CK => CLK, Q => 
                           n_1202, QN => n22251);
   REGISTERS_reg_14_63_inst : DFF_X1 port map( D => n7169, CK => CLK, Q => 
                           n_1203, QN => n21155);
   REGISTERS_reg_14_62_inst : DFF_X1 port map( D => n7168, CK => CLK, Q => 
                           n_1204, QN => n20772);
   REGISTERS_reg_14_61_inst : DFF_X1 port map( D => n7167, CK => CLK, Q => 
                           n_1205, QN => n20773);
   REGISTERS_reg_14_60_inst : DFF_X1 port map( D => n7166, CK => CLK, Q => 
                           n_1206, QN => n20774);
   REGISTERS_reg_11_63_inst : DFF_X1 port map( D => n7361, CK => CLK, Q => 
                           n_1207, QN => n21504);
   REGISTERS_reg_11_62_inst : DFF_X1 port map( D => n7360, CK => CLK, Q => 
                           n_1208, QN => n21505);
   REGISTERS_reg_11_61_inst : DFF_X1 port map( D => n7359, CK => CLK, Q => 
                           n_1209, QN => n21506);
   REGISTERS_reg_11_60_inst : DFF_X1 port map( D => n7358, CK => CLK, Q => 
                           n_1210, QN => n21507);
   REGISTERS_reg_8_63_inst : DFF_X1 port map( D => n7553, CK => CLK, Q => 
                           n_1211, QN => n22256);
   REGISTERS_reg_8_62_inst : DFF_X1 port map( D => n7552, CK => CLK, Q => 
                           n_1212, QN => n22257);
   REGISTERS_reg_8_61_inst : DFF_X1 port map( D => n7551, CK => CLK, Q => 
                           n_1213, QN => n22258);
   REGISTERS_reg_8_60_inst : DFF_X1 port map( D => n7550, CK => CLK, Q => 
                           n_1214, QN => n22259);
   REGISTERS_reg_3_63_inst : DFF_X1 port map( D => n7873, CK => CLK, Q => 
                           n_1215, QN => n21168);
   REGISTERS_reg_3_62_inst : DFF_X1 port map( D => n7872, CK => CLK, Q => 
                           n_1216, QN => n21169);
   REGISTERS_reg_3_61_inst : DFF_X1 port map( D => n7871, CK => CLK, Q => 
                           n_1217, QN => n21170);
   REGISTERS_reg_3_60_inst : DFF_X1 port map( D => n7870, CK => CLK, Q => 
                           n_1218, QN => n21171);
   REGISTERS_reg_26_59_inst : DFF_X1 port map( D => n6397, CK => CLK, Q => 
                           n_1219, QN => n21580);
   REGISTERS_reg_26_58_inst : DFF_X1 port map( D => n6396, CK => CLK, Q => 
                           n_1220, QN => n21581);
   REGISTERS_reg_26_57_inst : DFF_X1 port map( D => n6395, CK => CLK, Q => 
                           n_1221, QN => n21582);
   REGISTERS_reg_26_56_inst : DFF_X1 port map( D => n6394, CK => CLK, Q => 
                           n_1222, QN => n21583);
   REGISTERS_reg_26_55_inst : DFF_X1 port map( D => n6393, CK => CLK, Q => 
                           n_1223, QN => n21584);
   REGISTERS_reg_26_54_inst : DFF_X1 port map( D => n6392, CK => CLK, Q => 
                           n_1224, QN => n21585);
   REGISTERS_reg_26_53_inst : DFF_X1 port map( D => n6391, CK => CLK, Q => 
                           n_1225, QN => n21586);
   REGISTERS_reg_26_52_inst : DFF_X1 port map( D => n6390, CK => CLK, Q => 
                           n_1226, QN => n21587);
   REGISTERS_reg_26_51_inst : DFF_X1 port map( D => n6389, CK => CLK, Q => 
                           n_1227, QN => n21588);
   REGISTERS_reg_26_50_inst : DFF_X1 port map( D => n6388, CK => CLK, Q => 
                           n_1228, QN => n21589);
   REGISTERS_reg_26_49_inst : DFF_X1 port map( D => n6387, CK => CLK, Q => 
                           n_1229, QN => n21590);
   REGISTERS_reg_26_48_inst : DFF_X1 port map( D => n6386, CK => CLK, Q => 
                           n_1230, QN => n21591);
   REGISTERS_reg_26_47_inst : DFF_X1 port map( D => n6385, CK => CLK, Q => 
                           n_1231, QN => n21592);
   REGISTERS_reg_26_46_inst : DFF_X1 port map( D => n6384, CK => CLK, Q => 
                           n_1232, QN => n21593);
   REGISTERS_reg_26_45_inst : DFF_X1 port map( D => n6383, CK => CLK, Q => 
                           n_1233, QN => n21594);
   REGISTERS_reg_26_44_inst : DFF_X1 port map( D => n6382, CK => CLK, Q => 
                           n_1234, QN => n21595);
   REGISTERS_reg_26_43_inst : DFF_X1 port map( D => n6381, CK => CLK, Q => 
                           n_1235, QN => n21596);
   REGISTERS_reg_26_42_inst : DFF_X1 port map( D => n6380, CK => CLK, Q => 
                           n_1236, QN => n21597);
   REGISTERS_reg_26_41_inst : DFF_X1 port map( D => n6379, CK => CLK, Q => 
                           n_1237, QN => n21598);
   REGISTERS_reg_26_40_inst : DFF_X1 port map( D => n6378, CK => CLK, Q => 
                           n_1238, QN => n21599);
   REGISTERS_reg_26_39_inst : DFF_X1 port map( D => n6377, CK => CLK, Q => 
                           n_1239, QN => n21600);
   REGISTERS_reg_26_38_inst : DFF_X1 port map( D => n6376, CK => CLK, Q => 
                           n_1240, QN => n21601);
   REGISTERS_reg_26_37_inst : DFF_X1 port map( D => n6375, CK => CLK, Q => 
                           n_1241, QN => n21602);
   REGISTERS_reg_26_36_inst : DFF_X1 port map( D => n6374, CK => CLK, Q => 
                           n_1242, QN => n21603);
   REGISTERS_reg_26_35_inst : DFF_X1 port map( D => n6373, CK => CLK, Q => 
                           n_1243, QN => n21604);
   REGISTERS_reg_26_34_inst : DFF_X1 port map( D => n6372, CK => CLK, Q => 
                           n_1244, QN => n21605);
   REGISTERS_reg_26_33_inst : DFF_X1 port map( D => n6371, CK => CLK, Q => 
                           n_1245, QN => n21606);
   REGISTERS_reg_26_32_inst : DFF_X1 port map( D => n6370, CK => CLK, Q => 
                           n_1246, QN => n21607);
   REGISTERS_reg_26_31_inst : DFF_X1 port map( D => n6369, CK => CLK, Q => 
                           n_1247, QN => n21608);
   REGISTERS_reg_26_30_inst : DFF_X1 port map( D => n6368, CK => CLK, Q => 
                           n_1248, QN => n21609);
   REGISTERS_reg_26_29_inst : DFF_X1 port map( D => n6367, CK => CLK, Q => 
                           n_1249, QN => n21610);
   REGISTERS_reg_26_28_inst : DFF_X1 port map( D => n6366, CK => CLK, Q => 
                           n_1250, QN => n21611);
   REGISTERS_reg_26_27_inst : DFF_X1 port map( D => n6365, CK => CLK, Q => 
                           n_1251, QN => n21612);
   REGISTERS_reg_26_26_inst : DFF_X1 port map( D => n6364, CK => CLK, Q => 
                           n_1252, QN => n21613);
   REGISTERS_reg_26_25_inst : DFF_X1 port map( D => n6363, CK => CLK, Q => 
                           n_1253, QN => n21614);
   REGISTERS_reg_26_24_inst : DFF_X1 port map( D => n6362, CK => CLK, Q => 
                           n_1254, QN => n21615);
   REGISTERS_reg_26_23_inst : DFF_X1 port map( D => n6361, CK => CLK, Q => 
                           n_1255, QN => n21616);
   REGISTERS_reg_26_22_inst : DFF_X1 port map( D => n6360, CK => CLK, Q => 
                           n_1256, QN => n21617);
   REGISTERS_reg_26_21_inst : DFF_X1 port map( D => n6359, CK => CLK, Q => 
                           n_1257, QN => n21618);
   REGISTERS_reg_26_20_inst : DFF_X1 port map( D => n6358, CK => CLK, Q => 
                           n_1258, QN => n21619);
   REGISTERS_reg_26_19_inst : DFF_X1 port map( D => n6357, CK => CLK, Q => 
                           n_1259, QN => n21620);
   REGISTERS_reg_26_18_inst : DFF_X1 port map( D => n6356, CK => CLK, Q => 
                           n_1260, QN => n21621);
   REGISTERS_reg_26_17_inst : DFF_X1 port map( D => n6355, CK => CLK, Q => 
                           n_1261, QN => n21622);
   REGISTERS_reg_26_16_inst : DFF_X1 port map( D => n6354, CK => CLK, Q => 
                           n_1262, QN => n21623);
   REGISTERS_reg_26_15_inst : DFF_X1 port map( D => n6353, CK => CLK, Q => 
                           n_1263, QN => n21624);
   REGISTERS_reg_26_14_inst : DFF_X1 port map( D => n6352, CK => CLK, Q => 
                           n_1264, QN => n21625);
   REGISTERS_reg_26_13_inst : DFF_X1 port map( D => n6351, CK => CLK, Q => 
                           n_1265, QN => n21626);
   REGISTERS_reg_26_12_inst : DFF_X1 port map( D => n6350, CK => CLK, Q => 
                           n_1266, QN => n21627);
   REGISTERS_reg_26_11_inst : DFF_X1 port map( D => n6349, CK => CLK, Q => 
                           n_1267, QN => n21628);
   REGISTERS_reg_26_10_inst : DFF_X1 port map( D => n6348, CK => CLK, Q => 
                           n_1268, QN => n21629);
   REGISTERS_reg_26_9_inst : DFF_X1 port map( D => n6347, CK => CLK, Q => 
                           n_1269, QN => n21630);
   REGISTERS_reg_26_8_inst : DFF_X1 port map( D => n6346, CK => CLK, Q => 
                           n_1270, QN => n21631);
   REGISTERS_reg_26_7_inst : DFF_X1 port map( D => n6345, CK => CLK, Q => 
                           n_1271, QN => n21632);
   REGISTERS_reg_26_6_inst : DFF_X1 port map( D => n6344, CK => CLK, Q => 
                           n_1272, QN => n21633);
   REGISTERS_reg_26_5_inst : DFF_X1 port map( D => n6343, CK => CLK, Q => 
                           n_1273, QN => n21634);
   REGISTERS_reg_26_4_inst : DFF_X1 port map( D => n6342, CK => CLK, Q => 
                           n_1274, QN => n21635);
   REGISTERS_reg_26_3_inst : DFF_X1 port map( D => n6341, CK => CLK, Q => 
                           n_1275, QN => n21636);
   REGISTERS_reg_26_2_inst : DFF_X1 port map( D => n6340, CK => CLK, Q => 
                           n_1276, QN => n21637);
   REGISTERS_reg_26_1_inst : DFF_X1 port map( D => n6339, CK => CLK, Q => 
                           n_1277, QN => n21638);
   REGISTERS_reg_26_0_inst : DFF_X1 port map( D => n6338, CK => CLK, Q => 
                           n_1278, QN => n21639);
   REGISTERS_reg_25_59_inst : DFF_X1 port map( D => n6461, CK => CLK, Q => 
                           n_1279, QN => n21180);
   REGISTERS_reg_25_58_inst : DFF_X1 port map( D => n6460, CK => CLK, Q => 
                           n_1280, QN => n21181);
   REGISTERS_reg_25_57_inst : DFF_X1 port map( D => n6459, CK => CLK, Q => 
                           n_1281, QN => n21182);
   REGISTERS_reg_25_56_inst : DFF_X1 port map( D => n6458, CK => CLK, Q => 
                           n_1282, QN => n21183);
   REGISTERS_reg_25_55_inst : DFF_X1 port map( D => n6457, CK => CLK, Q => 
                           n_1283, QN => n21184);
   REGISTERS_reg_25_54_inst : DFF_X1 port map( D => n6456, CK => CLK, Q => 
                           n_1284, QN => n21185);
   REGISTERS_reg_25_53_inst : DFF_X1 port map( D => n6455, CK => CLK, Q => 
                           n_1285, QN => n21186);
   REGISTERS_reg_25_52_inst : DFF_X1 port map( D => n6454, CK => CLK, Q => 
                           n_1286, QN => n21187);
   REGISTERS_reg_25_51_inst : DFF_X1 port map( D => n6453, CK => CLK, Q => 
                           n_1287, QN => n21188);
   REGISTERS_reg_25_50_inst : DFF_X1 port map( D => n6452, CK => CLK, Q => 
                           n_1288, QN => n21189);
   REGISTERS_reg_25_49_inst : DFF_X1 port map( D => n6451, CK => CLK, Q => 
                           n_1289, QN => n21190);
   REGISTERS_reg_25_48_inst : DFF_X1 port map( D => n6450, CK => CLK, Q => 
                           n_1290, QN => n21191);
   REGISTERS_reg_25_47_inst : DFF_X1 port map( D => n6449, CK => CLK, Q => 
                           n_1291, QN => n21192);
   REGISTERS_reg_25_46_inst : DFF_X1 port map( D => n6448, CK => CLK, Q => 
                           n_1292, QN => n21193);
   REGISTERS_reg_25_45_inst : DFF_X1 port map( D => n6447, CK => CLK, Q => 
                           n_1293, QN => n21194);
   REGISTERS_reg_25_44_inst : DFF_X1 port map( D => n6446, CK => CLK, Q => 
                           n_1294, QN => n21195);
   REGISTERS_reg_25_43_inst : DFF_X1 port map( D => n6445, CK => CLK, Q => 
                           n_1295, QN => n21196);
   REGISTERS_reg_25_42_inst : DFF_X1 port map( D => n6444, CK => CLK, Q => 
                           n_1296, QN => n21197);
   REGISTERS_reg_25_41_inst : DFF_X1 port map( D => n6443, CK => CLK, Q => 
                           n_1297, QN => n21198);
   REGISTERS_reg_25_40_inst : DFF_X1 port map( D => n6442, CK => CLK, Q => 
                           n_1298, QN => n21199);
   REGISTERS_reg_25_39_inst : DFF_X1 port map( D => n6441, CK => CLK, Q => 
                           n_1299, QN => n21200);
   REGISTERS_reg_25_38_inst : DFF_X1 port map( D => n6440, CK => CLK, Q => 
                           n_1300, QN => n21201);
   REGISTERS_reg_25_37_inst : DFF_X1 port map( D => n6439, CK => CLK, Q => 
                           n_1301, QN => n21202);
   REGISTERS_reg_25_36_inst : DFF_X1 port map( D => n6438, CK => CLK, Q => 
                           n_1302, QN => n21203);
   REGISTERS_reg_25_35_inst : DFF_X1 port map( D => n6437, CK => CLK, Q => 
                           n_1303, QN => n21204);
   REGISTERS_reg_25_34_inst : DFF_X1 port map( D => n6436, CK => CLK, Q => 
                           n_1304, QN => n21205);
   REGISTERS_reg_25_33_inst : DFF_X1 port map( D => n6435, CK => CLK, Q => 
                           n_1305, QN => n21206);
   REGISTERS_reg_25_32_inst : DFF_X1 port map( D => n6434, CK => CLK, Q => 
                           n_1306, QN => n21207);
   REGISTERS_reg_25_31_inst : DFF_X1 port map( D => n6433, CK => CLK, Q => 
                           n_1307, QN => n21208);
   REGISTERS_reg_25_30_inst : DFF_X1 port map( D => n6432, CK => CLK, Q => 
                           n_1308, QN => n21209);
   REGISTERS_reg_25_29_inst : DFF_X1 port map( D => n6431, CK => CLK, Q => 
                           n_1309, QN => n21210);
   REGISTERS_reg_25_28_inst : DFF_X1 port map( D => n6430, CK => CLK, Q => 
                           n_1310, QN => n21211);
   REGISTERS_reg_25_27_inst : DFF_X1 port map( D => n6429, CK => CLK, Q => 
                           n_1311, QN => n21212);
   REGISTERS_reg_25_26_inst : DFF_X1 port map( D => n6428, CK => CLK, Q => 
                           n_1312, QN => n21213);
   REGISTERS_reg_25_25_inst : DFF_X1 port map( D => n6427, CK => CLK, Q => 
                           n_1313, QN => n21214);
   REGISTERS_reg_25_24_inst : DFF_X1 port map( D => n6426, CK => CLK, Q => 
                           n_1314, QN => n21215);
   REGISTERS_reg_25_23_inst : DFF_X1 port map( D => n6425, CK => CLK, Q => 
                           n_1315, QN => n21216);
   REGISTERS_reg_25_22_inst : DFF_X1 port map( D => n6424, CK => CLK, Q => 
                           n_1316, QN => n21217);
   REGISTERS_reg_25_21_inst : DFF_X1 port map( D => n6423, CK => CLK, Q => 
                           n_1317, QN => n21218);
   REGISTERS_reg_25_20_inst : DFF_X1 port map( D => n6422, CK => CLK, Q => 
                           n_1318, QN => n21219);
   REGISTERS_reg_25_19_inst : DFF_X1 port map( D => n6421, CK => CLK, Q => 
                           n_1319, QN => n21220);
   REGISTERS_reg_25_18_inst : DFF_X1 port map( D => n6420, CK => CLK, Q => 
                           n_1320, QN => n21221);
   REGISTERS_reg_25_17_inst : DFF_X1 port map( D => n6419, CK => CLK, Q => 
                           n_1321, QN => n21222);
   REGISTERS_reg_25_16_inst : DFF_X1 port map( D => n6418, CK => CLK, Q => 
                           n_1322, QN => n21223);
   REGISTERS_reg_25_15_inst : DFF_X1 port map( D => n6417, CK => CLK, Q => 
                           n_1323, QN => n21224);
   REGISTERS_reg_25_14_inst : DFF_X1 port map( D => n6416, CK => CLK, Q => 
                           n_1324, QN => n21225);
   REGISTERS_reg_25_13_inst : DFF_X1 port map( D => n6415, CK => CLK, Q => 
                           n_1325, QN => n21226);
   REGISTERS_reg_25_12_inst : DFF_X1 port map( D => n6414, CK => CLK, Q => 
                           n_1326, QN => n21227);
   REGISTERS_reg_25_11_inst : DFF_X1 port map( D => n6413, CK => CLK, Q => 
                           n_1327, QN => n21228);
   REGISTERS_reg_25_10_inst : DFF_X1 port map( D => n6412, CK => CLK, Q => 
                           n_1328, QN => n21229);
   REGISTERS_reg_25_9_inst : DFF_X1 port map( D => n6411, CK => CLK, Q => 
                           n_1329, QN => n21230);
   REGISTERS_reg_25_8_inst : DFF_X1 port map( D => n6410, CK => CLK, Q => 
                           n_1330, QN => n21231);
   REGISTERS_reg_25_7_inst : DFF_X1 port map( D => n6409, CK => CLK, Q => 
                           n_1331, QN => n21232);
   REGISTERS_reg_25_6_inst : DFF_X1 port map( D => n6408, CK => CLK, Q => 
                           n_1332, QN => n21233);
   REGISTERS_reg_25_5_inst : DFF_X1 port map( D => n6407, CK => CLK, Q => 
                           n_1333, QN => n21234);
   REGISTERS_reg_25_4_inst : DFF_X1 port map( D => n6406, CK => CLK, Q => 
                           n_1334, QN => n21235);
   REGISTERS_reg_25_3_inst : DFF_X1 port map( D => n6405, CK => CLK, Q => 
                           n_1335, QN => n21236);
   REGISTERS_reg_25_2_inst : DFF_X1 port map( D => n6404, CK => CLK, Q => 
                           n_1336, QN => n21237);
   REGISTERS_reg_25_1_inst : DFF_X1 port map( D => n6403, CK => CLK, Q => 
                           n_1337, QN => n21238);
   REGISTERS_reg_25_0_inst : DFF_X1 port map( D => n6402, CK => CLK, Q => 
                           n_1338, QN => n21239);
   REGISTERS_reg_19_59_inst : DFF_X1 port map( D => n6845, CK => CLK, Q => 
                           n_1339, QN => n22320);
   REGISTERS_reg_19_58_inst : DFF_X1 port map( D => n6844, CK => CLK, Q => 
                           n_1340, QN => n22321);
   REGISTERS_reg_19_57_inst : DFF_X1 port map( D => n6843, CK => CLK, Q => 
                           n_1341, QN => n22322);
   REGISTERS_reg_19_56_inst : DFF_X1 port map( D => n6842, CK => CLK, Q => 
                           n_1342, QN => n22323);
   REGISTERS_reg_19_55_inst : DFF_X1 port map( D => n6841, CK => CLK, Q => 
                           n_1343, QN => n22324);
   REGISTERS_reg_19_54_inst : DFF_X1 port map( D => n6840, CK => CLK, Q => 
                           n_1344, QN => n22325);
   REGISTERS_reg_19_53_inst : DFF_X1 port map( D => n6839, CK => CLK, Q => 
                           n_1345, QN => n22326);
   REGISTERS_reg_19_52_inst : DFF_X1 port map( D => n6838, CK => CLK, Q => 
                           n_1346, QN => n22327);
   REGISTERS_reg_19_51_inst : DFF_X1 port map( D => n6837, CK => CLK, Q => 
                           n_1347, QN => n22328);
   REGISTERS_reg_19_50_inst : DFF_X1 port map( D => n6836, CK => CLK, Q => 
                           n_1348, QN => n22329);
   REGISTERS_reg_19_49_inst : DFF_X1 port map( D => n6835, CK => CLK, Q => 
                           n_1349, QN => n22330);
   REGISTERS_reg_19_48_inst : DFF_X1 port map( D => n6834, CK => CLK, Q => 
                           n_1350, QN => n22331);
   REGISTERS_reg_19_47_inst : DFF_X1 port map( D => n6833, CK => CLK, Q => 
                           n_1351, QN => n22332);
   REGISTERS_reg_19_46_inst : DFF_X1 port map( D => n6832, CK => CLK, Q => 
                           n_1352, QN => n22333);
   REGISTERS_reg_19_45_inst : DFF_X1 port map( D => n6831, CK => CLK, Q => 
                           n_1353, QN => n22334);
   REGISTERS_reg_19_44_inst : DFF_X1 port map( D => n6830, CK => CLK, Q => 
                           n_1354, QN => n22335);
   REGISTERS_reg_19_43_inst : DFF_X1 port map( D => n6829, CK => CLK, Q => 
                           n_1355, QN => n22336);
   REGISTERS_reg_19_42_inst : DFF_X1 port map( D => n6828, CK => CLK, Q => 
                           n_1356, QN => n22337);
   REGISTERS_reg_19_41_inst : DFF_X1 port map( D => n6827, CK => CLK, Q => 
                           n_1357, QN => n22338);
   REGISTERS_reg_19_40_inst : DFF_X1 port map( D => n6826, CK => CLK, Q => 
                           n_1358, QN => n22339);
   REGISTERS_reg_19_39_inst : DFF_X1 port map( D => n6825, CK => CLK, Q => 
                           n_1359, QN => n22340);
   REGISTERS_reg_19_38_inst : DFF_X1 port map( D => n6824, CK => CLK, Q => 
                           n_1360, QN => n22341);
   REGISTERS_reg_19_37_inst : DFF_X1 port map( D => n6823, CK => CLK, Q => 
                           n_1361, QN => n22342);
   REGISTERS_reg_19_36_inst : DFF_X1 port map( D => n6822, CK => CLK, Q => 
                           n_1362, QN => n22343);
   REGISTERS_reg_19_35_inst : DFF_X1 port map( D => n6821, CK => CLK, Q => 
                           n_1363, QN => n22344);
   REGISTERS_reg_19_34_inst : DFF_X1 port map( D => n6820, CK => CLK, Q => 
                           n_1364, QN => n22345);
   REGISTERS_reg_19_33_inst : DFF_X1 port map( D => n6819, CK => CLK, Q => 
                           n_1365, QN => n22346);
   REGISTERS_reg_19_32_inst : DFF_X1 port map( D => n6818, CK => CLK, Q => 
                           n_1366, QN => n22347);
   REGISTERS_reg_19_31_inst : DFF_X1 port map( D => n6817, CK => CLK, Q => 
                           n_1367, QN => n22348);
   REGISTERS_reg_19_30_inst : DFF_X1 port map( D => n6816, CK => CLK, Q => 
                           n_1368, QN => n22349);
   REGISTERS_reg_19_29_inst : DFF_X1 port map( D => n6815, CK => CLK, Q => 
                           n_1369, QN => n22350);
   REGISTERS_reg_19_28_inst : DFF_X1 port map( D => n6814, CK => CLK, Q => 
                           n_1370, QN => n22351);
   REGISTERS_reg_19_27_inst : DFF_X1 port map( D => n6813, CK => CLK, Q => 
                           n_1371, QN => n22352);
   REGISTERS_reg_19_26_inst : DFF_X1 port map( D => n6812, CK => CLK, Q => 
                           n_1372, QN => n22353);
   REGISTERS_reg_19_25_inst : DFF_X1 port map( D => n6811, CK => CLK, Q => 
                           n_1373, QN => n22354);
   REGISTERS_reg_19_24_inst : DFF_X1 port map( D => n6810, CK => CLK, Q => 
                           n_1374, QN => n22355);
   REGISTERS_reg_19_23_inst : DFF_X1 port map( D => n6809, CK => CLK, Q => 
                           n_1375, QN => n22356);
   REGISTERS_reg_19_22_inst : DFF_X1 port map( D => n6808, CK => CLK, Q => 
                           n_1376, QN => n22357);
   REGISTERS_reg_19_21_inst : DFF_X1 port map( D => n6807, CK => CLK, Q => 
                           n_1377, QN => n22358);
   REGISTERS_reg_19_20_inst : DFF_X1 port map( D => n6806, CK => CLK, Q => 
                           n_1378, QN => n22359);
   REGISTERS_reg_19_19_inst : DFF_X1 port map( D => n6805, CK => CLK, Q => 
                           n_1379, QN => n22360);
   REGISTERS_reg_19_18_inst : DFF_X1 port map( D => n6804, CK => CLK, Q => 
                           n_1380, QN => n22361);
   REGISTERS_reg_19_17_inst : DFF_X1 port map( D => n6803, CK => CLK, Q => 
                           n_1381, QN => n22362);
   REGISTERS_reg_19_16_inst : DFF_X1 port map( D => n6802, CK => CLK, Q => 
                           n_1382, QN => n22363);
   REGISTERS_reg_19_15_inst : DFF_X1 port map( D => n6801, CK => CLK, Q => 
                           n_1383, QN => n22364);
   REGISTERS_reg_19_14_inst : DFF_X1 port map( D => n6800, CK => CLK, Q => 
                           n_1384, QN => n22365);
   REGISTERS_reg_19_13_inst : DFF_X1 port map( D => n6799, CK => CLK, Q => 
                           n_1385, QN => n22366);
   REGISTERS_reg_19_12_inst : DFF_X1 port map( D => n6798, CK => CLK, Q => 
                           n_1386, QN => n22367);
   REGISTERS_reg_19_11_inst : DFF_X1 port map( D => n6797, CK => CLK, Q => 
                           n_1387, QN => n22368);
   REGISTERS_reg_19_10_inst : DFF_X1 port map( D => n6796, CK => CLK, Q => 
                           n_1388, QN => n22369);
   REGISTERS_reg_19_9_inst : DFF_X1 port map( D => n6795, CK => CLK, Q => 
                           n_1389, QN => n22370);
   REGISTERS_reg_19_8_inst : DFF_X1 port map( D => n6794, CK => CLK, Q => 
                           n_1390, QN => n22371);
   REGISTERS_reg_19_7_inst : DFF_X1 port map( D => n6793, CK => CLK, Q => 
                           n_1391, QN => n22372);
   REGISTERS_reg_19_6_inst : DFF_X1 port map( D => n6792, CK => CLK, Q => 
                           n_1392, QN => n22373);
   REGISTERS_reg_19_5_inst : DFF_X1 port map( D => n6791, CK => CLK, Q => 
                           n_1393, QN => n22374);
   REGISTERS_reg_19_4_inst : DFF_X1 port map( D => n6790, CK => CLK, Q => 
                           n_1394, QN => n22375);
   REGISTERS_reg_19_3_inst : DFF_X1 port map( D => n6789, CK => CLK, Q => 
                           n_1395, QN => n22376);
   REGISTERS_reg_19_2_inst : DFF_X1 port map( D => n6788, CK => CLK, Q => 
                           n_1396, QN => n22377);
   REGISTERS_reg_19_1_inst : DFF_X1 port map( D => n6787, CK => CLK, Q => 
                           n_1397, QN => n22378);
   REGISTERS_reg_19_0_inst : DFF_X1 port map( D => n6786, CK => CLK, Q => 
                           n_1398, QN => n22379);
   REGISTERS_reg_14_59_inst : DFF_X1 port map( D => n7165, CK => CLK, Q => 
                           n_1399, QN => n20775);
   REGISTERS_reg_14_58_inst : DFF_X1 port map( D => n7164, CK => CLK, Q => 
                           n_1400, QN => n20776);
   REGISTERS_reg_14_57_inst : DFF_X1 port map( D => n7163, CK => CLK, Q => 
                           n_1401, QN => n20777);
   REGISTERS_reg_14_56_inst : DFF_X1 port map( D => n7162, CK => CLK, Q => 
                           n_1402, QN => n20778);
   REGISTERS_reg_14_55_inst : DFF_X1 port map( D => n7161, CK => CLK, Q => 
                           n_1403, QN => n20779);
   REGISTERS_reg_14_54_inst : DFF_X1 port map( D => n7160, CK => CLK, Q => 
                           n_1404, QN => n20780);
   REGISTERS_reg_14_53_inst : DFF_X1 port map( D => n7159, CK => CLK, Q => 
                           n_1405, QN => n20781);
   REGISTERS_reg_14_52_inst : DFF_X1 port map( D => n7158, CK => CLK, Q => 
                           n_1406, QN => n20782);
   REGISTERS_reg_14_51_inst : DFF_X1 port map( D => n7157, CK => CLK, Q => 
                           n_1407, QN => n20783);
   REGISTERS_reg_14_50_inst : DFF_X1 port map( D => n7156, CK => CLK, Q => 
                           n_1408, QN => n20784);
   REGISTERS_reg_14_49_inst : DFF_X1 port map( D => n7155, CK => CLK, Q => 
                           n_1409, QN => n20785);
   REGISTERS_reg_14_48_inst : DFF_X1 port map( D => n7154, CK => CLK, Q => 
                           n_1410, QN => n20786);
   REGISTERS_reg_14_47_inst : DFF_X1 port map( D => n7153, CK => CLK, Q => 
                           n_1411, QN => n20787);
   REGISTERS_reg_14_46_inst : DFF_X1 port map( D => n7152, CK => CLK, Q => 
                           n_1412, QN => n20788);
   REGISTERS_reg_14_45_inst : DFF_X1 port map( D => n7151, CK => CLK, Q => 
                           n_1413, QN => n20789);
   REGISTERS_reg_14_44_inst : DFF_X1 port map( D => n7150, CK => CLK, Q => 
                           n_1414, QN => n20790);
   REGISTERS_reg_14_43_inst : DFF_X1 port map( D => n7149, CK => CLK, Q => 
                           n_1415, QN => n20791);
   REGISTERS_reg_14_42_inst : DFF_X1 port map( D => n7148, CK => CLK, Q => 
                           n_1416, QN => n20792);
   REGISTERS_reg_14_41_inst : DFF_X1 port map( D => n7147, CK => CLK, Q => 
                           n_1417, QN => n20793);
   REGISTERS_reg_14_40_inst : DFF_X1 port map( D => n7146, CK => CLK, Q => 
                           n_1418, QN => n20794);
   REGISTERS_reg_14_39_inst : DFF_X1 port map( D => n7145, CK => CLK, Q => 
                           n_1419, QN => n20795);
   REGISTERS_reg_14_38_inst : DFF_X1 port map( D => n7144, CK => CLK, Q => 
                           n_1420, QN => n20796);
   REGISTERS_reg_14_37_inst : DFF_X1 port map( D => n7143, CK => CLK, Q => 
                           n_1421, QN => n20797);
   REGISTERS_reg_14_36_inst : DFF_X1 port map( D => n7142, CK => CLK, Q => 
                           n_1422, QN => n20798);
   REGISTERS_reg_14_35_inst : DFF_X1 port map( D => n7141, CK => CLK, Q => 
                           n_1423, QN => n20799);
   REGISTERS_reg_14_34_inst : DFF_X1 port map( D => n7140, CK => CLK, Q => 
                           n_1424, QN => n20800);
   REGISTERS_reg_14_33_inst : DFF_X1 port map( D => n7139, CK => CLK, Q => 
                           n_1425, QN => n20801);
   REGISTERS_reg_14_32_inst : DFF_X1 port map( D => n7138, CK => CLK, Q => 
                           n_1426, QN => n20802);
   REGISTERS_reg_14_31_inst : DFF_X1 port map( D => n7137, CK => CLK, Q => 
                           n_1427, QN => n20803);
   REGISTERS_reg_14_30_inst : DFF_X1 port map( D => n7136, CK => CLK, Q => 
                           n_1428, QN => n20804);
   REGISTERS_reg_14_29_inst : DFF_X1 port map( D => n7135, CK => CLK, Q => 
                           n_1429, QN => n20805);
   REGISTERS_reg_14_28_inst : DFF_X1 port map( D => n7134, CK => CLK, Q => 
                           n_1430, QN => n20806);
   REGISTERS_reg_14_27_inst : DFF_X1 port map( D => n7133, CK => CLK, Q => 
                           n_1431, QN => n20807);
   REGISTERS_reg_14_26_inst : DFF_X1 port map( D => n7132, CK => CLK, Q => 
                           n_1432, QN => n20808);
   REGISTERS_reg_14_25_inst : DFF_X1 port map( D => n7131, CK => CLK, Q => 
                           n_1433, QN => n20809);
   REGISTERS_reg_14_24_inst : DFF_X1 port map( D => n7130, CK => CLK, Q => 
                           n_1434, QN => n20810);
   REGISTERS_reg_14_23_inst : DFF_X1 port map( D => n7129, CK => CLK, Q => 
                           n_1435, QN => n20811);
   REGISTERS_reg_14_22_inst : DFF_X1 port map( D => n7128, CK => CLK, Q => 
                           n_1436, QN => n20812);
   REGISTERS_reg_14_21_inst : DFF_X1 port map( D => n7127, CK => CLK, Q => 
                           n_1437, QN => n20813);
   REGISTERS_reg_14_20_inst : DFF_X1 port map( D => n7126, CK => CLK, Q => 
                           n_1438, QN => n20814);
   REGISTERS_reg_14_19_inst : DFF_X1 port map( D => n7125, CK => CLK, Q => 
                           n_1439, QN => n20815);
   REGISTERS_reg_14_18_inst : DFF_X1 port map( D => n7124, CK => CLK, Q => 
                           n_1440, QN => n20816);
   REGISTERS_reg_14_17_inst : DFF_X1 port map( D => n7123, CK => CLK, Q => 
                           n_1441, QN => n20817);
   REGISTERS_reg_14_16_inst : DFF_X1 port map( D => n7122, CK => CLK, Q => 
                           n_1442, QN => n20818);
   REGISTERS_reg_14_15_inst : DFF_X1 port map( D => n7121, CK => CLK, Q => 
                           n_1443, QN => n20819);
   REGISTERS_reg_14_14_inst : DFF_X1 port map( D => n7120, CK => CLK, Q => 
                           n_1444, QN => n20820);
   REGISTERS_reg_14_13_inst : DFF_X1 port map( D => n7119, CK => CLK, Q => 
                           n_1445, QN => n20821);
   REGISTERS_reg_14_12_inst : DFF_X1 port map( D => n7118, CK => CLK, Q => 
                           n_1446, QN => n20822);
   REGISTERS_reg_14_11_inst : DFF_X1 port map( D => n7117, CK => CLK, Q => 
                           n_1447, QN => n20823);
   REGISTERS_reg_14_10_inst : DFF_X1 port map( D => n7116, CK => CLK, Q => 
                           n_1448, QN => n20824);
   REGISTERS_reg_14_9_inst : DFF_X1 port map( D => n7115, CK => CLK, Q => 
                           n_1449, QN => n20825);
   REGISTERS_reg_14_8_inst : DFF_X1 port map( D => n7114, CK => CLK, Q => 
                           n_1450, QN => n20826);
   REGISTERS_reg_14_7_inst : DFF_X1 port map( D => n7113, CK => CLK, Q => 
                           n_1451, QN => n20827);
   REGISTERS_reg_14_6_inst : DFF_X1 port map( D => n7112, CK => CLK, Q => 
                           n_1452, QN => n20828);
   REGISTERS_reg_14_5_inst : DFF_X1 port map( D => n7111, CK => CLK, Q => 
                           n_1453, QN => n20829);
   REGISTERS_reg_14_4_inst : DFF_X1 port map( D => n7110, CK => CLK, Q => 
                           n_1454, QN => n20830);
   REGISTERS_reg_14_3_inst : DFF_X1 port map( D => n7109, CK => CLK, Q => 
                           n_1455, QN => n20831);
   REGISTERS_reg_14_2_inst : DFF_X1 port map( D => n7108, CK => CLK, Q => 
                           n_1456, QN => n20832);
   REGISTERS_reg_14_1_inst : DFF_X1 port map( D => n7107, CK => CLK, Q => 
                           n_1457, QN => n20833);
   REGISTERS_reg_14_0_inst : DFF_X1 port map( D => n7106, CK => CLK, Q => 
                           n_1458, QN => n20834);
   REGISTERS_reg_11_59_inst : DFF_X1 port map( D => n7357, CK => CLK, Q => 
                           n_1459, QN => n21940);
   REGISTERS_reg_11_58_inst : DFF_X1 port map( D => n7356, CK => CLK, Q => 
                           n_1460, QN => n21941);
   REGISTERS_reg_11_57_inst : DFF_X1 port map( D => n7355, CK => CLK, Q => 
                           n_1461, QN => n21942);
   REGISTERS_reg_11_56_inst : DFF_X1 port map( D => n7354, CK => CLK, Q => 
                           n_1462, QN => n21943);
   REGISTERS_reg_11_55_inst : DFF_X1 port map( D => n7353, CK => CLK, Q => 
                           n_1463, QN => n21944);
   REGISTERS_reg_11_54_inst : DFF_X1 port map( D => n7352, CK => CLK, Q => 
                           n_1464, QN => n21945);
   REGISTERS_reg_11_53_inst : DFF_X1 port map( D => n7351, CK => CLK, Q => 
                           n_1465, QN => n21946);
   REGISTERS_reg_11_52_inst : DFF_X1 port map( D => n7350, CK => CLK, Q => 
                           n_1466, QN => n21947);
   REGISTERS_reg_11_51_inst : DFF_X1 port map( D => n7349, CK => CLK, Q => 
                           n_1467, QN => n21948);
   REGISTERS_reg_11_50_inst : DFF_X1 port map( D => n7348, CK => CLK, Q => 
                           n_1468, QN => n21949);
   REGISTERS_reg_11_49_inst : DFF_X1 port map( D => n7347, CK => CLK, Q => 
                           n_1469, QN => n21950);
   REGISTERS_reg_11_48_inst : DFF_X1 port map( D => n7346, CK => CLK, Q => 
                           n_1470, QN => n21951);
   REGISTERS_reg_11_47_inst : DFF_X1 port map( D => n7345, CK => CLK, Q => 
                           n_1471, QN => n21952);
   REGISTERS_reg_11_46_inst : DFF_X1 port map( D => n7344, CK => CLK, Q => 
                           n_1472, QN => n21953);
   REGISTERS_reg_11_45_inst : DFF_X1 port map( D => n7343, CK => CLK, Q => 
                           n_1473, QN => n21954);
   REGISTERS_reg_11_44_inst : DFF_X1 port map( D => n7342, CK => CLK, Q => 
                           n_1474, QN => n21955);
   REGISTERS_reg_11_43_inst : DFF_X1 port map( D => n7341, CK => CLK, Q => 
                           n_1475, QN => n21956);
   REGISTERS_reg_11_42_inst : DFF_X1 port map( D => n7340, CK => CLK, Q => 
                           n_1476, QN => n21957);
   REGISTERS_reg_11_41_inst : DFF_X1 port map( D => n7339, CK => CLK, Q => 
                           n_1477, QN => n21958);
   REGISTERS_reg_11_40_inst : DFF_X1 port map( D => n7338, CK => CLK, Q => 
                           n_1478, QN => n21959);
   REGISTERS_reg_11_39_inst : DFF_X1 port map( D => n7337, CK => CLK, Q => 
                           n_1479, QN => n21960);
   REGISTERS_reg_11_38_inst : DFF_X1 port map( D => n7336, CK => CLK, Q => 
                           n_1480, QN => n21961);
   REGISTERS_reg_11_37_inst : DFF_X1 port map( D => n7335, CK => CLK, Q => 
                           n_1481, QN => n21962);
   REGISTERS_reg_11_36_inst : DFF_X1 port map( D => n7334, CK => CLK, Q => 
                           n_1482, QN => n21963);
   REGISTERS_reg_11_35_inst : DFF_X1 port map( D => n7333, CK => CLK, Q => 
                           n_1483, QN => n21964);
   REGISTERS_reg_11_34_inst : DFF_X1 port map( D => n7332, CK => CLK, Q => 
                           n_1484, QN => n21965);
   REGISTERS_reg_11_33_inst : DFF_X1 port map( D => n7331, CK => CLK, Q => 
                           n_1485, QN => n21966);
   REGISTERS_reg_11_32_inst : DFF_X1 port map( D => n7330, CK => CLK, Q => 
                           n_1486, QN => n21967);
   REGISTERS_reg_11_31_inst : DFF_X1 port map( D => n7329, CK => CLK, Q => 
                           n_1487, QN => n21968);
   REGISTERS_reg_11_30_inst : DFF_X1 port map( D => n7328, CK => CLK, Q => 
                           n_1488, QN => n21969);
   REGISTERS_reg_11_29_inst : DFF_X1 port map( D => n7327, CK => CLK, Q => 
                           n_1489, QN => n21970);
   REGISTERS_reg_11_28_inst : DFF_X1 port map( D => n7326, CK => CLK, Q => 
                           n_1490, QN => n21971);
   REGISTERS_reg_11_27_inst : DFF_X1 port map( D => n7325, CK => CLK, Q => 
                           n_1491, QN => n21972);
   REGISTERS_reg_11_26_inst : DFF_X1 port map( D => n7324, CK => CLK, Q => 
                           n_1492, QN => n21973);
   REGISTERS_reg_11_25_inst : DFF_X1 port map( D => n7323, CK => CLK, Q => 
                           n_1493, QN => n21974);
   REGISTERS_reg_11_24_inst : DFF_X1 port map( D => n7322, CK => CLK, Q => 
                           n_1494, QN => n21975);
   REGISTERS_reg_11_23_inst : DFF_X1 port map( D => n7321, CK => CLK, Q => 
                           n_1495, QN => n21976);
   REGISTERS_reg_11_22_inst : DFF_X1 port map( D => n7320, CK => CLK, Q => 
                           n_1496, QN => n21977);
   REGISTERS_reg_11_21_inst : DFF_X1 port map( D => n7319, CK => CLK, Q => 
                           n_1497, QN => n21978);
   REGISTERS_reg_11_20_inst : DFF_X1 port map( D => n7318, CK => CLK, Q => 
                           n_1498, QN => n21979);
   REGISTERS_reg_11_19_inst : DFF_X1 port map( D => n7317, CK => CLK, Q => 
                           n_1499, QN => n21980);
   REGISTERS_reg_11_18_inst : DFF_X1 port map( D => n7316, CK => CLK, Q => 
                           n_1500, QN => n21981);
   REGISTERS_reg_11_17_inst : DFF_X1 port map( D => n7315, CK => CLK, Q => 
                           n_1501, QN => n21982);
   REGISTERS_reg_11_16_inst : DFF_X1 port map( D => n7314, CK => CLK, Q => 
                           n_1502, QN => n21983);
   REGISTERS_reg_11_15_inst : DFF_X1 port map( D => n7313, CK => CLK, Q => 
                           n_1503, QN => n21984);
   REGISTERS_reg_11_14_inst : DFF_X1 port map( D => n7312, CK => CLK, Q => 
                           n_1504, QN => n21985);
   REGISTERS_reg_11_13_inst : DFF_X1 port map( D => n7311, CK => CLK, Q => 
                           n_1505, QN => n21986);
   REGISTERS_reg_11_12_inst : DFF_X1 port map( D => n7310, CK => CLK, Q => 
                           n_1506, QN => n21987);
   REGISTERS_reg_11_11_inst : DFF_X1 port map( D => n7309, CK => CLK, Q => 
                           n_1507, QN => n21988);
   REGISTERS_reg_11_10_inst : DFF_X1 port map( D => n7308, CK => CLK, Q => 
                           n_1508, QN => n21989);
   REGISTERS_reg_11_9_inst : DFF_X1 port map( D => n7307, CK => CLK, Q => 
                           n_1509, QN => n21990);
   REGISTERS_reg_11_8_inst : DFF_X1 port map( D => n7306, CK => CLK, Q => 
                           n_1510, QN => n21991);
   REGISTERS_reg_11_7_inst : DFF_X1 port map( D => n7305, CK => CLK, Q => 
                           n_1511, QN => n21992);
   REGISTERS_reg_11_6_inst : DFF_X1 port map( D => n7304, CK => CLK, Q => 
                           n_1512, QN => n21993);
   REGISTERS_reg_11_5_inst : DFF_X1 port map( D => n7303, CK => CLK, Q => 
                           n_1513, QN => n21994);
   REGISTERS_reg_11_4_inst : DFF_X1 port map( D => n7302, CK => CLK, Q => 
                           n_1514, QN => n21995);
   REGISTERS_reg_11_3_inst : DFF_X1 port map( D => n7301, CK => CLK, Q => 
                           n_1515, QN => n21996);
   REGISTERS_reg_11_2_inst : DFF_X1 port map( D => n7300, CK => CLK, Q => 
                           n_1516, QN => n21997);
   REGISTERS_reg_11_1_inst : DFF_X1 port map( D => n7299, CK => CLK, Q => 
                           n_1517, QN => n21998);
   REGISTERS_reg_11_0_inst : DFF_X1 port map( D => n7298, CK => CLK, Q => 
                           n_1518, QN => n21999);
   REGISTERS_reg_8_59_inst : DFF_X1 port map( D => n7549, CK => CLK, Q => 
                           n_1519, QN => n22440);
   REGISTERS_reg_8_58_inst : DFF_X1 port map( D => n7548, CK => CLK, Q => 
                           n_1520, QN => n22441);
   REGISTERS_reg_8_57_inst : DFF_X1 port map( D => n7547, CK => CLK, Q => 
                           n_1521, QN => n22442);
   REGISTERS_reg_8_56_inst : DFF_X1 port map( D => n7546, CK => CLK, Q => 
                           n_1522, QN => n22443);
   REGISTERS_reg_8_55_inst : DFF_X1 port map( D => n7545, CK => CLK, Q => 
                           n_1523, QN => n22444);
   REGISTERS_reg_8_54_inst : DFF_X1 port map( D => n7544, CK => CLK, Q => 
                           n_1524, QN => n22445);
   REGISTERS_reg_8_53_inst : DFF_X1 port map( D => n7543, CK => CLK, Q => 
                           n_1525, QN => n22446);
   REGISTERS_reg_8_52_inst : DFF_X1 port map( D => n7542, CK => CLK, Q => 
                           n_1526, QN => n22447);
   REGISTERS_reg_8_51_inst : DFF_X1 port map( D => n7541, CK => CLK, Q => 
                           n_1527, QN => n22448);
   REGISTERS_reg_8_50_inst : DFF_X1 port map( D => n7540, CK => CLK, Q => 
                           n_1528, QN => n22449);
   REGISTERS_reg_8_49_inst : DFF_X1 port map( D => n7539, CK => CLK, Q => 
                           n_1529, QN => n22450);
   REGISTERS_reg_8_48_inst : DFF_X1 port map( D => n7538, CK => CLK, Q => 
                           n_1530, QN => n22451);
   REGISTERS_reg_8_47_inst : DFF_X1 port map( D => n7537, CK => CLK, Q => 
                           n_1531, QN => n22452);
   REGISTERS_reg_8_46_inst : DFF_X1 port map( D => n7536, CK => CLK, Q => 
                           n_1532, QN => n22453);
   REGISTERS_reg_8_45_inst : DFF_X1 port map( D => n7535, CK => CLK, Q => 
                           n_1533, QN => n22454);
   REGISTERS_reg_8_44_inst : DFF_X1 port map( D => n7534, CK => CLK, Q => 
                           n_1534, QN => n22455);
   REGISTERS_reg_8_43_inst : DFF_X1 port map( D => n7533, CK => CLK, Q => 
                           n_1535, QN => n22456);
   REGISTERS_reg_8_42_inst : DFF_X1 port map( D => n7532, CK => CLK, Q => 
                           n_1536, QN => n22457);
   REGISTERS_reg_8_41_inst : DFF_X1 port map( D => n7531, CK => CLK, Q => 
                           n_1537, QN => n22458);
   REGISTERS_reg_8_40_inst : DFF_X1 port map( D => n7530, CK => CLK, Q => 
                           n_1538, QN => n22459);
   REGISTERS_reg_8_39_inst : DFF_X1 port map( D => n7529, CK => CLK, Q => 
                           n_1539, QN => n22460);
   REGISTERS_reg_8_38_inst : DFF_X1 port map( D => n7528, CK => CLK, Q => 
                           n_1540, QN => n22461);
   REGISTERS_reg_8_37_inst : DFF_X1 port map( D => n7527, CK => CLK, Q => 
                           n_1541, QN => n22462);
   REGISTERS_reg_8_36_inst : DFF_X1 port map( D => n7526, CK => CLK, Q => 
                           n_1542, QN => n22463);
   REGISTERS_reg_8_35_inst : DFF_X1 port map( D => n7525, CK => CLK, Q => 
                           n_1543, QN => n22464);
   REGISTERS_reg_8_34_inst : DFF_X1 port map( D => n7524, CK => CLK, Q => 
                           n_1544, QN => n22465);
   REGISTERS_reg_8_33_inst : DFF_X1 port map( D => n7523, CK => CLK, Q => 
                           n_1545, QN => n22466);
   REGISTERS_reg_8_32_inst : DFF_X1 port map( D => n7522, CK => CLK, Q => 
                           n_1546, QN => n22467);
   REGISTERS_reg_8_31_inst : DFF_X1 port map( D => n7521, CK => CLK, Q => 
                           n_1547, QN => n22468);
   REGISTERS_reg_8_30_inst : DFF_X1 port map( D => n7520, CK => CLK, Q => 
                           n_1548, QN => n22469);
   REGISTERS_reg_8_29_inst : DFF_X1 port map( D => n7519, CK => CLK, Q => 
                           n_1549, QN => n22470);
   REGISTERS_reg_8_28_inst : DFF_X1 port map( D => n7518, CK => CLK, Q => 
                           n_1550, QN => n22471);
   REGISTERS_reg_8_27_inst : DFF_X1 port map( D => n7517, CK => CLK, Q => 
                           n_1551, QN => n22472);
   REGISTERS_reg_8_26_inst : DFF_X1 port map( D => n7516, CK => CLK, Q => 
                           n_1552, QN => n22473);
   REGISTERS_reg_8_25_inst : DFF_X1 port map( D => n7515, CK => CLK, Q => 
                           n_1553, QN => n22474);
   REGISTERS_reg_8_24_inst : DFF_X1 port map( D => n7514, CK => CLK, Q => 
                           n_1554, QN => n22475);
   REGISTERS_reg_8_23_inst : DFF_X1 port map( D => n7513, CK => CLK, Q => 
                           n_1555, QN => n22476);
   REGISTERS_reg_8_22_inst : DFF_X1 port map( D => n7512, CK => CLK, Q => 
                           n_1556, QN => n22477);
   REGISTERS_reg_8_21_inst : DFF_X1 port map( D => n7511, CK => CLK, Q => 
                           n_1557, QN => n22478);
   REGISTERS_reg_8_20_inst : DFF_X1 port map( D => n7510, CK => CLK, Q => 
                           n_1558, QN => n22479);
   REGISTERS_reg_8_19_inst : DFF_X1 port map( D => n7509, CK => CLK, Q => 
                           n_1559, QN => n22480);
   REGISTERS_reg_8_18_inst : DFF_X1 port map( D => n7508, CK => CLK, Q => 
                           n_1560, QN => n22481);
   REGISTERS_reg_8_17_inst : DFF_X1 port map( D => n7507, CK => CLK, Q => 
                           n_1561, QN => n22482);
   REGISTERS_reg_8_16_inst : DFF_X1 port map( D => n7506, CK => CLK, Q => 
                           n_1562, QN => n22483);
   REGISTERS_reg_8_15_inst : DFF_X1 port map( D => n7505, CK => CLK, Q => 
                           n_1563, QN => n22484);
   REGISTERS_reg_8_14_inst : DFF_X1 port map( D => n7504, CK => CLK, Q => 
                           n_1564, QN => n22485);
   REGISTERS_reg_8_13_inst : DFF_X1 port map( D => n7503, CK => CLK, Q => 
                           n_1565, QN => n22486);
   REGISTERS_reg_8_12_inst : DFF_X1 port map( D => n7502, CK => CLK, Q => 
                           n_1566, QN => n22487);
   REGISTERS_reg_8_11_inst : DFF_X1 port map( D => n7501, CK => CLK, Q => 
                           n_1567, QN => n22488);
   REGISTERS_reg_8_10_inst : DFF_X1 port map( D => n7500, CK => CLK, Q => 
                           n_1568, QN => n22489);
   REGISTERS_reg_8_9_inst : DFF_X1 port map( D => n7499, CK => CLK, Q => n_1569
                           , QN => n22490);
   REGISTERS_reg_8_8_inst : DFF_X1 port map( D => n7498, CK => CLK, Q => n_1570
                           , QN => n22491);
   REGISTERS_reg_8_7_inst : DFF_X1 port map( D => n7497, CK => CLK, Q => n_1571
                           , QN => n22492);
   REGISTERS_reg_8_6_inst : DFF_X1 port map( D => n7496, CK => CLK, Q => n_1572
                           , QN => n22493);
   REGISTERS_reg_8_5_inst : DFF_X1 port map( D => n7495, CK => CLK, Q => n_1573
                           , QN => n22494);
   REGISTERS_reg_8_4_inst : DFF_X1 port map( D => n7494, CK => CLK, Q => n_1574
                           , QN => n22495);
   REGISTERS_reg_8_3_inst : DFF_X1 port map( D => n7493, CK => CLK, Q => n_1575
                           , QN => n22496);
   REGISTERS_reg_8_2_inst : DFF_X1 port map( D => n7492, CK => CLK, Q => n_1576
                           , QN => n22497);
   REGISTERS_reg_8_1_inst : DFF_X1 port map( D => n7491, CK => CLK, Q => n_1577
                           , QN => n22498);
   REGISTERS_reg_8_0_inst : DFF_X1 port map( D => n7490, CK => CLK, Q => n_1578
                           , QN => n22499);
   REGISTERS_reg_3_59_inst : DFF_X1 port map( D => n7869, CK => CLK, Q => 
                           n_1579, QN => n21360);
   REGISTERS_reg_3_58_inst : DFF_X1 port map( D => n7868, CK => CLK, Q => 
                           n_1580, QN => n21361);
   REGISTERS_reg_3_57_inst : DFF_X1 port map( D => n7867, CK => CLK, Q => 
                           n_1581, QN => n21362);
   REGISTERS_reg_3_56_inst : DFF_X1 port map( D => n7866, CK => CLK, Q => 
                           n_1582, QN => n21363);
   REGISTERS_reg_3_55_inst : DFF_X1 port map( D => n7865, CK => CLK, Q => 
                           n_1583, QN => n21364);
   REGISTERS_reg_3_54_inst : DFF_X1 port map( D => n7864, CK => CLK, Q => 
                           n_1584, QN => n21365);
   REGISTERS_reg_3_53_inst : DFF_X1 port map( D => n7863, CK => CLK, Q => 
                           n_1585, QN => n21366);
   REGISTERS_reg_3_52_inst : DFF_X1 port map( D => n7862, CK => CLK, Q => 
                           n_1586, QN => n21367);
   REGISTERS_reg_3_51_inst : DFF_X1 port map( D => n7861, CK => CLK, Q => 
                           n_1587, QN => n21368);
   REGISTERS_reg_3_50_inst : DFF_X1 port map( D => n7860, CK => CLK, Q => 
                           n_1588, QN => n21369);
   REGISTERS_reg_3_49_inst : DFF_X1 port map( D => n7859, CK => CLK, Q => 
                           n_1589, QN => n21370);
   REGISTERS_reg_3_48_inst : DFF_X1 port map( D => n7858, CK => CLK, Q => 
                           n_1590, QN => n21371);
   REGISTERS_reg_3_47_inst : DFF_X1 port map( D => n7857, CK => CLK, Q => 
                           n_1591, QN => n21372);
   REGISTERS_reg_3_46_inst : DFF_X1 port map( D => n7856, CK => CLK, Q => 
                           n_1592, QN => n21373);
   REGISTERS_reg_3_45_inst : DFF_X1 port map( D => n7855, CK => CLK, Q => 
                           n_1593, QN => n21374);
   REGISTERS_reg_3_44_inst : DFF_X1 port map( D => n7854, CK => CLK, Q => 
                           n_1594, QN => n21375);
   REGISTERS_reg_3_43_inst : DFF_X1 port map( D => n7853, CK => CLK, Q => 
                           n_1595, QN => n21376);
   REGISTERS_reg_3_42_inst : DFF_X1 port map( D => n7852, CK => CLK, Q => 
                           n_1596, QN => n21377);
   REGISTERS_reg_3_41_inst : DFF_X1 port map( D => n7851, CK => CLK, Q => 
                           n_1597, QN => n21378);
   REGISTERS_reg_3_40_inst : DFF_X1 port map( D => n7850, CK => CLK, Q => 
                           n_1598, QN => n21379);
   REGISTERS_reg_3_39_inst : DFF_X1 port map( D => n7849, CK => CLK, Q => 
                           n_1599, QN => n21380);
   REGISTERS_reg_3_38_inst : DFF_X1 port map( D => n7848, CK => CLK, Q => 
                           n_1600, QN => n21381);
   REGISTERS_reg_3_37_inst : DFF_X1 port map( D => n7847, CK => CLK, Q => 
                           n_1601, QN => n21382);
   REGISTERS_reg_3_36_inst : DFF_X1 port map( D => n7846, CK => CLK, Q => 
                           n_1602, QN => n21383);
   REGISTERS_reg_3_35_inst : DFF_X1 port map( D => n7845, CK => CLK, Q => 
                           n_1603, QN => n21384);
   REGISTERS_reg_3_34_inst : DFF_X1 port map( D => n7844, CK => CLK, Q => 
                           n_1604, QN => n21385);
   REGISTERS_reg_3_33_inst : DFF_X1 port map( D => n7843, CK => CLK, Q => 
                           n_1605, QN => n21386);
   REGISTERS_reg_3_32_inst : DFF_X1 port map( D => n7842, CK => CLK, Q => 
                           n_1606, QN => n21387);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n7841, CK => CLK, Q => 
                           n_1607, QN => n21388);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n7840, CK => CLK, Q => 
                           n_1608, QN => n21389);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n7839, CK => CLK, Q => 
                           n_1609, QN => n21390);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n7838, CK => CLK, Q => 
                           n_1610, QN => n21391);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n7837, CK => CLK, Q => 
                           n_1611, QN => n21392);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n7836, CK => CLK, Q => 
                           n_1612, QN => n21393);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n7835, CK => CLK, Q => 
                           n_1613, QN => n21394);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n7834, CK => CLK, Q => 
                           n_1614, QN => n21395);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n7833, CK => CLK, Q => 
                           n_1615, QN => n21396);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n7832, CK => CLK, Q => 
                           n_1616, QN => n21397);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n7831, CK => CLK, Q => 
                           n_1617, QN => n21398);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n7830, CK => CLK, Q => 
                           n_1618, QN => n21399);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n7829, CK => CLK, Q => 
                           n_1619, QN => n21400);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n7828, CK => CLK, Q => 
                           n_1620, QN => n21401);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n7827, CK => CLK, Q => 
                           n_1621, QN => n21402);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n7826, CK => CLK, Q => 
                           n_1622, QN => n21403);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n7825, CK => CLK, Q => 
                           n_1623, QN => n21404);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n7824, CK => CLK, Q => 
                           n_1624, QN => n21405);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n7823, CK => CLK, Q => 
                           n_1625, QN => n21406);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n7822, CK => CLK, Q => 
                           n_1626, QN => n21407);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n7821, CK => CLK, Q => 
                           n_1627, QN => n21408);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n7820, CK => CLK, Q => 
                           n_1628, QN => n21409);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n7819, CK => CLK, Q => n_1629
                           , QN => n21410);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n7818, CK => CLK, Q => n_1630
                           , QN => n21411);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n7817, CK => CLK, Q => n_1631
                           , QN => n21412);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n7816, CK => CLK, Q => n_1632
                           , QN => n21413);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n7815, CK => CLK, Q => n_1633
                           , QN => n21414);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n7814, CK => CLK, Q => n_1634
                           , QN => n21415);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n7813, CK => CLK, Q => n_1635
                           , QN => n21416);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n7812, CK => CLK, Q => n_1636
                           , QN => n21417);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n7811, CK => CLK, Q => n_1637
                           , QN => n21418);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n7810, CK => CLK, Q => n_1638
                           , QN => n21419);
   REGISTERS_reg_24_63_inst : DFF_X1 port map( D => n6529, CK => CLK, Q => 
                           n_1639, QN => n22500);
   REGISTERS_reg_24_62_inst : DFF_X1 port map( D => n6528, CK => CLK, Q => 
                           n_1640, QN => n22501);
   REGISTERS_reg_24_61_inst : DFF_X1 port map( D => n6527, CK => CLK, Q => 
                           n_1641, QN => n22502);
   REGISTERS_reg_24_60_inst : DFF_X1 port map( D => n6526, CK => CLK, Q => 
                           n_1642, QN => n22503);
   REGISTERS_reg_23_63_inst : DFF_X1 port map( D => n6593, CK => CLK, Q => 
                           n_1643, QN => n21164);
   REGISTERS_reg_23_62_inst : DFF_X1 port map( D => n6592, CK => CLK, Q => 
                           n_1644, QN => n21165);
   REGISTERS_reg_23_61_inst : DFF_X1 port map( D => n6591, CK => CLK, Q => 
                           n_1645, QN => n21166);
   REGISTERS_reg_23_60_inst : DFF_X1 port map( D => n6590, CK => CLK, Q => 
                           n_1646, QN => n21167);
   REGISTERS_reg_17_63_inst : DFF_X1 port map( D => n6977, CK => CLK, Q => 
                           n_1647, QN => n21488);
   REGISTERS_reg_17_62_inst : DFF_X1 port map( D => n6976, CK => CLK, Q => 
                           n_1648, QN => n21489);
   REGISTERS_reg_17_61_inst : DFF_X1 port map( D => n6975, CK => CLK, Q => 
                           n_1649, QN => n21490);
   REGISTERS_reg_17_60_inst : DFF_X1 port map( D => n6974, CK => CLK, Q => 
                           n_1650, QN => n21491);
   REGISTERS_reg_12_63_inst : DFF_X1 port map( D => n7297, CK => CLK, Q => 
                           n_1651, QN => n20708);
   REGISTERS_reg_12_62_inst : DFF_X1 port map( D => n7296, CK => CLK, Q => 
                           n_1652, QN => n20709);
   REGISTERS_reg_12_61_inst : DFF_X1 port map( D => n7295, CK => CLK, Q => 
                           n_1653, QN => n20710);
   REGISTERS_reg_12_60_inst : DFF_X1 port map( D => n7294, CK => CLK, Q => 
                           n_1654, QN => n20711);
   REGISTERS_reg_9_63_inst : DFF_X1 port map( D => n7489, CK => CLK, Q => 
                           n_1655, QN => n22508);
   REGISTERS_reg_9_62_inst : DFF_X1 port map( D => n7488, CK => CLK, Q => 
                           n_1656, QN => n22509);
   REGISTERS_reg_9_61_inst : DFF_X1 port map( D => n7487, CK => CLK, Q => 
                           n_1657, QN => n22510);
   REGISTERS_reg_9_60_inst : DFF_X1 port map( D => n7486, CK => CLK, Q => 
                           n_1658, QN => n22511);
   REGISTERS_reg_7_63_inst : DFF_X1 port map( D => n7617, CK => CLK, Q => 
                           n_1659, QN => n21508);
   REGISTERS_reg_7_62_inst : DFF_X1 port map( D => n7616, CK => CLK, Q => 
                           n_1660, QN => n21509);
   REGISTERS_reg_7_61_inst : DFF_X1 port map( D => n7615, CK => CLK, Q => 
                           n_1661, QN => n21510);
   REGISTERS_reg_7_60_inst : DFF_X1 port map( D => n7614, CK => CLK, Q => 
                           n_1662, QN => n21511);
   REGISTERS_reg_5_63_inst : DFF_X1 port map( D => n7745, CK => CLK, Q => 
                           n_1663, QN => n21176);
   REGISTERS_reg_5_62_inst : DFF_X1 port map( D => n7744, CK => CLK, Q => 
                           n_1664, QN => n21177);
   REGISTERS_reg_5_61_inst : DFF_X1 port map( D => n7743, CK => CLK, Q => 
                           n_1665, QN => n21178);
   REGISTERS_reg_5_60_inst : DFF_X1 port map( D => n7742, CK => CLK, Q => 
                           n_1666, QN => n21179);
   REGISTERS_reg_24_59_inst : DFF_X1 port map( D => n6525, CK => CLK, Q => 
                           n_1667, QN => n22512);
   REGISTERS_reg_24_58_inst : DFF_X1 port map( D => n6524, CK => CLK, Q => 
                           n_1668, QN => n22513);
   REGISTERS_reg_24_57_inst : DFF_X1 port map( D => n6523, CK => CLK, Q => 
                           n_1669, QN => n22514);
   REGISTERS_reg_24_56_inst : DFF_X1 port map( D => n6522, CK => CLK, Q => 
                           n_1670, QN => n22515);
   REGISTERS_reg_24_55_inst : DFF_X1 port map( D => n6521, CK => CLK, Q => 
                           n_1671, QN => n22516);
   REGISTERS_reg_24_54_inst : DFF_X1 port map( D => n6520, CK => CLK, Q => 
                           n_1672, QN => n22517);
   REGISTERS_reg_24_53_inst : DFF_X1 port map( D => n6519, CK => CLK, Q => 
                           n_1673, QN => n22518);
   REGISTERS_reg_24_52_inst : DFF_X1 port map( D => n6518, CK => CLK, Q => 
                           n_1674, QN => n22519);
   REGISTERS_reg_24_51_inst : DFF_X1 port map( D => n6517, CK => CLK, Q => 
                           n_1675, QN => n22520);
   REGISTERS_reg_24_50_inst : DFF_X1 port map( D => n6516, CK => CLK, Q => 
                           n_1676, QN => n22521);
   REGISTERS_reg_24_49_inst : DFF_X1 port map( D => n6515, CK => CLK, Q => 
                           n_1677, QN => n22522);
   REGISTERS_reg_24_48_inst : DFF_X1 port map( D => n6514, CK => CLK, Q => 
                           n_1678, QN => n22523);
   REGISTERS_reg_24_47_inst : DFF_X1 port map( D => n6513, CK => CLK, Q => 
                           n_1679, QN => n22524);
   REGISTERS_reg_24_46_inst : DFF_X1 port map( D => n6512, CK => CLK, Q => 
                           n_1680, QN => n22525);
   REGISTERS_reg_24_45_inst : DFF_X1 port map( D => n6511, CK => CLK, Q => 
                           n_1681, QN => n22526);
   REGISTERS_reg_24_44_inst : DFF_X1 port map( D => n6510, CK => CLK, Q => 
                           n_1682, QN => n22527);
   REGISTERS_reg_24_43_inst : DFF_X1 port map( D => n6509, CK => CLK, Q => 
                           n_1683, QN => n22528);
   REGISTERS_reg_24_42_inst : DFF_X1 port map( D => n6508, CK => CLK, Q => 
                           n_1684, QN => n22529);
   REGISTERS_reg_24_41_inst : DFF_X1 port map( D => n6507, CK => CLK, Q => 
                           n_1685, QN => n22530);
   REGISTERS_reg_24_40_inst : DFF_X1 port map( D => n6506, CK => CLK, Q => 
                           n_1686, QN => n22531);
   REGISTERS_reg_24_39_inst : DFF_X1 port map( D => n6505, CK => CLK, Q => 
                           n_1687, QN => n22532);
   REGISTERS_reg_24_38_inst : DFF_X1 port map( D => n6504, CK => CLK, Q => 
                           n_1688, QN => n22533);
   REGISTERS_reg_24_37_inst : DFF_X1 port map( D => n6503, CK => CLK, Q => 
                           n_1689, QN => n22534);
   REGISTERS_reg_24_36_inst : DFF_X1 port map( D => n6502, CK => CLK, Q => 
                           n_1690, QN => n22535);
   REGISTERS_reg_24_35_inst : DFF_X1 port map( D => n6501, CK => CLK, Q => 
                           n_1691, QN => n22536);
   REGISTERS_reg_24_34_inst : DFF_X1 port map( D => n6500, CK => CLK, Q => 
                           n_1692, QN => n22537);
   REGISTERS_reg_24_33_inst : DFF_X1 port map( D => n6499, CK => CLK, Q => 
                           n_1693, QN => n22538);
   REGISTERS_reg_24_32_inst : DFF_X1 port map( D => n6498, CK => CLK, Q => 
                           n_1694, QN => n22539);
   REGISTERS_reg_24_31_inst : DFF_X1 port map( D => n6497, CK => CLK, Q => 
                           n_1695, QN => n22540);
   REGISTERS_reg_24_30_inst : DFF_X1 port map( D => n6496, CK => CLK, Q => 
                           n_1696, QN => n22541);
   REGISTERS_reg_24_29_inst : DFF_X1 port map( D => n6495, CK => CLK, Q => 
                           n_1697, QN => n22542);
   REGISTERS_reg_24_28_inst : DFF_X1 port map( D => n6494, CK => CLK, Q => 
                           n_1698, QN => n22543);
   REGISTERS_reg_24_27_inst : DFF_X1 port map( D => n6493, CK => CLK, Q => 
                           n_1699, QN => n22544);
   REGISTERS_reg_24_26_inst : DFF_X1 port map( D => n6492, CK => CLK, Q => 
                           n_1700, QN => n22545);
   REGISTERS_reg_24_25_inst : DFF_X1 port map( D => n6491, CK => CLK, Q => 
                           n_1701, QN => n22546);
   REGISTERS_reg_24_24_inst : DFF_X1 port map( D => n6490, CK => CLK, Q => 
                           n_1702, QN => n22547);
   REGISTERS_reg_24_23_inst : DFF_X1 port map( D => n6489, CK => CLK, Q => 
                           n_1703, QN => n22548);
   REGISTERS_reg_24_22_inst : DFF_X1 port map( D => n6488, CK => CLK, Q => 
                           n_1704, QN => n22549);
   REGISTERS_reg_24_21_inst : DFF_X1 port map( D => n6487, CK => CLK, Q => 
                           n_1705, QN => n22550);
   REGISTERS_reg_24_20_inst : DFF_X1 port map( D => n6486, CK => CLK, Q => 
                           n_1706, QN => n22551);
   REGISTERS_reg_24_19_inst : DFF_X1 port map( D => n6485, CK => CLK, Q => 
                           n_1707, QN => n22552);
   REGISTERS_reg_24_18_inst : DFF_X1 port map( D => n6484, CK => CLK, Q => 
                           n_1708, QN => n22553);
   REGISTERS_reg_24_17_inst : DFF_X1 port map( D => n6483, CK => CLK, Q => 
                           n_1709, QN => n22554);
   REGISTERS_reg_24_16_inst : DFF_X1 port map( D => n6482, CK => CLK, Q => 
                           n_1710, QN => n22555);
   REGISTERS_reg_24_15_inst : DFF_X1 port map( D => n6481, CK => CLK, Q => 
                           n_1711, QN => n22556);
   REGISTERS_reg_24_14_inst : DFF_X1 port map( D => n6480, CK => CLK, Q => 
                           n_1712, QN => n22557);
   REGISTERS_reg_24_13_inst : DFF_X1 port map( D => n6479, CK => CLK, Q => 
                           n_1713, QN => n22558);
   REGISTERS_reg_24_12_inst : DFF_X1 port map( D => n6478, CK => CLK, Q => 
                           n_1714, QN => n22559);
   REGISTERS_reg_24_11_inst : DFF_X1 port map( D => n6477, CK => CLK, Q => 
                           n_1715, QN => n22560);
   REGISTERS_reg_24_10_inst : DFF_X1 port map( D => n6476, CK => CLK, Q => 
                           n_1716, QN => n22561);
   REGISTERS_reg_24_9_inst : DFF_X1 port map( D => n6475, CK => CLK, Q => 
                           n_1717, QN => n22562);
   REGISTERS_reg_24_8_inst : DFF_X1 port map( D => n6474, CK => CLK, Q => 
                           n_1718, QN => n22563);
   REGISTERS_reg_24_7_inst : DFF_X1 port map( D => n6473, CK => CLK, Q => 
                           n_1719, QN => n22564);
   REGISTERS_reg_24_6_inst : DFF_X1 port map( D => n6472, CK => CLK, Q => 
                           n_1720, QN => n22565);
   REGISTERS_reg_24_5_inst : DFF_X1 port map( D => n6471, CK => CLK, Q => 
                           n_1721, QN => n22566);
   REGISTERS_reg_24_4_inst : DFF_X1 port map( D => n6470, CK => CLK, Q => 
                           n_1722, QN => n22567);
   REGISTERS_reg_24_3_inst : DFF_X1 port map( D => n6469, CK => CLK, Q => 
                           n_1723, QN => n22568);
   REGISTERS_reg_24_2_inst : DFF_X1 port map( D => n6468, CK => CLK, Q => 
                           n_1724, QN => n22569);
   REGISTERS_reg_24_1_inst : DFF_X1 port map( D => n6467, CK => CLK, Q => 
                           n_1725, QN => n22570);
   REGISTERS_reg_24_0_inst : DFF_X1 port map( D => n6466, CK => CLK, Q => 
                           n_1726, QN => n22571);
   REGISTERS_reg_23_59_inst : DFF_X1 port map( D => n6589, CK => CLK, Q => 
                           n_1727, QN => n21300);
   REGISTERS_reg_23_58_inst : DFF_X1 port map( D => n6588, CK => CLK, Q => 
                           n_1728, QN => n21301);
   REGISTERS_reg_23_57_inst : DFF_X1 port map( D => n6587, CK => CLK, Q => 
                           n_1729, QN => n21302);
   REGISTERS_reg_23_56_inst : DFF_X1 port map( D => n6586, CK => CLK, Q => 
                           n_1730, QN => n21303);
   REGISTERS_reg_23_55_inst : DFF_X1 port map( D => n6585, CK => CLK, Q => 
                           n_1731, QN => n21304);
   REGISTERS_reg_23_54_inst : DFF_X1 port map( D => n6584, CK => CLK, Q => 
                           n_1732, QN => n21305);
   REGISTERS_reg_23_53_inst : DFF_X1 port map( D => n6583, CK => CLK, Q => 
                           n_1733, QN => n21306);
   REGISTERS_reg_23_52_inst : DFF_X1 port map( D => n6582, CK => CLK, Q => 
                           n_1734, QN => n21307);
   REGISTERS_reg_23_51_inst : DFF_X1 port map( D => n6581, CK => CLK, Q => 
                           n_1735, QN => n21308);
   REGISTERS_reg_23_50_inst : DFF_X1 port map( D => n6580, CK => CLK, Q => 
                           n_1736, QN => n21309);
   REGISTERS_reg_23_49_inst : DFF_X1 port map( D => n6579, CK => CLK, Q => 
                           n_1737, QN => n21310);
   REGISTERS_reg_23_48_inst : DFF_X1 port map( D => n6578, CK => CLK, Q => 
                           n_1738, QN => n21311);
   REGISTERS_reg_23_47_inst : DFF_X1 port map( D => n6577, CK => CLK, Q => 
                           n_1739, QN => n21312);
   REGISTERS_reg_23_46_inst : DFF_X1 port map( D => n6576, CK => CLK, Q => 
                           n_1740, QN => n21313);
   REGISTERS_reg_23_45_inst : DFF_X1 port map( D => n6575, CK => CLK, Q => 
                           n_1741, QN => n21314);
   REGISTERS_reg_23_44_inst : DFF_X1 port map( D => n6574, CK => CLK, Q => 
                           n_1742, QN => n21315);
   REGISTERS_reg_23_43_inst : DFF_X1 port map( D => n6573, CK => CLK, Q => 
                           n_1743, QN => n21316);
   REGISTERS_reg_23_42_inst : DFF_X1 port map( D => n6572, CK => CLK, Q => 
                           n_1744, QN => n21317);
   REGISTERS_reg_23_41_inst : DFF_X1 port map( D => n6571, CK => CLK, Q => 
                           n_1745, QN => n21318);
   REGISTERS_reg_23_40_inst : DFF_X1 port map( D => n6570, CK => CLK, Q => 
                           n_1746, QN => n21319);
   REGISTERS_reg_23_39_inst : DFF_X1 port map( D => n6569, CK => CLK, Q => 
                           n_1747, QN => n21320);
   REGISTERS_reg_23_38_inst : DFF_X1 port map( D => n6568, CK => CLK, Q => 
                           n_1748, QN => n21321);
   REGISTERS_reg_23_37_inst : DFF_X1 port map( D => n6567, CK => CLK, Q => 
                           n_1749, QN => n21322);
   REGISTERS_reg_23_36_inst : DFF_X1 port map( D => n6566, CK => CLK, Q => 
                           n_1750, QN => n21323);
   REGISTERS_reg_23_35_inst : DFF_X1 port map( D => n6565, CK => CLK, Q => 
                           n_1751, QN => n21324);
   REGISTERS_reg_23_34_inst : DFF_X1 port map( D => n6564, CK => CLK, Q => 
                           n_1752, QN => n21325);
   REGISTERS_reg_23_33_inst : DFF_X1 port map( D => n6563, CK => CLK, Q => 
                           n_1753, QN => n21326);
   REGISTERS_reg_23_32_inst : DFF_X1 port map( D => n6562, CK => CLK, Q => 
                           n_1754, QN => n21327);
   REGISTERS_reg_23_31_inst : DFF_X1 port map( D => n6561, CK => CLK, Q => 
                           n_1755, QN => n21328);
   REGISTERS_reg_23_30_inst : DFF_X1 port map( D => n6560, CK => CLK, Q => 
                           n_1756, QN => n21329);
   REGISTERS_reg_23_29_inst : DFF_X1 port map( D => n6559, CK => CLK, Q => 
                           n_1757, QN => n21330);
   REGISTERS_reg_23_28_inst : DFF_X1 port map( D => n6558, CK => CLK, Q => 
                           n_1758, QN => n21331);
   REGISTERS_reg_23_27_inst : DFF_X1 port map( D => n6557, CK => CLK, Q => 
                           n_1759, QN => n21332);
   REGISTERS_reg_23_26_inst : DFF_X1 port map( D => n6556, CK => CLK, Q => 
                           n_1760, QN => n21333);
   REGISTERS_reg_23_25_inst : DFF_X1 port map( D => n6555, CK => CLK, Q => 
                           n_1761, QN => n21334);
   REGISTERS_reg_23_24_inst : DFF_X1 port map( D => n6554, CK => CLK, Q => 
                           n_1762, QN => n21335);
   REGISTERS_reg_23_23_inst : DFF_X1 port map( D => n6553, CK => CLK, Q => 
                           n_1763, QN => n21336);
   REGISTERS_reg_23_22_inst : DFF_X1 port map( D => n6552, CK => CLK, Q => 
                           n_1764, QN => n21337);
   REGISTERS_reg_23_21_inst : DFF_X1 port map( D => n6551, CK => CLK, Q => 
                           n_1765, QN => n21338);
   REGISTERS_reg_23_20_inst : DFF_X1 port map( D => n6550, CK => CLK, Q => 
                           n_1766, QN => n21339);
   REGISTERS_reg_23_19_inst : DFF_X1 port map( D => n6549, CK => CLK, Q => 
                           n_1767, QN => n21340);
   REGISTERS_reg_23_18_inst : DFF_X1 port map( D => n6548, CK => CLK, Q => 
                           n_1768, QN => n21341);
   REGISTERS_reg_23_17_inst : DFF_X1 port map( D => n6547, CK => CLK, Q => 
                           n_1769, QN => n21342);
   REGISTERS_reg_23_16_inst : DFF_X1 port map( D => n6546, CK => CLK, Q => 
                           n_1770, QN => n21343);
   REGISTERS_reg_23_15_inst : DFF_X1 port map( D => n6545, CK => CLK, Q => 
                           n_1771, QN => n21344);
   REGISTERS_reg_23_14_inst : DFF_X1 port map( D => n6544, CK => CLK, Q => 
                           n_1772, QN => n21345);
   REGISTERS_reg_23_13_inst : DFF_X1 port map( D => n6543, CK => CLK, Q => 
                           n_1773, QN => n21346);
   REGISTERS_reg_23_12_inst : DFF_X1 port map( D => n6542, CK => CLK, Q => 
                           n_1774, QN => n21347);
   REGISTERS_reg_23_11_inst : DFF_X1 port map( D => n6541, CK => CLK, Q => 
                           n_1775, QN => n21348);
   REGISTERS_reg_23_10_inst : DFF_X1 port map( D => n6540, CK => CLK, Q => 
                           n_1776, QN => n21349);
   REGISTERS_reg_23_9_inst : DFF_X1 port map( D => n6539, CK => CLK, Q => 
                           n_1777, QN => n21350);
   REGISTERS_reg_23_8_inst : DFF_X1 port map( D => n6538, CK => CLK, Q => 
                           n_1778, QN => n21351);
   REGISTERS_reg_23_7_inst : DFF_X1 port map( D => n6537, CK => CLK, Q => 
                           n_1779, QN => n21352);
   REGISTERS_reg_23_6_inst : DFF_X1 port map( D => n6536, CK => CLK, Q => 
                           n_1780, QN => n21353);
   REGISTERS_reg_23_5_inst : DFF_X1 port map( D => n6535, CK => CLK, Q => 
                           n_1781, QN => n21354);
   REGISTERS_reg_23_4_inst : DFF_X1 port map( D => n6534, CK => CLK, Q => 
                           n_1782, QN => n21355);
   REGISTERS_reg_23_3_inst : DFF_X1 port map( D => n6533, CK => CLK, Q => 
                           n_1783, QN => n21356);
   REGISTERS_reg_23_2_inst : DFF_X1 port map( D => n6532, CK => CLK, Q => 
                           n_1784, QN => n21357);
   REGISTERS_reg_23_1_inst : DFF_X1 port map( D => n6531, CK => CLK, Q => 
                           n_1785, QN => n21358);
   REGISTERS_reg_23_0_inst : DFF_X1 port map( D => n6530, CK => CLK, Q => 
                           n_1786, QN => n21359);
   REGISTERS_reg_17_59_inst : DFF_X1 port map( D => n6973, CK => CLK, Q => 
                           n_1787, QN => n21700);
   REGISTERS_reg_17_58_inst : DFF_X1 port map( D => n6972, CK => CLK, Q => 
                           n_1788, QN => n21701);
   REGISTERS_reg_17_57_inst : DFF_X1 port map( D => n6971, CK => CLK, Q => 
                           n_1789, QN => n21702);
   REGISTERS_reg_17_56_inst : DFF_X1 port map( D => n6970, CK => CLK, Q => 
                           n_1790, QN => n21703);
   REGISTERS_reg_17_55_inst : DFF_X1 port map( D => n6969, CK => CLK, Q => 
                           n_1791, QN => n21704);
   REGISTERS_reg_17_54_inst : DFF_X1 port map( D => n6968, CK => CLK, Q => 
                           n_1792, QN => n21705);
   REGISTERS_reg_17_53_inst : DFF_X1 port map( D => n6967, CK => CLK, Q => 
                           n_1793, QN => n21706);
   REGISTERS_reg_17_52_inst : DFF_X1 port map( D => n6966, CK => CLK, Q => 
                           n_1794, QN => n21707);
   REGISTERS_reg_17_51_inst : DFF_X1 port map( D => n6965, CK => CLK, Q => 
                           n_1795, QN => n21708);
   REGISTERS_reg_17_50_inst : DFF_X1 port map( D => n6964, CK => CLK, Q => 
                           n_1796, QN => n21709);
   REGISTERS_reg_17_49_inst : DFF_X1 port map( D => n6963, CK => CLK, Q => 
                           n_1797, QN => n21710);
   REGISTERS_reg_17_48_inst : DFF_X1 port map( D => n6962, CK => CLK, Q => 
                           n_1798, QN => n21711);
   REGISTERS_reg_17_47_inst : DFF_X1 port map( D => n6961, CK => CLK, Q => 
                           n_1799, QN => n21712);
   REGISTERS_reg_17_46_inst : DFF_X1 port map( D => n6960, CK => CLK, Q => 
                           n_1800, QN => n21713);
   REGISTERS_reg_17_45_inst : DFF_X1 port map( D => n6959, CK => CLK, Q => 
                           n_1801, QN => n21714);
   REGISTERS_reg_17_44_inst : DFF_X1 port map( D => n6958, CK => CLK, Q => 
                           n_1802, QN => n21715);
   REGISTERS_reg_17_43_inst : DFF_X1 port map( D => n6957, CK => CLK, Q => 
                           n_1803, QN => n21716);
   REGISTERS_reg_17_42_inst : DFF_X1 port map( D => n6956, CK => CLK, Q => 
                           n_1804, QN => n21717);
   REGISTERS_reg_17_41_inst : DFF_X1 port map( D => n6955, CK => CLK, Q => 
                           n_1805, QN => n21718);
   REGISTERS_reg_17_40_inst : DFF_X1 port map( D => n6954, CK => CLK, Q => 
                           n_1806, QN => n21719);
   REGISTERS_reg_17_39_inst : DFF_X1 port map( D => n6953, CK => CLK, Q => 
                           n_1807, QN => n21720);
   REGISTERS_reg_17_38_inst : DFF_X1 port map( D => n6952, CK => CLK, Q => 
                           n_1808, QN => n21721);
   REGISTERS_reg_17_37_inst : DFF_X1 port map( D => n6951, CK => CLK, Q => 
                           n_1809, QN => n21722);
   REGISTERS_reg_17_36_inst : DFF_X1 port map( D => n6950, CK => CLK, Q => 
                           n_1810, QN => n21723);
   REGISTERS_reg_17_35_inst : DFF_X1 port map( D => n6949, CK => CLK, Q => 
                           n_1811, QN => n21724);
   REGISTERS_reg_17_34_inst : DFF_X1 port map( D => n6948, CK => CLK, Q => 
                           n_1812, QN => n21725);
   REGISTERS_reg_17_33_inst : DFF_X1 port map( D => n6947, CK => CLK, Q => 
                           n_1813, QN => n21726);
   REGISTERS_reg_17_32_inst : DFF_X1 port map( D => n6946, CK => CLK, Q => 
                           n_1814, QN => n21727);
   REGISTERS_reg_17_31_inst : DFF_X1 port map( D => n6945, CK => CLK, Q => 
                           n_1815, QN => n21728);
   REGISTERS_reg_17_30_inst : DFF_X1 port map( D => n6944, CK => CLK, Q => 
                           n_1816, QN => n21729);
   REGISTERS_reg_17_29_inst : DFF_X1 port map( D => n6943, CK => CLK, Q => 
                           n_1817, QN => n21730);
   REGISTERS_reg_17_28_inst : DFF_X1 port map( D => n6942, CK => CLK, Q => 
                           n_1818, QN => n21731);
   REGISTERS_reg_17_27_inst : DFF_X1 port map( D => n6941, CK => CLK, Q => 
                           n_1819, QN => n21732);
   REGISTERS_reg_17_26_inst : DFF_X1 port map( D => n6940, CK => CLK, Q => 
                           n_1820, QN => n21733);
   REGISTERS_reg_17_25_inst : DFF_X1 port map( D => n6939, CK => CLK, Q => 
                           n_1821, QN => n21734);
   REGISTERS_reg_17_24_inst : DFF_X1 port map( D => n6938, CK => CLK, Q => 
                           n_1822, QN => n21735);
   REGISTERS_reg_17_23_inst : DFF_X1 port map( D => n6937, CK => CLK, Q => 
                           n_1823, QN => n21736);
   REGISTERS_reg_17_22_inst : DFF_X1 port map( D => n6936, CK => CLK, Q => 
                           n_1824, QN => n21737);
   REGISTERS_reg_17_21_inst : DFF_X1 port map( D => n6935, CK => CLK, Q => 
                           n_1825, QN => n21738);
   REGISTERS_reg_17_20_inst : DFF_X1 port map( D => n6934, CK => CLK, Q => 
                           n_1826, QN => n21739);
   REGISTERS_reg_17_19_inst : DFF_X1 port map( D => n6933, CK => CLK, Q => 
                           n_1827, QN => n21740);
   REGISTERS_reg_17_18_inst : DFF_X1 port map( D => n6932, CK => CLK, Q => 
                           n_1828, QN => n21741);
   REGISTERS_reg_17_17_inst : DFF_X1 port map( D => n6931, CK => CLK, Q => 
                           n_1829, QN => n21742);
   REGISTERS_reg_17_16_inst : DFF_X1 port map( D => n6930, CK => CLK, Q => 
                           n_1830, QN => n21743);
   REGISTERS_reg_17_15_inst : DFF_X1 port map( D => n6929, CK => CLK, Q => 
                           n_1831, QN => n21744);
   REGISTERS_reg_17_14_inst : DFF_X1 port map( D => n6928, CK => CLK, Q => 
                           n_1832, QN => n21745);
   REGISTERS_reg_17_13_inst : DFF_X1 port map( D => n6927, CK => CLK, Q => 
                           n_1833, QN => n21746);
   REGISTERS_reg_17_12_inst : DFF_X1 port map( D => n6926, CK => CLK, Q => 
                           n_1834, QN => n21747);
   REGISTERS_reg_17_11_inst : DFF_X1 port map( D => n6925, CK => CLK, Q => 
                           n_1835, QN => n21748);
   REGISTERS_reg_17_10_inst : DFF_X1 port map( D => n6924, CK => CLK, Q => 
                           n_1836, QN => n21749);
   REGISTERS_reg_17_9_inst : DFF_X1 port map( D => n6923, CK => CLK, Q => 
                           n_1837, QN => n21750);
   REGISTERS_reg_17_8_inst : DFF_X1 port map( D => n6922, CK => CLK, Q => 
                           n_1838, QN => n21751);
   REGISTERS_reg_17_7_inst : DFF_X1 port map( D => n6921, CK => CLK, Q => 
                           n_1839, QN => n21752);
   REGISTERS_reg_17_6_inst : DFF_X1 port map( D => n6920, CK => CLK, Q => 
                           n_1840, QN => n21753);
   REGISTERS_reg_17_5_inst : DFF_X1 port map( D => n6919, CK => CLK, Q => 
                           n_1841, QN => n21754);
   REGISTERS_reg_17_4_inst : DFF_X1 port map( D => n6918, CK => CLK, Q => 
                           n_1842, QN => n21755);
   REGISTERS_reg_17_3_inst : DFF_X1 port map( D => n6917, CK => CLK, Q => 
                           n_1843, QN => n21756);
   REGISTERS_reg_17_2_inst : DFF_X1 port map( D => n6916, CK => CLK, Q => 
                           n_1844, QN => n21757);
   REGISTERS_reg_17_1_inst : DFF_X1 port map( D => n6915, CK => CLK, Q => 
                           n_1845, QN => n21758);
   REGISTERS_reg_17_0_inst : DFF_X1 port map( D => n6914, CK => CLK, Q => 
                           n_1846, QN => n21759);
   REGISTERS_reg_12_59_inst : DFF_X1 port map( D => n7293, CK => CLK, Q => 
                           n_1847, QN => n20712);
   REGISTERS_reg_12_58_inst : DFF_X1 port map( D => n7292, CK => CLK, Q => 
                           n_1848, QN => n20713);
   REGISTERS_reg_12_57_inst : DFF_X1 port map( D => n7291, CK => CLK, Q => 
                           n_1849, QN => n20714);
   REGISTERS_reg_12_56_inst : DFF_X1 port map( D => n7290, CK => CLK, Q => 
                           n_1850, QN => n20715);
   REGISTERS_reg_12_55_inst : DFF_X1 port map( D => n7289, CK => CLK, Q => 
                           n_1851, QN => n20716);
   REGISTERS_reg_12_54_inst : DFF_X1 port map( D => n7288, CK => CLK, Q => 
                           n_1852, QN => n20717);
   REGISTERS_reg_12_53_inst : DFF_X1 port map( D => n7287, CK => CLK, Q => 
                           n_1853, QN => n20718);
   REGISTERS_reg_12_52_inst : DFF_X1 port map( D => n7286, CK => CLK, Q => 
                           n_1854, QN => n20719);
   REGISTERS_reg_12_51_inst : DFF_X1 port map( D => n7285, CK => CLK, Q => 
                           n_1855, QN => n20720);
   REGISTERS_reg_12_50_inst : DFF_X1 port map( D => n7284, CK => CLK, Q => 
                           n_1856, QN => n20721);
   REGISTERS_reg_12_49_inst : DFF_X1 port map( D => n7283, CK => CLK, Q => 
                           n_1857, QN => n20722);
   REGISTERS_reg_12_48_inst : DFF_X1 port map( D => n7282, CK => CLK, Q => 
                           n_1858, QN => n20723);
   REGISTERS_reg_12_47_inst : DFF_X1 port map( D => n7281, CK => CLK, Q => 
                           n_1859, QN => n20724);
   REGISTERS_reg_12_46_inst : DFF_X1 port map( D => n7280, CK => CLK, Q => 
                           n_1860, QN => n20725);
   REGISTERS_reg_12_45_inst : DFF_X1 port map( D => n7279, CK => CLK, Q => 
                           n_1861, QN => n20726);
   REGISTERS_reg_12_44_inst : DFF_X1 port map( D => n7278, CK => CLK, Q => 
                           n_1862, QN => n20727);
   REGISTERS_reg_12_43_inst : DFF_X1 port map( D => n7277, CK => CLK, Q => 
                           n_1863, QN => n20728);
   REGISTERS_reg_12_42_inst : DFF_X1 port map( D => n7276, CK => CLK, Q => 
                           n_1864, QN => n20729);
   REGISTERS_reg_12_41_inst : DFF_X1 port map( D => n7275, CK => CLK, Q => 
                           n_1865, QN => n20730);
   REGISTERS_reg_12_40_inst : DFF_X1 port map( D => n7274, CK => CLK, Q => 
                           n_1866, QN => n20731);
   REGISTERS_reg_12_39_inst : DFF_X1 port map( D => n7273, CK => CLK, Q => 
                           n_1867, QN => n20732);
   REGISTERS_reg_12_38_inst : DFF_X1 port map( D => n7272, CK => CLK, Q => 
                           n_1868, QN => n20733);
   REGISTERS_reg_12_37_inst : DFF_X1 port map( D => n7271, CK => CLK, Q => 
                           n_1869, QN => n20734);
   REGISTERS_reg_12_36_inst : DFF_X1 port map( D => n7270, CK => CLK, Q => 
                           n_1870, QN => n20735);
   REGISTERS_reg_12_35_inst : DFF_X1 port map( D => n7269, CK => CLK, Q => 
                           n_1871, QN => n20736);
   REGISTERS_reg_12_34_inst : DFF_X1 port map( D => n7268, CK => CLK, Q => 
                           n_1872, QN => n20737);
   REGISTERS_reg_12_33_inst : DFF_X1 port map( D => n7267, CK => CLK, Q => 
                           n_1873, QN => n20738);
   REGISTERS_reg_12_32_inst : DFF_X1 port map( D => n7266, CK => CLK, Q => 
                           n_1874, QN => n20739);
   REGISTERS_reg_12_31_inst : DFF_X1 port map( D => n7265, CK => CLK, Q => 
                           n_1875, QN => n20740);
   REGISTERS_reg_12_30_inst : DFF_X1 port map( D => n7264, CK => CLK, Q => 
                           n_1876, QN => n20741);
   REGISTERS_reg_12_29_inst : DFF_X1 port map( D => n7263, CK => CLK, Q => 
                           n_1877, QN => n20742);
   REGISTERS_reg_12_28_inst : DFF_X1 port map( D => n7262, CK => CLK, Q => 
                           n_1878, QN => n20743);
   REGISTERS_reg_12_27_inst : DFF_X1 port map( D => n7261, CK => CLK, Q => 
                           n_1879, QN => n20744);
   REGISTERS_reg_12_26_inst : DFF_X1 port map( D => n7260, CK => CLK, Q => 
                           n_1880, QN => n20745);
   REGISTERS_reg_12_25_inst : DFF_X1 port map( D => n7259, CK => CLK, Q => 
                           n_1881, QN => n20746);
   REGISTERS_reg_12_24_inst : DFF_X1 port map( D => n7258, CK => CLK, Q => 
                           n_1882, QN => n20747);
   REGISTERS_reg_12_23_inst : DFF_X1 port map( D => n7257, CK => CLK, Q => 
                           n_1883, QN => n20748);
   REGISTERS_reg_12_22_inst : DFF_X1 port map( D => n7256, CK => CLK, Q => 
                           n_1884, QN => n20749);
   REGISTERS_reg_12_21_inst : DFF_X1 port map( D => n7255, CK => CLK, Q => 
                           n_1885, QN => n20750);
   REGISTERS_reg_12_20_inst : DFF_X1 port map( D => n7254, CK => CLK, Q => 
                           n_1886, QN => n20751);
   REGISTERS_reg_12_19_inst : DFF_X1 port map( D => n7253, CK => CLK, Q => 
                           n_1887, QN => n20752);
   REGISTERS_reg_12_18_inst : DFF_X1 port map( D => n7252, CK => CLK, Q => 
                           n_1888, QN => n20753);
   REGISTERS_reg_12_17_inst : DFF_X1 port map( D => n7251, CK => CLK, Q => 
                           n_1889, QN => n20754);
   REGISTERS_reg_12_16_inst : DFF_X1 port map( D => n7250, CK => CLK, Q => 
                           n_1890, QN => n20755);
   REGISTERS_reg_12_15_inst : DFF_X1 port map( D => n7249, CK => CLK, Q => 
                           n_1891, QN => n20756);
   REGISTERS_reg_12_14_inst : DFF_X1 port map( D => n7248, CK => CLK, Q => 
                           n_1892, QN => n20757);
   REGISTERS_reg_12_13_inst : DFF_X1 port map( D => n7247, CK => CLK, Q => 
                           n_1893, QN => n20758);
   REGISTERS_reg_12_12_inst : DFF_X1 port map( D => n7246, CK => CLK, Q => 
                           n_1894, QN => n20759);
   REGISTERS_reg_12_11_inst : DFF_X1 port map( D => n7245, CK => CLK, Q => 
                           n_1895, QN => n20760);
   REGISTERS_reg_12_10_inst : DFF_X1 port map( D => n7244, CK => CLK, Q => 
                           n_1896, QN => n20761);
   REGISTERS_reg_12_9_inst : DFF_X1 port map( D => n7243, CK => CLK, Q => 
                           n_1897, QN => n20762);
   REGISTERS_reg_12_8_inst : DFF_X1 port map( D => n7242, CK => CLK, Q => 
                           n_1898, QN => n20763);
   REGISTERS_reg_12_7_inst : DFF_X1 port map( D => n7241, CK => CLK, Q => 
                           n_1899, QN => n20764);
   REGISTERS_reg_12_6_inst : DFF_X1 port map( D => n7240, CK => CLK, Q => 
                           n_1900, QN => n20765);
   REGISTERS_reg_12_5_inst : DFF_X1 port map( D => n7239, CK => CLK, Q => 
                           n_1901, QN => n20766);
   REGISTERS_reg_12_4_inst : DFF_X1 port map( D => n7238, CK => CLK, Q => 
                           n_1902, QN => n20767);
   REGISTERS_reg_12_3_inst : DFF_X1 port map( D => n7237, CK => CLK, Q => 
                           n_1903, QN => n20768);
   REGISTERS_reg_12_2_inst : DFF_X1 port map( D => n7236, CK => CLK, Q => 
                           n_1904, QN => n20769);
   REGISTERS_reg_12_1_inst : DFF_X1 port map( D => n7235, CK => CLK, Q => 
                           n_1905, QN => n20770);
   REGISTERS_reg_12_0_inst : DFF_X1 port map( D => n7234, CK => CLK, Q => 
                           n_1906, QN => n20771);
   REGISTERS_reg_9_59_inst : DFF_X1 port map( D => n7485, CK => CLK, Q => 
                           n_1907, QN => n22632);
   REGISTERS_reg_9_58_inst : DFF_X1 port map( D => n7484, CK => CLK, Q => 
                           n_1908, QN => n22633);
   REGISTERS_reg_9_57_inst : DFF_X1 port map( D => n7483, CK => CLK, Q => 
                           n_1909, QN => n22634);
   REGISTERS_reg_9_56_inst : DFF_X1 port map( D => n7482, CK => CLK, Q => 
                           n_1910, QN => n22635);
   REGISTERS_reg_9_55_inst : DFF_X1 port map( D => n7481, CK => CLK, Q => 
                           n_1911, QN => n22636);
   REGISTERS_reg_9_54_inst : DFF_X1 port map( D => n7480, CK => CLK, Q => 
                           n_1912, QN => n22637);
   REGISTERS_reg_9_53_inst : DFF_X1 port map( D => n7479, CK => CLK, Q => 
                           n_1913, QN => n22638);
   REGISTERS_reg_9_52_inst : DFF_X1 port map( D => n7478, CK => CLK, Q => 
                           n_1914, QN => n22639);
   REGISTERS_reg_9_51_inst : DFF_X1 port map( D => n7477, CK => CLK, Q => 
                           n_1915, QN => n22640);
   REGISTERS_reg_9_50_inst : DFF_X1 port map( D => n7476, CK => CLK, Q => 
                           n_1916, QN => n22641);
   REGISTERS_reg_9_49_inst : DFF_X1 port map( D => n7475, CK => CLK, Q => 
                           n_1917, QN => n22642);
   REGISTERS_reg_9_48_inst : DFF_X1 port map( D => n7474, CK => CLK, Q => 
                           n_1918, QN => n22643);
   REGISTERS_reg_9_47_inst : DFF_X1 port map( D => n7473, CK => CLK, Q => 
                           n_1919, QN => n22644);
   REGISTERS_reg_9_46_inst : DFF_X1 port map( D => n7472, CK => CLK, Q => 
                           n_1920, QN => n22645);
   REGISTERS_reg_9_45_inst : DFF_X1 port map( D => n7471, CK => CLK, Q => 
                           n_1921, QN => n22646);
   REGISTERS_reg_9_44_inst : DFF_X1 port map( D => n7470, CK => CLK, Q => 
                           n_1922, QN => n22647);
   REGISTERS_reg_9_43_inst : DFF_X1 port map( D => n7469, CK => CLK, Q => 
                           n_1923, QN => n22648);
   REGISTERS_reg_9_42_inst : DFF_X1 port map( D => n7468, CK => CLK, Q => 
                           n_1924, QN => n22649);
   REGISTERS_reg_9_41_inst : DFF_X1 port map( D => n7467, CK => CLK, Q => 
                           n_1925, QN => n22650);
   REGISTERS_reg_9_40_inst : DFF_X1 port map( D => n7466, CK => CLK, Q => 
                           n_1926, QN => n22651);
   REGISTERS_reg_9_39_inst : DFF_X1 port map( D => n7465, CK => CLK, Q => 
                           n_1927, QN => n22652);
   REGISTERS_reg_9_38_inst : DFF_X1 port map( D => n7464, CK => CLK, Q => 
                           n_1928, QN => n22653);
   REGISTERS_reg_9_37_inst : DFF_X1 port map( D => n7463, CK => CLK, Q => 
                           n_1929, QN => n22654);
   REGISTERS_reg_9_36_inst : DFF_X1 port map( D => n7462, CK => CLK, Q => 
                           n_1930, QN => n22655);
   REGISTERS_reg_9_35_inst : DFF_X1 port map( D => n7461, CK => CLK, Q => 
                           n_1931, QN => n22656);
   REGISTERS_reg_9_34_inst : DFF_X1 port map( D => n7460, CK => CLK, Q => 
                           n_1932, QN => n22657);
   REGISTERS_reg_9_33_inst : DFF_X1 port map( D => n7459, CK => CLK, Q => 
                           n_1933, QN => n22658);
   REGISTERS_reg_9_32_inst : DFF_X1 port map( D => n7458, CK => CLK, Q => 
                           n_1934, QN => n22659);
   REGISTERS_reg_9_31_inst : DFF_X1 port map( D => n7457, CK => CLK, Q => 
                           n_1935, QN => n22660);
   REGISTERS_reg_9_30_inst : DFF_X1 port map( D => n7456, CK => CLK, Q => 
                           n_1936, QN => n22661);
   REGISTERS_reg_9_29_inst : DFF_X1 port map( D => n7455, CK => CLK, Q => 
                           n_1937, QN => n22662);
   REGISTERS_reg_9_28_inst : DFF_X1 port map( D => n7454, CK => CLK, Q => 
                           n_1938, QN => n22663);
   REGISTERS_reg_9_27_inst : DFF_X1 port map( D => n7453, CK => CLK, Q => 
                           n_1939, QN => n22664);
   REGISTERS_reg_9_26_inst : DFF_X1 port map( D => n7452, CK => CLK, Q => 
                           n_1940, QN => n22665);
   REGISTERS_reg_9_25_inst : DFF_X1 port map( D => n7451, CK => CLK, Q => 
                           n_1941, QN => n22666);
   REGISTERS_reg_9_24_inst : DFF_X1 port map( D => n7450, CK => CLK, Q => 
                           n_1942, QN => n22667);
   REGISTERS_reg_9_23_inst : DFF_X1 port map( D => n7449, CK => CLK, Q => 
                           n_1943, QN => n22668);
   REGISTERS_reg_9_22_inst : DFF_X1 port map( D => n7448, CK => CLK, Q => 
                           n_1944, QN => n22669);
   REGISTERS_reg_9_21_inst : DFF_X1 port map( D => n7447, CK => CLK, Q => 
                           n_1945, QN => n22670);
   REGISTERS_reg_9_20_inst : DFF_X1 port map( D => n7446, CK => CLK, Q => 
                           n_1946, QN => n22671);
   REGISTERS_reg_9_19_inst : DFF_X1 port map( D => n7445, CK => CLK, Q => 
                           n_1947, QN => n22672);
   REGISTERS_reg_9_18_inst : DFF_X1 port map( D => n7444, CK => CLK, Q => 
                           n_1948, QN => n22673);
   REGISTERS_reg_9_17_inst : DFF_X1 port map( D => n7443, CK => CLK, Q => 
                           n_1949, QN => n22674);
   REGISTERS_reg_9_16_inst : DFF_X1 port map( D => n7442, CK => CLK, Q => 
                           n_1950, QN => n22675);
   REGISTERS_reg_9_15_inst : DFF_X1 port map( D => n7441, CK => CLK, Q => 
                           n_1951, QN => n22676);
   REGISTERS_reg_9_14_inst : DFF_X1 port map( D => n7440, CK => CLK, Q => 
                           n_1952, QN => n22677);
   REGISTERS_reg_9_13_inst : DFF_X1 port map( D => n7439, CK => CLK, Q => 
                           n_1953, QN => n22678);
   REGISTERS_reg_9_12_inst : DFF_X1 port map( D => n7438, CK => CLK, Q => 
                           n_1954, QN => n22679);
   REGISTERS_reg_9_11_inst : DFF_X1 port map( D => n7437, CK => CLK, Q => 
                           n_1955, QN => n22680);
   REGISTERS_reg_9_10_inst : DFF_X1 port map( D => n7436, CK => CLK, Q => 
                           n_1956, QN => n22681);
   REGISTERS_reg_9_9_inst : DFF_X1 port map( D => n7435, CK => CLK, Q => n_1957
                           , QN => n22682);
   REGISTERS_reg_9_8_inst : DFF_X1 port map( D => n7434, CK => CLK, Q => n_1958
                           , QN => n22683);
   REGISTERS_reg_9_7_inst : DFF_X1 port map( D => n7433, CK => CLK, Q => n_1959
                           , QN => n22684);
   REGISTERS_reg_9_6_inst : DFF_X1 port map( D => n7432, CK => CLK, Q => n_1960
                           , QN => n22685);
   REGISTERS_reg_9_5_inst : DFF_X1 port map( D => n7431, CK => CLK, Q => n_1961
                           , QN => n22686);
   REGISTERS_reg_9_4_inst : DFF_X1 port map( D => n7430, CK => CLK, Q => n_1962
                           , QN => n22687);
   REGISTERS_reg_9_3_inst : DFF_X1 port map( D => n7429, CK => CLK, Q => n_1963
                           , QN => n22688);
   REGISTERS_reg_9_2_inst : DFF_X1 port map( D => n7428, CK => CLK, Q => n_1964
                           , QN => n22689);
   REGISTERS_reg_9_1_inst : DFF_X1 port map( D => n7427, CK => CLK, Q => n_1965
                           , QN => n22690);
   REGISTERS_reg_9_0_inst : DFF_X1 port map( D => n7426, CK => CLK, Q => n_1966
                           , QN => n22691);
   REGISTERS_reg_7_59_inst : DFF_X1 port map( D => n7613, CK => CLK, Q => 
                           n_1967, QN => n22000);
   REGISTERS_reg_7_58_inst : DFF_X1 port map( D => n7612, CK => CLK, Q => 
                           n_1968, QN => n22001);
   REGISTERS_reg_7_57_inst : DFF_X1 port map( D => n7611, CK => CLK, Q => 
                           n_1969, QN => n22002);
   REGISTERS_reg_7_56_inst : DFF_X1 port map( D => n7610, CK => CLK, Q => 
                           n_1970, QN => n22003);
   REGISTERS_reg_7_55_inst : DFF_X1 port map( D => n7609, CK => CLK, Q => 
                           n_1971, QN => n22004);
   REGISTERS_reg_7_54_inst : DFF_X1 port map( D => n7608, CK => CLK, Q => 
                           n_1972, QN => n22005);
   REGISTERS_reg_7_53_inst : DFF_X1 port map( D => n7607, CK => CLK, Q => 
                           n_1973, QN => n22006);
   REGISTERS_reg_7_52_inst : DFF_X1 port map( D => n7606, CK => CLK, Q => 
                           n_1974, QN => n22007);
   REGISTERS_reg_7_51_inst : DFF_X1 port map( D => n7605, CK => CLK, Q => 
                           n_1975, QN => n22008);
   REGISTERS_reg_7_50_inst : DFF_X1 port map( D => n7604, CK => CLK, Q => 
                           n_1976, QN => n22009);
   REGISTERS_reg_7_49_inst : DFF_X1 port map( D => n7603, CK => CLK, Q => 
                           n_1977, QN => n22010);
   REGISTERS_reg_7_48_inst : DFF_X1 port map( D => n7602, CK => CLK, Q => 
                           n_1978, QN => n22011);
   REGISTERS_reg_7_47_inst : DFF_X1 port map( D => n7601, CK => CLK, Q => 
                           n_1979, QN => n22012);
   REGISTERS_reg_7_46_inst : DFF_X1 port map( D => n7600, CK => CLK, Q => 
                           n_1980, QN => n22013);
   REGISTERS_reg_7_45_inst : DFF_X1 port map( D => n7599, CK => CLK, Q => 
                           n_1981, QN => n22014);
   REGISTERS_reg_7_44_inst : DFF_X1 port map( D => n7598, CK => CLK, Q => 
                           n_1982, QN => n22015);
   REGISTERS_reg_7_43_inst : DFF_X1 port map( D => n7597, CK => CLK, Q => 
                           n_1983, QN => n22016);
   REGISTERS_reg_7_42_inst : DFF_X1 port map( D => n7596, CK => CLK, Q => 
                           n_1984, QN => n22017);
   REGISTERS_reg_7_41_inst : DFF_X1 port map( D => n7595, CK => CLK, Q => 
                           n_1985, QN => n22018);
   REGISTERS_reg_7_40_inst : DFF_X1 port map( D => n7594, CK => CLK, Q => 
                           n_1986, QN => n22019);
   REGISTERS_reg_7_39_inst : DFF_X1 port map( D => n7593, CK => CLK, Q => 
                           n_1987, QN => n22020);
   REGISTERS_reg_7_38_inst : DFF_X1 port map( D => n7592, CK => CLK, Q => 
                           n_1988, QN => n22021);
   REGISTERS_reg_7_37_inst : DFF_X1 port map( D => n7591, CK => CLK, Q => 
                           n_1989, QN => n22022);
   REGISTERS_reg_7_36_inst : DFF_X1 port map( D => n7590, CK => CLK, Q => 
                           n_1990, QN => n22023);
   REGISTERS_reg_7_35_inst : DFF_X1 port map( D => n7589, CK => CLK, Q => 
                           n_1991, QN => n22024);
   REGISTERS_reg_7_34_inst : DFF_X1 port map( D => n7588, CK => CLK, Q => 
                           n_1992, QN => n22025);
   REGISTERS_reg_7_33_inst : DFF_X1 port map( D => n7587, CK => CLK, Q => 
                           n_1993, QN => n22026);
   REGISTERS_reg_7_32_inst : DFF_X1 port map( D => n7586, CK => CLK, Q => 
                           n_1994, QN => n22027);
   REGISTERS_reg_7_31_inst : DFF_X1 port map( D => n7585, CK => CLK, Q => 
                           n_1995, QN => n22028);
   REGISTERS_reg_7_30_inst : DFF_X1 port map( D => n7584, CK => CLK, Q => 
                           n_1996, QN => n22029);
   REGISTERS_reg_7_29_inst : DFF_X1 port map( D => n7583, CK => CLK, Q => 
                           n_1997, QN => n22030);
   REGISTERS_reg_7_28_inst : DFF_X1 port map( D => n7582, CK => CLK, Q => 
                           n_1998, QN => n22031);
   REGISTERS_reg_7_27_inst : DFF_X1 port map( D => n7581, CK => CLK, Q => 
                           n_1999, QN => n22032);
   REGISTERS_reg_7_26_inst : DFF_X1 port map( D => n7580, CK => CLK, Q => 
                           n_2000, QN => n22033);
   REGISTERS_reg_7_25_inst : DFF_X1 port map( D => n7579, CK => CLK, Q => 
                           n_2001, QN => n22034);
   REGISTERS_reg_7_24_inst : DFF_X1 port map( D => n7578, CK => CLK, Q => 
                           n_2002, QN => n22035);
   REGISTERS_reg_7_23_inst : DFF_X1 port map( D => n7577, CK => CLK, Q => 
                           n_2003, QN => n22036);
   REGISTERS_reg_7_22_inst : DFF_X1 port map( D => n7576, CK => CLK, Q => 
                           n_2004, QN => n22037);
   REGISTERS_reg_7_21_inst : DFF_X1 port map( D => n7575, CK => CLK, Q => 
                           n_2005, QN => n22038);
   REGISTERS_reg_7_20_inst : DFF_X1 port map( D => n7574, CK => CLK, Q => 
                           n_2006, QN => n22039);
   REGISTERS_reg_7_19_inst : DFF_X1 port map( D => n7573, CK => CLK, Q => 
                           n_2007, QN => n22040);
   REGISTERS_reg_7_18_inst : DFF_X1 port map( D => n7572, CK => CLK, Q => 
                           n_2008, QN => n22041);
   REGISTERS_reg_7_17_inst : DFF_X1 port map( D => n7571, CK => CLK, Q => 
                           n_2009, QN => n22042);
   REGISTERS_reg_7_16_inst : DFF_X1 port map( D => n7570, CK => CLK, Q => 
                           n_2010, QN => n22043);
   REGISTERS_reg_7_15_inst : DFF_X1 port map( D => n7569, CK => CLK, Q => 
                           n_2011, QN => n22044);
   REGISTERS_reg_7_14_inst : DFF_X1 port map( D => n7568, CK => CLK, Q => 
                           n_2012, QN => n22045);
   REGISTERS_reg_7_13_inst : DFF_X1 port map( D => n7567, CK => CLK, Q => 
                           n_2013, QN => n22046);
   REGISTERS_reg_7_12_inst : DFF_X1 port map( D => n7566, CK => CLK, Q => 
                           n_2014, QN => n22047);
   REGISTERS_reg_7_11_inst : DFF_X1 port map( D => n7565, CK => CLK, Q => 
                           n_2015, QN => n22048);
   REGISTERS_reg_7_10_inst : DFF_X1 port map( D => n7564, CK => CLK, Q => 
                           n_2016, QN => n22049);
   REGISTERS_reg_7_9_inst : DFF_X1 port map( D => n7563, CK => CLK, Q => n_2017
                           , QN => n22050);
   REGISTERS_reg_7_8_inst : DFF_X1 port map( D => n7562, CK => CLK, Q => n_2018
                           , QN => n22051);
   REGISTERS_reg_7_7_inst : DFF_X1 port map( D => n7561, CK => CLK, Q => n_2019
                           , QN => n22052);
   REGISTERS_reg_7_6_inst : DFF_X1 port map( D => n7560, CK => CLK, Q => n_2020
                           , QN => n22053);
   REGISTERS_reg_7_5_inst : DFF_X1 port map( D => n7559, CK => CLK, Q => n_2021
                           , QN => n22054);
   REGISTERS_reg_7_4_inst : DFF_X1 port map( D => n7558, CK => CLK, Q => n_2022
                           , QN => n22055);
   REGISTERS_reg_7_3_inst : DFF_X1 port map( D => n7557, CK => CLK, Q => n_2023
                           , QN => n22056);
   REGISTERS_reg_7_2_inst : DFF_X1 port map( D => n7556, CK => CLK, Q => n_2024
                           , QN => n22057);
   REGISTERS_reg_7_1_inst : DFF_X1 port map( D => n7555, CK => CLK, Q => n_2025
                           , QN => n22058);
   REGISTERS_reg_7_0_inst : DFF_X1 port map( D => n7554, CK => CLK, Q => n_2026
                           , QN => n22059);
   REGISTERS_reg_5_59_inst : DFF_X1 port map( D => n7741, CK => CLK, Q => 
                           n_2027, QN => n21520);
   REGISTERS_reg_5_58_inst : DFF_X1 port map( D => n7740, CK => CLK, Q => 
                           n_2028, QN => n21521);
   REGISTERS_reg_5_57_inst : DFF_X1 port map( D => n7739, CK => CLK, Q => 
                           n_2029, QN => n21522);
   REGISTERS_reg_5_56_inst : DFF_X1 port map( D => n7738, CK => CLK, Q => 
                           n_2030, QN => n21523);
   REGISTERS_reg_5_55_inst : DFF_X1 port map( D => n7737, CK => CLK, Q => 
                           n_2031, QN => n21524);
   REGISTERS_reg_5_54_inst : DFF_X1 port map( D => n7736, CK => CLK, Q => 
                           n_2032, QN => n21525);
   REGISTERS_reg_5_53_inst : DFF_X1 port map( D => n7735, CK => CLK, Q => 
                           n_2033, QN => n21526);
   REGISTERS_reg_5_52_inst : DFF_X1 port map( D => n7734, CK => CLK, Q => 
                           n_2034, QN => n21527);
   REGISTERS_reg_5_51_inst : DFF_X1 port map( D => n7733, CK => CLK, Q => 
                           n_2035, QN => n21528);
   REGISTERS_reg_5_50_inst : DFF_X1 port map( D => n7732, CK => CLK, Q => 
                           n_2036, QN => n21529);
   REGISTERS_reg_5_49_inst : DFF_X1 port map( D => n7731, CK => CLK, Q => 
                           n_2037, QN => n21530);
   REGISTERS_reg_5_48_inst : DFF_X1 port map( D => n7730, CK => CLK, Q => 
                           n_2038, QN => n21531);
   REGISTERS_reg_5_47_inst : DFF_X1 port map( D => n7729, CK => CLK, Q => 
                           n_2039, QN => n21532);
   REGISTERS_reg_5_46_inst : DFF_X1 port map( D => n7728, CK => CLK, Q => 
                           n_2040, QN => n21533);
   REGISTERS_reg_5_45_inst : DFF_X1 port map( D => n7727, CK => CLK, Q => 
                           n_2041, QN => n21534);
   REGISTERS_reg_5_44_inst : DFF_X1 port map( D => n7726, CK => CLK, Q => 
                           n_2042, QN => n21535);
   REGISTERS_reg_5_43_inst : DFF_X1 port map( D => n7725, CK => CLK, Q => 
                           n_2043, QN => n21536);
   REGISTERS_reg_5_42_inst : DFF_X1 port map( D => n7724, CK => CLK, Q => 
                           n_2044, QN => n21537);
   REGISTERS_reg_5_41_inst : DFF_X1 port map( D => n7723, CK => CLK, Q => 
                           n_2045, QN => n21538);
   REGISTERS_reg_5_40_inst : DFF_X1 port map( D => n7722, CK => CLK, Q => 
                           n_2046, QN => n21539);
   REGISTERS_reg_5_39_inst : DFF_X1 port map( D => n7721, CK => CLK, Q => 
                           n_2047, QN => n21540);
   REGISTERS_reg_5_38_inst : DFF_X1 port map( D => n7720, CK => CLK, Q => 
                           n_2048, QN => n21541);
   REGISTERS_reg_5_37_inst : DFF_X1 port map( D => n7719, CK => CLK, Q => 
                           n_2049, QN => n21542);
   REGISTERS_reg_5_36_inst : DFF_X1 port map( D => n7718, CK => CLK, Q => 
                           n_2050, QN => n21543);
   REGISTERS_reg_5_35_inst : DFF_X1 port map( D => n7717, CK => CLK, Q => 
                           n_2051, QN => n21544);
   REGISTERS_reg_5_34_inst : DFF_X1 port map( D => n7716, CK => CLK, Q => 
                           n_2052, QN => n21545);
   REGISTERS_reg_5_33_inst : DFF_X1 port map( D => n7715, CK => CLK, Q => 
                           n_2053, QN => n21546);
   REGISTERS_reg_5_32_inst : DFF_X1 port map( D => n7714, CK => CLK, Q => 
                           n_2054, QN => n21547);
   REGISTERS_reg_5_31_inst : DFF_X1 port map( D => n7713, CK => CLK, Q => 
                           n_2055, QN => n21548);
   REGISTERS_reg_5_30_inst : DFF_X1 port map( D => n7712, CK => CLK, Q => 
                           n_2056, QN => n21549);
   REGISTERS_reg_5_29_inst : DFF_X1 port map( D => n7711, CK => CLK, Q => 
                           n_2057, QN => n21550);
   REGISTERS_reg_5_28_inst : DFF_X1 port map( D => n7710, CK => CLK, Q => 
                           n_2058, QN => n21551);
   REGISTERS_reg_5_27_inst : DFF_X1 port map( D => n7709, CK => CLK, Q => 
                           n_2059, QN => n21552);
   REGISTERS_reg_5_26_inst : DFF_X1 port map( D => n7708, CK => CLK, Q => 
                           n_2060, QN => n21553);
   REGISTERS_reg_5_25_inst : DFF_X1 port map( D => n7707, CK => CLK, Q => 
                           n_2061, QN => n21554);
   REGISTERS_reg_5_24_inst : DFF_X1 port map( D => n7706, CK => CLK, Q => 
                           n_2062, QN => n21555);
   REGISTERS_reg_5_23_inst : DFF_X1 port map( D => n7705, CK => CLK, Q => 
                           n_2063, QN => n21556);
   REGISTERS_reg_5_22_inst : DFF_X1 port map( D => n7704, CK => CLK, Q => 
                           n_2064, QN => n21557);
   REGISTERS_reg_5_21_inst : DFF_X1 port map( D => n7703, CK => CLK, Q => 
                           n_2065, QN => n21558);
   REGISTERS_reg_5_20_inst : DFF_X1 port map( D => n7702, CK => CLK, Q => 
                           n_2066, QN => n21559);
   REGISTERS_reg_5_19_inst : DFF_X1 port map( D => n7701, CK => CLK, Q => 
                           n_2067, QN => n21560);
   REGISTERS_reg_5_18_inst : DFF_X1 port map( D => n7700, CK => CLK, Q => 
                           n_2068, QN => n21561);
   REGISTERS_reg_5_17_inst : DFF_X1 port map( D => n7699, CK => CLK, Q => 
                           n_2069, QN => n21562);
   REGISTERS_reg_5_16_inst : DFF_X1 port map( D => n7698, CK => CLK, Q => 
                           n_2070, QN => n21563);
   REGISTERS_reg_5_15_inst : DFF_X1 port map( D => n7697, CK => CLK, Q => 
                           n_2071, QN => n21564);
   REGISTERS_reg_5_14_inst : DFF_X1 port map( D => n7696, CK => CLK, Q => 
                           n_2072, QN => n21565);
   REGISTERS_reg_5_13_inst : DFF_X1 port map( D => n7695, CK => CLK, Q => 
                           n_2073, QN => n21566);
   REGISTERS_reg_5_12_inst : DFF_X1 port map( D => n7694, CK => CLK, Q => 
                           n_2074, QN => n21567);
   REGISTERS_reg_5_11_inst : DFF_X1 port map( D => n7693, CK => CLK, Q => 
                           n_2075, QN => n21568);
   REGISTERS_reg_5_10_inst : DFF_X1 port map( D => n7692, CK => CLK, Q => 
                           n_2076, QN => n21569);
   REGISTERS_reg_5_9_inst : DFF_X1 port map( D => n7691, CK => CLK, Q => n_2077
                           , QN => n21570);
   REGISTERS_reg_5_8_inst : DFF_X1 port map( D => n7690, CK => CLK, Q => n_2078
                           , QN => n21571);
   REGISTERS_reg_5_7_inst : DFF_X1 port map( D => n7689, CK => CLK, Q => n_2079
                           , QN => n21572);
   REGISTERS_reg_5_6_inst : DFF_X1 port map( D => n7688, CK => CLK, Q => n_2080
                           , QN => n21573);
   REGISTERS_reg_5_5_inst : DFF_X1 port map( D => n7687, CK => CLK, Q => n_2081
                           , QN => n21574);
   REGISTERS_reg_5_4_inst : DFF_X1 port map( D => n7686, CK => CLK, Q => n_2082
                           , QN => n21575);
   REGISTERS_reg_5_3_inst : DFF_X1 port map( D => n7685, CK => CLK, Q => n_2083
                           , QN => n21576);
   REGISTERS_reg_5_2_inst : DFF_X1 port map( D => n7684, CK => CLK, Q => n_2084
                           , QN => n21577);
   REGISTERS_reg_5_1_inst : DFF_X1 port map( D => n7683, CK => CLK, Q => n_2085
                           , QN => n21578);
   REGISTERS_reg_5_0_inst : DFF_X1 port map( D => n7682, CK => CLK, Q => n_2086
                           , QN => n21579);
   REGISTERS_reg_0_63_inst : DFF_X1 port map( D => n8065, CK => CLK, Q => 
                           n25582, QN => n21516);
   REGISTERS_reg_0_62_inst : DFF_X1 port map( D => n8064, CK => CLK, Q => 
                           n25581, QN => n21517);
   REGISTERS_reg_0_61_inst : DFF_X1 port map( D => n8063, CK => CLK, Q => 
                           n25580, QN => n21518);
   REGISTERS_reg_0_60_inst : DFF_X1 port map( D => n8062, CK => CLK, Q => 
                           n25579, QN => n21519);
   REGISTERS_reg_0_59_inst : DFF_X1 port map( D => n8061, CK => CLK, Q => 
                           n25550, QN => n22120);
   REGISTERS_reg_0_58_inst : DFF_X1 port map( D => n8060, CK => CLK, Q => 
                           n25549, QN => n22121);
   REGISTERS_reg_0_57_inst : DFF_X1 port map( D => n8059, CK => CLK, Q => 
                           n25548, QN => n22122);
   REGISTERS_reg_0_56_inst : DFF_X1 port map( D => n8058, CK => CLK, Q => 
                           n25547, QN => n22123);
   REGISTERS_reg_0_55_inst : DFF_X1 port map( D => n8057, CK => CLK, Q => 
                           n25546, QN => n22124);
   REGISTERS_reg_0_54_inst : DFF_X1 port map( D => n8056, CK => CLK, Q => 
                           n25545, QN => n22125);
   REGISTERS_reg_0_53_inst : DFF_X1 port map( D => n8055, CK => CLK, Q => 
                           n25544, QN => n22126);
   REGISTERS_reg_0_52_inst : DFF_X1 port map( D => n8054, CK => CLK, Q => 
                           n25543, QN => n22127);
   REGISTERS_reg_0_51_inst : DFF_X1 port map( D => n8053, CK => CLK, Q => 
                           n25542, QN => n22128);
   REGISTERS_reg_0_50_inst : DFF_X1 port map( D => n8052, CK => CLK, Q => 
                           n25541, QN => n22129);
   REGISTERS_reg_0_49_inst : DFF_X1 port map( D => n8051, CK => CLK, Q => 
                           n25540, QN => n22130);
   REGISTERS_reg_0_48_inst : DFF_X1 port map( D => n8050, CK => CLK, Q => 
                           n25539, QN => n22131);
   REGISTERS_reg_0_47_inst : DFF_X1 port map( D => n8049, CK => CLK, Q => 
                           n25538, QN => n22132);
   REGISTERS_reg_0_46_inst : DFF_X1 port map( D => n8048, CK => CLK, Q => 
                           n25537, QN => n22133);
   REGISTERS_reg_0_45_inst : DFF_X1 port map( D => n8047, CK => CLK, Q => 
                           n25536, QN => n22134);
   REGISTERS_reg_0_44_inst : DFF_X1 port map( D => n8046, CK => CLK, Q => 
                           n25535, QN => n22135);
   REGISTERS_reg_0_43_inst : DFF_X1 port map( D => n8045, CK => CLK, Q => 
                           n25534, QN => n22136);
   REGISTERS_reg_0_42_inst : DFF_X1 port map( D => n8044, CK => CLK, Q => 
                           n25533, QN => n22137);
   REGISTERS_reg_0_41_inst : DFF_X1 port map( D => n8043, CK => CLK, Q => 
                           n25532, QN => n22138);
   REGISTERS_reg_0_40_inst : DFF_X1 port map( D => n8042, CK => CLK, Q => 
                           n25531, QN => n22139);
   REGISTERS_reg_0_39_inst : DFF_X1 port map( D => n8041, CK => CLK, Q => 
                           n25530, QN => n22140);
   REGISTERS_reg_0_38_inst : DFF_X1 port map( D => n8040, CK => CLK, Q => 
                           n25529, QN => n22141);
   REGISTERS_reg_0_37_inst : DFF_X1 port map( D => n8039, CK => CLK, Q => 
                           n25528, QN => n22142);
   REGISTERS_reg_0_36_inst : DFF_X1 port map( D => n8038, CK => CLK, Q => 
                           n25527, QN => n22143);
   REGISTERS_reg_0_35_inst : DFF_X1 port map( D => n8037, CK => CLK, Q => 
                           n25526, QN => n22144);
   REGISTERS_reg_0_34_inst : DFF_X1 port map( D => n8036, CK => CLK, Q => 
                           n25525, QN => n22145);
   REGISTERS_reg_0_33_inst : DFF_X1 port map( D => n8035, CK => CLK, Q => 
                           n25524, QN => n22146);
   REGISTERS_reg_0_32_inst : DFF_X1 port map( D => n8034, CK => CLK, Q => 
                           n25523, QN => n22147);
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n8033, CK => CLK, Q => 
                           n25522, QN => n22148);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n8032, CK => CLK, Q => 
                           n25521, QN => n22149);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n8031, CK => CLK, Q => 
                           n25520, QN => n22150);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n8030, CK => CLK, Q => 
                           n25519, QN => n22151);
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n8029, CK => CLK, Q => 
                           n25518, QN => n22152);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n8028, CK => CLK, Q => 
                           n25517, QN => n22153);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n8027, CK => CLK, Q => 
                           n25516, QN => n22154);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n8026, CK => CLK, Q => 
                           n25515, QN => n22155);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n8025, CK => CLK, Q => 
                           n25514, QN => n22156);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n8024, CK => CLK, Q => 
                           n25513, QN => n22157);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n8023, CK => CLK, Q => 
                           n25512, QN => n22158);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n8022, CK => CLK, Q => 
                           n25511, QN => n22159);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n8021, CK => CLK, Q => 
                           n25510, QN => n22160);
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n8020, CK => CLK, Q => 
                           n25509, QN => n22161);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n8019, CK => CLK, Q => 
                           n25508, QN => n22162);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n8018, CK => CLK, Q => 
                           n25507, QN => n22163);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n8017, CK => CLK, Q => 
                           n25506, QN => n22164);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n8016, CK => CLK, Q => 
                           n25505, QN => n22165);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n8015, CK => CLK, Q => 
                           n25504, QN => n22166);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n8014, CK => CLK, Q => 
                           n25503, QN => n22167);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n8013, CK => CLK, Q => 
                           n25678, QN => n22168);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n8012, CK => CLK, Q => 
                           n25677, QN => n22169);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n8011, CK => CLK, Q => n25676
                           , QN => n22170);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n8010, CK => CLK, Q => n25675
                           , QN => n22171);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n8009, CK => CLK, Q => n25674
                           , QN => n22172);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n8008, CK => CLK, Q => n25673
                           , QN => n22173);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n8007, CK => CLK, Q => n25672
                           , QN => n22174);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n8006, CK => CLK, Q => n25671
                           , QN => n22175);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n8005, CK => CLK, Q => n25670
                           , QN => n22176);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n8004, CK => CLK, Q => n25669
                           , QN => n22177);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n8003, CK => CLK, Q => n25668
                           , QN => n22178);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n8002, CK => CLK, Q => n25667
                           , QN => n22179);
   REGISTERS_reg_4_63_inst : DFF_X1 port map( D => n7809, CK => CLK, Q => 
                           n25574, QN => n21500);
   REGISTERS_reg_4_62_inst : DFF_X1 port map( D => n7808, CK => CLK, Q => 
                           n25573, QN => n21501);
   REGISTERS_reg_4_61_inst : DFF_X1 port map( D => n7807, CK => CLK, Q => 
                           n25572, QN => n21502);
   REGISTERS_reg_4_60_inst : DFF_X1 port map( D => n7806, CK => CLK, Q => 
                           n25571, QN => n21503);
   REGISTERS_reg_30_63_inst : DFF_X1 port map( D => n6145, CK => CLK, Q => 
                           n26198, QN => n20835);
   REGISTERS_reg_30_62_inst : DFF_X1 port map( D => n6144, CK => CLK, Q => 
                           n26197, QN => n20836);
   REGISTERS_reg_30_61_inst : DFF_X1 port map( D => n6143, CK => CLK, Q => 
                           n26196, QN => n20837);
   REGISTERS_reg_30_60_inst : DFF_X1 port map( D => n6142, CK => CLK, Q => 
                           n26195, QN => n20838);
   REGISTERS_reg_28_63_inst : DFF_X1 port map( D => n6273, CK => CLK, Q => 
                           n8450, QN => n22180);
   REGISTERS_reg_28_62_inst : DFF_X1 port map( D => n6272, CK => CLK, Q => 
                           n8453, QN => n22181);
   REGISTERS_reg_28_61_inst : DFF_X1 port map( D => n6271, CK => CLK, Q => 
                           n8456, QN => n22182);
   REGISTERS_reg_28_60_inst : DFF_X1 port map( D => n6270, CK => CLK, Q => 
                           n8459, QN => n22183);
   REGISTERS_reg_27_63_inst : DFF_X1 port map( D => n6337, CK => CLK, Q => 
                           n18367, QN => n22504);
   REGISTERS_reg_27_62_inst : DFF_X1 port map( D => n6336, CK => CLK, Q => 
                           n18384, QN => n22505);
   REGISTERS_reg_27_61_inst : DFF_X1 port map( D => n6335, CK => CLK, Q => 
                           n18401, QN => n22506);
   REGISTERS_reg_27_60_inst : DFF_X1 port map( D => n6334, CK => CLK, Q => 
                           n18418, QN => n22507);
   REGISTERS_reg_2_63_inst : DFF_X1 port map( D => n7937, CK => CLK, Q => 
                           n25566, QN => n21172);
   REGISTERS_reg_2_62_inst : DFF_X1 port map( D => n7936, CK => CLK, Q => 
                           n25565, QN => n21173);
   REGISTERS_reg_2_61_inst : DFF_X1 port map( D => n7935, CK => CLK, Q => 
                           n25564, QN => n21174);
   REGISTERS_reg_2_60_inst : DFF_X1 port map( D => n7934, CK => CLK, Q => 
                           n25563, QN => n21175);
   REGISTERS_reg_4_59_inst : DFF_X1 port map( D => n7805, CK => CLK, Q => 
                           n25454, QN => n21880);
   REGISTERS_reg_4_58_inst : DFF_X1 port map( D => n7804, CK => CLK, Q => 
                           n25453, QN => n21881);
   REGISTERS_reg_4_57_inst : DFF_X1 port map( D => n7803, CK => CLK, Q => 
                           n25452, QN => n21882);
   REGISTERS_reg_4_56_inst : DFF_X1 port map( D => n7802, CK => CLK, Q => 
                           n25451, QN => n21883);
   REGISTERS_reg_4_55_inst : DFF_X1 port map( D => n7801, CK => CLK, Q => 
                           n25450, QN => n21884);
   REGISTERS_reg_4_54_inst : DFF_X1 port map( D => n7800, CK => CLK, Q => 
                           n25449, QN => n21885);
   REGISTERS_reg_4_53_inst : DFF_X1 port map( D => n7799, CK => CLK, Q => 
                           n25448, QN => n21886);
   REGISTERS_reg_4_52_inst : DFF_X1 port map( D => n7798, CK => CLK, Q => 
                           n25447, QN => n21887);
   REGISTERS_reg_4_51_inst : DFF_X1 port map( D => n7797, CK => CLK, Q => 
                           n25446, QN => n21888);
   REGISTERS_reg_4_50_inst : DFF_X1 port map( D => n7796, CK => CLK, Q => 
                           n25445, QN => n21889);
   REGISTERS_reg_4_49_inst : DFF_X1 port map( D => n7795, CK => CLK, Q => 
                           n25444, QN => n21890);
   REGISTERS_reg_4_48_inst : DFF_X1 port map( D => n7794, CK => CLK, Q => 
                           n25443, QN => n21891);
   REGISTERS_reg_4_47_inst : DFF_X1 port map( D => n7793, CK => CLK, Q => 
                           n25442, QN => n21892);
   REGISTERS_reg_4_46_inst : DFF_X1 port map( D => n7792, CK => CLK, Q => 
                           n25441, QN => n21893);
   REGISTERS_reg_4_45_inst : DFF_X1 port map( D => n7791, CK => CLK, Q => 
                           n25440, QN => n21894);
   REGISTERS_reg_4_44_inst : DFF_X1 port map( D => n7790, CK => CLK, Q => 
                           n25439, QN => n21895);
   REGISTERS_reg_4_43_inst : DFF_X1 port map( D => n7789, CK => CLK, Q => 
                           n25438, QN => n21896);
   REGISTERS_reg_4_42_inst : DFF_X1 port map( D => n7788, CK => CLK, Q => 
                           n25437, QN => n21897);
   REGISTERS_reg_4_41_inst : DFF_X1 port map( D => n7787, CK => CLK, Q => 
                           n25436, QN => n21898);
   REGISTERS_reg_4_40_inst : DFF_X1 port map( D => n7786, CK => CLK, Q => 
                           n25435, QN => n21899);
   REGISTERS_reg_4_39_inst : DFF_X1 port map( D => n7785, CK => CLK, Q => 
                           n25434, QN => n21900);
   REGISTERS_reg_4_38_inst : DFF_X1 port map( D => n7784, CK => CLK, Q => 
                           n25433, QN => n21901);
   REGISTERS_reg_4_37_inst : DFF_X1 port map( D => n7783, CK => CLK, Q => 
                           n25432, QN => n21902);
   REGISTERS_reg_4_36_inst : DFF_X1 port map( D => n7782, CK => CLK, Q => 
                           n25431, QN => n21903);
   REGISTERS_reg_4_35_inst : DFF_X1 port map( D => n7781, CK => CLK, Q => 
                           n25430, QN => n21904);
   REGISTERS_reg_4_34_inst : DFF_X1 port map( D => n7780, CK => CLK, Q => 
                           n25429, QN => n21905);
   REGISTERS_reg_4_33_inst : DFF_X1 port map( D => n7779, CK => CLK, Q => 
                           n25428, QN => n21906);
   REGISTERS_reg_4_32_inst : DFF_X1 port map( D => n7778, CK => CLK, Q => 
                           n25427, QN => n21907);
   REGISTERS_reg_4_31_inst : DFF_X1 port map( D => n7777, CK => CLK, Q => 
                           n25426, QN => n21908);
   REGISTERS_reg_4_30_inst : DFF_X1 port map( D => n7776, CK => CLK, Q => 
                           n25425, QN => n21909);
   REGISTERS_reg_4_29_inst : DFF_X1 port map( D => n7775, CK => CLK, Q => 
                           n25424, QN => n21910);
   REGISTERS_reg_4_28_inst : DFF_X1 port map( D => n7774, CK => CLK, Q => 
                           n25423, QN => n21911);
   REGISTERS_reg_4_27_inst : DFF_X1 port map( D => n7773, CK => CLK, Q => 
                           n25422, QN => n21912);
   REGISTERS_reg_4_26_inst : DFF_X1 port map( D => n7772, CK => CLK, Q => 
                           n25421, QN => n21913);
   REGISTERS_reg_4_25_inst : DFF_X1 port map( D => n7771, CK => CLK, Q => 
                           n25420, QN => n21914);
   REGISTERS_reg_4_24_inst : DFF_X1 port map( D => n7770, CK => CLK, Q => 
                           n25419, QN => n21915);
   REGISTERS_reg_4_23_inst : DFF_X1 port map( D => n7769, CK => CLK, Q => 
                           n25418, QN => n21916);
   REGISTERS_reg_4_22_inst : DFF_X1 port map( D => n7768, CK => CLK, Q => 
                           n25417, QN => n21917);
   REGISTERS_reg_4_21_inst : DFF_X1 port map( D => n7767, CK => CLK, Q => 
                           n25416, QN => n21918);
   REGISTERS_reg_4_20_inst : DFF_X1 port map( D => n7766, CK => CLK, Q => 
                           n25415, QN => n21919);
   REGISTERS_reg_4_19_inst : DFF_X1 port map( D => n7765, CK => CLK, Q => 
                           n25414, QN => n21920);
   REGISTERS_reg_4_18_inst : DFF_X1 port map( D => n7764, CK => CLK, Q => 
                           n25413, QN => n21921);
   REGISTERS_reg_4_17_inst : DFF_X1 port map( D => n7763, CK => CLK, Q => 
                           n25412, QN => n21922);
   REGISTERS_reg_4_16_inst : DFF_X1 port map( D => n7762, CK => CLK, Q => 
                           n25411, QN => n21923);
   REGISTERS_reg_4_15_inst : DFF_X1 port map( D => n7761, CK => CLK, Q => 
                           n25410, QN => n21924);
   REGISTERS_reg_4_14_inst : DFF_X1 port map( D => n7760, CK => CLK, Q => 
                           n25409, QN => n21925);
   REGISTERS_reg_4_13_inst : DFF_X1 port map( D => n7759, CK => CLK, Q => 
                           n25408, QN => n21926);
   REGISTERS_reg_4_12_inst : DFF_X1 port map( D => n7758, CK => CLK, Q => 
                           n25407, QN => n21927);
   REGISTERS_reg_4_11_inst : DFF_X1 port map( D => n7757, CK => CLK, Q => 
                           n25630, QN => n21928);
   REGISTERS_reg_4_10_inst : DFF_X1 port map( D => n7756, CK => CLK, Q => 
                           n25629, QN => n21929);
   REGISTERS_reg_4_9_inst : DFF_X1 port map( D => n7755, CK => CLK, Q => n25628
                           , QN => n21930);
   REGISTERS_reg_4_8_inst : DFF_X1 port map( D => n7754, CK => CLK, Q => n25627
                           , QN => n21931);
   REGISTERS_reg_4_7_inst : DFF_X1 port map( D => n7753, CK => CLK, Q => n25626
                           , QN => n21932);
   REGISTERS_reg_4_6_inst : DFF_X1 port map( D => n7752, CK => CLK, Q => n25625
                           , QN => n21933);
   REGISTERS_reg_4_5_inst : DFF_X1 port map( D => n7751, CK => CLK, Q => n25624
                           , QN => n21934);
   REGISTERS_reg_4_4_inst : DFF_X1 port map( D => n7750, CK => CLK, Q => n25623
                           , QN => n21935);
   REGISTERS_reg_4_3_inst : DFF_X1 port map( D => n7749, CK => CLK, Q => n25622
                           , QN => n21936);
   REGISTERS_reg_4_2_inst : DFF_X1 port map( D => n7748, CK => CLK, Q => n25621
                           , QN => n21937);
   REGISTERS_reg_4_1_inst : DFF_X1 port map( D => n7747, CK => CLK, Q => n25620
                           , QN => n21938);
   REGISTERS_reg_4_0_inst : DFF_X1 port map( D => n7746, CK => CLK, Q => n25619
                           , QN => n21939);
   REGISTERS_reg_30_59_inst : DFF_X1 port map( D => n6141, CK => CLK, Q => 
                           n26386, QN => n20839);
   REGISTERS_reg_30_58_inst : DFF_X1 port map( D => n6140, CK => CLK, Q => 
                           n26385, QN => n20840);
   REGISTERS_reg_30_57_inst : DFF_X1 port map( D => n6139, CK => CLK, Q => 
                           n26384, QN => n20841);
   REGISTERS_reg_30_56_inst : DFF_X1 port map( D => n6138, CK => CLK, Q => 
                           n26383, QN => n20842);
   REGISTERS_reg_30_55_inst : DFF_X1 port map( D => n6137, CK => CLK, Q => 
                           n26382, QN => n20843);
   REGISTERS_reg_30_54_inst : DFF_X1 port map( D => n6136, CK => CLK, Q => 
                           n26381, QN => n20844);
   REGISTERS_reg_30_53_inst : DFF_X1 port map( D => n6135, CK => CLK, Q => 
                           n26380, QN => n20845);
   REGISTERS_reg_30_52_inst : DFF_X1 port map( D => n6134, CK => CLK, Q => 
                           n26379, QN => n20846);
   REGISTERS_reg_30_51_inst : DFF_X1 port map( D => n6133, CK => CLK, Q => 
                           n26378, QN => n20847);
   REGISTERS_reg_30_50_inst : DFF_X1 port map( D => n6132, CK => CLK, Q => 
                           n26377, QN => n20848);
   REGISTERS_reg_30_49_inst : DFF_X1 port map( D => n6131, CK => CLK, Q => 
                           n26376, QN => n20849);
   REGISTERS_reg_30_48_inst : DFF_X1 port map( D => n6130, CK => CLK, Q => 
                           n26375, QN => n20850);
   REGISTERS_reg_30_47_inst : DFF_X1 port map( D => n6129, CK => CLK, Q => 
                           n26374, QN => n20851);
   REGISTERS_reg_30_46_inst : DFF_X1 port map( D => n6128, CK => CLK, Q => 
                           n26373, QN => n20852);
   REGISTERS_reg_30_45_inst : DFF_X1 port map( D => n6127, CK => CLK, Q => 
                           n26372, QN => n20853);
   REGISTERS_reg_30_44_inst : DFF_X1 port map( D => n6126, CK => CLK, Q => 
                           n26371, QN => n20854);
   REGISTERS_reg_30_43_inst : DFF_X1 port map( D => n6125, CK => CLK, Q => 
                           n26370, QN => n20855);
   REGISTERS_reg_30_42_inst : DFF_X1 port map( D => n6124, CK => CLK, Q => 
                           n26369, QN => n20856);
   REGISTERS_reg_30_41_inst : DFF_X1 port map( D => n6123, CK => CLK, Q => 
                           n26368, QN => n20857);
   REGISTERS_reg_30_40_inst : DFF_X1 port map( D => n6122, CK => CLK, Q => 
                           n26367, QN => n20858);
   REGISTERS_reg_30_39_inst : DFF_X1 port map( D => n6121, CK => CLK, Q => 
                           n26366, QN => n20859);
   REGISTERS_reg_30_38_inst : DFF_X1 port map( D => n6120, CK => CLK, Q => 
                           n26365, QN => n20860);
   REGISTERS_reg_30_37_inst : DFF_X1 port map( D => n6119, CK => CLK, Q => 
                           n26364, QN => n20861);
   REGISTERS_reg_30_36_inst : DFF_X1 port map( D => n6118, CK => CLK, Q => 
                           n26363, QN => n20862);
   REGISTERS_reg_30_35_inst : DFF_X1 port map( D => n6117, CK => CLK, Q => 
                           n26362, QN => n20863);
   REGISTERS_reg_30_34_inst : DFF_X1 port map( D => n6116, CK => CLK, Q => 
                           n26361, QN => n20864);
   REGISTERS_reg_30_33_inst : DFF_X1 port map( D => n6115, CK => CLK, Q => 
                           n26360, QN => n20865);
   REGISTERS_reg_30_32_inst : DFF_X1 port map( D => n6114, CK => CLK, Q => 
                           n26359, QN => n20866);
   REGISTERS_reg_30_31_inst : DFF_X1 port map( D => n6113, CK => CLK, Q => 
                           n26358, QN => n20867);
   REGISTERS_reg_30_30_inst : DFF_X1 port map( D => n6112, CK => CLK, Q => 
                           n26357, QN => n20868);
   REGISTERS_reg_30_29_inst : DFF_X1 port map( D => n6111, CK => CLK, Q => 
                           n26356, QN => n20869);
   REGISTERS_reg_30_28_inst : DFF_X1 port map( D => n6110, CK => CLK, Q => 
                           n26355, QN => n20870);
   REGISTERS_reg_30_27_inst : DFF_X1 port map( D => n6109, CK => CLK, Q => 
                           n26354, QN => n20871);
   REGISTERS_reg_30_26_inst : DFF_X1 port map( D => n6108, CK => CLK, Q => 
                           n26353, QN => n20872);
   REGISTERS_reg_30_25_inst : DFF_X1 port map( D => n6107, CK => CLK, Q => 
                           n26352, QN => n20873);
   REGISTERS_reg_30_24_inst : DFF_X1 port map( D => n6106, CK => CLK, Q => 
                           n26351, QN => n20874);
   REGISTERS_reg_30_23_inst : DFF_X1 port map( D => n6105, CK => CLK, Q => 
                           n26350, QN => n20875);
   REGISTERS_reg_30_22_inst : DFF_X1 port map( D => n6104, CK => CLK, Q => 
                           n26349, QN => n20876);
   REGISTERS_reg_30_21_inst : DFF_X1 port map( D => n6103, CK => CLK, Q => 
                           n26348, QN => n20877);
   REGISTERS_reg_30_20_inst : DFF_X1 port map( D => n6102, CK => CLK, Q => 
                           n26347, QN => n20878);
   REGISTERS_reg_30_19_inst : DFF_X1 port map( D => n6101, CK => CLK, Q => 
                           n26346, QN => n20879);
   REGISTERS_reg_30_18_inst : DFF_X1 port map( D => n6100, CK => CLK, Q => 
                           n26345, QN => n20880);
   REGISTERS_reg_30_17_inst : DFF_X1 port map( D => n6099, CK => CLK, Q => 
                           n26344, QN => n20881);
   REGISTERS_reg_30_16_inst : DFF_X1 port map( D => n6098, CK => CLK, Q => 
                           n26343, QN => n20882);
   REGISTERS_reg_30_15_inst : DFF_X1 port map( D => n6097, CK => CLK, Q => 
                           n26342, QN => n20883);
   REGISTERS_reg_30_14_inst : DFF_X1 port map( D => n6096, CK => CLK, Q => 
                           n26341, QN => n20884);
   REGISTERS_reg_30_13_inst : DFF_X1 port map( D => n6095, CK => CLK, Q => 
                           n26340, QN => n20885);
   REGISTERS_reg_30_12_inst : DFF_X1 port map( D => n6094, CK => CLK, Q => 
                           n26339, QN => n20886);
   REGISTERS_reg_30_11_inst : DFF_X1 port map( D => n6093, CK => CLK, Q => 
                           n26338, QN => n20887);
   REGISTERS_reg_30_10_inst : DFF_X1 port map( D => n6092, CK => CLK, Q => 
                           n26337, QN => n20888);
   REGISTERS_reg_30_9_inst : DFF_X1 port map( D => n6091, CK => CLK, Q => 
                           n26336, QN => n20889);
   REGISTERS_reg_30_8_inst : DFF_X1 port map( D => n6090, CK => CLK, Q => 
                           n26335, QN => n20890);
   REGISTERS_reg_30_7_inst : DFF_X1 port map( D => n6089, CK => CLK, Q => 
                           n26334, QN => n20891);
   REGISTERS_reg_30_6_inst : DFF_X1 port map( D => n6088, CK => CLK, Q => 
                           n26333, QN => n20892);
   REGISTERS_reg_30_5_inst : DFF_X1 port map( D => n6087, CK => CLK, Q => 
                           n26332, QN => n20893);
   REGISTERS_reg_30_4_inst : DFF_X1 port map( D => n6086, CK => CLK, Q => 
                           n26331, QN => n20894);
   REGISTERS_reg_30_3_inst : DFF_X1 port map( D => n6085, CK => CLK, Q => 
                           n26330, QN => n20895);
   REGISTERS_reg_30_2_inst : DFF_X1 port map( D => n6084, CK => CLK, Q => 
                           n26329, QN => n20896);
   REGISTERS_reg_30_1_inst : DFF_X1 port map( D => n6083, CK => CLK, Q => 
                           n26328, QN => n20897);
   REGISTERS_reg_30_0_inst : DFF_X1 port map( D => n6082, CK => CLK, Q => 
                           n26327, QN => n20898);
   REGISTERS_reg_28_59_inst : DFF_X1 port map( D => n6269, CK => CLK, Q => 
                           n8462, QN => n22184);
   REGISTERS_reg_28_58_inst : DFF_X1 port map( D => n6268, CK => CLK, Q => 
                           n8465, QN => n22185);
   REGISTERS_reg_28_57_inst : DFF_X1 port map( D => n6267, CK => CLK, Q => 
                           n8468, QN => n22186);
   REGISTERS_reg_28_56_inst : DFF_X1 port map( D => n6266, CK => CLK, Q => 
                           n8471, QN => n22187);
   REGISTERS_reg_28_55_inst : DFF_X1 port map( D => n6265, CK => CLK, Q => 
                           n8474, QN => n22188);
   REGISTERS_reg_28_54_inst : DFF_X1 port map( D => n6264, CK => CLK, Q => 
                           n8477, QN => n22189);
   REGISTERS_reg_28_53_inst : DFF_X1 port map( D => n6263, CK => CLK, Q => 
                           n8480, QN => n22190);
   REGISTERS_reg_28_52_inst : DFF_X1 port map( D => n6262, CK => CLK, Q => 
                           n8483, QN => n22191);
   REGISTERS_reg_28_51_inst : DFF_X1 port map( D => n6261, CK => CLK, Q => 
                           n8486, QN => n22192);
   REGISTERS_reg_28_50_inst : DFF_X1 port map( D => n6260, CK => CLK, Q => 
                           n8489, QN => n22193);
   REGISTERS_reg_28_49_inst : DFF_X1 port map( D => n6259, CK => CLK, Q => 
                           n8492, QN => n22194);
   REGISTERS_reg_28_48_inst : DFF_X1 port map( D => n6258, CK => CLK, Q => 
                           n8495, QN => n22195);
   REGISTERS_reg_28_47_inst : DFF_X1 port map( D => n6257, CK => CLK, Q => 
                           n8498, QN => n22196);
   REGISTERS_reg_28_46_inst : DFF_X1 port map( D => n6256, CK => CLK, Q => 
                           n8501, QN => n22197);
   REGISTERS_reg_28_45_inst : DFF_X1 port map( D => n6255, CK => CLK, Q => 
                           n8504, QN => n22198);
   REGISTERS_reg_28_44_inst : DFF_X1 port map( D => n6254, CK => CLK, Q => 
                           n8507, QN => n22199);
   REGISTERS_reg_28_43_inst : DFF_X1 port map( D => n6253, CK => CLK, Q => 
                           n8510, QN => n22200);
   REGISTERS_reg_28_42_inst : DFF_X1 port map( D => n6252, CK => CLK, Q => 
                           n8513, QN => n22201);
   REGISTERS_reg_28_41_inst : DFF_X1 port map( D => n6251, CK => CLK, Q => 
                           n8516, QN => n22202);
   REGISTERS_reg_28_40_inst : DFF_X1 port map( D => n6250, CK => CLK, Q => 
                           n8519, QN => n22203);
   REGISTERS_reg_28_39_inst : DFF_X1 port map( D => n6249, CK => CLK, Q => 
                           n8522, QN => n22204);
   REGISTERS_reg_28_38_inst : DFF_X1 port map( D => n6248, CK => CLK, Q => 
                           n8525, QN => n22205);
   REGISTERS_reg_28_37_inst : DFF_X1 port map( D => n6247, CK => CLK, Q => 
                           n8528, QN => n22206);
   REGISTERS_reg_28_36_inst : DFF_X1 port map( D => n6246, CK => CLK, Q => 
                           n8531, QN => n22207);
   REGISTERS_reg_28_35_inst : DFF_X1 port map( D => n6245, CK => CLK, Q => 
                           n8534, QN => n22208);
   REGISTERS_reg_28_34_inst : DFF_X1 port map( D => n6244, CK => CLK, Q => 
                           n8537, QN => n22209);
   REGISTERS_reg_28_33_inst : DFF_X1 port map( D => n6243, CK => CLK, Q => 
                           n8540, QN => n22210);
   REGISTERS_reg_28_32_inst : DFF_X1 port map( D => n6242, CK => CLK, Q => 
                           n8543, QN => n22211);
   REGISTERS_reg_28_31_inst : DFF_X1 port map( D => n6241, CK => CLK, Q => 
                           n8546, QN => n22212);
   REGISTERS_reg_28_30_inst : DFF_X1 port map( D => n6240, CK => CLK, Q => 
                           n8549, QN => n22213);
   REGISTERS_reg_28_29_inst : DFF_X1 port map( D => n6239, CK => CLK, Q => 
                           n8552, QN => n22214);
   REGISTERS_reg_28_28_inst : DFF_X1 port map( D => n6238, CK => CLK, Q => 
                           n8555, QN => n22215);
   REGISTERS_reg_28_27_inst : DFF_X1 port map( D => n6237, CK => CLK, Q => 
                           n8558, QN => n22216);
   REGISTERS_reg_28_26_inst : DFF_X1 port map( D => n6236, CK => CLK, Q => 
                           n8561, QN => n22217);
   REGISTERS_reg_28_25_inst : DFF_X1 port map( D => n6235, CK => CLK, Q => 
                           n8564, QN => n22218);
   REGISTERS_reg_28_24_inst : DFF_X1 port map( D => n6234, CK => CLK, Q => 
                           n8567, QN => n22219);
   REGISTERS_reg_28_23_inst : DFF_X1 port map( D => n6233, CK => CLK, Q => 
                           n8570, QN => n22220);
   REGISTERS_reg_28_22_inst : DFF_X1 port map( D => n6232, CK => CLK, Q => 
                           n8573, QN => n22221);
   REGISTERS_reg_28_21_inst : DFF_X1 port map( D => n6231, CK => CLK, Q => 
                           n8576, QN => n22222);
   REGISTERS_reg_28_20_inst : DFF_X1 port map( D => n6230, CK => CLK, Q => 
                           n8579, QN => n22223);
   REGISTERS_reg_28_19_inst : DFF_X1 port map( D => n6229, CK => CLK, Q => 
                           n8582, QN => n22224);
   REGISTERS_reg_28_18_inst : DFF_X1 port map( D => n6228, CK => CLK, Q => 
                           n8585, QN => n22225);
   REGISTERS_reg_28_17_inst : DFF_X1 port map( D => n6227, CK => CLK, Q => 
                           n8588, QN => n22226);
   REGISTERS_reg_28_16_inst : DFF_X1 port map( D => n6226, CK => CLK, Q => 
                           n8591, QN => n22227);
   REGISTERS_reg_28_15_inst : DFF_X1 port map( D => n6225, CK => CLK, Q => 
                           n8594, QN => n22228);
   REGISTERS_reg_28_14_inst : DFF_X1 port map( D => n6224, CK => CLK, Q => 
                           n8597, QN => n22229);
   REGISTERS_reg_28_13_inst : DFF_X1 port map( D => n6223, CK => CLK, Q => 
                           n8600, QN => n22230);
   REGISTERS_reg_28_12_inst : DFF_X1 port map( D => n6222, CK => CLK, Q => 
                           n8603, QN => n22231);
   REGISTERS_reg_28_11_inst : DFF_X1 port map( D => n6221, CK => CLK, Q => 
                           n8606, QN => n22232);
   REGISTERS_reg_28_10_inst : DFF_X1 port map( D => n6220, CK => CLK, Q => 
                           n8609, QN => n22233);
   REGISTERS_reg_28_9_inst : DFF_X1 port map( D => n6219, CK => CLK, Q => n8612
                           , QN => n22234);
   REGISTERS_reg_28_8_inst : DFF_X1 port map( D => n6218, CK => CLK, Q => n8615
                           , QN => n22235);
   REGISTERS_reg_28_7_inst : DFF_X1 port map( D => n6217, CK => CLK, Q => n8618
                           , QN => n22236);
   REGISTERS_reg_28_6_inst : DFF_X1 port map( D => n6216, CK => CLK, Q => n8621
                           , QN => n22237);
   REGISTERS_reg_28_5_inst : DFF_X1 port map( D => n6215, CK => CLK, Q => n8624
                           , QN => n22238);
   REGISTERS_reg_28_4_inst : DFF_X1 port map( D => n6214, CK => CLK, Q => n8627
                           , QN => n22239);
   REGISTERS_reg_28_3_inst : DFF_X1 port map( D => n6213, CK => CLK, Q => n8630
                           , QN => n22240);
   REGISTERS_reg_28_2_inst : DFF_X1 port map( D => n6212, CK => CLK, Q => n8633
                           , QN => n22241);
   REGISTERS_reg_28_1_inst : DFF_X1 port map( D => n6211, CK => CLK, Q => n8636
                           , QN => n22242);
   REGISTERS_reg_28_0_inst : DFF_X1 port map( D => n6210, CK => CLK, Q => n8639
                           , QN => n22243);
   REGISTERS_reg_27_59_inst : DFF_X1 port map( D => n6333, CK => CLK, Q => 
                           n18435, QN => n22572);
   REGISTERS_reg_27_58_inst : DFF_X1 port map( D => n6332, CK => CLK, Q => 
                           n18452, QN => n22573);
   REGISTERS_reg_27_57_inst : DFF_X1 port map( D => n6331, CK => CLK, Q => 
                           n18469, QN => n22574);
   REGISTERS_reg_27_56_inst : DFF_X1 port map( D => n6330, CK => CLK, Q => 
                           n18486, QN => n22575);
   REGISTERS_reg_27_55_inst : DFF_X1 port map( D => n6329, CK => CLK, Q => 
                           n18503, QN => n22576);
   REGISTERS_reg_27_54_inst : DFF_X1 port map( D => n6328, CK => CLK, Q => 
                           n18520, QN => n22577);
   REGISTERS_reg_27_53_inst : DFF_X1 port map( D => n6327, CK => CLK, Q => 
                           n18537, QN => n22578);
   REGISTERS_reg_27_52_inst : DFF_X1 port map( D => n6326, CK => CLK, Q => 
                           n18554, QN => n22579);
   REGISTERS_reg_27_51_inst : DFF_X1 port map( D => n6325, CK => CLK, Q => 
                           n18571, QN => n22580);
   REGISTERS_reg_27_50_inst : DFF_X1 port map( D => n6324, CK => CLK, Q => 
                           n18588, QN => n22581);
   REGISTERS_reg_27_49_inst : DFF_X1 port map( D => n6323, CK => CLK, Q => 
                           n18605, QN => n22582);
   REGISTERS_reg_27_48_inst : DFF_X1 port map( D => n6322, CK => CLK, Q => 
                           n18622, QN => n22583);
   REGISTERS_reg_27_47_inst : DFF_X1 port map( D => n6321, CK => CLK, Q => 
                           n18639, QN => n22584);
   REGISTERS_reg_27_46_inst : DFF_X1 port map( D => n6320, CK => CLK, Q => 
                           n18656, QN => n22585);
   REGISTERS_reg_27_45_inst : DFF_X1 port map( D => n6319, CK => CLK, Q => 
                           n18673, QN => n22586);
   REGISTERS_reg_27_44_inst : DFF_X1 port map( D => n6318, CK => CLK, Q => 
                           n18690, QN => n22587);
   REGISTERS_reg_27_43_inst : DFF_X1 port map( D => n6317, CK => CLK, Q => 
                           n18707, QN => n22588);
   REGISTERS_reg_27_42_inst : DFF_X1 port map( D => n6316, CK => CLK, Q => 
                           n18724, QN => n22589);
   REGISTERS_reg_27_41_inst : DFF_X1 port map( D => n6315, CK => CLK, Q => 
                           n18741, QN => n22590);
   REGISTERS_reg_27_40_inst : DFF_X1 port map( D => n6314, CK => CLK, Q => 
                           n18758, QN => n22591);
   REGISTERS_reg_27_39_inst : DFF_X1 port map( D => n6313, CK => CLK, Q => 
                           n18775, QN => n22592);
   REGISTERS_reg_27_38_inst : DFF_X1 port map( D => n6312, CK => CLK, Q => 
                           n18792, QN => n22593);
   REGISTERS_reg_27_37_inst : DFF_X1 port map( D => n6311, CK => CLK, Q => 
                           n18809, QN => n22594);
   REGISTERS_reg_27_36_inst : DFF_X1 port map( D => n6310, CK => CLK, Q => 
                           n18826, QN => n22595);
   REGISTERS_reg_27_35_inst : DFF_X1 port map( D => n6309, CK => CLK, Q => 
                           n18843, QN => n22596);
   REGISTERS_reg_27_34_inst : DFF_X1 port map( D => n6308, CK => CLK, Q => 
                           n18860, QN => n22597);
   REGISTERS_reg_27_33_inst : DFF_X1 port map( D => n6307, CK => CLK, Q => 
                           n18877, QN => n22598);
   REGISTERS_reg_27_32_inst : DFF_X1 port map( D => n6306, CK => CLK, Q => 
                           n18894, QN => n22599);
   REGISTERS_reg_27_31_inst : DFF_X1 port map( D => n6305, CK => CLK, Q => 
                           n18911, QN => n22600);
   REGISTERS_reg_27_30_inst : DFF_X1 port map( D => n6304, CK => CLK, Q => 
                           n18928, QN => n22601);
   REGISTERS_reg_27_29_inst : DFF_X1 port map( D => n6303, CK => CLK, Q => 
                           n18945, QN => n22602);
   REGISTERS_reg_27_28_inst : DFF_X1 port map( D => n6302, CK => CLK, Q => 
                           n18962, QN => n22603);
   REGISTERS_reg_27_27_inst : DFF_X1 port map( D => n6301, CK => CLK, Q => 
                           n18979, QN => n22604);
   REGISTERS_reg_27_26_inst : DFF_X1 port map( D => n6300, CK => CLK, Q => 
                           n18996, QN => n22605);
   REGISTERS_reg_27_25_inst : DFF_X1 port map( D => n6299, CK => CLK, Q => 
                           n19013, QN => n22606);
   REGISTERS_reg_27_24_inst : DFF_X1 port map( D => n6298, CK => CLK, Q => 
                           n19030, QN => n22607);
   REGISTERS_reg_27_23_inst : DFF_X1 port map( D => n6297, CK => CLK, Q => 
                           n19047, QN => n22608);
   REGISTERS_reg_27_22_inst : DFF_X1 port map( D => n6296, CK => CLK, Q => 
                           n19064, QN => n22609);
   REGISTERS_reg_27_21_inst : DFF_X1 port map( D => n6295, CK => CLK, Q => 
                           n19081, QN => n22610);
   REGISTERS_reg_27_20_inst : DFF_X1 port map( D => n6294, CK => CLK, Q => 
                           n19098, QN => n22611);
   REGISTERS_reg_27_19_inst : DFF_X1 port map( D => n6293, CK => CLK, Q => 
                           n19115, QN => n22612);
   REGISTERS_reg_27_18_inst : DFF_X1 port map( D => n6292, CK => CLK, Q => 
                           n19132, QN => n22613);
   REGISTERS_reg_27_17_inst : DFF_X1 port map( D => n6291, CK => CLK, Q => 
                           n19149, QN => n22614);
   REGISTERS_reg_27_16_inst : DFF_X1 port map( D => n6290, CK => CLK, Q => 
                           n19166, QN => n22615);
   REGISTERS_reg_27_15_inst : DFF_X1 port map( D => n6289, CK => CLK, Q => 
                           n19183, QN => n22616);
   REGISTERS_reg_27_14_inst : DFF_X1 port map( D => n6288, CK => CLK, Q => 
                           n19200, QN => n22617);
   REGISTERS_reg_27_13_inst : DFF_X1 port map( D => n6287, CK => CLK, Q => 
                           n19217, QN => n22618);
   REGISTERS_reg_27_12_inst : DFF_X1 port map( D => n6286, CK => CLK, Q => 
                           n19234, QN => n22619);
   REGISTERS_reg_27_11_inst : DFF_X1 port map( D => n6285, CK => CLK, Q => 
                           n19251, QN => n22620);
   REGISTERS_reg_27_10_inst : DFF_X1 port map( D => n6284, CK => CLK, Q => 
                           n19268, QN => n22621);
   REGISTERS_reg_27_9_inst : DFF_X1 port map( D => n6283, CK => CLK, Q => 
                           n19285, QN => n22622);
   REGISTERS_reg_27_8_inst : DFF_X1 port map( D => n6282, CK => CLK, Q => 
                           n19302, QN => n22623);
   REGISTERS_reg_27_7_inst : DFF_X1 port map( D => n6281, CK => CLK, Q => 
                           n19319, QN => n22624);
   REGISTERS_reg_27_6_inst : DFF_X1 port map( D => n6280, CK => CLK, Q => 
                           n19336, QN => n22625);
   REGISTERS_reg_27_5_inst : DFF_X1 port map( D => n6279, CK => CLK, Q => 
                           n19353, QN => n22626);
   REGISTERS_reg_27_4_inst : DFF_X1 port map( D => n6278, CK => CLK, Q => 
                           n19370, QN => n22627);
   REGISTERS_reg_27_3_inst : DFF_X1 port map( D => n6277, CK => CLK, Q => 
                           n19387, QN => n22628);
   REGISTERS_reg_27_2_inst : DFF_X1 port map( D => n6276, CK => CLK, Q => 
                           n19404, QN => n22629);
   REGISTERS_reg_27_1_inst : DFF_X1 port map( D => n6275, CK => CLK, Q => 
                           n19421, QN => n22630);
   REGISTERS_reg_27_0_inst : DFF_X1 port map( D => n6274, CK => CLK, Q => 
                           n19438, QN => n22631);
   REGISTERS_reg_2_59_inst : DFF_X1 port map( D => n7933, CK => CLK, Q => 
                           n25358, QN => n21420);
   REGISTERS_reg_2_58_inst : DFF_X1 port map( D => n7932, CK => CLK, Q => 
                           n25357, QN => n21421);
   REGISTERS_reg_2_57_inst : DFF_X1 port map( D => n7931, CK => CLK, Q => 
                           n25356, QN => n21422);
   REGISTERS_reg_2_56_inst : DFF_X1 port map( D => n7930, CK => CLK, Q => 
                           n25355, QN => n21423);
   REGISTERS_reg_2_55_inst : DFF_X1 port map( D => n7929, CK => CLK, Q => 
                           n25354, QN => n21424);
   REGISTERS_reg_2_54_inst : DFF_X1 port map( D => n7928, CK => CLK, Q => 
                           n25353, QN => n21425);
   REGISTERS_reg_2_53_inst : DFF_X1 port map( D => n7927, CK => CLK, Q => 
                           n25352, QN => n21426);
   REGISTERS_reg_2_52_inst : DFF_X1 port map( D => n7926, CK => CLK, Q => 
                           n25351, QN => n21427);
   REGISTERS_reg_2_51_inst : DFF_X1 port map( D => n7925, CK => CLK, Q => 
                           n25350, QN => n21428);
   REGISTERS_reg_2_50_inst : DFF_X1 port map( D => n7924, CK => CLK, Q => 
                           n25349, QN => n21429);
   REGISTERS_reg_2_49_inst : DFF_X1 port map( D => n7923, CK => CLK, Q => 
                           n25348, QN => n21430);
   REGISTERS_reg_2_48_inst : DFF_X1 port map( D => n7922, CK => CLK, Q => 
                           n25347, QN => n21431);
   REGISTERS_reg_2_47_inst : DFF_X1 port map( D => n7921, CK => CLK, Q => 
                           n25346, QN => n21432);
   REGISTERS_reg_2_46_inst : DFF_X1 port map( D => n7920, CK => CLK, Q => 
                           n25345, QN => n21433);
   REGISTERS_reg_2_45_inst : DFF_X1 port map( D => n7919, CK => CLK, Q => 
                           n25344, QN => n21434);
   REGISTERS_reg_2_44_inst : DFF_X1 port map( D => n7918, CK => CLK, Q => 
                           n25343, QN => n21435);
   REGISTERS_reg_2_43_inst : DFF_X1 port map( D => n7917, CK => CLK, Q => 
                           n25342, QN => n21436);
   REGISTERS_reg_2_42_inst : DFF_X1 port map( D => n7916, CK => CLK, Q => 
                           n25341, QN => n21437);
   REGISTERS_reg_2_41_inst : DFF_X1 port map( D => n7915, CK => CLK, Q => 
                           n25340, QN => n21438);
   REGISTERS_reg_2_40_inst : DFF_X1 port map( D => n7914, CK => CLK, Q => 
                           n25339, QN => n21439);
   REGISTERS_reg_2_39_inst : DFF_X1 port map( D => n7913, CK => CLK, Q => 
                           n25338, QN => n21440);
   REGISTERS_reg_2_38_inst : DFF_X1 port map( D => n7912, CK => CLK, Q => 
                           n25337, QN => n21441);
   REGISTERS_reg_2_37_inst : DFF_X1 port map( D => n7911, CK => CLK, Q => 
                           n25336, QN => n21442);
   REGISTERS_reg_2_36_inst : DFF_X1 port map( D => n7910, CK => CLK, Q => 
                           n25335, QN => n21443);
   REGISTERS_reg_2_35_inst : DFF_X1 port map( D => n7909, CK => CLK, Q => 
                           n25334, QN => n21444);
   REGISTERS_reg_2_34_inst : DFF_X1 port map( D => n7908, CK => CLK, Q => 
                           n25333, QN => n21445);
   REGISTERS_reg_2_33_inst : DFF_X1 port map( D => n7907, CK => CLK, Q => 
                           n25332, QN => n21446);
   REGISTERS_reg_2_32_inst : DFF_X1 port map( D => n7906, CK => CLK, Q => 
                           n25331, QN => n21447);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n7905, CK => CLK, Q => 
                           n25330, QN => n21448);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n7904, CK => CLK, Q => 
                           n25329, QN => n21449);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n7903, CK => CLK, Q => 
                           n25328, QN => n21450);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n7902, CK => CLK, Q => 
                           n25327, QN => n21451);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n7901, CK => CLK, Q => 
                           n25326, QN => n21452);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n7900, CK => CLK, Q => 
                           n25325, QN => n21453);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n7899, CK => CLK, Q => 
                           n25324, QN => n21454);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n7898, CK => CLK, Q => 
                           n25323, QN => n21455);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n7897, CK => CLK, Q => 
                           n25322, QN => n21456);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n7896, CK => CLK, Q => 
                           n25321, QN => n21457);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n7895, CK => CLK, Q => 
                           n25320, QN => n21458);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n7894, CK => CLK, Q => 
                           n25319, QN => n21459);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n7893, CK => CLK, Q => 
                           n25318, QN => n21460);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n7892, CK => CLK, Q => 
                           n25317, QN => n21461);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n7891, CK => CLK, Q => 
                           n25316, QN => n21462);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n7890, CK => CLK, Q => 
                           n25315, QN => n21463);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n7889, CK => CLK, Q => 
                           n25314, QN => n21464);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n7888, CK => CLK, Q => 
                           n25313, QN => n21465);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n7887, CK => CLK, Q => 
                           n25312, QN => n21466);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n7886, CK => CLK, Q => 
                           n25311, QN => n21467);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n7885, CK => CLK, Q => 
                           n25654, QN => n21468);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n7884, CK => CLK, Q => 
                           n25653, QN => n21469);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n7883, CK => CLK, Q => n25652
                           , QN => n21470);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n7882, CK => CLK, Q => n25651
                           , QN => n21471);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n7881, CK => CLK, Q => n25650
                           , QN => n21472);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n7880, CK => CLK, Q => n25649
                           , QN => n21473);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n7879, CK => CLK, Q => n25648
                           , QN => n21474);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n7878, CK => CLK, Q => n25647
                           , QN => n21475);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n7877, CK => CLK, Q => n25646
                           , QN => n21476);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n7876, CK => CLK, Q => n25645
                           , QN => n21477);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n7875, CK => CLK, Q => n25644
                           , QN => n21478);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n7874, CK => CLK, Q => n25643
                           , QN => n21479);
   REGISTERS_reg_31_63_inst : DFF_X1 port map( D => n6081, CK => CLK, Q => 
                           n26194, QN => n20899);
   REGISTERS_reg_31_62_inst : DFF_X1 port map( D => n6080, CK => CLK, Q => 
                           n26193, QN => n20900);
   REGISTERS_reg_31_61_inst : DFF_X1 port map( D => n6079, CK => CLK, Q => 
                           n26192, QN => n20901);
   REGISTERS_reg_31_60_inst : DFF_X1 port map( D => n6078, CK => CLK, Q => 
                           n26191, QN => n20902);
   REGISTERS_reg_29_63_inst : DFF_X1 port map( D => n6209, CK => CLK, Q => 
                           n9249, QN => n22244);
   REGISTERS_reg_29_62_inst : DFF_X1 port map( D => n6208, CK => CLK, Q => 
                           n9252, QN => n22245);
   REGISTERS_reg_29_61_inst : DFF_X1 port map( D => n6207, CK => CLK, Q => 
                           n9255, QN => n22246);
   REGISTERS_reg_29_60_inst : DFF_X1 port map( D => n6206, CK => CLK, Q => 
                           n9258, QN => n22247);
   REGISTERS_reg_22_63_inst : DFF_X1 port map( D => n6657, CK => CLK, Q => 
                           n25695, QN => n21492);
   REGISTERS_reg_22_62_inst : DFF_X1 port map( D => n6656, CK => CLK, Q => 
                           n25690, QN => n21493);
   REGISTERS_reg_22_61_inst : DFF_X1 port map( D => n6655, CK => CLK, Q => 
                           n25685, QN => n21494);
   REGISTERS_reg_22_60_inst : DFF_X1 port map( D => n6654, CK => CLK, Q => 
                           n25680, QN => n21495);
   REGISTERS_reg_18_63_inst : DFF_X1 port map( D => n6913, CK => CLK, Q => 
                           n25696, QN => n21484);
   REGISTERS_reg_18_62_inst : DFF_X1 port map( D => n6912, CK => CLK, Q => 
                           n25691, QN => n21485);
   REGISTERS_reg_18_61_inst : DFF_X1 port map( D => n6911, CK => CLK, Q => 
                           n25686, QN => n21486);
   REGISTERS_reg_18_60_inst : DFF_X1 port map( D => n6910, CK => CLK, Q => 
                           n25681, QN => n21487);
   REGISTERS_reg_10_63_inst : DFF_X1 port map( D => n7425, CK => CLK, Q => 
                           n18382, QN => n22252);
   REGISTERS_reg_10_62_inst : DFF_X1 port map( D => n7424, CK => CLK, Q => 
                           n18399, QN => n22253);
   REGISTERS_reg_10_61_inst : DFF_X1 port map( D => n7423, CK => CLK, Q => 
                           n18416, QN => n22254);
   REGISTERS_reg_10_60_inst : DFF_X1 port map( D => n7422, CK => CLK, Q => 
                           n18433, QN => n22255);
   REGISTERS_reg_1_63_inst : DFF_X1 port map( D => n8001, CK => CLK, Q => 
                           n25578, QN => n21512);
   REGISTERS_reg_1_62_inst : DFF_X1 port map( D => n8000, CK => CLK, Q => 
                           n25577, QN => n21513);
   REGISTERS_reg_1_61_inst : DFF_X1 port map( D => n7999, CK => CLK, Q => 
                           n25576, QN => n21514);
   REGISTERS_reg_1_60_inst : DFF_X1 port map( D => n7998, CK => CLK, Q => 
                           n25575, QN => n21515);
   REGISTERS_reg_16_63_inst : DFF_X1 port map( D => n7041, CK => CLK, Q => 
                           n25697, QN => n21160);
   REGISTERS_reg_16_62_inst : DFF_X1 port map( D => n7040, CK => CLK, Q => 
                           n25692, QN => n21161);
   REGISTERS_reg_16_61_inst : DFF_X1 port map( D => n7039, CK => CLK, Q => 
                           n25687, QN => n21162);
   REGISTERS_reg_16_60_inst : DFF_X1 port map( D => n7038, CK => CLK, Q => 
                           n25682, QN => n21163);
   REGISTERS_reg_6_63_inst : DFF_X1 port map( D => n7681, CK => CLK, Q => 
                           n25558, QN => n21496);
   REGISTERS_reg_6_62_inst : DFF_X1 port map( D => n7680, CK => CLK, Q => 
                           n25557, QN => n21497);
   REGISTERS_reg_6_61_inst : DFF_X1 port map( D => n7679, CK => CLK, Q => 
                           n25556, QN => n21498);
   REGISTERS_reg_6_60_inst : DFF_X1 port map( D => n7678, CK => CLK, Q => 
                           n25555, QN => n21499);
   REGISTERS_reg_31_59_inst : DFF_X1 port map( D => n6077, CK => CLK, Q => 
                           n26266, QN => n20903);
   REGISTERS_reg_31_58_inst : DFF_X1 port map( D => n6076, CK => CLK, Q => 
                           n26265, QN => n20904);
   REGISTERS_reg_31_57_inst : DFF_X1 port map( D => n6075, CK => CLK, Q => 
                           n26264, QN => n20905);
   REGISTERS_reg_31_56_inst : DFF_X1 port map( D => n6074, CK => CLK, Q => 
                           n26263, QN => n20906);
   REGISTERS_reg_31_55_inst : DFF_X1 port map( D => n6073, CK => CLK, Q => 
                           n26262, QN => n20907);
   REGISTERS_reg_31_54_inst : DFF_X1 port map( D => n6072, CK => CLK, Q => 
                           n26261, QN => n20908);
   REGISTERS_reg_31_53_inst : DFF_X1 port map( D => n6071, CK => CLK, Q => 
                           n26260, QN => n20909);
   REGISTERS_reg_31_52_inst : DFF_X1 port map( D => n6070, CK => CLK, Q => 
                           n26259, QN => n20910);
   REGISTERS_reg_31_51_inst : DFF_X1 port map( D => n6069, CK => CLK, Q => 
                           n26258, QN => n20911);
   REGISTERS_reg_31_50_inst : DFF_X1 port map( D => n6068, CK => CLK, Q => 
                           n26257, QN => n20912);
   REGISTERS_reg_31_49_inst : DFF_X1 port map( D => n6067, CK => CLK, Q => 
                           n26256, QN => n20913);
   REGISTERS_reg_31_48_inst : DFF_X1 port map( D => n6066, CK => CLK, Q => 
                           n26255, QN => n20914);
   REGISTERS_reg_31_47_inst : DFF_X1 port map( D => n6065, CK => CLK, Q => 
                           n26254, QN => n20915);
   REGISTERS_reg_31_46_inst : DFF_X1 port map( D => n6064, CK => CLK, Q => 
                           n26253, QN => n20916);
   REGISTERS_reg_31_45_inst : DFF_X1 port map( D => n6063, CK => CLK, Q => 
                           n26252, QN => n20917);
   REGISTERS_reg_31_44_inst : DFF_X1 port map( D => n6062, CK => CLK, Q => 
                           n26251, QN => n20918);
   REGISTERS_reg_31_43_inst : DFF_X1 port map( D => n6061, CK => CLK, Q => 
                           n26250, QN => n20919);
   REGISTERS_reg_31_42_inst : DFF_X1 port map( D => n6060, CK => CLK, Q => 
                           n26249, QN => n20920);
   REGISTERS_reg_31_41_inst : DFF_X1 port map( D => n6059, CK => CLK, Q => 
                           n26248, QN => n20921);
   REGISTERS_reg_31_40_inst : DFF_X1 port map( D => n6058, CK => CLK, Q => 
                           n26247, QN => n20922);
   REGISTERS_reg_31_39_inst : DFF_X1 port map( D => n6057, CK => CLK, Q => 
                           n26246, QN => n20923);
   REGISTERS_reg_31_38_inst : DFF_X1 port map( D => n6056, CK => CLK, Q => 
                           n26245, QN => n20924);
   REGISTERS_reg_31_37_inst : DFF_X1 port map( D => n6055, CK => CLK, Q => 
                           n26244, QN => n20925);
   REGISTERS_reg_31_36_inst : DFF_X1 port map( D => n6054, CK => CLK, Q => 
                           n26243, QN => n20926);
   REGISTERS_reg_31_35_inst : DFF_X1 port map( D => n6053, CK => CLK, Q => 
                           n26242, QN => n20927);
   REGISTERS_reg_31_34_inst : DFF_X1 port map( D => n6052, CK => CLK, Q => 
                           n26241, QN => n20928);
   REGISTERS_reg_31_33_inst : DFF_X1 port map( D => n6051, CK => CLK, Q => 
                           n26240, QN => n20929);
   REGISTERS_reg_31_32_inst : DFF_X1 port map( D => n6050, CK => CLK, Q => 
                           n26239, QN => n20930);
   REGISTERS_reg_31_31_inst : DFF_X1 port map( D => n6049, CK => CLK, Q => 
                           n26238, QN => n20931);
   REGISTERS_reg_31_30_inst : DFF_X1 port map( D => n6048, CK => CLK, Q => 
                           n26237, QN => n20932);
   REGISTERS_reg_31_29_inst : DFF_X1 port map( D => n6047, CK => CLK, Q => 
                           n26236, QN => n20933);
   REGISTERS_reg_31_28_inst : DFF_X1 port map( D => n6046, CK => CLK, Q => 
                           n26235, QN => n20934);
   REGISTERS_reg_31_27_inst : DFF_X1 port map( D => n6045, CK => CLK, Q => 
                           n26234, QN => n20935);
   REGISTERS_reg_31_26_inst : DFF_X1 port map( D => n6044, CK => CLK, Q => 
                           n26233, QN => n20936);
   REGISTERS_reg_31_25_inst : DFF_X1 port map( D => n6043, CK => CLK, Q => 
                           n26232, QN => n20937);
   REGISTERS_reg_31_24_inst : DFF_X1 port map( D => n6042, CK => CLK, Q => 
                           n26231, QN => n20938);
   REGISTERS_reg_31_23_inst : DFF_X1 port map( D => n6041, CK => CLK, Q => 
                           n26230, QN => n20939);
   REGISTERS_reg_31_22_inst : DFF_X1 port map( D => n6040, CK => CLK, Q => 
                           n26229, QN => n20940);
   REGISTERS_reg_31_21_inst : DFF_X1 port map( D => n6039, CK => CLK, Q => 
                           n26228, QN => n20941);
   REGISTERS_reg_31_20_inst : DFF_X1 port map( D => n6038, CK => CLK, Q => 
                           n26227, QN => n20942);
   REGISTERS_reg_31_19_inst : DFF_X1 port map( D => n6037, CK => CLK, Q => 
                           n26226, QN => n20943);
   REGISTERS_reg_31_18_inst : DFF_X1 port map( D => n6036, CK => CLK, Q => 
                           n26225, QN => n20944);
   REGISTERS_reg_31_17_inst : DFF_X1 port map( D => n6035, CK => CLK, Q => 
                           n26224, QN => n20945);
   REGISTERS_reg_31_16_inst : DFF_X1 port map( D => n6034, CK => CLK, Q => 
                           n26223, QN => n20946);
   REGISTERS_reg_31_15_inst : DFF_X1 port map( D => n6033, CK => CLK, Q => 
                           n26222, QN => n20947);
   REGISTERS_reg_31_14_inst : DFF_X1 port map( D => n6032, CK => CLK, Q => 
                           n26221, QN => n20948);
   REGISTERS_reg_31_13_inst : DFF_X1 port map( D => n6031, CK => CLK, Q => 
                           n26220, QN => n20949);
   REGISTERS_reg_31_12_inst : DFF_X1 port map( D => n6030, CK => CLK, Q => 
                           n26219, QN => n20950);
   REGISTERS_reg_31_11_inst : DFF_X1 port map( D => n6029, CK => CLK, Q => 
                           n26218, QN => n20951);
   REGISTERS_reg_31_10_inst : DFF_X1 port map( D => n6028, CK => CLK, Q => 
                           n26217, QN => n20952);
   REGISTERS_reg_31_9_inst : DFF_X1 port map( D => n6027, CK => CLK, Q => 
                           n26216, QN => n20953);
   REGISTERS_reg_31_8_inst : DFF_X1 port map( D => n6026, CK => CLK, Q => 
                           n26215, QN => n20954);
   REGISTERS_reg_31_7_inst : DFF_X1 port map( D => n6025, CK => CLK, Q => 
                           n26214, QN => n20955);
   REGISTERS_reg_31_6_inst : DFF_X1 port map( D => n6024, CK => CLK, Q => 
                           n26213, QN => n20956);
   REGISTERS_reg_31_5_inst : DFF_X1 port map( D => n6023, CK => CLK, Q => 
                           n26212, QN => n20957);
   REGISTERS_reg_31_4_inst : DFF_X1 port map( D => n6022, CK => CLK, Q => 
                           n26211, QN => n20958);
   REGISTERS_reg_31_3_inst : DFF_X1 port map( D => n6021, CK => CLK, Q => 
                           n26210, QN => n20959);
   REGISTERS_reg_31_2_inst : DFF_X1 port map( D => n6020, CK => CLK, Q => 
                           n26209, QN => n20960);
   REGISTERS_reg_31_1_inst : DFF_X1 port map( D => n6019, CK => CLK, Q => 
                           n26208, QN => n20961);
   REGISTERS_reg_31_0_inst : DFF_X1 port map( D => n6018, CK => CLK, Q => 
                           n26207, QN => n20962);
   REGISTERS_reg_29_59_inst : DFF_X1 port map( D => n6205, CK => CLK, Q => 
                           n9261, QN => n22260);
   REGISTERS_reg_29_58_inst : DFF_X1 port map( D => n6204, CK => CLK, Q => 
                           n9264, QN => n22261);
   REGISTERS_reg_29_57_inst : DFF_X1 port map( D => n6203, CK => CLK, Q => 
                           n9267, QN => n22262);
   REGISTERS_reg_29_56_inst : DFF_X1 port map( D => n6202, CK => CLK, Q => 
                           n9270, QN => n22263);
   REGISTERS_reg_29_55_inst : DFF_X1 port map( D => n6201, CK => CLK, Q => 
                           n9273, QN => n22264);
   REGISTERS_reg_29_54_inst : DFF_X1 port map( D => n6200, CK => CLK, Q => 
                           n9276, QN => n22265);
   REGISTERS_reg_29_53_inst : DFF_X1 port map( D => n6199, CK => CLK, Q => 
                           n9279, QN => n22266);
   REGISTERS_reg_29_52_inst : DFF_X1 port map( D => n6198, CK => CLK, Q => 
                           n9282, QN => n22267);
   REGISTERS_reg_29_51_inst : DFF_X1 port map( D => n6197, CK => CLK, Q => 
                           n9285, QN => n22268);
   REGISTERS_reg_29_50_inst : DFF_X1 port map( D => n6196, CK => CLK, Q => 
                           n9288, QN => n22269);
   REGISTERS_reg_29_49_inst : DFF_X1 port map( D => n6195, CK => CLK, Q => 
                           n9291, QN => n22270);
   REGISTERS_reg_29_48_inst : DFF_X1 port map( D => n6194, CK => CLK, Q => 
                           n9294, QN => n22271);
   REGISTERS_reg_29_47_inst : DFF_X1 port map( D => n6193, CK => CLK, Q => 
                           n9297, QN => n22272);
   REGISTERS_reg_29_46_inst : DFF_X1 port map( D => n6192, CK => CLK, Q => 
                           n9300, QN => n22273);
   REGISTERS_reg_29_45_inst : DFF_X1 port map( D => n6191, CK => CLK, Q => 
                           n9303, QN => n22274);
   REGISTERS_reg_29_44_inst : DFF_X1 port map( D => n6190, CK => CLK, Q => 
                           n9306, QN => n22275);
   REGISTERS_reg_29_43_inst : DFF_X1 port map( D => n6189, CK => CLK, Q => 
                           n9309, QN => n22276);
   REGISTERS_reg_29_42_inst : DFF_X1 port map( D => n6188, CK => CLK, Q => 
                           n9312, QN => n22277);
   REGISTERS_reg_29_41_inst : DFF_X1 port map( D => n6187, CK => CLK, Q => 
                           n9315, QN => n22278);
   REGISTERS_reg_29_40_inst : DFF_X1 port map( D => n6186, CK => CLK, Q => 
                           n9318, QN => n22279);
   REGISTERS_reg_29_39_inst : DFF_X1 port map( D => n6185, CK => CLK, Q => 
                           n9321, QN => n22280);
   REGISTERS_reg_29_38_inst : DFF_X1 port map( D => n6184, CK => CLK, Q => 
                           n9324, QN => n22281);
   REGISTERS_reg_29_37_inst : DFF_X1 port map( D => n6183, CK => CLK, Q => 
                           n9327, QN => n22282);
   REGISTERS_reg_29_36_inst : DFF_X1 port map( D => n6182, CK => CLK, Q => 
                           n9330, QN => n22283);
   REGISTERS_reg_29_35_inst : DFF_X1 port map( D => n6181, CK => CLK, Q => 
                           n9333, QN => n22284);
   REGISTERS_reg_29_34_inst : DFF_X1 port map( D => n6180, CK => CLK, Q => 
                           n9336, QN => n22285);
   REGISTERS_reg_29_33_inst : DFF_X1 port map( D => n6179, CK => CLK, Q => 
                           n9339, QN => n22286);
   REGISTERS_reg_29_32_inst : DFF_X1 port map( D => n6178, CK => CLK, Q => 
                           n9342, QN => n22287);
   REGISTERS_reg_29_31_inst : DFF_X1 port map( D => n6177, CK => CLK, Q => 
                           n9345, QN => n22288);
   REGISTERS_reg_29_30_inst : DFF_X1 port map( D => n6176, CK => CLK, Q => 
                           n9348, QN => n22289);
   REGISTERS_reg_29_29_inst : DFF_X1 port map( D => n6175, CK => CLK, Q => 
                           n9351, QN => n22290);
   REGISTERS_reg_29_28_inst : DFF_X1 port map( D => n6174, CK => CLK, Q => 
                           n9354, QN => n22291);
   REGISTERS_reg_29_27_inst : DFF_X1 port map( D => n6173, CK => CLK, Q => 
                           n9357, QN => n22292);
   REGISTERS_reg_29_26_inst : DFF_X1 port map( D => n6172, CK => CLK, Q => 
                           n9360, QN => n22293);
   REGISTERS_reg_29_25_inst : DFF_X1 port map( D => n6171, CK => CLK, Q => 
                           n9363, QN => n22294);
   REGISTERS_reg_29_24_inst : DFF_X1 port map( D => n6170, CK => CLK, Q => 
                           n9366, QN => n22295);
   REGISTERS_reg_29_23_inst : DFF_X1 port map( D => n6169, CK => CLK, Q => 
                           n9369, QN => n22296);
   REGISTERS_reg_29_22_inst : DFF_X1 port map( D => n6168, CK => CLK, Q => 
                           n9372, QN => n22297);
   REGISTERS_reg_29_21_inst : DFF_X1 port map( D => n6167, CK => CLK, Q => 
                           n9375, QN => n22298);
   REGISTERS_reg_29_20_inst : DFF_X1 port map( D => n6166, CK => CLK, Q => 
                           n9378, QN => n22299);
   REGISTERS_reg_29_19_inst : DFF_X1 port map( D => n6165, CK => CLK, Q => 
                           n9381, QN => n22300);
   REGISTERS_reg_29_18_inst : DFF_X1 port map( D => n6164, CK => CLK, Q => 
                           n9384, QN => n22301);
   REGISTERS_reg_29_17_inst : DFF_X1 port map( D => n6163, CK => CLK, Q => 
                           n9387, QN => n22302);
   REGISTERS_reg_29_16_inst : DFF_X1 port map( D => n6162, CK => CLK, Q => 
                           n9390, QN => n22303);
   REGISTERS_reg_29_15_inst : DFF_X1 port map( D => n6161, CK => CLK, Q => 
                           n9393, QN => n22304);
   REGISTERS_reg_29_14_inst : DFF_X1 port map( D => n6160, CK => CLK, Q => 
                           n9396, QN => n22305);
   REGISTERS_reg_29_13_inst : DFF_X1 port map( D => n6159, CK => CLK, Q => 
                           n9399, QN => n22306);
   REGISTERS_reg_29_12_inst : DFF_X1 port map( D => n6158, CK => CLK, Q => 
                           n9402, QN => n22307);
   REGISTERS_reg_29_11_inst : DFF_X1 port map( D => n6157, CK => CLK, Q => 
                           n9405, QN => n22308);
   REGISTERS_reg_29_10_inst : DFF_X1 port map( D => n6156, CK => CLK, Q => 
                           n9408, QN => n22309);
   REGISTERS_reg_29_9_inst : DFF_X1 port map( D => n6155, CK => CLK, Q => n9411
                           , QN => n22310);
   REGISTERS_reg_29_8_inst : DFF_X1 port map( D => n6154, CK => CLK, Q => n9414
                           , QN => n22311);
   REGISTERS_reg_29_7_inst : DFF_X1 port map( D => n6153, CK => CLK, Q => n9417
                           , QN => n22312);
   REGISTERS_reg_29_6_inst : DFF_X1 port map( D => n6152, CK => CLK, Q => n9420
                           , QN => n22313);
   REGISTERS_reg_29_5_inst : DFF_X1 port map( D => n6151, CK => CLK, Q => n9423
                           , QN => n22314);
   REGISTERS_reg_29_4_inst : DFF_X1 port map( D => n6150, CK => CLK, Q => n9426
                           , QN => n22315);
   REGISTERS_reg_29_3_inst : DFF_X1 port map( D => n6149, CK => CLK, Q => n9429
                           , QN => n22316);
   REGISTERS_reg_29_2_inst : DFF_X1 port map( D => n6148, CK => CLK, Q => n9432
                           , QN => n22317);
   REGISTERS_reg_29_1_inst : DFF_X1 port map( D => n6147, CK => CLK, Q => n9435
                           , QN => n22318);
   REGISTERS_reg_29_0_inst : DFF_X1 port map( D => n6146, CK => CLK, Q => n9438
                           , QN => n22319);
   REGISTERS_reg_22_59_inst : DFF_X1 port map( D => n6653, CK => CLK, Q => 
                           n25995, QN => n21760);
   REGISTERS_reg_22_58_inst : DFF_X1 port map( D => n6652, CK => CLK, Q => 
                           n25990, QN => n21761);
   REGISTERS_reg_22_57_inst : DFF_X1 port map( D => n6651, CK => CLK, Q => 
                           n25985, QN => n21762);
   REGISTERS_reg_22_56_inst : DFF_X1 port map( D => n6650, CK => CLK, Q => 
                           n25980, QN => n21763);
   REGISTERS_reg_22_55_inst : DFF_X1 port map( D => n6649, CK => CLK, Q => 
                           n25975, QN => n21764);
   REGISTERS_reg_22_54_inst : DFF_X1 port map( D => n6648, CK => CLK, Q => 
                           n25970, QN => n21765);
   REGISTERS_reg_22_53_inst : DFF_X1 port map( D => n6647, CK => CLK, Q => 
                           n25965, QN => n21766);
   REGISTERS_reg_22_52_inst : DFF_X1 port map( D => n6646, CK => CLK, Q => 
                           n25960, QN => n21767);
   REGISTERS_reg_22_51_inst : DFF_X1 port map( D => n6645, CK => CLK, Q => 
                           n25955, QN => n21768);
   REGISTERS_reg_22_50_inst : DFF_X1 port map( D => n6644, CK => CLK, Q => 
                           n25950, QN => n21769);
   REGISTERS_reg_22_49_inst : DFF_X1 port map( D => n6643, CK => CLK, Q => 
                           n25945, QN => n21770);
   REGISTERS_reg_22_48_inst : DFF_X1 port map( D => n6642, CK => CLK, Q => 
                           n25940, QN => n21771);
   REGISTERS_reg_22_47_inst : DFF_X1 port map( D => n6641, CK => CLK, Q => 
                           n25935, QN => n21772);
   REGISTERS_reg_22_46_inst : DFF_X1 port map( D => n6640, CK => CLK, Q => 
                           n25930, QN => n21773);
   REGISTERS_reg_22_45_inst : DFF_X1 port map( D => n6639, CK => CLK, Q => 
                           n25925, QN => n21774);
   REGISTERS_reg_22_44_inst : DFF_X1 port map( D => n6638, CK => CLK, Q => 
                           n25920, QN => n21775);
   REGISTERS_reg_22_43_inst : DFF_X1 port map( D => n6637, CK => CLK, Q => 
                           n25915, QN => n21776);
   REGISTERS_reg_22_42_inst : DFF_X1 port map( D => n6636, CK => CLK, Q => 
                           n25910, QN => n21777);
   REGISTERS_reg_22_41_inst : DFF_X1 port map( D => n6635, CK => CLK, Q => 
                           n25905, QN => n21778);
   REGISTERS_reg_22_40_inst : DFF_X1 port map( D => n6634, CK => CLK, Q => 
                           n25900, QN => n21779);
   REGISTERS_reg_22_39_inst : DFF_X1 port map( D => n6633, CK => CLK, Q => 
                           n25895, QN => n21780);
   REGISTERS_reg_22_38_inst : DFF_X1 port map( D => n6632, CK => CLK, Q => 
                           n25890, QN => n21781);
   REGISTERS_reg_22_37_inst : DFF_X1 port map( D => n6631, CK => CLK, Q => 
                           n25885, QN => n21782);
   REGISTERS_reg_22_36_inst : DFF_X1 port map( D => n6630, CK => CLK, Q => 
                           n25880, QN => n21783);
   REGISTERS_reg_22_35_inst : DFF_X1 port map( D => n6629, CK => CLK, Q => 
                           n25875, QN => n21784);
   REGISTERS_reg_22_34_inst : DFF_X1 port map( D => n6628, CK => CLK, Q => 
                           n25870, QN => n21785);
   REGISTERS_reg_22_33_inst : DFF_X1 port map( D => n6627, CK => CLK, Q => 
                           n25865, QN => n21786);
   REGISTERS_reg_22_32_inst : DFF_X1 port map( D => n6626, CK => CLK, Q => 
                           n25860, QN => n21787);
   REGISTERS_reg_22_31_inst : DFF_X1 port map( D => n6625, CK => CLK, Q => 
                           n25855, QN => n21788);
   REGISTERS_reg_22_30_inst : DFF_X1 port map( D => n6624, CK => CLK, Q => 
                           n25850, QN => n21789);
   REGISTERS_reg_22_29_inst : DFF_X1 port map( D => n6623, CK => CLK, Q => 
                           n25845, QN => n21790);
   REGISTERS_reg_22_28_inst : DFF_X1 port map( D => n6622, CK => CLK, Q => 
                           n25840, QN => n21791);
   REGISTERS_reg_22_27_inst : DFF_X1 port map( D => n6621, CK => CLK, Q => 
                           n25835, QN => n21792);
   REGISTERS_reg_22_26_inst : DFF_X1 port map( D => n6620, CK => CLK, Q => 
                           n25830, QN => n21793);
   REGISTERS_reg_22_25_inst : DFF_X1 port map( D => n6619, CK => CLK, Q => 
                           n25825, QN => n21794);
   REGISTERS_reg_22_24_inst : DFF_X1 port map( D => n6618, CK => CLK, Q => 
                           n25820, QN => n21795);
   REGISTERS_reg_22_23_inst : DFF_X1 port map( D => n6617, CK => CLK, Q => 
                           n25815, QN => n21796);
   REGISTERS_reg_22_22_inst : DFF_X1 port map( D => n6616, CK => CLK, Q => 
                           n25810, QN => n21797);
   REGISTERS_reg_22_21_inst : DFF_X1 port map( D => n6615, CK => CLK, Q => 
                           n25805, QN => n21798);
   REGISTERS_reg_22_20_inst : DFF_X1 port map( D => n6614, CK => CLK, Q => 
                           n25800, QN => n21799);
   REGISTERS_reg_22_19_inst : DFF_X1 port map( D => n6613, CK => CLK, Q => 
                           n25795, QN => n21800);
   REGISTERS_reg_22_18_inst : DFF_X1 port map( D => n6612, CK => CLK, Q => 
                           n25790, QN => n21801);
   REGISTERS_reg_22_17_inst : DFF_X1 port map( D => n6611, CK => CLK, Q => 
                           n25785, QN => n21802);
   REGISTERS_reg_22_16_inst : DFF_X1 port map( D => n6610, CK => CLK, Q => 
                           n25780, QN => n21803);
   REGISTERS_reg_22_15_inst : DFF_X1 port map( D => n6609, CK => CLK, Q => 
                           n25775, QN => n21804);
   REGISTERS_reg_22_14_inst : DFF_X1 port map( D => n6608, CK => CLK, Q => 
                           n25770, QN => n21805);
   REGISTERS_reg_22_13_inst : DFF_X1 port map( D => n6607, CK => CLK, Q => 
                           n25765, QN => n21806);
   REGISTERS_reg_22_12_inst : DFF_X1 port map( D => n6606, CK => CLK, Q => 
                           n25760, QN => n21807);
   REGISTERS_reg_22_11_inst : DFF_X1 port map( D => n6605, CK => CLK, Q => 
                           n25755, QN => n21808);
   REGISTERS_reg_22_10_inst : DFF_X1 port map( D => n6604, CK => CLK, Q => 
                           n25750, QN => n21809);
   REGISTERS_reg_22_9_inst : DFF_X1 port map( D => n6603, CK => CLK, Q => 
                           n25745, QN => n21810);
   REGISTERS_reg_22_8_inst : DFF_X1 port map( D => n6602, CK => CLK, Q => 
                           n25740, QN => n21811);
   REGISTERS_reg_22_7_inst : DFF_X1 port map( D => n6601, CK => CLK, Q => 
                           n25735, QN => n21812);
   REGISTERS_reg_22_6_inst : DFF_X1 port map( D => n6600, CK => CLK, Q => 
                           n25730, QN => n21813);
   REGISTERS_reg_22_5_inst : DFF_X1 port map( D => n6599, CK => CLK, Q => 
                           n25725, QN => n21814);
   REGISTERS_reg_22_4_inst : DFF_X1 port map( D => n6598, CK => CLK, Q => 
                           n25720, QN => n21815);
   REGISTERS_reg_22_3_inst : DFF_X1 port map( D => n6597, CK => CLK, Q => 
                           n25715, QN => n21816);
   REGISTERS_reg_22_2_inst : DFF_X1 port map( D => n6596, CK => CLK, Q => 
                           n25710, QN => n21817);
   REGISTERS_reg_22_1_inst : DFF_X1 port map( D => n6595, CK => CLK, Q => 
                           n25705, QN => n21818);
   REGISTERS_reg_22_0_inst : DFF_X1 port map( D => n6594, CK => CLK, Q => 
                           n25700, QN => n21819);
   REGISTERS_reg_18_59_inst : DFF_X1 port map( D => n6909, CK => CLK, Q => 
                           n25996, QN => n21640);
   REGISTERS_reg_18_58_inst : DFF_X1 port map( D => n6908, CK => CLK, Q => 
                           n25991, QN => n21641);
   REGISTERS_reg_18_57_inst : DFF_X1 port map( D => n6907, CK => CLK, Q => 
                           n25986, QN => n21642);
   REGISTERS_reg_18_56_inst : DFF_X1 port map( D => n6906, CK => CLK, Q => 
                           n25981, QN => n21643);
   REGISTERS_reg_18_55_inst : DFF_X1 port map( D => n6905, CK => CLK, Q => 
                           n25976, QN => n21644);
   REGISTERS_reg_18_54_inst : DFF_X1 port map( D => n6904, CK => CLK, Q => 
                           n25971, QN => n21645);
   REGISTERS_reg_18_53_inst : DFF_X1 port map( D => n6903, CK => CLK, Q => 
                           n25966, QN => n21646);
   REGISTERS_reg_18_52_inst : DFF_X1 port map( D => n6902, CK => CLK, Q => 
                           n25961, QN => n21647);
   REGISTERS_reg_18_51_inst : DFF_X1 port map( D => n6901, CK => CLK, Q => 
                           n25956, QN => n21648);
   REGISTERS_reg_18_50_inst : DFF_X1 port map( D => n6900, CK => CLK, Q => 
                           n25951, QN => n21649);
   REGISTERS_reg_18_49_inst : DFF_X1 port map( D => n6899, CK => CLK, Q => 
                           n25946, QN => n21650);
   REGISTERS_reg_18_48_inst : DFF_X1 port map( D => n6898, CK => CLK, Q => 
                           n25941, QN => n21651);
   REGISTERS_reg_18_47_inst : DFF_X1 port map( D => n6897, CK => CLK, Q => 
                           n25936, QN => n21652);
   REGISTERS_reg_18_46_inst : DFF_X1 port map( D => n6896, CK => CLK, Q => 
                           n25931, QN => n21653);
   REGISTERS_reg_18_45_inst : DFF_X1 port map( D => n6895, CK => CLK, Q => 
                           n25926, QN => n21654);
   REGISTERS_reg_18_44_inst : DFF_X1 port map( D => n6894, CK => CLK, Q => 
                           n25921, QN => n21655);
   REGISTERS_reg_18_43_inst : DFF_X1 port map( D => n6893, CK => CLK, Q => 
                           n25916, QN => n21656);
   REGISTERS_reg_18_42_inst : DFF_X1 port map( D => n6892, CK => CLK, Q => 
                           n25911, QN => n21657);
   REGISTERS_reg_18_41_inst : DFF_X1 port map( D => n6891, CK => CLK, Q => 
                           n25906, QN => n21658);
   REGISTERS_reg_18_40_inst : DFF_X1 port map( D => n6890, CK => CLK, Q => 
                           n25901, QN => n21659);
   REGISTERS_reg_18_39_inst : DFF_X1 port map( D => n6889, CK => CLK, Q => 
                           n25896, QN => n21660);
   REGISTERS_reg_18_38_inst : DFF_X1 port map( D => n6888, CK => CLK, Q => 
                           n25891, QN => n21661);
   REGISTERS_reg_18_37_inst : DFF_X1 port map( D => n6887, CK => CLK, Q => 
                           n25886, QN => n21662);
   REGISTERS_reg_18_36_inst : DFF_X1 port map( D => n6886, CK => CLK, Q => 
                           n25881, QN => n21663);
   REGISTERS_reg_18_35_inst : DFF_X1 port map( D => n6885, CK => CLK, Q => 
                           n25876, QN => n21664);
   REGISTERS_reg_18_34_inst : DFF_X1 port map( D => n6884, CK => CLK, Q => 
                           n25871, QN => n21665);
   REGISTERS_reg_18_33_inst : DFF_X1 port map( D => n6883, CK => CLK, Q => 
                           n25866, QN => n21666);
   REGISTERS_reg_18_32_inst : DFF_X1 port map( D => n6882, CK => CLK, Q => 
                           n25861, QN => n21667);
   REGISTERS_reg_18_31_inst : DFF_X1 port map( D => n6881, CK => CLK, Q => 
                           n25856, QN => n21668);
   REGISTERS_reg_18_30_inst : DFF_X1 port map( D => n6880, CK => CLK, Q => 
                           n25851, QN => n21669);
   REGISTERS_reg_18_29_inst : DFF_X1 port map( D => n6879, CK => CLK, Q => 
                           n25846, QN => n21670);
   REGISTERS_reg_18_28_inst : DFF_X1 port map( D => n6878, CK => CLK, Q => 
                           n25841, QN => n21671);
   REGISTERS_reg_18_27_inst : DFF_X1 port map( D => n6877, CK => CLK, Q => 
                           n25836, QN => n21672);
   REGISTERS_reg_18_26_inst : DFF_X1 port map( D => n6876, CK => CLK, Q => 
                           n25831, QN => n21673);
   REGISTERS_reg_18_25_inst : DFF_X1 port map( D => n6875, CK => CLK, Q => 
                           n25826, QN => n21674);
   REGISTERS_reg_18_24_inst : DFF_X1 port map( D => n6874, CK => CLK, Q => 
                           n25821, QN => n21675);
   REGISTERS_reg_18_23_inst : DFF_X1 port map( D => n6873, CK => CLK, Q => 
                           n25816, QN => n21676);
   REGISTERS_reg_18_22_inst : DFF_X1 port map( D => n6872, CK => CLK, Q => 
                           n25811, QN => n21677);
   REGISTERS_reg_18_21_inst : DFF_X1 port map( D => n6871, CK => CLK, Q => 
                           n25806, QN => n21678);
   REGISTERS_reg_18_20_inst : DFF_X1 port map( D => n6870, CK => CLK, Q => 
                           n25801, QN => n21679);
   REGISTERS_reg_18_19_inst : DFF_X1 port map( D => n6869, CK => CLK, Q => 
                           n25796, QN => n21680);
   REGISTERS_reg_18_18_inst : DFF_X1 port map( D => n6868, CK => CLK, Q => 
                           n25791, QN => n21681);
   REGISTERS_reg_18_17_inst : DFF_X1 port map( D => n6867, CK => CLK, Q => 
                           n25786, QN => n21682);
   REGISTERS_reg_18_16_inst : DFF_X1 port map( D => n6866, CK => CLK, Q => 
                           n25781, QN => n21683);
   REGISTERS_reg_18_15_inst : DFF_X1 port map( D => n6865, CK => CLK, Q => 
                           n25776, QN => n21684);
   REGISTERS_reg_18_14_inst : DFF_X1 port map( D => n6864, CK => CLK, Q => 
                           n25771, QN => n21685);
   REGISTERS_reg_18_13_inst : DFF_X1 port map( D => n6863, CK => CLK, Q => 
                           n25766, QN => n21686);
   REGISTERS_reg_18_12_inst : DFF_X1 port map( D => n6862, CK => CLK, Q => 
                           n25761, QN => n21687);
   REGISTERS_reg_18_11_inst : DFF_X1 port map( D => n6861, CK => CLK, Q => 
                           n25756, QN => n21688);
   REGISTERS_reg_18_10_inst : DFF_X1 port map( D => n6860, CK => CLK, Q => 
                           n25751, QN => n21689);
   REGISTERS_reg_18_9_inst : DFF_X1 port map( D => n6859, CK => CLK, Q => 
                           n25746, QN => n21690);
   REGISTERS_reg_18_8_inst : DFF_X1 port map( D => n6858, CK => CLK, Q => 
                           n25741, QN => n21691);
   REGISTERS_reg_18_7_inst : DFF_X1 port map( D => n6857, CK => CLK, Q => 
                           n25736, QN => n21692);
   REGISTERS_reg_18_6_inst : DFF_X1 port map( D => n6856, CK => CLK, Q => 
                           n25731, QN => n21693);
   REGISTERS_reg_18_5_inst : DFF_X1 port map( D => n6855, CK => CLK, Q => 
                           n25726, QN => n21694);
   REGISTERS_reg_18_4_inst : DFF_X1 port map( D => n6854, CK => CLK, Q => 
                           n25721, QN => n21695);
   REGISTERS_reg_18_3_inst : DFF_X1 port map( D => n6853, CK => CLK, Q => 
                           n25716, QN => n21696);
   REGISTERS_reg_18_2_inst : DFF_X1 port map( D => n6852, CK => CLK, Q => 
                           n25711, QN => n21697);
   REGISTERS_reg_18_1_inst : DFF_X1 port map( D => n6851, CK => CLK, Q => 
                           n25706, QN => n21698);
   REGISTERS_reg_18_0_inst : DFF_X1 port map( D => n6850, CK => CLK, Q => 
                           n25701, QN => n21699);
   REGISTERS_reg_10_59_inst : DFF_X1 port map( D => n7421, CK => CLK, Q => 
                           n18450, QN => n22380);
   REGISTERS_reg_10_58_inst : DFF_X1 port map( D => n7420, CK => CLK, Q => 
                           n18467, QN => n22381);
   REGISTERS_reg_10_57_inst : DFF_X1 port map( D => n7419, CK => CLK, Q => 
                           n18484, QN => n22382);
   REGISTERS_reg_10_56_inst : DFF_X1 port map( D => n7418, CK => CLK, Q => 
                           n18501, QN => n22383);
   REGISTERS_reg_10_55_inst : DFF_X1 port map( D => n7417, CK => CLK, Q => 
                           n18518, QN => n22384);
   REGISTERS_reg_10_54_inst : DFF_X1 port map( D => n7416, CK => CLK, Q => 
                           n18535, QN => n22385);
   REGISTERS_reg_10_53_inst : DFF_X1 port map( D => n7415, CK => CLK, Q => 
                           n18552, QN => n22386);
   REGISTERS_reg_10_52_inst : DFF_X1 port map( D => n7414, CK => CLK, Q => 
                           n18569, QN => n22387);
   REGISTERS_reg_10_51_inst : DFF_X1 port map( D => n7413, CK => CLK, Q => 
                           n18586, QN => n22388);
   REGISTERS_reg_10_50_inst : DFF_X1 port map( D => n7412, CK => CLK, Q => 
                           n18603, QN => n22389);
   REGISTERS_reg_10_49_inst : DFF_X1 port map( D => n7411, CK => CLK, Q => 
                           n18620, QN => n22390);
   REGISTERS_reg_10_48_inst : DFF_X1 port map( D => n7410, CK => CLK, Q => 
                           n18637, QN => n22391);
   REGISTERS_reg_10_47_inst : DFF_X1 port map( D => n7409, CK => CLK, Q => 
                           n18654, QN => n22392);
   REGISTERS_reg_10_46_inst : DFF_X1 port map( D => n7408, CK => CLK, Q => 
                           n18671, QN => n22393);
   REGISTERS_reg_10_45_inst : DFF_X1 port map( D => n7407, CK => CLK, Q => 
                           n18688, QN => n22394);
   REGISTERS_reg_10_44_inst : DFF_X1 port map( D => n7406, CK => CLK, Q => 
                           n18705, QN => n22395);
   REGISTERS_reg_10_43_inst : DFF_X1 port map( D => n7405, CK => CLK, Q => 
                           n18722, QN => n22396);
   REGISTERS_reg_10_42_inst : DFF_X1 port map( D => n7404, CK => CLK, Q => 
                           n18739, QN => n22397);
   REGISTERS_reg_10_41_inst : DFF_X1 port map( D => n7403, CK => CLK, Q => 
                           n18756, QN => n22398);
   REGISTERS_reg_10_40_inst : DFF_X1 port map( D => n7402, CK => CLK, Q => 
                           n18773, QN => n22399);
   REGISTERS_reg_10_39_inst : DFF_X1 port map( D => n7401, CK => CLK, Q => 
                           n18790, QN => n22400);
   REGISTERS_reg_10_38_inst : DFF_X1 port map( D => n7400, CK => CLK, Q => 
                           n18807, QN => n22401);
   REGISTERS_reg_10_37_inst : DFF_X1 port map( D => n7399, CK => CLK, Q => 
                           n18824, QN => n22402);
   REGISTERS_reg_10_36_inst : DFF_X1 port map( D => n7398, CK => CLK, Q => 
                           n18841, QN => n22403);
   REGISTERS_reg_10_35_inst : DFF_X1 port map( D => n7397, CK => CLK, Q => 
                           n18858, QN => n22404);
   REGISTERS_reg_10_34_inst : DFF_X1 port map( D => n7396, CK => CLK, Q => 
                           n18875, QN => n22405);
   REGISTERS_reg_10_33_inst : DFF_X1 port map( D => n7395, CK => CLK, Q => 
                           n18892, QN => n22406);
   REGISTERS_reg_10_32_inst : DFF_X1 port map( D => n7394, CK => CLK, Q => 
                           n18909, QN => n22407);
   REGISTERS_reg_10_31_inst : DFF_X1 port map( D => n7393, CK => CLK, Q => 
                           n18926, QN => n22408);
   REGISTERS_reg_10_30_inst : DFF_X1 port map( D => n7392, CK => CLK, Q => 
                           n18943, QN => n22409);
   REGISTERS_reg_10_29_inst : DFF_X1 port map( D => n7391, CK => CLK, Q => 
                           n18960, QN => n22410);
   REGISTERS_reg_10_28_inst : DFF_X1 port map( D => n7390, CK => CLK, Q => 
                           n18977, QN => n22411);
   REGISTERS_reg_10_27_inst : DFF_X1 port map( D => n7389, CK => CLK, Q => 
                           n18994, QN => n22412);
   REGISTERS_reg_10_26_inst : DFF_X1 port map( D => n7388, CK => CLK, Q => 
                           n19011, QN => n22413);
   REGISTERS_reg_10_25_inst : DFF_X1 port map( D => n7387, CK => CLK, Q => 
                           n19028, QN => n22414);
   REGISTERS_reg_10_24_inst : DFF_X1 port map( D => n7386, CK => CLK, Q => 
                           n19045, QN => n22415);
   REGISTERS_reg_10_23_inst : DFF_X1 port map( D => n7385, CK => CLK, Q => 
                           n19062, QN => n22416);
   REGISTERS_reg_10_22_inst : DFF_X1 port map( D => n7384, CK => CLK, Q => 
                           n19079, QN => n22417);
   REGISTERS_reg_10_21_inst : DFF_X1 port map( D => n7383, CK => CLK, Q => 
                           n19096, QN => n22418);
   REGISTERS_reg_10_20_inst : DFF_X1 port map( D => n7382, CK => CLK, Q => 
                           n19113, QN => n22419);
   REGISTERS_reg_10_19_inst : DFF_X1 port map( D => n7381, CK => CLK, Q => 
                           n19130, QN => n22420);
   REGISTERS_reg_10_18_inst : DFF_X1 port map( D => n7380, CK => CLK, Q => 
                           n19147, QN => n22421);
   REGISTERS_reg_10_17_inst : DFF_X1 port map( D => n7379, CK => CLK, Q => 
                           n19164, QN => n22422);
   REGISTERS_reg_10_16_inst : DFF_X1 port map( D => n7378, CK => CLK, Q => 
                           n19181, QN => n22423);
   REGISTERS_reg_10_15_inst : DFF_X1 port map( D => n7377, CK => CLK, Q => 
                           n19198, QN => n22424);
   REGISTERS_reg_10_14_inst : DFF_X1 port map( D => n7376, CK => CLK, Q => 
                           n19215, QN => n22425);
   REGISTERS_reg_10_13_inst : DFF_X1 port map( D => n7375, CK => CLK, Q => 
                           n19232, QN => n22426);
   REGISTERS_reg_10_12_inst : DFF_X1 port map( D => n7374, CK => CLK, Q => 
                           n19249, QN => n22427);
   REGISTERS_reg_10_11_inst : DFF_X1 port map( D => n7373, CK => CLK, Q => 
                           n19266, QN => n22428);
   REGISTERS_reg_10_10_inst : DFF_X1 port map( D => n7372, CK => CLK, Q => 
                           n19283, QN => n22429);
   REGISTERS_reg_10_9_inst : DFF_X1 port map( D => n7371, CK => CLK, Q => 
                           n19300, QN => n22430);
   REGISTERS_reg_10_8_inst : DFF_X1 port map( D => n7370, CK => CLK, Q => 
                           n19317, QN => n22431);
   REGISTERS_reg_10_7_inst : DFF_X1 port map( D => n7369, CK => CLK, Q => 
                           n19334, QN => n22432);
   REGISTERS_reg_10_6_inst : DFF_X1 port map( D => n7368, CK => CLK, Q => 
                           n19351, QN => n22433);
   REGISTERS_reg_10_5_inst : DFF_X1 port map( D => n7367, CK => CLK, Q => 
                           n19368, QN => n22434);
   REGISTERS_reg_10_4_inst : DFF_X1 port map( D => n7366, CK => CLK, Q => 
                           n19385, QN => n22435);
   REGISTERS_reg_10_3_inst : DFF_X1 port map( D => n7365, CK => CLK, Q => 
                           n19402, QN => n22436);
   REGISTERS_reg_10_2_inst : DFF_X1 port map( D => n7364, CK => CLK, Q => 
                           n19419, QN => n22437);
   REGISTERS_reg_10_1_inst : DFF_X1 port map( D => n7363, CK => CLK, Q => 
                           n19436, QN => n22438);
   REGISTERS_reg_10_0_inst : DFF_X1 port map( D => n7362, CK => CLK, Q => 
                           n19453, QN => n22439);
   REGISTERS_reg_1_59_inst : DFF_X1 port map( D => n7997, CK => CLK, Q => 
                           n25502, QN => n22060);
   REGISTERS_reg_1_58_inst : DFF_X1 port map( D => n7996, CK => CLK, Q => 
                           n25501, QN => n22061);
   REGISTERS_reg_1_57_inst : DFF_X1 port map( D => n7995, CK => CLK, Q => 
                           n25500, QN => n22062);
   REGISTERS_reg_1_56_inst : DFF_X1 port map( D => n7994, CK => CLK, Q => 
                           n25499, QN => n22063);
   REGISTERS_reg_1_55_inst : DFF_X1 port map( D => n7993, CK => CLK, Q => 
                           n25498, QN => n22064);
   REGISTERS_reg_1_54_inst : DFF_X1 port map( D => n7992, CK => CLK, Q => 
                           n25497, QN => n22065);
   REGISTERS_reg_1_53_inst : DFF_X1 port map( D => n7991, CK => CLK, Q => 
                           n25496, QN => n22066);
   REGISTERS_reg_1_52_inst : DFF_X1 port map( D => n7990, CK => CLK, Q => 
                           n25495, QN => n22067);
   REGISTERS_reg_1_51_inst : DFF_X1 port map( D => n7989, CK => CLK, Q => 
                           n25494, QN => n22068);
   REGISTERS_reg_1_50_inst : DFF_X1 port map( D => n7988, CK => CLK, Q => 
                           n25493, QN => n22069);
   REGISTERS_reg_1_49_inst : DFF_X1 port map( D => n7987, CK => CLK, Q => 
                           n25492, QN => n22070);
   REGISTERS_reg_1_48_inst : DFF_X1 port map( D => n7986, CK => CLK, Q => 
                           n25491, QN => n22071);
   REGISTERS_reg_1_47_inst : DFF_X1 port map( D => n7985, CK => CLK, Q => 
                           n25490, QN => n22072);
   REGISTERS_reg_1_46_inst : DFF_X1 port map( D => n7984, CK => CLK, Q => 
                           n25489, QN => n22073);
   REGISTERS_reg_1_45_inst : DFF_X1 port map( D => n7983, CK => CLK, Q => 
                           n25488, QN => n22074);
   REGISTERS_reg_1_44_inst : DFF_X1 port map( D => n7982, CK => CLK, Q => 
                           n25487, QN => n22075);
   REGISTERS_reg_1_43_inst : DFF_X1 port map( D => n7981, CK => CLK, Q => 
                           n25486, QN => n22076);
   REGISTERS_reg_1_42_inst : DFF_X1 port map( D => n7980, CK => CLK, Q => 
                           n25485, QN => n22077);
   REGISTERS_reg_1_41_inst : DFF_X1 port map( D => n7979, CK => CLK, Q => 
                           n25484, QN => n22078);
   REGISTERS_reg_1_40_inst : DFF_X1 port map( D => n7978, CK => CLK, Q => 
                           n25483, QN => n22079);
   REGISTERS_reg_1_39_inst : DFF_X1 port map( D => n7977, CK => CLK, Q => 
                           n25482, QN => n22080);
   REGISTERS_reg_1_38_inst : DFF_X1 port map( D => n7976, CK => CLK, Q => 
                           n25481, QN => n22081);
   REGISTERS_reg_1_37_inst : DFF_X1 port map( D => n7975, CK => CLK, Q => 
                           n25480, QN => n22082);
   REGISTERS_reg_1_36_inst : DFF_X1 port map( D => n7974, CK => CLK, Q => 
                           n25479, QN => n22083);
   REGISTERS_reg_1_35_inst : DFF_X1 port map( D => n7973, CK => CLK, Q => 
                           n25478, QN => n22084);
   REGISTERS_reg_1_34_inst : DFF_X1 port map( D => n7972, CK => CLK, Q => 
                           n25477, QN => n22085);
   REGISTERS_reg_1_33_inst : DFF_X1 port map( D => n7971, CK => CLK, Q => 
                           n25476, QN => n22086);
   REGISTERS_reg_1_32_inst : DFF_X1 port map( D => n7970, CK => CLK, Q => 
                           n25475, QN => n22087);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n7969, CK => CLK, Q => 
                           n25474, QN => n22088);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n7968, CK => CLK, Q => 
                           n25473, QN => n22089);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n7967, CK => CLK, Q => 
                           n25472, QN => n22090);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n7966, CK => CLK, Q => 
                           n25471, QN => n22091);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n7965, CK => CLK, Q => 
                           n25470, QN => n22092);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n7964, CK => CLK, Q => 
                           n25469, QN => n22093);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n7963, CK => CLK, Q => 
                           n25468, QN => n22094);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n7962, CK => CLK, Q => 
                           n25467, QN => n22095);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n7961, CK => CLK, Q => 
                           n25466, QN => n22096);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n7960, CK => CLK, Q => 
                           n25465, QN => n22097);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n7959, CK => CLK, Q => 
                           n25464, QN => n22098);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n7958, CK => CLK, Q => 
                           n25463, QN => n22099);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n7957, CK => CLK, Q => 
                           n25462, QN => n22100);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n7956, CK => CLK, Q => 
                           n25461, QN => n22101);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n7955, CK => CLK, Q => 
                           n25460, QN => n22102);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n7954, CK => CLK, Q => 
                           n25459, QN => n22103);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n7953, CK => CLK, Q => 
                           n25458, QN => n22104);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n7952, CK => CLK, Q => 
                           n25457, QN => n22105);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n7951, CK => CLK, Q => 
                           n25456, QN => n22106);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n7950, CK => CLK, Q => 
                           n25455, QN => n22107);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n7949, CK => CLK, Q => 
                           n25666, QN => n22108);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n7948, CK => CLK, Q => 
                           n25665, QN => n22109);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n7947, CK => CLK, Q => n25664
                           , QN => n22110);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n7946, CK => CLK, Q => n25663
                           , QN => n22111);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n7945, CK => CLK, Q => n25662
                           , QN => n22112);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n7944, CK => CLK, Q => n25661
                           , QN => n22113);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n7943, CK => CLK, Q => n25660
                           , QN => n22114);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n7942, CK => CLK, Q => n25659
                           , QN => n22115);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n7941, CK => CLK, Q => n25658
                           , QN => n22116);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n7940, CK => CLK, Q => n25657
                           , QN => n22117);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n7939, CK => CLK, Q => n25656
                           , QN => n22118);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n7938, CK => CLK, Q => n25655
                           , QN => n22119);
   REGISTERS_reg_16_59_inst : DFF_X1 port map( D => n7037, CK => CLK, Q => 
                           n25997, QN => n21240);
   REGISTERS_reg_16_58_inst : DFF_X1 port map( D => n7036, CK => CLK, Q => 
                           n25992, QN => n21241);
   REGISTERS_reg_16_57_inst : DFF_X1 port map( D => n7035, CK => CLK, Q => 
                           n25987, QN => n21242);
   REGISTERS_reg_16_56_inst : DFF_X1 port map( D => n7034, CK => CLK, Q => 
                           n25982, QN => n21243);
   REGISTERS_reg_16_55_inst : DFF_X1 port map( D => n7033, CK => CLK, Q => 
                           n25977, QN => n21244);
   REGISTERS_reg_16_54_inst : DFF_X1 port map( D => n7032, CK => CLK, Q => 
                           n25972, QN => n21245);
   REGISTERS_reg_16_53_inst : DFF_X1 port map( D => n7031, CK => CLK, Q => 
                           n25967, QN => n21246);
   REGISTERS_reg_16_52_inst : DFF_X1 port map( D => n7030, CK => CLK, Q => 
                           n25962, QN => n21247);
   REGISTERS_reg_16_51_inst : DFF_X1 port map( D => n7029, CK => CLK, Q => 
                           n25957, QN => n21248);
   REGISTERS_reg_16_50_inst : DFF_X1 port map( D => n7028, CK => CLK, Q => 
                           n25952, QN => n21249);
   REGISTERS_reg_16_49_inst : DFF_X1 port map( D => n7027, CK => CLK, Q => 
                           n25947, QN => n21250);
   REGISTERS_reg_16_48_inst : DFF_X1 port map( D => n7026, CK => CLK, Q => 
                           n25942, QN => n21251);
   REGISTERS_reg_16_47_inst : DFF_X1 port map( D => n7025, CK => CLK, Q => 
                           n25937, QN => n21252);
   REGISTERS_reg_16_46_inst : DFF_X1 port map( D => n7024, CK => CLK, Q => 
                           n25932, QN => n21253);
   REGISTERS_reg_16_45_inst : DFF_X1 port map( D => n7023, CK => CLK, Q => 
                           n25927, QN => n21254);
   REGISTERS_reg_16_44_inst : DFF_X1 port map( D => n7022, CK => CLK, Q => 
                           n25922, QN => n21255);
   REGISTERS_reg_16_43_inst : DFF_X1 port map( D => n7021, CK => CLK, Q => 
                           n25917, QN => n21256);
   REGISTERS_reg_16_42_inst : DFF_X1 port map( D => n7020, CK => CLK, Q => 
                           n25912, QN => n21257);
   REGISTERS_reg_16_41_inst : DFF_X1 port map( D => n7019, CK => CLK, Q => 
                           n25907, QN => n21258);
   REGISTERS_reg_16_40_inst : DFF_X1 port map( D => n7018, CK => CLK, Q => 
                           n25902, QN => n21259);
   REGISTERS_reg_16_39_inst : DFF_X1 port map( D => n7017, CK => CLK, Q => 
                           n25897, QN => n21260);
   REGISTERS_reg_16_38_inst : DFF_X1 port map( D => n7016, CK => CLK, Q => 
                           n25892, QN => n21261);
   REGISTERS_reg_16_37_inst : DFF_X1 port map( D => n7015, CK => CLK, Q => 
                           n25887, QN => n21262);
   REGISTERS_reg_16_36_inst : DFF_X1 port map( D => n7014, CK => CLK, Q => 
                           n25882, QN => n21263);
   REGISTERS_reg_16_35_inst : DFF_X1 port map( D => n7013, CK => CLK, Q => 
                           n25877, QN => n21264);
   REGISTERS_reg_16_34_inst : DFF_X1 port map( D => n7012, CK => CLK, Q => 
                           n25872, QN => n21265);
   REGISTERS_reg_16_33_inst : DFF_X1 port map( D => n7011, CK => CLK, Q => 
                           n25867, QN => n21266);
   REGISTERS_reg_16_32_inst : DFF_X1 port map( D => n7010, CK => CLK, Q => 
                           n25862, QN => n21267);
   REGISTERS_reg_16_31_inst : DFF_X1 port map( D => n7009, CK => CLK, Q => 
                           n25857, QN => n21268);
   REGISTERS_reg_16_30_inst : DFF_X1 port map( D => n7008, CK => CLK, Q => 
                           n25852, QN => n21269);
   REGISTERS_reg_16_29_inst : DFF_X1 port map( D => n7007, CK => CLK, Q => 
                           n25847, QN => n21270);
   REGISTERS_reg_16_28_inst : DFF_X1 port map( D => n7006, CK => CLK, Q => 
                           n25842, QN => n21271);
   REGISTERS_reg_16_27_inst : DFF_X1 port map( D => n7005, CK => CLK, Q => 
                           n25837, QN => n21272);
   REGISTERS_reg_16_26_inst : DFF_X1 port map( D => n7004, CK => CLK, Q => 
                           n25832, QN => n21273);
   REGISTERS_reg_16_25_inst : DFF_X1 port map( D => n7003, CK => CLK, Q => 
                           n25827, QN => n21274);
   REGISTERS_reg_16_24_inst : DFF_X1 port map( D => n7002, CK => CLK, Q => 
                           n25822, QN => n21275);
   REGISTERS_reg_16_23_inst : DFF_X1 port map( D => n7001, CK => CLK, Q => 
                           n25817, QN => n21276);
   REGISTERS_reg_16_22_inst : DFF_X1 port map( D => n7000, CK => CLK, Q => 
                           n25812, QN => n21277);
   REGISTERS_reg_16_21_inst : DFF_X1 port map( D => n6999, CK => CLK, Q => 
                           n25807, QN => n21278);
   REGISTERS_reg_16_20_inst : DFF_X1 port map( D => n6998, CK => CLK, Q => 
                           n25802, QN => n21279);
   REGISTERS_reg_16_19_inst : DFF_X1 port map( D => n6997, CK => CLK, Q => 
                           n25797, QN => n21280);
   REGISTERS_reg_16_18_inst : DFF_X1 port map( D => n6996, CK => CLK, Q => 
                           n25792, QN => n21281);
   REGISTERS_reg_16_17_inst : DFF_X1 port map( D => n6995, CK => CLK, Q => 
                           n25787, QN => n21282);
   REGISTERS_reg_16_16_inst : DFF_X1 port map( D => n6994, CK => CLK, Q => 
                           n25782, QN => n21283);
   REGISTERS_reg_16_15_inst : DFF_X1 port map( D => n6993, CK => CLK, Q => 
                           n25777, QN => n21284);
   REGISTERS_reg_16_14_inst : DFF_X1 port map( D => n6992, CK => CLK, Q => 
                           n25772, QN => n21285);
   REGISTERS_reg_16_13_inst : DFF_X1 port map( D => n6991, CK => CLK, Q => 
                           n25767, QN => n21286);
   REGISTERS_reg_16_12_inst : DFF_X1 port map( D => n6990, CK => CLK, Q => 
                           n25762, QN => n21287);
   REGISTERS_reg_16_11_inst : DFF_X1 port map( D => n6989, CK => CLK, Q => 
                           n25757, QN => n21288);
   REGISTERS_reg_16_10_inst : DFF_X1 port map( D => n6988, CK => CLK, Q => 
                           n25752, QN => n21289);
   REGISTERS_reg_16_9_inst : DFF_X1 port map( D => n6987, CK => CLK, Q => 
                           n25747, QN => n21290);
   REGISTERS_reg_16_8_inst : DFF_X1 port map( D => n6986, CK => CLK, Q => 
                           n25742, QN => n21291);
   REGISTERS_reg_16_7_inst : DFF_X1 port map( D => n6985, CK => CLK, Q => 
                           n25737, QN => n21292);
   REGISTERS_reg_16_6_inst : DFF_X1 port map( D => n6984, CK => CLK, Q => 
                           n25732, QN => n21293);
   REGISTERS_reg_16_5_inst : DFF_X1 port map( D => n6983, CK => CLK, Q => 
                           n25727, QN => n21294);
   REGISTERS_reg_16_4_inst : DFF_X1 port map( D => n6982, CK => CLK, Q => 
                           n25722, QN => n21295);
   REGISTERS_reg_16_3_inst : DFF_X1 port map( D => n6981, CK => CLK, Q => 
                           n25717, QN => n21296);
   REGISTERS_reg_16_2_inst : DFF_X1 port map( D => n6980, CK => CLK, Q => 
                           n25712, QN => n21297);
   REGISTERS_reg_16_1_inst : DFF_X1 port map( D => n6979, CK => CLK, Q => 
                           n25707, QN => n21298);
   REGISTERS_reg_16_0_inst : DFF_X1 port map( D => n6978, CK => CLK, Q => 
                           n25702, QN => n21299);
   REGISTERS_reg_6_59_inst : DFF_X1 port map( D => n7677, CK => CLK, Q => 
                           n25262, QN => n21820);
   REGISTERS_reg_6_58_inst : DFF_X1 port map( D => n7676, CK => CLK, Q => 
                           n25261, QN => n21821);
   REGISTERS_reg_6_57_inst : DFF_X1 port map( D => n7675, CK => CLK, Q => 
                           n25260, QN => n21822);
   REGISTERS_reg_6_56_inst : DFF_X1 port map( D => n7674, CK => CLK, Q => 
                           n25259, QN => n21823);
   REGISTERS_reg_6_55_inst : DFF_X1 port map( D => n7673, CK => CLK, Q => 
                           n25258, QN => n21824);
   REGISTERS_reg_6_54_inst : DFF_X1 port map( D => n7672, CK => CLK, Q => 
                           n25257, QN => n21825);
   REGISTERS_reg_6_53_inst : DFF_X1 port map( D => n7671, CK => CLK, Q => 
                           n25256, QN => n21826);
   REGISTERS_reg_6_52_inst : DFF_X1 port map( D => n7670, CK => CLK, Q => 
                           n25255, QN => n21827);
   REGISTERS_reg_6_51_inst : DFF_X1 port map( D => n7669, CK => CLK, Q => 
                           n25254, QN => n21828);
   REGISTERS_reg_6_50_inst : DFF_X1 port map( D => n7668, CK => CLK, Q => 
                           n25253, QN => n21829);
   REGISTERS_reg_6_49_inst : DFF_X1 port map( D => n7667, CK => CLK, Q => 
                           n25252, QN => n21830);
   REGISTERS_reg_6_48_inst : DFF_X1 port map( D => n7666, CK => CLK, Q => 
                           n25251, QN => n21831);
   REGISTERS_reg_6_47_inst : DFF_X1 port map( D => n7665, CK => CLK, Q => 
                           n25250, QN => n21832);
   REGISTERS_reg_6_46_inst : DFF_X1 port map( D => n7664, CK => CLK, Q => 
                           n25249, QN => n21833);
   REGISTERS_reg_6_45_inst : DFF_X1 port map( D => n7663, CK => CLK, Q => 
                           n25248, QN => n21834);
   REGISTERS_reg_6_44_inst : DFF_X1 port map( D => n7662, CK => CLK, Q => 
                           n25247, QN => n21835);
   REGISTERS_reg_6_43_inst : DFF_X1 port map( D => n7661, CK => CLK, Q => 
                           n25246, QN => n21836);
   REGISTERS_reg_6_42_inst : DFF_X1 port map( D => n7660, CK => CLK, Q => 
                           n25245, QN => n21837);
   REGISTERS_reg_6_41_inst : DFF_X1 port map( D => n7659, CK => CLK, Q => 
                           n25244, QN => n21838);
   REGISTERS_reg_6_40_inst : DFF_X1 port map( D => n7658, CK => CLK, Q => 
                           n25243, QN => n21839);
   REGISTERS_reg_6_39_inst : DFF_X1 port map( D => n7657, CK => CLK, Q => 
                           n25242, QN => n21840);
   REGISTERS_reg_6_38_inst : DFF_X1 port map( D => n7656, CK => CLK, Q => 
                           n25241, QN => n21841);
   REGISTERS_reg_6_37_inst : DFF_X1 port map( D => n7655, CK => CLK, Q => 
                           n25240, QN => n21842);
   REGISTERS_reg_6_36_inst : DFF_X1 port map( D => n7654, CK => CLK, Q => 
                           n25239, QN => n21843);
   REGISTERS_reg_6_35_inst : DFF_X1 port map( D => n7653, CK => CLK, Q => 
                           n25238, QN => n21844);
   REGISTERS_reg_6_34_inst : DFF_X1 port map( D => n7652, CK => CLK, Q => 
                           n25237, QN => n21845);
   REGISTERS_reg_6_33_inst : DFF_X1 port map( D => n7651, CK => CLK, Q => 
                           n25236, QN => n21846);
   REGISTERS_reg_6_32_inst : DFF_X1 port map( D => n7650, CK => CLK, Q => 
                           n25235, QN => n21847);
   REGISTERS_reg_6_31_inst : DFF_X1 port map( D => n7649, CK => CLK, Q => 
                           n25234, QN => n21848);
   REGISTERS_reg_6_30_inst : DFF_X1 port map( D => n7648, CK => CLK, Q => 
                           n25233, QN => n21849);
   REGISTERS_reg_6_29_inst : DFF_X1 port map( D => n7647, CK => CLK, Q => 
                           n25232, QN => n21850);
   REGISTERS_reg_6_28_inst : DFF_X1 port map( D => n7646, CK => CLK, Q => 
                           n25231, QN => n21851);
   REGISTERS_reg_6_27_inst : DFF_X1 port map( D => n7645, CK => CLK, Q => 
                           n25230, QN => n21852);
   REGISTERS_reg_6_26_inst : DFF_X1 port map( D => n7644, CK => CLK, Q => 
                           n25229, QN => n21853);
   REGISTERS_reg_6_25_inst : DFF_X1 port map( D => n7643, CK => CLK, Q => 
                           n25228, QN => n21854);
   REGISTERS_reg_6_24_inst : DFF_X1 port map( D => n7642, CK => CLK, Q => 
                           n25227, QN => n21855);
   REGISTERS_reg_6_23_inst : DFF_X1 port map( D => n7641, CK => CLK, Q => 
                           n25226, QN => n21856);
   REGISTERS_reg_6_22_inst : DFF_X1 port map( D => n7640, CK => CLK, Q => 
                           n25225, QN => n21857);
   REGISTERS_reg_6_21_inst : DFF_X1 port map( D => n7639, CK => CLK, Q => 
                           n25224, QN => n21858);
   REGISTERS_reg_6_20_inst : DFF_X1 port map( D => n7638, CK => CLK, Q => 
                           n25223, QN => n21859);
   REGISTERS_reg_6_19_inst : DFF_X1 port map( D => n7637, CK => CLK, Q => 
                           n25222, QN => n21860);
   REGISTERS_reg_6_18_inst : DFF_X1 port map( D => n7636, CK => CLK, Q => 
                           n25221, QN => n21861);
   REGISTERS_reg_6_17_inst : DFF_X1 port map( D => n7635, CK => CLK, Q => 
                           n25220, QN => n21862);
   REGISTERS_reg_6_16_inst : DFF_X1 port map( D => n7634, CK => CLK, Q => 
                           n25219, QN => n21863);
   REGISTERS_reg_6_15_inst : DFF_X1 port map( D => n7633, CK => CLK, Q => 
                           n25218, QN => n21864);
   REGISTERS_reg_6_14_inst : DFF_X1 port map( D => n7632, CK => CLK, Q => 
                           n25217, QN => n21865);
   REGISTERS_reg_6_13_inst : DFF_X1 port map( D => n7631, CK => CLK, Q => 
                           n25216, QN => n21866);
   REGISTERS_reg_6_12_inst : DFF_X1 port map( D => n7630, CK => CLK, Q => 
                           n25215, QN => n21867);
   REGISTERS_reg_6_11_inst : DFF_X1 port map( D => n7629, CK => CLK, Q => 
                           n25606, QN => n21868);
   REGISTERS_reg_6_10_inst : DFF_X1 port map( D => n7628, CK => CLK, Q => 
                           n25605, QN => n21869);
   REGISTERS_reg_6_9_inst : DFF_X1 port map( D => n7627, CK => CLK, Q => n25604
                           , QN => n21870);
   REGISTERS_reg_6_8_inst : DFF_X1 port map( D => n7626, CK => CLK, Q => n25603
                           , QN => n21871);
   REGISTERS_reg_6_7_inst : DFF_X1 port map( D => n7625, CK => CLK, Q => n25602
                           , QN => n21872);
   REGISTERS_reg_6_6_inst : DFF_X1 port map( D => n7624, CK => CLK, Q => n25601
                           , QN => n21873);
   REGISTERS_reg_6_5_inst : DFF_X1 port map( D => n7623, CK => CLK, Q => n25600
                           , QN => n21874);
   REGISTERS_reg_6_4_inst : DFF_X1 port map( D => n7622, CK => CLK, Q => n25599
                           , QN => n21875);
   REGISTERS_reg_6_3_inst : DFF_X1 port map( D => n7621, CK => CLK, Q => n25598
                           , QN => n21876);
   REGISTERS_reg_6_2_inst : DFF_X1 port map( D => n7620, CK => CLK, Q => n25597
                           , QN => n21877);
   REGISTERS_reg_6_1_inst : DFF_X1 port map( D => n7619, CK => CLK, Q => n25596
                           , QN => n21878);
   REGISTERS_reg_6_0_inst : DFF_X1 port map( D => n7618, CK => CLK, Q => n25595
                           , QN => n21879);
   OUT2_reg_63_inst : DFF_X1 port map( D => n5889, CK => CLK, Q => n4226, QN =>
                           n_2087);
   U19266 : INV_X1 port map( A => n26537, ZN => n26533);
   U19267 : INV_X1 port map( A => n26762, ZN => n26758);
   U19268 : INV_X1 port map( A => n26541, ZN => n26535);
   U19269 : INV_X1 port map( A => n26540, ZN => n26534);
   U19270 : INV_X1 port map( A => n26765, ZN => n26760);
   U19271 : INV_X1 port map( A => n26763, ZN => n26759);
   U19272 : BUF_X1 port map( A => n22722, Z => n27162);
   U19273 : BUF_X1 port map( A => n22722, Z => n27163);
   U19274 : BUF_X1 port map( A => n22722, Z => n27164);
   U19275 : BUF_X1 port map( A => n22722, Z => n27165);
   U19276 : BUF_X1 port map( A => n22760, Z => n26946);
   U19277 : BUF_X1 port map( A => n22760, Z => n26947);
   U19278 : BUF_X1 port map( A => n22760, Z => n26948);
   U19279 : BUF_X1 port map( A => n22760, Z => n26949);
   U19280 : BUF_X1 port map( A => n22753, Z => n26982);
   U19281 : BUF_X1 port map( A => n22753, Z => n26983);
   U19282 : BUF_X1 port map( A => n22753, Z => n26984);
   U19283 : BUF_X1 port map( A => n22753, Z => n26985);
   U19284 : BUF_X1 port map( A => n22719, Z => n27174);
   U19285 : BUF_X1 port map( A => n22719, Z => n27175);
   U19286 : BUF_X1 port map( A => n22719, Z => n27176);
   U19287 : BUF_X1 port map( A => n22719, Z => n27177);
   U19288 : BUF_X1 port map( A => n22724, Z => n27150);
   U19289 : BUF_X1 port map( A => n22724, Z => n27151);
   U19290 : BUF_X1 port map( A => n22724, Z => n27152);
   U19291 : BUF_X1 port map( A => n22724, Z => n27153);
   U19292 : BUF_X1 port map( A => n22743, Z => n27042);
   U19293 : BUF_X1 port map( A => n22743, Z => n27043);
   U19294 : BUF_X1 port map( A => n22743, Z => n27044);
   U19295 : BUF_X1 port map( A => n22743, Z => n27045);
   U19296 : BUF_X1 port map( A => n22764, Z => n26922);
   U19297 : BUF_X1 port map( A => n22764, Z => n26923);
   U19298 : BUF_X1 port map( A => n22764, Z => n26924);
   U19299 : BUF_X1 port map( A => n22764, Z => n26925);
   U19300 : BUF_X1 port map( A => n22762, Z => n26934);
   U19301 : BUF_X1 port map( A => n22762, Z => n26935);
   U19302 : BUF_X1 port map( A => n22762, Z => n26936);
   U19303 : BUF_X1 port map( A => n22762, Z => n26937);
   U19304 : BUF_X1 port map( A => n22693, Z => n27270);
   U19305 : BUF_X1 port map( A => n22693, Z => n27271);
   U19306 : BUF_X1 port map( A => n22693, Z => n27272);
   U19307 : BUF_X1 port map( A => n22693, Z => n27273);
   U19308 : BUF_X1 port map( A => n22697, Z => n27258);
   U19309 : BUF_X1 port map( A => n22697, Z => n27259);
   U19310 : BUF_X1 port map( A => n22697, Z => n27260);
   U19311 : BUF_X1 port map( A => n22697, Z => n27261);
   U19312 : BUF_X1 port map( A => n22715, Z => n27186);
   U19313 : BUF_X1 port map( A => n22715, Z => n27187);
   U19314 : BUF_X1 port map( A => n22715, Z => n27188);
   U19315 : BUF_X1 port map( A => n22715, Z => n27189);
   U19316 : BUF_X1 port map( A => n22726, Z => n27138);
   U19317 : BUF_X1 port map( A => n22726, Z => n27139);
   U19318 : BUF_X1 port map( A => n22726, Z => n27140);
   U19319 : BUF_X1 port map( A => n22726, Z => n27141);
   U19320 : BUF_X1 port map( A => n22706, Z => n27222);
   U19321 : BUF_X1 port map( A => n22706, Z => n27223);
   U19322 : BUF_X1 port map( A => n22706, Z => n27224);
   U19323 : BUF_X1 port map( A => n22706, Z => n27225);
   U19324 : BUF_X1 port map( A => n22712, Z => n27198);
   U19325 : BUF_X1 port map( A => n22712, Z => n27199);
   U19326 : BUF_X1 port map( A => n22712, Z => n27200);
   U19327 : BUF_X1 port map( A => n22712, Z => n27201);
   U19328 : BUF_X1 port map( A => n22749, Z => n27006);
   U19329 : BUF_X1 port map( A => n22749, Z => n27007);
   U19330 : BUF_X1 port map( A => n22749, Z => n27008);
   U19331 : BUF_X1 port map( A => n22749, Z => n27009);
   U19332 : BUF_X1 port map( A => n22739, Z => n27066);
   U19333 : BUF_X1 port map( A => n22739, Z => n27067);
   U19334 : BUF_X1 port map( A => n22739, Z => n27068);
   U19335 : BUF_X1 port map( A => n22739, Z => n27069);
   U19336 : BUF_X1 port map( A => n22741, Z => n27054);
   U19337 : BUF_X1 port map( A => n22741, Z => n27055);
   U19338 : BUF_X1 port map( A => n22741, Z => n27056);
   U19339 : BUF_X1 port map( A => n22741, Z => n27057);
   U19340 : BUF_X1 port map( A => n22758, Z => n26958);
   U19341 : BUF_X1 port map( A => n22758, Z => n26959);
   U19342 : BUF_X1 port map( A => n22758, Z => n26960);
   U19343 : BUF_X1 port map( A => n22758, Z => n26961);
   U19344 : BUF_X1 port map( A => n22709, Z => n27210);
   U19345 : BUF_X1 port map( A => n22709, Z => n27211);
   U19346 : BUF_X1 port map( A => n22709, Z => n27212);
   U19347 : BUF_X1 port map( A => n22709, Z => n27213);
   U19348 : BUF_X1 port map( A => n22700, Z => n27246);
   U19349 : BUF_X1 port map( A => n22700, Z => n27247);
   U19350 : BUF_X1 port map( A => n22700, Z => n27248);
   U19351 : BUF_X1 port map( A => n22700, Z => n27249);
   U19352 : BUF_X1 port map( A => n22703, Z => n27234);
   U19353 : BUF_X1 port map( A => n22703, Z => n27235);
   U19354 : BUF_X1 port map( A => n22703, Z => n27236);
   U19355 : BUF_X1 port map( A => n22703, Z => n27237);
   U19356 : BUF_X1 port map( A => n22751, Z => n26994);
   U19357 : BUF_X1 port map( A => n22751, Z => n26995);
   U19358 : BUF_X1 port map( A => n22751, Z => n26996);
   U19359 : BUF_X1 port map( A => n22751, Z => n26997);
   U19360 : BUF_X1 port map( A => n22736, Z => n27078);
   U19361 : BUF_X1 port map( A => n22736, Z => n27079);
   U19362 : BUF_X1 port map( A => n22736, Z => n27080);
   U19363 : BUF_X1 port map( A => n22736, Z => n27081);
   U19364 : BUF_X1 port map( A => n22756, Z => n26970);
   U19365 : BUF_X1 port map( A => n22756, Z => n26971);
   U19366 : BUF_X1 port map( A => n22756, Z => n26972);
   U19367 : BUF_X1 port map( A => n22756, Z => n26973);
   U19368 : BUF_X1 port map( A => n22768, Z => n26898);
   U19369 : BUF_X1 port map( A => n22768, Z => n26899);
   U19370 : BUF_X1 port map( A => n22768, Z => n26900);
   U19371 : BUF_X1 port map( A => n22768, Z => n26901);
   U19372 : BUF_X1 port map( A => n22766, Z => n26910);
   U19373 : BUF_X1 port map( A => n22766, Z => n26911);
   U19374 : BUF_X1 port map( A => n22766, Z => n26912);
   U19375 : BUF_X1 port map( A => n22766, Z => n26913);
   U19376 : BUF_X1 port map( A => n22732, Z => n27102);
   U19377 : BUF_X1 port map( A => n22732, Z => n27103);
   U19378 : BUF_X1 port map( A => n22732, Z => n27104);
   U19379 : BUF_X1 port map( A => n22732, Z => n27105);
   U19380 : BUF_X1 port map( A => n22728, Z => n27126);
   U19381 : BUF_X1 port map( A => n22728, Z => n27127);
   U19382 : BUF_X1 port map( A => n22728, Z => n27128);
   U19383 : BUF_X1 port map( A => n22728, Z => n27129);
   U19384 : BUF_X1 port map( A => n27275, Z => n27277);
   U19385 : BUF_X1 port map( A => n27275, Z => n27278);
   U19386 : BUF_X1 port map( A => n27275, Z => n27279);
   U19387 : BUF_X1 port map( A => n27276, Z => n27280);
   U19388 : BUF_X1 port map( A => n27276, Z => n27281);
   U19389 : BUF_X1 port map( A => n22730, Z => n27113);
   U19390 : BUF_X1 port map( A => n22730, Z => n27114);
   U19391 : BUF_X1 port map( A => n22730, Z => n27115);
   U19392 : BUF_X1 port map( A => n22730, Z => n27116);
   U19393 : BUF_X1 port map( A => n22730, Z => n27117);
   U19394 : BUF_X1 port map( A => n22734, Z => n27089);
   U19395 : BUF_X1 port map( A => n22734, Z => n27090);
   U19396 : BUF_X1 port map( A => n22734, Z => n27091);
   U19397 : BUF_X1 port map( A => n22734, Z => n27092);
   U19398 : BUF_X1 port map( A => n22734, Z => n27093);
   U19399 : BUF_X1 port map( A => n22745, Z => n27029);
   U19400 : BUF_X1 port map( A => n22745, Z => n27030);
   U19401 : BUF_X1 port map( A => n22745, Z => n27031);
   U19402 : BUF_X1 port map( A => n22745, Z => n27032);
   U19403 : BUF_X1 port map( A => n22745, Z => n27033);
   U19404 : BUF_X1 port map( A => n22747, Z => n27017);
   U19405 : BUF_X1 port map( A => n22747, Z => n27018);
   U19406 : BUF_X1 port map( A => n22747, Z => n27019);
   U19407 : BUF_X1 port map( A => n22747, Z => n27020);
   U19408 : BUF_X1 port map( A => n22747, Z => n27021);
   U19409 : BUF_X1 port map( A => n23980, Z => n26636);
   U19410 : BUF_X1 port map( A => n23980, Z => n26637);
   U19411 : BUF_X1 port map( A => n23980, Z => n26638);
   U19412 : BUF_X1 port map( A => n23980, Z => n26639);
   U19413 : BUF_X1 port map( A => n23980, Z => n26640);
   U19414 : BUF_X1 port map( A => n22781, Z => n26861);
   U19415 : BUF_X1 port map( A => n22781, Z => n26862);
   U19416 : BUF_X1 port map( A => n22781, Z => n26863);
   U19417 : BUF_X1 port map( A => n22781, Z => n26864);
   U19418 : BUF_X1 port map( A => n22781, Z => n26865);
   U19419 : BUF_X1 port map( A => n22760, Z => n26945);
   U19420 : BUF_X1 port map( A => n22753, Z => n26981);
   U19421 : BUF_X1 port map( A => n22764, Z => n26921);
   U19422 : BUF_X1 port map( A => n22762, Z => n26933);
   U19423 : BUF_X1 port map( A => n22758, Z => n26957);
   U19424 : BUF_X1 port map( A => n22756, Z => n26969);
   U19425 : BUF_X1 port map( A => n22768, Z => n26897);
   U19426 : BUF_X1 port map( A => n22766, Z => n26909);
   U19427 : BUF_X1 port map( A => n22722, Z => n27161);
   U19428 : BUF_X1 port map( A => n22719, Z => n27173);
   U19429 : BUF_X1 port map( A => n22724, Z => n27149);
   U19430 : BUF_X1 port map( A => n22743, Z => n27041);
   U19431 : BUF_X1 port map( A => n22693, Z => n27269);
   U19432 : BUF_X1 port map( A => n22697, Z => n27257);
   U19433 : BUF_X1 port map( A => n22715, Z => n27185);
   U19434 : BUF_X1 port map( A => n22726, Z => n27137);
   U19435 : BUF_X1 port map( A => n22706, Z => n27221);
   U19436 : BUF_X1 port map( A => n22712, Z => n27197);
   U19437 : BUF_X1 port map( A => n22749, Z => n27005);
   U19438 : BUF_X1 port map( A => n22739, Z => n27065);
   U19439 : BUF_X1 port map( A => n22741, Z => n27053);
   U19440 : BUF_X1 port map( A => n22709, Z => n27209);
   U19441 : BUF_X1 port map( A => n22700, Z => n27245);
   U19442 : BUF_X1 port map( A => n22703, Z => n27233);
   U19443 : BUF_X1 port map( A => n22751, Z => n26993);
   U19444 : BUF_X1 port map( A => n22736, Z => n27077);
   U19445 : BUF_X1 port map( A => n22732, Z => n27101);
   U19446 : BUF_X1 port map( A => n22728, Z => n27125);
   U19447 : BUF_X1 port map( A => n26526, Z => n26541);
   U19448 : BUF_X1 port map( A => n26526, Z => n26540);
   U19449 : BUF_X1 port map( A => n26526, Z => n26539);
   U19450 : BUF_X1 port map( A => n26525, Z => n26538);
   U19451 : BUF_X1 port map( A => n26525, Z => n26537);
   U19452 : BUF_X1 port map( A => n26751, Z => n26766);
   U19453 : BUF_X1 port map( A => n26751, Z => n26765);
   U19454 : BUF_X1 port map( A => n26751, Z => n26764);
   U19455 : BUF_X1 port map( A => n26750, Z => n26763);
   U19456 : BUF_X1 port map( A => n26750, Z => n26762);
   U19457 : BUF_X1 port map( A => n26525, Z => n26536);
   U19458 : BUF_X1 port map( A => n26750, Z => n26761);
   U19459 : BUF_X1 port map( A => n26529, Z => n26550);
   U19460 : BUF_X1 port map( A => n26529, Z => n26549);
   U19461 : BUF_X1 port map( A => n26529, Z => n26548);
   U19462 : BUF_X1 port map( A => n26528, Z => n26547);
   U19463 : BUF_X1 port map( A => n26528, Z => n26546);
   U19464 : BUF_X1 port map( A => n26528, Z => n26545);
   U19465 : BUF_X1 port map( A => n26527, Z => n26544);
   U19466 : BUF_X1 port map( A => n26527, Z => n26543);
   U19467 : BUF_X1 port map( A => n26527, Z => n26542);
   U19468 : BUF_X1 port map( A => n26754, Z => n26775);
   U19469 : BUF_X1 port map( A => n26754, Z => n26774);
   U19470 : BUF_X1 port map( A => n26754, Z => n26773);
   U19471 : BUF_X1 port map( A => n26753, Z => n26772);
   U19472 : BUF_X1 port map( A => n26753, Z => n26771);
   U19473 : BUF_X1 port map( A => n26753, Z => n26770);
   U19474 : BUF_X1 port map( A => n26752, Z => n26768);
   U19475 : BUF_X1 port map( A => n26752, Z => n26767);
   U19476 : BUF_X1 port map( A => n26752, Z => n26769);
   U19477 : BUF_X1 port map( A => n26530, Z => n26551);
   U19478 : BUF_X1 port map( A => n26755, Z => n26776);
   U19479 : BUF_X1 port map( A => n23992, Z => n26582);
   U19480 : BUF_X1 port map( A => n24017, Z => n26459);
   U19481 : BUF_X1 port map( A => n23992, Z => n26583);
   U19482 : BUF_X1 port map( A => n24017, Z => n26460);
   U19483 : BUF_X1 port map( A => n23992, Z => n26584);
   U19484 : BUF_X1 port map( A => n24017, Z => n26461);
   U19485 : BUF_X1 port map( A => n23992, Z => n26585);
   U19486 : BUF_X1 port map( A => n24017, Z => n26462);
   U19487 : BUF_X1 port map( A => n23992, Z => n26586);
   U19488 : BUF_X1 port map( A => n24017, Z => n26463);
   U19489 : BUF_X1 port map( A => n22793, Z => n26807);
   U19490 : BUF_X1 port map( A => n22818, Z => n26684);
   U19491 : BUF_X1 port map( A => n22793, Z => n26808);
   U19492 : BUF_X1 port map( A => n22818, Z => n26685);
   U19493 : BUF_X1 port map( A => n22793, Z => n26809);
   U19494 : BUF_X1 port map( A => n22818, Z => n26686);
   U19495 : BUF_X1 port map( A => n22793, Z => n26810);
   U19496 : BUF_X1 port map( A => n22818, Z => n26687);
   U19497 : BUF_X1 port map( A => n22793, Z => n26811);
   U19498 : BUF_X1 port map( A => n22818, Z => n26688);
   U19499 : BUF_X1 port map( A => n24012, Z => n26483);
   U19500 : BUF_X1 port map( A => n24012, Z => n26484);
   U19501 : BUF_X1 port map( A => n24012, Z => n26485);
   U19502 : BUF_X1 port map( A => n24012, Z => n26486);
   U19503 : BUF_X1 port map( A => n24012, Z => n26487);
   U19504 : BUF_X1 port map( A => n22813, Z => n26708);
   U19505 : BUF_X1 port map( A => n22813, Z => n26709);
   U19506 : BUF_X1 port map( A => n22813, Z => n26710);
   U19507 : BUF_X1 port map( A => n22813, Z => n26711);
   U19508 : BUF_X1 port map( A => n22813, Z => n26712);
   U19509 : BUF_X1 port map( A => n23987, Z => n26606);
   U19510 : BUF_X1 port map( A => n23977, Z => n26654);
   U19511 : BUF_X1 port map( A => n23982, Z => n26630);
   U19512 : BUF_X1 port map( A => n24007, Z => n26507);
   U19513 : BUF_X1 port map( A => n24002, Z => n26552);
   U19514 : BUF_X1 port map( A => n23987, Z => n26607);
   U19515 : BUF_X1 port map( A => n23977, Z => n26655);
   U19516 : BUF_X1 port map( A => n23982, Z => n26631);
   U19517 : BUF_X1 port map( A => n24007, Z => n26508);
   U19518 : BUF_X1 port map( A => n24002, Z => n26553);
   U19519 : BUF_X1 port map( A => n23987, Z => n26608);
   U19520 : BUF_X1 port map( A => n23977, Z => n26656);
   U19521 : BUF_X1 port map( A => n23982, Z => n26632);
   U19522 : BUF_X1 port map( A => n24007, Z => n26509);
   U19523 : BUF_X1 port map( A => n24002, Z => n26554);
   U19524 : BUF_X1 port map( A => n23987, Z => n26609);
   U19525 : BUF_X1 port map( A => n23977, Z => n26657);
   U19526 : BUF_X1 port map( A => n23982, Z => n26633);
   U19527 : BUF_X1 port map( A => n24007, Z => n26510);
   U19528 : BUF_X1 port map( A => n24002, Z => n26555);
   U19529 : BUF_X1 port map( A => n23987, Z => n26610);
   U19530 : BUF_X1 port map( A => n23977, Z => n26658);
   U19531 : BUF_X1 port map( A => n23982, Z => n26634);
   U19532 : BUF_X1 port map( A => n24007, Z => n26511);
   U19533 : BUF_X1 port map( A => n24002, Z => n26556);
   U19534 : BUF_X1 port map( A => n22788, Z => n26831);
   U19535 : BUF_X1 port map( A => n22778, Z => n26879);
   U19536 : BUF_X1 port map( A => n22783, Z => n26855);
   U19537 : BUF_X1 port map( A => n22808, Z => n26732);
   U19538 : BUF_X1 port map( A => n22803, Z => n26777);
   U19539 : BUF_X1 port map( A => n22788, Z => n26832);
   U19540 : BUF_X1 port map( A => n22778, Z => n26880);
   U19541 : BUF_X1 port map( A => n22783, Z => n26856);
   U19542 : BUF_X1 port map( A => n22808, Z => n26733);
   U19543 : BUF_X1 port map( A => n22803, Z => n26778);
   U19544 : BUF_X1 port map( A => n22788, Z => n26833);
   U19545 : BUF_X1 port map( A => n22778, Z => n26881);
   U19546 : BUF_X1 port map( A => n22783, Z => n26857);
   U19547 : BUF_X1 port map( A => n22808, Z => n26734);
   U19548 : BUF_X1 port map( A => n22803, Z => n26779);
   U19549 : BUF_X1 port map( A => n22788, Z => n26834);
   U19550 : BUF_X1 port map( A => n22778, Z => n26882);
   U19551 : BUF_X1 port map( A => n22783, Z => n26858);
   U19552 : BUF_X1 port map( A => n22808, Z => n26735);
   U19553 : BUF_X1 port map( A => n22803, Z => n26780);
   U19554 : BUF_X1 port map( A => n22788, Z => n26835);
   U19555 : BUF_X1 port map( A => n22778, Z => n26883);
   U19556 : BUF_X1 port map( A => n22783, Z => n26859);
   U19557 : BUF_X1 port map( A => n22808, Z => n26736);
   U19558 : BUF_X1 port map( A => n22803, Z => n26781);
   U19559 : BUF_X1 port map( A => n23989, Z => n26595);
   U19560 : BUF_X1 port map( A => n23984, Z => n26619);
   U19561 : BUF_X1 port map( A => n23974, Z => n26667);
   U19562 : BUF_X1 port map( A => n23979, Z => n26643);
   U19563 : BUF_X1 port map( A => n24004, Z => n26520);
   U19564 : BUF_X1 port map( A => n23999, Z => n26565);
   U19565 : BUF_X1 port map( A => n23989, Z => n26596);
   U19566 : BUF_X1 port map( A => n23984, Z => n26620);
   U19567 : BUF_X1 port map( A => n23974, Z => n26668);
   U19568 : BUF_X1 port map( A => n23979, Z => n26644);
   U19569 : BUF_X1 port map( A => n24004, Z => n26521);
   U19570 : BUF_X1 port map( A => n23999, Z => n26566);
   U19571 : BUF_X1 port map( A => n23989, Z => n26597);
   U19572 : BUF_X1 port map( A => n23984, Z => n26621);
   U19573 : BUF_X1 port map( A => n23974, Z => n26669);
   U19574 : BUF_X1 port map( A => n23979, Z => n26645);
   U19575 : BUF_X1 port map( A => n24004, Z => n26522);
   U19576 : BUF_X1 port map( A => n23999, Z => n26567);
   U19577 : BUF_X1 port map( A => n23989, Z => n26598);
   U19578 : BUF_X1 port map( A => n23984, Z => n26622);
   U19579 : BUF_X1 port map( A => n23974, Z => n26670);
   U19580 : BUF_X1 port map( A => n23979, Z => n26646);
   U19581 : BUF_X1 port map( A => n24004, Z => n26523);
   U19582 : BUF_X1 port map( A => n23999, Z => n26568);
   U19583 : BUF_X1 port map( A => n22790, Z => n26820);
   U19584 : BUF_X1 port map( A => n22785, Z => n26844);
   U19585 : BUF_X1 port map( A => n22775, Z => n26892);
   U19586 : BUF_X1 port map( A => n22780, Z => n26868);
   U19587 : BUF_X1 port map( A => n22805, Z => n26745);
   U19588 : BUF_X1 port map( A => n22800, Z => n26790);
   U19589 : BUF_X1 port map( A => n22790, Z => n26821);
   U19590 : BUF_X1 port map( A => n22785, Z => n26845);
   U19591 : BUF_X1 port map( A => n22775, Z => n26893);
   U19592 : BUF_X1 port map( A => n22780, Z => n26869);
   U19593 : BUF_X1 port map( A => n22805, Z => n26746);
   U19594 : BUF_X1 port map( A => n22800, Z => n26791);
   U19595 : BUF_X1 port map( A => n22790, Z => n26822);
   U19596 : BUF_X1 port map( A => n22785, Z => n26846);
   U19597 : BUF_X1 port map( A => n22775, Z => n26894);
   U19598 : BUF_X1 port map( A => n22780, Z => n26870);
   U19599 : BUF_X1 port map( A => n22805, Z => n26747);
   U19600 : BUF_X1 port map( A => n22800, Z => n26792);
   U19601 : BUF_X1 port map( A => n22790, Z => n26823);
   U19602 : BUF_X1 port map( A => n22785, Z => n26847);
   U19603 : BUF_X1 port map( A => n22775, Z => n26895);
   U19604 : BUF_X1 port map( A => n22780, Z => n26871);
   U19605 : BUF_X1 port map( A => n22805, Z => n26748);
   U19606 : BUF_X1 port map( A => n22800, Z => n26793);
   U19607 : BUF_X1 port map( A => n23993, Z => n26576);
   U19608 : BUF_X1 port map( A => n24018, Z => n26453);
   U19609 : BUF_X1 port map( A => n23993, Z => n26577);
   U19610 : BUF_X1 port map( A => n24018, Z => n26454);
   U19611 : BUF_X1 port map( A => n23993, Z => n26578);
   U19612 : BUF_X1 port map( A => n24018, Z => n26455);
   U19613 : BUF_X1 port map( A => n23993, Z => n26579);
   U19614 : BUF_X1 port map( A => n24018, Z => n26456);
   U19615 : BUF_X1 port map( A => n23993, Z => n26580);
   U19616 : BUF_X1 port map( A => n24018, Z => n26457);
   U19617 : BUF_X1 port map( A => n22794, Z => n26801);
   U19618 : BUF_X1 port map( A => n22819, Z => n26678);
   U19619 : BUF_X1 port map( A => n22794, Z => n26802);
   U19620 : BUF_X1 port map( A => n22819, Z => n26679);
   U19621 : BUF_X1 port map( A => n22794, Z => n26803);
   U19622 : BUF_X1 port map( A => n22819, Z => n26680);
   U19623 : BUF_X1 port map( A => n22794, Z => n26804);
   U19624 : BUF_X1 port map( A => n22819, Z => n26681);
   U19625 : BUF_X1 port map( A => n22794, Z => n26805);
   U19626 : BUF_X1 port map( A => n22819, Z => n26682);
   U19627 : BUF_X1 port map( A => n23988, Z => n26600);
   U19628 : BUF_X1 port map( A => n23978, Z => n26648);
   U19629 : BUF_X1 port map( A => n23983, Z => n26624);
   U19630 : BUF_X1 port map( A => n24008, Z => n26501);
   U19631 : BUF_X1 port map( A => n24013, Z => n26477);
   U19632 : BUF_X1 port map( A => n23988, Z => n26601);
   U19633 : BUF_X1 port map( A => n23978, Z => n26649);
   U19634 : BUF_X1 port map( A => n23983, Z => n26625);
   U19635 : BUF_X1 port map( A => n24008, Z => n26502);
   U19636 : BUF_X1 port map( A => n24013, Z => n26478);
   U19637 : BUF_X1 port map( A => n23988, Z => n26602);
   U19638 : BUF_X1 port map( A => n23978, Z => n26650);
   U19639 : BUF_X1 port map( A => n23983, Z => n26626);
   U19640 : BUF_X1 port map( A => n24008, Z => n26503);
   U19641 : BUF_X1 port map( A => n24013, Z => n26479);
   U19642 : BUF_X1 port map( A => n23988, Z => n26603);
   U19643 : BUF_X1 port map( A => n23978, Z => n26651);
   U19644 : BUF_X1 port map( A => n23983, Z => n26627);
   U19645 : BUF_X1 port map( A => n24008, Z => n26504);
   U19646 : BUF_X1 port map( A => n24013, Z => n26480);
   U19647 : BUF_X1 port map( A => n23988, Z => n26604);
   U19648 : BUF_X1 port map( A => n23978, Z => n26652);
   U19649 : BUF_X1 port map( A => n23983, Z => n26628);
   U19650 : BUF_X1 port map( A => n24008, Z => n26505);
   U19651 : BUF_X1 port map( A => n24013, Z => n26481);
   U19652 : BUF_X1 port map( A => n22789, Z => n26825);
   U19653 : BUF_X1 port map( A => n22779, Z => n26873);
   U19654 : BUF_X1 port map( A => n22784, Z => n26849);
   U19655 : BUF_X1 port map( A => n22809, Z => n26726);
   U19656 : BUF_X1 port map( A => n22814, Z => n26702);
   U19657 : BUF_X1 port map( A => n22789, Z => n26826);
   U19658 : BUF_X1 port map( A => n22779, Z => n26874);
   U19659 : BUF_X1 port map( A => n22784, Z => n26850);
   U19660 : BUF_X1 port map( A => n22809, Z => n26727);
   U19661 : BUF_X1 port map( A => n22814, Z => n26703);
   U19662 : BUF_X1 port map( A => n22789, Z => n26827);
   U19663 : BUF_X1 port map( A => n22779, Z => n26875);
   U19664 : BUF_X1 port map( A => n22784, Z => n26851);
   U19665 : BUF_X1 port map( A => n22809, Z => n26728);
   U19666 : BUF_X1 port map( A => n22814, Z => n26704);
   U19667 : BUF_X1 port map( A => n22789, Z => n26828);
   U19668 : BUF_X1 port map( A => n22779, Z => n26876);
   U19669 : BUF_X1 port map( A => n22784, Z => n26852);
   U19670 : BUF_X1 port map( A => n22809, Z => n26729);
   U19671 : BUF_X1 port map( A => n22814, Z => n26705);
   U19672 : BUF_X1 port map( A => n22789, Z => n26829);
   U19673 : BUF_X1 port map( A => n22779, Z => n26877);
   U19674 : BUF_X1 port map( A => n22784, Z => n26853);
   U19675 : BUF_X1 port map( A => n22809, Z => n26730);
   U19676 : BUF_X1 port map( A => n22814, Z => n26706);
   U19677 : BUF_X1 port map( A => n23994, Z => n26570);
   U19678 : BUF_X1 port map( A => n24019, Z => n26447);
   U19679 : BUF_X1 port map( A => n23994, Z => n26571);
   U19680 : BUF_X1 port map( A => n24019, Z => n26448);
   U19681 : BUF_X1 port map( A => n23994, Z => n26572);
   U19682 : BUF_X1 port map( A => n24019, Z => n26449);
   U19683 : BUF_X1 port map( A => n23994, Z => n26573);
   U19684 : BUF_X1 port map( A => n24019, Z => n26450);
   U19685 : BUF_X1 port map( A => n23994, Z => n26574);
   U19686 : BUF_X1 port map( A => n24019, Z => n26451);
   U19687 : BUF_X1 port map( A => n22795, Z => n26795);
   U19688 : BUF_X1 port map( A => n22820, Z => n26672);
   U19689 : BUF_X1 port map( A => n22795, Z => n26796);
   U19690 : BUF_X1 port map( A => n22820, Z => n26673);
   U19691 : BUF_X1 port map( A => n22795, Z => n26797);
   U19692 : BUF_X1 port map( A => n22820, Z => n26674);
   U19693 : BUF_X1 port map( A => n22795, Z => n26798);
   U19694 : BUF_X1 port map( A => n22820, Z => n26675);
   U19695 : BUF_X1 port map( A => n22795, Z => n26799);
   U19696 : BUF_X1 port map( A => n22820, Z => n26676);
   U19697 : BUF_X1 port map( A => n22696, Z => n27263);
   U19698 : BUF_X1 port map( A => n22714, Z => n27191);
   U19699 : BUF_X1 port map( A => n22705, Z => n27227);
   U19700 : BUF_X1 port map( A => n22711, Z => n27203);
   U19701 : BUF_X1 port map( A => n22708, Z => n27215);
   U19702 : BUF_X1 port map( A => n22699, Z => n27251);
   U19703 : BUF_X1 port map( A => n22702, Z => n27239);
   U19704 : BUF_X1 port map( A => n22721, Z => n27167);
   U19705 : BUF_X1 port map( A => n22759, Z => n26951);
   U19706 : BUF_X1 port map( A => n22752, Z => n26987);
   U19707 : BUF_X1 port map( A => n22718, Z => n27179);
   U19708 : BUF_X1 port map( A => n22723, Z => n27155);
   U19709 : BUF_X1 port map( A => n22742, Z => n27047);
   U19710 : BUF_X1 port map( A => n22763, Z => n26927);
   U19711 : BUF_X1 port map( A => n22761, Z => n26939);
   U19712 : BUF_X1 port map( A => n22725, Z => n27143);
   U19713 : BUF_X1 port map( A => n22748, Z => n27011);
   U19714 : BUF_X1 port map( A => n22738, Z => n27071);
   U19715 : BUF_X1 port map( A => n22740, Z => n27059);
   U19716 : BUF_X1 port map( A => n22757, Z => n26963);
   U19717 : BUF_X1 port map( A => n22750, Z => n26999);
   U19718 : BUF_X1 port map( A => n22735, Z => n27083);
   U19719 : BUF_X1 port map( A => n22755, Z => n26975);
   U19720 : BUF_X1 port map( A => n22729, Z => n27119);
   U19721 : BUF_X1 port map( A => n22733, Z => n27095);
   U19722 : BUF_X1 port map( A => n22744, Z => n27035);
   U19723 : BUF_X1 port map( A => n22746, Z => n27023);
   U19724 : BUF_X1 port map( A => n22767, Z => n26903);
   U19725 : BUF_X1 port map( A => n22765, Z => n26915);
   U19726 : BUF_X1 port map( A => n22731, Z => n27107);
   U19727 : BUF_X1 port map( A => n22727, Z => n27131);
   U19728 : BUF_X1 port map( A => n22696, Z => n27264);
   U19729 : BUF_X1 port map( A => n22696, Z => n27265);
   U19730 : BUF_X1 port map( A => n22696, Z => n27266);
   U19731 : BUF_X1 port map( A => n22696, Z => n27267);
   U19732 : BUF_X1 port map( A => n22714, Z => n27192);
   U19733 : BUF_X1 port map( A => n22714, Z => n27193);
   U19734 : BUF_X1 port map( A => n22714, Z => n27194);
   U19735 : BUF_X1 port map( A => n22714, Z => n27195);
   U19736 : BUF_X1 port map( A => n22705, Z => n27228);
   U19737 : BUF_X1 port map( A => n22705, Z => n27229);
   U19738 : BUF_X1 port map( A => n22705, Z => n27230);
   U19739 : BUF_X1 port map( A => n22705, Z => n27231);
   U19740 : BUF_X1 port map( A => n22711, Z => n27204);
   U19741 : BUF_X1 port map( A => n22711, Z => n27205);
   U19742 : BUF_X1 port map( A => n22711, Z => n27206);
   U19743 : BUF_X1 port map( A => n22711, Z => n27207);
   U19744 : BUF_X1 port map( A => n22708, Z => n27216);
   U19745 : BUF_X1 port map( A => n22708, Z => n27217);
   U19746 : BUF_X1 port map( A => n22708, Z => n27218);
   U19747 : BUF_X1 port map( A => n22708, Z => n27219);
   U19748 : BUF_X1 port map( A => n22699, Z => n27252);
   U19749 : BUF_X1 port map( A => n22699, Z => n27253);
   U19750 : BUF_X1 port map( A => n22699, Z => n27254);
   U19751 : BUF_X1 port map( A => n22699, Z => n27255);
   U19752 : BUF_X1 port map( A => n22702, Z => n27240);
   U19753 : BUF_X1 port map( A => n22702, Z => n27241);
   U19754 : BUF_X1 port map( A => n22702, Z => n27242);
   U19755 : BUF_X1 port map( A => n22702, Z => n27243);
   U19756 : BUF_X1 port map( A => n22721, Z => n27168);
   U19757 : BUF_X1 port map( A => n22721, Z => n27169);
   U19758 : BUF_X1 port map( A => n22721, Z => n27170);
   U19759 : BUF_X1 port map( A => n22721, Z => n27171);
   U19760 : BUF_X1 port map( A => n22759, Z => n26952);
   U19761 : BUF_X1 port map( A => n22759, Z => n26953);
   U19762 : BUF_X1 port map( A => n22759, Z => n26954);
   U19763 : BUF_X1 port map( A => n22759, Z => n26955);
   U19764 : BUF_X1 port map( A => n22752, Z => n26988);
   U19765 : BUF_X1 port map( A => n22752, Z => n26989);
   U19766 : BUF_X1 port map( A => n22752, Z => n26990);
   U19767 : BUF_X1 port map( A => n22752, Z => n26991);
   U19768 : BUF_X1 port map( A => n22718, Z => n27180);
   U19769 : BUF_X1 port map( A => n22718, Z => n27181);
   U19770 : BUF_X1 port map( A => n22718, Z => n27182);
   U19771 : BUF_X1 port map( A => n22718, Z => n27183);
   U19772 : BUF_X1 port map( A => n22723, Z => n27156);
   U19773 : BUF_X1 port map( A => n22723, Z => n27157);
   U19774 : BUF_X1 port map( A => n22723, Z => n27158);
   U19775 : BUF_X1 port map( A => n22723, Z => n27159);
   U19776 : BUF_X1 port map( A => n22742, Z => n27048);
   U19777 : BUF_X1 port map( A => n22742, Z => n27049);
   U19778 : BUF_X1 port map( A => n22742, Z => n27050);
   U19779 : BUF_X1 port map( A => n22742, Z => n27051);
   U19780 : BUF_X1 port map( A => n22763, Z => n26928);
   U19781 : BUF_X1 port map( A => n22763, Z => n26929);
   U19782 : BUF_X1 port map( A => n22763, Z => n26930);
   U19783 : BUF_X1 port map( A => n22763, Z => n26931);
   U19784 : BUF_X1 port map( A => n22761, Z => n26940);
   U19785 : BUF_X1 port map( A => n22761, Z => n26941);
   U19786 : BUF_X1 port map( A => n22761, Z => n26942);
   U19787 : BUF_X1 port map( A => n22761, Z => n26943);
   U19788 : BUF_X1 port map( A => n22725, Z => n27144);
   U19789 : BUF_X1 port map( A => n22725, Z => n27145);
   U19790 : BUF_X1 port map( A => n22725, Z => n27146);
   U19791 : BUF_X1 port map( A => n22725, Z => n27147);
   U19792 : BUF_X1 port map( A => n22748, Z => n27012);
   U19793 : BUF_X1 port map( A => n22748, Z => n27013);
   U19794 : BUF_X1 port map( A => n22748, Z => n27014);
   U19795 : BUF_X1 port map( A => n22748, Z => n27015);
   U19796 : BUF_X1 port map( A => n22738, Z => n27072);
   U19797 : BUF_X1 port map( A => n22738, Z => n27073);
   U19798 : BUF_X1 port map( A => n22738, Z => n27074);
   U19799 : BUF_X1 port map( A => n22738, Z => n27075);
   U19800 : BUF_X1 port map( A => n22740, Z => n27060);
   U19801 : BUF_X1 port map( A => n22740, Z => n27061);
   U19802 : BUF_X1 port map( A => n22740, Z => n27062);
   U19803 : BUF_X1 port map( A => n22740, Z => n27063);
   U19804 : BUF_X1 port map( A => n22757, Z => n26964);
   U19805 : BUF_X1 port map( A => n22757, Z => n26965);
   U19806 : BUF_X1 port map( A => n22757, Z => n26966);
   U19807 : BUF_X1 port map( A => n22757, Z => n26967);
   U19808 : BUF_X1 port map( A => n22750, Z => n27000);
   U19809 : BUF_X1 port map( A => n22750, Z => n27001);
   U19810 : BUF_X1 port map( A => n22750, Z => n27002);
   U19811 : BUF_X1 port map( A => n22750, Z => n27003);
   U19812 : BUF_X1 port map( A => n22735, Z => n27084);
   U19813 : BUF_X1 port map( A => n22735, Z => n27085);
   U19814 : BUF_X1 port map( A => n22735, Z => n27086);
   U19815 : BUF_X1 port map( A => n22735, Z => n27087);
   U19816 : BUF_X1 port map( A => n22755, Z => n26976);
   U19817 : BUF_X1 port map( A => n22755, Z => n26977);
   U19818 : BUF_X1 port map( A => n22755, Z => n26978);
   U19819 : BUF_X1 port map( A => n22755, Z => n26979);
   U19820 : BUF_X1 port map( A => n22729, Z => n27120);
   U19821 : BUF_X1 port map( A => n22729, Z => n27121);
   U19822 : BUF_X1 port map( A => n22729, Z => n27122);
   U19823 : BUF_X1 port map( A => n22729, Z => n27123);
   U19824 : BUF_X1 port map( A => n22733, Z => n27096);
   U19825 : BUF_X1 port map( A => n22733, Z => n27097);
   U19826 : BUF_X1 port map( A => n22733, Z => n27098);
   U19827 : BUF_X1 port map( A => n22733, Z => n27099);
   U19828 : BUF_X1 port map( A => n22744, Z => n27036);
   U19829 : BUF_X1 port map( A => n22744, Z => n27037);
   U19830 : BUF_X1 port map( A => n22744, Z => n27038);
   U19831 : BUF_X1 port map( A => n22744, Z => n27039);
   U19832 : BUF_X1 port map( A => n22746, Z => n27024);
   U19833 : BUF_X1 port map( A => n22746, Z => n27025);
   U19834 : BUF_X1 port map( A => n22746, Z => n27026);
   U19835 : BUF_X1 port map( A => n22746, Z => n27027);
   U19836 : BUF_X1 port map( A => n22767, Z => n26904);
   U19837 : BUF_X1 port map( A => n22767, Z => n26905);
   U19838 : BUF_X1 port map( A => n22767, Z => n26906);
   U19839 : BUF_X1 port map( A => n22767, Z => n26907);
   U19840 : BUF_X1 port map( A => n22765, Z => n26916);
   U19841 : BUF_X1 port map( A => n22765, Z => n26917);
   U19842 : BUF_X1 port map( A => n22765, Z => n26918);
   U19843 : BUF_X1 port map( A => n22765, Z => n26919);
   U19844 : BUF_X1 port map( A => n22731, Z => n27108);
   U19845 : BUF_X1 port map( A => n22731, Z => n27109);
   U19846 : BUF_X1 port map( A => n22731, Z => n27110);
   U19847 : BUF_X1 port map( A => n22731, Z => n27111);
   U19848 : BUF_X1 port map( A => n22727, Z => n27132);
   U19849 : BUF_X1 port map( A => n22727, Z => n27133);
   U19850 : BUF_X1 port map( A => n22727, Z => n27134);
   U19851 : BUF_X1 port map( A => n22727, Z => n27135);
   U19852 : NAND2_X1 port map( A1 => n25143, A2 => n25151, ZN => n23980);
   U19853 : NAND2_X1 port map( A1 => n23944, A2 => n23952, ZN => n22781);
   U19854 : NAND2_X1 port map( A1 => n27475, A2 => n27119, ZN => n22730);
   U19855 : NAND2_X1 port map( A1 => n27475, A2 => n27095, ZN => n22734);
   U19856 : NAND2_X1 port map( A1 => n27475, A2 => n27035, ZN => n22745);
   U19857 : NAND2_X1 port map( A1 => n27475, A2 => n27023, ZN => n22747);
   U19858 : BUF_X1 port map( A => n23990, Z => n26588);
   U19859 : BUF_X1 port map( A => n23985, Z => n26612);
   U19860 : BUF_X1 port map( A => n23975, Z => n26660);
   U19861 : BUF_X1 port map( A => n24005, Z => n26513);
   U19862 : BUF_X1 port map( A => n24000, Z => n26558);
   U19863 : BUF_X1 port map( A => n23990, Z => n26589);
   U19864 : BUF_X1 port map( A => n23985, Z => n26613);
   U19865 : BUF_X1 port map( A => n23975, Z => n26661);
   U19866 : BUF_X1 port map( A => n24005, Z => n26514);
   U19867 : BUF_X1 port map( A => n24000, Z => n26559);
   U19868 : BUF_X1 port map( A => n23990, Z => n26590);
   U19869 : BUF_X1 port map( A => n23985, Z => n26614);
   U19870 : BUF_X1 port map( A => n23975, Z => n26662);
   U19871 : BUF_X1 port map( A => n24005, Z => n26515);
   U19872 : BUF_X1 port map( A => n24000, Z => n26560);
   U19873 : BUF_X1 port map( A => n23990, Z => n26591);
   U19874 : BUF_X1 port map( A => n23985, Z => n26615);
   U19875 : BUF_X1 port map( A => n23975, Z => n26663);
   U19876 : BUF_X1 port map( A => n24005, Z => n26516);
   U19877 : BUF_X1 port map( A => n24000, Z => n26561);
   U19878 : BUF_X1 port map( A => n23990, Z => n26592);
   U19879 : BUF_X1 port map( A => n23985, Z => n26616);
   U19880 : BUF_X1 port map( A => n23975, Z => n26664);
   U19881 : BUF_X1 port map( A => n24005, Z => n26517);
   U19882 : BUF_X1 port map( A => n24000, Z => n26562);
   U19883 : BUF_X1 port map( A => n22791, Z => n26813);
   U19884 : BUF_X1 port map( A => n22786, Z => n26837);
   U19885 : BUF_X1 port map( A => n22776, Z => n26885);
   U19886 : BUF_X1 port map( A => n22806, Z => n26738);
   U19887 : BUF_X1 port map( A => n22801, Z => n26783);
   U19888 : BUF_X1 port map( A => n22791, Z => n26814);
   U19889 : BUF_X1 port map( A => n22786, Z => n26838);
   U19890 : BUF_X1 port map( A => n22776, Z => n26886);
   U19891 : BUF_X1 port map( A => n22806, Z => n26739);
   U19892 : BUF_X1 port map( A => n22801, Z => n26784);
   U19893 : BUF_X1 port map( A => n22791, Z => n26815);
   U19894 : BUF_X1 port map( A => n22786, Z => n26839);
   U19895 : BUF_X1 port map( A => n22776, Z => n26887);
   U19896 : BUF_X1 port map( A => n22806, Z => n26740);
   U19897 : BUF_X1 port map( A => n22801, Z => n26785);
   U19898 : BUF_X1 port map( A => n22791, Z => n26816);
   U19899 : BUF_X1 port map( A => n22786, Z => n26840);
   U19900 : BUF_X1 port map( A => n22776, Z => n26888);
   U19901 : BUF_X1 port map( A => n22806, Z => n26741);
   U19902 : BUF_X1 port map( A => n22801, Z => n26786);
   U19903 : BUF_X1 port map( A => n22791, Z => n26817);
   U19904 : BUF_X1 port map( A => n22786, Z => n26841);
   U19905 : BUF_X1 port map( A => n22776, Z => n26889);
   U19906 : BUF_X1 port map( A => n22806, Z => n26742);
   U19907 : BUF_X1 port map( A => n22801, Z => n26787);
   U19908 : BUF_X1 port map( A => n23989, Z => n26594);
   U19909 : BUF_X1 port map( A => n23984, Z => n26618);
   U19910 : BUF_X1 port map( A => n23974, Z => n26666);
   U19911 : BUF_X1 port map( A => n23979, Z => n26642);
   U19912 : BUF_X1 port map( A => n24004, Z => n26519);
   U19913 : BUF_X1 port map( A => n23999, Z => n26564);
   U19914 : BUF_X1 port map( A => n22790, Z => n26819);
   U19915 : BUF_X1 port map( A => n22785, Z => n26843);
   U19916 : BUF_X1 port map( A => n22775, Z => n26891);
   U19917 : BUF_X1 port map( A => n22780, Z => n26867);
   U19918 : BUF_X1 port map( A => n22805, Z => n26744);
   U19919 : BUF_X1 port map( A => n22800, Z => n26789);
   U19920 : NAND2_X1 port map( A1 => n27476, A2 => n26951, ZN => n22760);
   U19921 : NAND2_X1 port map( A1 => n27476, A2 => n26987, ZN => n22753);
   U19922 : NAND2_X1 port map( A1 => n27476, A2 => n26927, ZN => n22764);
   U19923 : NAND2_X1 port map( A1 => n27476, A2 => n26939, ZN => n22762);
   U19924 : NAND2_X1 port map( A1 => n27476, A2 => n26963, ZN => n22758);
   U19925 : NAND2_X1 port map( A1 => n27476, A2 => n26975, ZN => n22756);
   U19926 : NAND2_X1 port map( A1 => n27476, A2 => n26903, ZN => n22768);
   U19927 : NAND2_X1 port map( A1 => n27476, A2 => n26915, ZN => n22766);
   U19928 : NAND2_X1 port map( A1 => n27474, A2 => n27263, ZN => n22697);
   U19929 : NAND2_X1 port map( A1 => n27474, A2 => n27251, ZN => n22700);
   U19930 : NAND2_X1 port map( A1 => n27474, A2 => n27239, ZN => n22703);
   U19931 : NAND2_X1 port map( A1 => n27474, A2 => n27167, ZN => n22722);
   U19932 : NAND2_X1 port map( A1 => n27474, A2 => n27179, ZN => n22719);
   U19933 : NAND2_X1 port map( A1 => n27474, A2 => n27155, ZN => n22724);
   U19934 : NAND2_X1 port map( A1 => n27475, A2 => n27047, ZN => n22743);
   U19935 : NAND2_X1 port map( A1 => n27474, A2 => n27277, ZN => n22693);
   U19936 : NAND2_X1 port map( A1 => n27474, A2 => n27143, ZN => n22726);
   U19937 : NAND2_X1 port map( A1 => n27475, A2 => n27011, ZN => n22749);
   U19938 : NAND2_X1 port map( A1 => n27475, A2 => n27071, ZN => n22739);
   U19939 : NAND2_X1 port map( A1 => n27475, A2 => n27059, ZN => n22741);
   U19940 : NAND2_X1 port map( A1 => n27475, A2 => n26999, ZN => n22751);
   U19941 : NAND2_X1 port map( A1 => n27475, A2 => n27083, ZN => n22736);
   U19942 : NAND2_X1 port map( A1 => n27474, A2 => n27191, ZN => n22715);
   U19943 : NAND2_X1 port map( A1 => n27474, A2 => n27227, ZN => n22706);
   U19944 : NAND2_X1 port map( A1 => n27474, A2 => n27203, ZN => n22712);
   U19945 : NAND2_X1 port map( A1 => n27474, A2 => n27215, ZN => n22709);
   U19946 : NAND2_X1 port map( A1 => n27475, A2 => n27107, ZN => n22732);
   U19947 : NAND2_X1 port map( A1 => n27475, A2 => n27131, ZN => n22728);
   U19948 : BUF_X1 port map( A => n22692, Z => n27275);
   U19949 : BUF_X1 port map( A => n22692, Z => n27276);
   U19950 : BUF_X1 port map( A => n26531, Z => n26529);
   U19951 : BUF_X1 port map( A => n26531, Z => n26528);
   U19952 : BUF_X1 port map( A => n26532, Z => n26527);
   U19953 : BUF_X1 port map( A => n26532, Z => n26526);
   U19954 : BUF_X1 port map( A => n26532, Z => n26525);
   U19955 : BUF_X1 port map( A => n26756, Z => n26754);
   U19956 : BUF_X1 port map( A => n26756, Z => n26753);
   U19957 : BUF_X1 port map( A => n26757, Z => n26751);
   U19958 : BUF_X1 port map( A => n26757, Z => n26750);
   U19959 : BUF_X1 port map( A => n26757, Z => n26752);
   U19960 : BUF_X1 port map( A => n26531, Z => n26530);
   U19961 : BUF_X1 port map( A => n26756, Z => n26755);
   U19962 : OAI22_X1 port map( A1 => n27318, A2 => n27168, B1 => n27162, B2 => 
                           n22679, ZN => n7438);
   U19963 : OAI22_X1 port map( A1 => n27321, A2 => n27168, B1 => n27162, B2 => 
                           n22678, ZN => n7439);
   U19964 : OAI22_X1 port map( A1 => n27324, A2 => n27168, B1 => n27162, B2 => 
                           n22677, ZN => n7440);
   U19965 : OAI22_X1 port map( A1 => n27327, A2 => n27168, B1 => n27162, B2 => 
                           n22676, ZN => n7441);
   U19966 : OAI22_X1 port map( A1 => n27330, A2 => n27168, B1 => n27162, B2 => 
                           n22675, ZN => n7442);
   U19967 : OAI22_X1 port map( A1 => n27333, A2 => n27168, B1 => n27162, B2 => 
                           n22674, ZN => n7443);
   U19968 : OAI22_X1 port map( A1 => n27336, A2 => n27168, B1 => n27162, B2 => 
                           n22673, ZN => n7444);
   U19969 : OAI22_X1 port map( A1 => n27339, A2 => n27168, B1 => n27162, B2 => 
                           n22672, ZN => n7445);
   U19970 : OAI22_X1 port map( A1 => n27342, A2 => n27168, B1 => n27162, B2 => 
                           n22671, ZN => n7446);
   U19971 : OAI22_X1 port map( A1 => n27345, A2 => n27168, B1 => n27162, B2 => 
                           n22670, ZN => n7447);
   U19972 : OAI22_X1 port map( A1 => n27348, A2 => n27168, B1 => n27162, B2 => 
                           n22669, ZN => n7448);
   U19973 : OAI22_X1 port map( A1 => n27351, A2 => n27169, B1 => n27162, B2 => 
                           n22668, ZN => n7449);
   U19974 : OAI22_X1 port map( A1 => n27354, A2 => n27169, B1 => n27163, B2 => 
                           n22667, ZN => n7450);
   U19975 : OAI22_X1 port map( A1 => n27357, A2 => n27169, B1 => n27163, B2 => 
                           n22666, ZN => n7451);
   U19976 : OAI22_X1 port map( A1 => n27360, A2 => n27169, B1 => n27163, B2 => 
                           n22665, ZN => n7452);
   U19977 : OAI22_X1 port map( A1 => n27363, A2 => n27169, B1 => n27163, B2 => 
                           n22664, ZN => n7453);
   U19978 : OAI22_X1 port map( A1 => n27366, A2 => n27169, B1 => n27163, B2 => 
                           n22663, ZN => n7454);
   U19979 : OAI22_X1 port map( A1 => n27369, A2 => n27169, B1 => n27163, B2 => 
                           n22662, ZN => n7455);
   U19980 : OAI22_X1 port map( A1 => n27372, A2 => n27169, B1 => n27163, B2 => 
                           n22661, ZN => n7456);
   U19981 : OAI22_X1 port map( A1 => n27375, A2 => n27169, B1 => n27163, B2 => 
                           n22660, ZN => n7457);
   U19982 : OAI22_X1 port map( A1 => n27378, A2 => n27169, B1 => n27163, B2 => 
                           n22659, ZN => n7458);
   U19983 : OAI22_X1 port map( A1 => n27381, A2 => n27169, B1 => n27163, B2 => 
                           n22658, ZN => n7459);
   U19984 : OAI22_X1 port map( A1 => n27384, A2 => n27169, B1 => n27163, B2 => 
                           n22657, ZN => n7460);
   U19985 : OAI22_X1 port map( A1 => n27387, A2 => n27170, B1 => n27163, B2 => 
                           n22656, ZN => n7461);
   U19986 : OAI22_X1 port map( A1 => n27390, A2 => n27170, B1 => n27164, B2 => 
                           n22655, ZN => n7462);
   U19987 : OAI22_X1 port map( A1 => n27393, A2 => n27170, B1 => n27164, B2 => 
                           n22654, ZN => n7463);
   U19988 : OAI22_X1 port map( A1 => n27396, A2 => n27170, B1 => n27164, B2 => 
                           n22653, ZN => n7464);
   U19989 : OAI22_X1 port map( A1 => n27399, A2 => n27170, B1 => n27164, B2 => 
                           n22652, ZN => n7465);
   U19990 : OAI22_X1 port map( A1 => n27402, A2 => n27170, B1 => n27164, B2 => 
                           n22651, ZN => n7466);
   U19991 : OAI22_X1 port map( A1 => n27405, A2 => n27170, B1 => n27164, B2 => 
                           n22650, ZN => n7467);
   U19992 : OAI22_X1 port map( A1 => n27408, A2 => n27170, B1 => n27164, B2 => 
                           n22649, ZN => n7468);
   U19993 : OAI22_X1 port map( A1 => n27411, A2 => n27170, B1 => n27164, B2 => 
                           n22648, ZN => n7469);
   U19994 : OAI22_X1 port map( A1 => n27414, A2 => n27170, B1 => n27164, B2 => 
                           n22647, ZN => n7470);
   U19995 : OAI22_X1 port map( A1 => n27417, A2 => n27170, B1 => n27164, B2 => 
                           n22646, ZN => n7471);
   U19996 : OAI22_X1 port map( A1 => n27420, A2 => n27170, B1 => n27164, B2 => 
                           n22645, ZN => n7472);
   U19997 : OAI22_X1 port map( A1 => n27423, A2 => n27171, B1 => n27164, B2 => 
                           n22644, ZN => n7473);
   U19998 : OAI22_X1 port map( A1 => n27426, A2 => n27171, B1 => n27165, B2 => 
                           n22643, ZN => n7474);
   U19999 : OAI22_X1 port map( A1 => n27429, A2 => n27171, B1 => n27165, B2 => 
                           n22642, ZN => n7475);
   U20000 : OAI22_X1 port map( A1 => n27432, A2 => n27171, B1 => n27165, B2 => 
                           n22641, ZN => n7476);
   U20001 : OAI22_X1 port map( A1 => n27435, A2 => n27171, B1 => n27165, B2 => 
                           n22640, ZN => n7477);
   U20002 : OAI22_X1 port map( A1 => n27438, A2 => n27171, B1 => n27165, B2 => 
                           n22639, ZN => n7478);
   U20003 : OAI22_X1 port map( A1 => n27441, A2 => n27171, B1 => n27165, B2 => 
                           n22638, ZN => n7479);
   U20004 : OAI22_X1 port map( A1 => n27444, A2 => n27171, B1 => n27165, B2 => 
                           n22637, ZN => n7480);
   U20005 : OAI22_X1 port map( A1 => n27447, A2 => n27171, B1 => n27165, B2 => 
                           n22636, ZN => n7481);
   U20006 : OAI22_X1 port map( A1 => n27450, A2 => n27171, B1 => n27165, B2 => 
                           n22635, ZN => n7482);
   U20007 : OAI22_X1 port map( A1 => n27453, A2 => n27171, B1 => n27165, B2 => 
                           n22634, ZN => n7483);
   U20008 : OAI22_X1 port map( A1 => n27456, A2 => n27171, B1 => n27165, B2 => 
                           n22633, ZN => n7484);
   U20009 : OAI22_X1 port map( A1 => n27459, A2 => n27172, B1 => n27165, B2 => 
                           n22632, ZN => n7485);
   U20010 : OAI22_X1 port map( A1 => n27319, A2 => n26988, B1 => n26982, B2 => 
                           n22559, ZN => n6478);
   U20011 : OAI22_X1 port map( A1 => n27322, A2 => n26988, B1 => n26982, B2 => 
                           n22558, ZN => n6479);
   U20012 : OAI22_X1 port map( A1 => n27325, A2 => n26988, B1 => n26982, B2 => 
                           n22557, ZN => n6480);
   U20013 : OAI22_X1 port map( A1 => n27328, A2 => n26988, B1 => n26982, B2 => 
                           n22556, ZN => n6481);
   U20014 : OAI22_X1 port map( A1 => n27331, A2 => n26988, B1 => n26982, B2 => 
                           n22555, ZN => n6482);
   U20015 : OAI22_X1 port map( A1 => n27334, A2 => n26988, B1 => n26982, B2 => 
                           n22554, ZN => n6483);
   U20016 : OAI22_X1 port map( A1 => n27337, A2 => n26988, B1 => n26982, B2 => 
                           n22553, ZN => n6484);
   U20017 : OAI22_X1 port map( A1 => n27340, A2 => n26988, B1 => n26982, B2 => 
                           n22552, ZN => n6485);
   U20018 : OAI22_X1 port map( A1 => n27343, A2 => n26988, B1 => n26982, B2 => 
                           n22551, ZN => n6486);
   U20019 : OAI22_X1 port map( A1 => n27346, A2 => n26988, B1 => n26982, B2 => 
                           n22550, ZN => n6487);
   U20020 : OAI22_X1 port map( A1 => n27349, A2 => n26988, B1 => n26982, B2 => 
                           n22549, ZN => n6488);
   U20021 : OAI22_X1 port map( A1 => n27352, A2 => n26989, B1 => n26982, B2 => 
                           n22548, ZN => n6489);
   U20022 : OAI22_X1 port map( A1 => n27355, A2 => n26989, B1 => n26983, B2 => 
                           n22547, ZN => n6490);
   U20023 : OAI22_X1 port map( A1 => n27358, A2 => n26989, B1 => n26983, B2 => 
                           n22546, ZN => n6491);
   U20024 : OAI22_X1 port map( A1 => n27361, A2 => n26989, B1 => n26983, B2 => 
                           n22545, ZN => n6492);
   U20025 : OAI22_X1 port map( A1 => n27364, A2 => n26989, B1 => n26983, B2 => 
                           n22544, ZN => n6493);
   U20026 : OAI22_X1 port map( A1 => n27367, A2 => n26989, B1 => n26983, B2 => 
                           n22543, ZN => n6494);
   U20027 : OAI22_X1 port map( A1 => n27370, A2 => n26989, B1 => n26983, B2 => 
                           n22542, ZN => n6495);
   U20028 : OAI22_X1 port map( A1 => n27373, A2 => n26989, B1 => n26983, B2 => 
                           n22541, ZN => n6496);
   U20029 : OAI22_X1 port map( A1 => n27376, A2 => n26989, B1 => n26983, B2 => 
                           n22540, ZN => n6497);
   U20030 : OAI22_X1 port map( A1 => n27379, A2 => n26989, B1 => n26983, B2 => 
                           n22539, ZN => n6498);
   U20031 : OAI22_X1 port map( A1 => n27382, A2 => n26989, B1 => n26983, B2 => 
                           n22538, ZN => n6499);
   U20032 : OAI22_X1 port map( A1 => n27385, A2 => n26989, B1 => n26983, B2 => 
                           n22537, ZN => n6500);
   U20033 : OAI22_X1 port map( A1 => n27388, A2 => n26990, B1 => n26983, B2 => 
                           n22536, ZN => n6501);
   U20034 : OAI22_X1 port map( A1 => n27391, A2 => n26990, B1 => n26984, B2 => 
                           n22535, ZN => n6502);
   U20035 : OAI22_X1 port map( A1 => n27394, A2 => n26990, B1 => n26984, B2 => 
                           n22534, ZN => n6503);
   U20036 : OAI22_X1 port map( A1 => n27397, A2 => n26990, B1 => n26984, B2 => 
                           n22533, ZN => n6504);
   U20037 : OAI22_X1 port map( A1 => n27400, A2 => n26990, B1 => n26984, B2 => 
                           n22532, ZN => n6505);
   U20038 : OAI22_X1 port map( A1 => n27403, A2 => n26990, B1 => n26984, B2 => 
                           n22531, ZN => n6506);
   U20039 : OAI22_X1 port map( A1 => n27406, A2 => n26990, B1 => n26984, B2 => 
                           n22530, ZN => n6507);
   U20040 : OAI22_X1 port map( A1 => n27409, A2 => n26990, B1 => n26984, B2 => 
                           n22529, ZN => n6508);
   U20041 : OAI22_X1 port map( A1 => n27412, A2 => n26990, B1 => n26984, B2 => 
                           n22528, ZN => n6509);
   U20042 : OAI22_X1 port map( A1 => n27415, A2 => n26990, B1 => n26984, B2 => 
                           n22527, ZN => n6510);
   U20043 : OAI22_X1 port map( A1 => n27418, A2 => n26990, B1 => n26984, B2 => 
                           n22526, ZN => n6511);
   U20044 : OAI22_X1 port map( A1 => n27421, A2 => n26990, B1 => n26984, B2 => 
                           n22525, ZN => n6512);
   U20045 : OAI22_X1 port map( A1 => n27424, A2 => n26991, B1 => n26984, B2 => 
                           n22524, ZN => n6513);
   U20046 : OAI22_X1 port map( A1 => n27427, A2 => n26991, B1 => n26985, B2 => 
                           n22523, ZN => n6514);
   U20047 : OAI22_X1 port map( A1 => n27430, A2 => n26991, B1 => n26985, B2 => 
                           n22522, ZN => n6515);
   U20048 : OAI22_X1 port map( A1 => n27433, A2 => n26991, B1 => n26985, B2 => 
                           n22521, ZN => n6516);
   U20049 : OAI22_X1 port map( A1 => n27436, A2 => n26991, B1 => n26985, B2 => 
                           n22520, ZN => n6517);
   U20050 : OAI22_X1 port map( A1 => n27439, A2 => n26991, B1 => n26985, B2 => 
                           n22519, ZN => n6518);
   U20051 : OAI22_X1 port map( A1 => n27442, A2 => n26991, B1 => n26985, B2 => 
                           n22518, ZN => n6519);
   U20052 : OAI22_X1 port map( A1 => n27445, A2 => n26991, B1 => n26985, B2 => 
                           n22517, ZN => n6520);
   U20053 : OAI22_X1 port map( A1 => n27448, A2 => n26991, B1 => n26985, B2 => 
                           n22516, ZN => n6521);
   U20054 : OAI22_X1 port map( A1 => n27451, A2 => n26991, B1 => n26985, B2 => 
                           n22515, ZN => n6522);
   U20055 : OAI22_X1 port map( A1 => n27454, A2 => n26991, B1 => n26985, B2 => 
                           n22514, ZN => n6523);
   U20056 : OAI22_X1 port map( A1 => n27457, A2 => n26991, B1 => n26985, B2 => 
                           n22513, ZN => n6524);
   U20057 : OAI22_X1 port map( A1 => n27460, A2 => n26992, B1 => n26985, B2 => 
                           n22512, ZN => n6525);
   U20058 : OAI22_X1 port map( A1 => n27318, A2 => n27180, B1 => n27174, B2 => 
                           n22487, ZN => n7502);
   U20059 : OAI22_X1 port map( A1 => n27321, A2 => n27180, B1 => n27174, B2 => 
                           n22486, ZN => n7503);
   U20060 : OAI22_X1 port map( A1 => n27324, A2 => n27180, B1 => n27174, B2 => 
                           n22485, ZN => n7504);
   U20061 : OAI22_X1 port map( A1 => n27327, A2 => n27180, B1 => n27174, B2 => 
                           n22484, ZN => n7505);
   U20062 : OAI22_X1 port map( A1 => n27330, A2 => n27180, B1 => n27174, B2 => 
                           n22483, ZN => n7506);
   U20063 : OAI22_X1 port map( A1 => n27333, A2 => n27180, B1 => n27174, B2 => 
                           n22482, ZN => n7507);
   U20064 : OAI22_X1 port map( A1 => n27336, A2 => n27180, B1 => n27174, B2 => 
                           n22481, ZN => n7508);
   U20065 : OAI22_X1 port map( A1 => n27339, A2 => n27180, B1 => n27174, B2 => 
                           n22480, ZN => n7509);
   U20066 : OAI22_X1 port map( A1 => n27342, A2 => n27180, B1 => n27174, B2 => 
                           n22479, ZN => n7510);
   U20067 : OAI22_X1 port map( A1 => n27345, A2 => n27180, B1 => n27174, B2 => 
                           n22478, ZN => n7511);
   U20068 : OAI22_X1 port map( A1 => n27348, A2 => n27180, B1 => n27174, B2 => 
                           n22477, ZN => n7512);
   U20069 : OAI22_X1 port map( A1 => n27351, A2 => n27181, B1 => n27174, B2 => 
                           n22476, ZN => n7513);
   U20070 : OAI22_X1 port map( A1 => n27354, A2 => n27181, B1 => n27175, B2 => 
                           n22475, ZN => n7514);
   U20071 : OAI22_X1 port map( A1 => n27357, A2 => n27181, B1 => n27175, B2 => 
                           n22474, ZN => n7515);
   U20072 : OAI22_X1 port map( A1 => n27360, A2 => n27181, B1 => n27175, B2 => 
                           n22473, ZN => n7516);
   U20073 : OAI22_X1 port map( A1 => n27363, A2 => n27181, B1 => n27175, B2 => 
                           n22472, ZN => n7517);
   U20074 : OAI22_X1 port map( A1 => n27366, A2 => n27181, B1 => n27175, B2 => 
                           n22471, ZN => n7518);
   U20075 : OAI22_X1 port map( A1 => n27369, A2 => n27181, B1 => n27175, B2 => 
                           n22470, ZN => n7519);
   U20076 : OAI22_X1 port map( A1 => n27372, A2 => n27181, B1 => n27175, B2 => 
                           n22469, ZN => n7520);
   U20077 : OAI22_X1 port map( A1 => n27375, A2 => n27181, B1 => n27175, B2 => 
                           n22468, ZN => n7521);
   U20078 : OAI22_X1 port map( A1 => n27378, A2 => n27181, B1 => n27175, B2 => 
                           n22467, ZN => n7522);
   U20079 : OAI22_X1 port map( A1 => n27381, A2 => n27181, B1 => n27175, B2 => 
                           n22466, ZN => n7523);
   U20080 : OAI22_X1 port map( A1 => n27384, A2 => n27181, B1 => n27175, B2 => 
                           n22465, ZN => n7524);
   U20081 : OAI22_X1 port map( A1 => n27387, A2 => n27182, B1 => n27175, B2 => 
                           n22464, ZN => n7525);
   U20082 : OAI22_X1 port map( A1 => n27390, A2 => n27182, B1 => n27176, B2 => 
                           n22463, ZN => n7526);
   U20083 : OAI22_X1 port map( A1 => n27393, A2 => n27182, B1 => n27176, B2 => 
                           n22462, ZN => n7527);
   U20084 : OAI22_X1 port map( A1 => n27396, A2 => n27182, B1 => n27176, B2 => 
                           n22461, ZN => n7528);
   U20085 : OAI22_X1 port map( A1 => n27399, A2 => n27182, B1 => n27176, B2 => 
                           n22460, ZN => n7529);
   U20086 : OAI22_X1 port map( A1 => n27402, A2 => n27182, B1 => n27176, B2 => 
                           n22459, ZN => n7530);
   U20087 : OAI22_X1 port map( A1 => n27405, A2 => n27182, B1 => n27176, B2 => 
                           n22458, ZN => n7531);
   U20088 : OAI22_X1 port map( A1 => n27408, A2 => n27182, B1 => n27176, B2 => 
                           n22457, ZN => n7532);
   U20089 : OAI22_X1 port map( A1 => n27411, A2 => n27182, B1 => n27176, B2 => 
                           n22456, ZN => n7533);
   U20090 : OAI22_X1 port map( A1 => n27414, A2 => n27182, B1 => n27176, B2 => 
                           n22455, ZN => n7534);
   U20091 : OAI22_X1 port map( A1 => n27417, A2 => n27182, B1 => n27176, B2 => 
                           n22454, ZN => n7535);
   U20092 : OAI22_X1 port map( A1 => n27420, A2 => n27182, B1 => n27176, B2 => 
                           n22453, ZN => n7536);
   U20093 : OAI22_X1 port map( A1 => n27423, A2 => n27183, B1 => n27176, B2 => 
                           n22452, ZN => n7537);
   U20094 : OAI22_X1 port map( A1 => n27426, A2 => n27183, B1 => n27177, B2 => 
                           n22451, ZN => n7538);
   U20095 : OAI22_X1 port map( A1 => n27429, A2 => n27183, B1 => n27177, B2 => 
                           n22450, ZN => n7539);
   U20096 : OAI22_X1 port map( A1 => n27432, A2 => n27183, B1 => n27177, B2 => 
                           n22449, ZN => n7540);
   U20097 : OAI22_X1 port map( A1 => n27435, A2 => n27183, B1 => n27177, B2 => 
                           n22448, ZN => n7541);
   U20098 : OAI22_X1 port map( A1 => n27438, A2 => n27183, B1 => n27177, B2 => 
                           n22447, ZN => n7542);
   U20099 : OAI22_X1 port map( A1 => n27441, A2 => n27183, B1 => n27177, B2 => 
                           n22446, ZN => n7543);
   U20100 : OAI22_X1 port map( A1 => n27444, A2 => n27183, B1 => n27177, B2 => 
                           n22445, ZN => n7544);
   U20101 : OAI22_X1 port map( A1 => n27447, A2 => n27183, B1 => n27177, B2 => 
                           n22444, ZN => n7545);
   U20102 : OAI22_X1 port map( A1 => n27450, A2 => n27183, B1 => n27177, B2 => 
                           n22443, ZN => n7546);
   U20103 : OAI22_X1 port map( A1 => n27453, A2 => n27183, B1 => n27177, B2 => 
                           n22442, ZN => n7547);
   U20104 : OAI22_X1 port map( A1 => n27456, A2 => n27183, B1 => n27177, B2 => 
                           n22441, ZN => n7548);
   U20105 : OAI22_X1 port map( A1 => n27459, A2 => n27184, B1 => n27177, B2 => 
                           n22440, ZN => n7549);
   U20106 : OAI22_X1 port map( A1 => n27319, A2 => n27048, B1 => n27042, B2 => 
                           n22367, ZN => n6798);
   U20107 : OAI22_X1 port map( A1 => n27322, A2 => n27048, B1 => n27042, B2 => 
                           n22366, ZN => n6799);
   U20108 : OAI22_X1 port map( A1 => n27325, A2 => n27048, B1 => n27042, B2 => 
                           n22365, ZN => n6800);
   U20109 : OAI22_X1 port map( A1 => n27328, A2 => n27048, B1 => n27042, B2 => 
                           n22364, ZN => n6801);
   U20110 : OAI22_X1 port map( A1 => n27331, A2 => n27048, B1 => n27042, B2 => 
                           n22363, ZN => n6802);
   U20111 : OAI22_X1 port map( A1 => n27334, A2 => n27048, B1 => n27042, B2 => 
                           n22362, ZN => n6803);
   U20112 : OAI22_X1 port map( A1 => n27337, A2 => n27048, B1 => n27042, B2 => 
                           n22361, ZN => n6804);
   U20113 : OAI22_X1 port map( A1 => n27340, A2 => n27048, B1 => n27042, B2 => 
                           n22360, ZN => n6805);
   U20114 : OAI22_X1 port map( A1 => n27343, A2 => n27048, B1 => n27042, B2 => 
                           n22359, ZN => n6806);
   U20115 : OAI22_X1 port map( A1 => n27346, A2 => n27048, B1 => n27042, B2 => 
                           n22358, ZN => n6807);
   U20116 : OAI22_X1 port map( A1 => n27349, A2 => n27048, B1 => n27042, B2 => 
                           n22357, ZN => n6808);
   U20117 : OAI22_X1 port map( A1 => n27352, A2 => n27049, B1 => n27042, B2 => 
                           n22356, ZN => n6809);
   U20118 : OAI22_X1 port map( A1 => n27355, A2 => n27049, B1 => n27043, B2 => 
                           n22355, ZN => n6810);
   U20119 : OAI22_X1 port map( A1 => n27358, A2 => n27049, B1 => n27043, B2 => 
                           n22354, ZN => n6811);
   U20120 : OAI22_X1 port map( A1 => n27361, A2 => n27049, B1 => n27043, B2 => 
                           n22353, ZN => n6812);
   U20121 : OAI22_X1 port map( A1 => n27364, A2 => n27049, B1 => n27043, B2 => 
                           n22352, ZN => n6813);
   U20122 : OAI22_X1 port map( A1 => n27367, A2 => n27049, B1 => n27043, B2 => 
                           n22351, ZN => n6814);
   U20123 : OAI22_X1 port map( A1 => n27370, A2 => n27049, B1 => n27043, B2 => 
                           n22350, ZN => n6815);
   U20124 : OAI22_X1 port map( A1 => n27373, A2 => n27049, B1 => n27043, B2 => 
                           n22349, ZN => n6816);
   U20125 : OAI22_X1 port map( A1 => n27376, A2 => n27049, B1 => n27043, B2 => 
                           n22348, ZN => n6817);
   U20126 : OAI22_X1 port map( A1 => n27379, A2 => n27049, B1 => n27043, B2 => 
                           n22347, ZN => n6818);
   U20127 : OAI22_X1 port map( A1 => n27382, A2 => n27049, B1 => n27043, B2 => 
                           n22346, ZN => n6819);
   U20128 : OAI22_X1 port map( A1 => n27385, A2 => n27049, B1 => n27043, B2 => 
                           n22345, ZN => n6820);
   U20129 : OAI22_X1 port map( A1 => n27388, A2 => n27050, B1 => n27043, B2 => 
                           n22344, ZN => n6821);
   U20130 : OAI22_X1 port map( A1 => n27391, A2 => n27050, B1 => n27044, B2 => 
                           n22343, ZN => n6822);
   U20131 : OAI22_X1 port map( A1 => n27394, A2 => n27050, B1 => n27044, B2 => 
                           n22342, ZN => n6823);
   U20132 : OAI22_X1 port map( A1 => n27397, A2 => n27050, B1 => n27044, B2 => 
                           n22341, ZN => n6824);
   U20133 : OAI22_X1 port map( A1 => n27400, A2 => n27050, B1 => n27044, B2 => 
                           n22340, ZN => n6825);
   U20134 : OAI22_X1 port map( A1 => n27403, A2 => n27050, B1 => n27044, B2 => 
                           n22339, ZN => n6826);
   U20135 : OAI22_X1 port map( A1 => n27406, A2 => n27050, B1 => n27044, B2 => 
                           n22338, ZN => n6827);
   U20136 : OAI22_X1 port map( A1 => n27409, A2 => n27050, B1 => n27044, B2 => 
                           n22337, ZN => n6828);
   U20137 : OAI22_X1 port map( A1 => n27412, A2 => n27050, B1 => n27044, B2 => 
                           n22336, ZN => n6829);
   U20138 : OAI22_X1 port map( A1 => n27415, A2 => n27050, B1 => n27044, B2 => 
                           n22335, ZN => n6830);
   U20139 : OAI22_X1 port map( A1 => n27418, A2 => n27050, B1 => n27044, B2 => 
                           n22334, ZN => n6831);
   U20140 : OAI22_X1 port map( A1 => n27421, A2 => n27050, B1 => n27044, B2 => 
                           n22333, ZN => n6832);
   U20141 : OAI22_X1 port map( A1 => n27424, A2 => n27051, B1 => n27044, B2 => 
                           n22332, ZN => n6833);
   U20142 : OAI22_X1 port map( A1 => n27427, A2 => n27051, B1 => n27045, B2 => 
                           n22331, ZN => n6834);
   U20143 : OAI22_X1 port map( A1 => n27430, A2 => n27051, B1 => n27045, B2 => 
                           n22330, ZN => n6835);
   U20144 : OAI22_X1 port map( A1 => n27433, A2 => n27051, B1 => n27045, B2 => 
                           n22329, ZN => n6836);
   U20145 : OAI22_X1 port map( A1 => n27436, A2 => n27051, B1 => n27045, B2 => 
                           n22328, ZN => n6837);
   U20146 : OAI22_X1 port map( A1 => n27439, A2 => n27051, B1 => n27045, B2 => 
                           n22327, ZN => n6838);
   U20147 : OAI22_X1 port map( A1 => n27442, A2 => n27051, B1 => n27045, B2 => 
                           n22326, ZN => n6839);
   U20148 : OAI22_X1 port map( A1 => n27445, A2 => n27051, B1 => n27045, B2 => 
                           n22325, ZN => n6840);
   U20149 : OAI22_X1 port map( A1 => n27448, A2 => n27051, B1 => n27045, B2 => 
                           n22324, ZN => n6841);
   U20150 : OAI22_X1 port map( A1 => n27451, A2 => n27051, B1 => n27045, B2 => 
                           n22323, ZN => n6842);
   U20151 : OAI22_X1 port map( A1 => n27454, A2 => n27051, B1 => n27045, B2 => 
                           n22322, ZN => n6843);
   U20152 : OAI22_X1 port map( A1 => n27457, A2 => n27051, B1 => n27045, B2 => 
                           n22321, ZN => n6844);
   U20153 : OAI22_X1 port map( A1 => n27460, A2 => n27052, B1 => n27045, B2 => 
                           n22320, ZN => n6845);
   U20154 : OAI22_X1 port map( A1 => n27318, A2 => n27192, B1 => n27186, B2 => 
                           n22047, ZN => n7566);
   U20155 : OAI22_X1 port map( A1 => n27321, A2 => n27192, B1 => n27186, B2 => 
                           n22046, ZN => n7567);
   U20156 : OAI22_X1 port map( A1 => n27324, A2 => n27192, B1 => n27186, B2 => 
                           n22045, ZN => n7568);
   U20157 : OAI22_X1 port map( A1 => n27327, A2 => n27192, B1 => n27186, B2 => 
                           n22044, ZN => n7569);
   U20158 : OAI22_X1 port map( A1 => n27330, A2 => n27192, B1 => n27186, B2 => 
                           n22043, ZN => n7570);
   U20159 : OAI22_X1 port map( A1 => n27333, A2 => n27192, B1 => n27186, B2 => 
                           n22042, ZN => n7571);
   U20160 : OAI22_X1 port map( A1 => n27336, A2 => n27192, B1 => n27186, B2 => 
                           n22041, ZN => n7572);
   U20161 : OAI22_X1 port map( A1 => n27339, A2 => n27192, B1 => n27186, B2 => 
                           n22040, ZN => n7573);
   U20162 : OAI22_X1 port map( A1 => n27342, A2 => n27192, B1 => n27186, B2 => 
                           n22039, ZN => n7574);
   U20163 : OAI22_X1 port map( A1 => n27345, A2 => n27192, B1 => n27186, B2 => 
                           n22038, ZN => n7575);
   U20164 : OAI22_X1 port map( A1 => n27348, A2 => n27192, B1 => n27186, B2 => 
                           n22037, ZN => n7576);
   U20165 : OAI22_X1 port map( A1 => n27351, A2 => n27193, B1 => n27186, B2 => 
                           n22036, ZN => n7577);
   U20166 : OAI22_X1 port map( A1 => n27354, A2 => n27193, B1 => n27187, B2 => 
                           n22035, ZN => n7578);
   U20167 : OAI22_X1 port map( A1 => n27357, A2 => n27193, B1 => n27187, B2 => 
                           n22034, ZN => n7579);
   U20168 : OAI22_X1 port map( A1 => n27360, A2 => n27193, B1 => n27187, B2 => 
                           n22033, ZN => n7580);
   U20169 : OAI22_X1 port map( A1 => n27363, A2 => n27193, B1 => n27187, B2 => 
                           n22032, ZN => n7581);
   U20170 : OAI22_X1 port map( A1 => n27366, A2 => n27193, B1 => n27187, B2 => 
                           n22031, ZN => n7582);
   U20171 : OAI22_X1 port map( A1 => n27369, A2 => n27193, B1 => n27187, B2 => 
                           n22030, ZN => n7583);
   U20172 : OAI22_X1 port map( A1 => n27372, A2 => n27193, B1 => n27187, B2 => 
                           n22029, ZN => n7584);
   U20173 : OAI22_X1 port map( A1 => n27375, A2 => n27193, B1 => n27187, B2 => 
                           n22028, ZN => n7585);
   U20174 : OAI22_X1 port map( A1 => n27378, A2 => n27193, B1 => n27187, B2 => 
                           n22027, ZN => n7586);
   U20175 : OAI22_X1 port map( A1 => n27381, A2 => n27193, B1 => n27187, B2 => 
                           n22026, ZN => n7587);
   U20176 : OAI22_X1 port map( A1 => n27384, A2 => n27193, B1 => n27187, B2 => 
                           n22025, ZN => n7588);
   U20177 : OAI22_X1 port map( A1 => n27387, A2 => n27194, B1 => n27187, B2 => 
                           n22024, ZN => n7589);
   U20178 : OAI22_X1 port map( A1 => n27390, A2 => n27194, B1 => n27188, B2 => 
                           n22023, ZN => n7590);
   U20179 : OAI22_X1 port map( A1 => n27393, A2 => n27194, B1 => n27188, B2 => 
                           n22022, ZN => n7591);
   U20180 : OAI22_X1 port map( A1 => n27396, A2 => n27194, B1 => n27188, B2 => 
                           n22021, ZN => n7592);
   U20181 : OAI22_X1 port map( A1 => n27399, A2 => n27194, B1 => n27188, B2 => 
                           n22020, ZN => n7593);
   U20182 : OAI22_X1 port map( A1 => n27402, A2 => n27194, B1 => n27188, B2 => 
                           n22019, ZN => n7594);
   U20183 : OAI22_X1 port map( A1 => n27405, A2 => n27194, B1 => n27188, B2 => 
                           n22018, ZN => n7595);
   U20184 : OAI22_X1 port map( A1 => n27408, A2 => n27194, B1 => n27188, B2 => 
                           n22017, ZN => n7596);
   U20185 : OAI22_X1 port map( A1 => n27411, A2 => n27194, B1 => n27188, B2 => 
                           n22016, ZN => n7597);
   U20186 : OAI22_X1 port map( A1 => n27414, A2 => n27194, B1 => n27188, B2 => 
                           n22015, ZN => n7598);
   U20187 : OAI22_X1 port map( A1 => n27417, A2 => n27194, B1 => n27188, B2 => 
                           n22014, ZN => n7599);
   U20188 : OAI22_X1 port map( A1 => n27420, A2 => n27194, B1 => n27188, B2 => 
                           n22013, ZN => n7600);
   U20189 : OAI22_X1 port map( A1 => n27423, A2 => n27195, B1 => n27188, B2 => 
                           n22012, ZN => n7601);
   U20190 : OAI22_X1 port map( A1 => n27426, A2 => n27195, B1 => n27189, B2 => 
                           n22011, ZN => n7602);
   U20191 : OAI22_X1 port map( A1 => n27429, A2 => n27195, B1 => n27189, B2 => 
                           n22010, ZN => n7603);
   U20192 : OAI22_X1 port map( A1 => n27432, A2 => n27195, B1 => n27189, B2 => 
                           n22009, ZN => n7604);
   U20193 : OAI22_X1 port map( A1 => n27435, A2 => n27195, B1 => n27189, B2 => 
                           n22008, ZN => n7605);
   U20194 : OAI22_X1 port map( A1 => n27438, A2 => n27195, B1 => n27189, B2 => 
                           n22007, ZN => n7606);
   U20195 : OAI22_X1 port map( A1 => n27441, A2 => n27195, B1 => n27189, B2 => 
                           n22006, ZN => n7607);
   U20196 : OAI22_X1 port map( A1 => n27444, A2 => n27195, B1 => n27189, B2 => 
                           n22005, ZN => n7608);
   U20197 : OAI22_X1 port map( A1 => n27447, A2 => n27195, B1 => n27189, B2 => 
                           n22004, ZN => n7609);
   U20198 : OAI22_X1 port map( A1 => n27450, A2 => n27195, B1 => n27189, B2 => 
                           n22003, ZN => n7610);
   U20199 : OAI22_X1 port map( A1 => n27453, A2 => n27195, B1 => n27189, B2 => 
                           n22002, ZN => n7611);
   U20200 : OAI22_X1 port map( A1 => n27456, A2 => n27195, B1 => n27189, B2 => 
                           n22001, ZN => n7612);
   U20201 : OAI22_X1 port map( A1 => n27459, A2 => n27196, B1 => n27189, B2 => 
                           n22000, ZN => n7613);
   U20202 : OAI22_X1 port map( A1 => n27318, A2 => n27144, B1 => n27138, B2 => 
                           n21987, ZN => n7310);
   U20203 : OAI22_X1 port map( A1 => n27321, A2 => n27144, B1 => n27138, B2 => 
                           n21986, ZN => n7311);
   U20204 : OAI22_X1 port map( A1 => n27324, A2 => n27144, B1 => n27138, B2 => 
                           n21985, ZN => n7312);
   U20205 : OAI22_X1 port map( A1 => n27327, A2 => n27144, B1 => n27138, B2 => 
                           n21984, ZN => n7313);
   U20206 : OAI22_X1 port map( A1 => n27330, A2 => n27144, B1 => n27138, B2 => 
                           n21983, ZN => n7314);
   U20207 : OAI22_X1 port map( A1 => n27333, A2 => n27144, B1 => n27138, B2 => 
                           n21982, ZN => n7315);
   U20208 : OAI22_X1 port map( A1 => n27336, A2 => n27144, B1 => n27138, B2 => 
                           n21981, ZN => n7316);
   U20209 : OAI22_X1 port map( A1 => n27339, A2 => n27144, B1 => n27138, B2 => 
                           n21980, ZN => n7317);
   U20210 : OAI22_X1 port map( A1 => n27342, A2 => n27144, B1 => n27138, B2 => 
                           n21979, ZN => n7318);
   U20211 : OAI22_X1 port map( A1 => n27345, A2 => n27144, B1 => n27138, B2 => 
                           n21978, ZN => n7319);
   U20212 : OAI22_X1 port map( A1 => n27348, A2 => n27144, B1 => n27138, B2 => 
                           n21977, ZN => n7320);
   U20213 : OAI22_X1 port map( A1 => n27351, A2 => n27145, B1 => n27138, B2 => 
                           n21976, ZN => n7321);
   U20214 : OAI22_X1 port map( A1 => n27354, A2 => n27145, B1 => n27139, B2 => 
                           n21975, ZN => n7322);
   U20215 : OAI22_X1 port map( A1 => n27357, A2 => n27145, B1 => n27139, B2 => 
                           n21974, ZN => n7323);
   U20216 : OAI22_X1 port map( A1 => n27360, A2 => n27145, B1 => n27139, B2 => 
                           n21973, ZN => n7324);
   U20217 : OAI22_X1 port map( A1 => n27363, A2 => n27145, B1 => n27139, B2 => 
                           n21972, ZN => n7325);
   U20218 : OAI22_X1 port map( A1 => n27366, A2 => n27145, B1 => n27139, B2 => 
                           n21971, ZN => n7326);
   U20219 : OAI22_X1 port map( A1 => n27369, A2 => n27145, B1 => n27139, B2 => 
                           n21970, ZN => n7327);
   U20220 : OAI22_X1 port map( A1 => n27372, A2 => n27145, B1 => n27139, B2 => 
                           n21969, ZN => n7328);
   U20221 : OAI22_X1 port map( A1 => n27375, A2 => n27145, B1 => n27139, B2 => 
                           n21968, ZN => n7329);
   U20222 : OAI22_X1 port map( A1 => n27378, A2 => n27145, B1 => n27139, B2 => 
                           n21967, ZN => n7330);
   U20223 : OAI22_X1 port map( A1 => n27381, A2 => n27145, B1 => n27139, B2 => 
                           n21966, ZN => n7331);
   U20224 : OAI22_X1 port map( A1 => n27384, A2 => n27145, B1 => n27139, B2 => 
                           n21965, ZN => n7332);
   U20225 : OAI22_X1 port map( A1 => n27387, A2 => n27146, B1 => n27139, B2 => 
                           n21964, ZN => n7333);
   U20226 : OAI22_X1 port map( A1 => n27390, A2 => n27146, B1 => n27140, B2 => 
                           n21963, ZN => n7334);
   U20227 : OAI22_X1 port map( A1 => n27393, A2 => n27146, B1 => n27140, B2 => 
                           n21962, ZN => n7335);
   U20228 : OAI22_X1 port map( A1 => n27396, A2 => n27146, B1 => n27140, B2 => 
                           n21961, ZN => n7336);
   U20229 : OAI22_X1 port map( A1 => n27399, A2 => n27146, B1 => n27140, B2 => 
                           n21960, ZN => n7337);
   U20230 : OAI22_X1 port map( A1 => n27402, A2 => n27146, B1 => n27140, B2 => 
                           n21959, ZN => n7338);
   U20231 : OAI22_X1 port map( A1 => n27405, A2 => n27146, B1 => n27140, B2 => 
                           n21958, ZN => n7339);
   U20232 : OAI22_X1 port map( A1 => n27408, A2 => n27146, B1 => n27140, B2 => 
                           n21957, ZN => n7340);
   U20233 : OAI22_X1 port map( A1 => n27411, A2 => n27146, B1 => n27140, B2 => 
                           n21956, ZN => n7341);
   U20234 : OAI22_X1 port map( A1 => n27414, A2 => n27146, B1 => n27140, B2 => 
                           n21955, ZN => n7342);
   U20235 : OAI22_X1 port map( A1 => n27417, A2 => n27146, B1 => n27140, B2 => 
                           n21954, ZN => n7343);
   U20236 : OAI22_X1 port map( A1 => n27420, A2 => n27146, B1 => n27140, B2 => 
                           n21953, ZN => n7344);
   U20237 : OAI22_X1 port map( A1 => n27423, A2 => n27147, B1 => n27140, B2 => 
                           n21952, ZN => n7345);
   U20238 : OAI22_X1 port map( A1 => n27426, A2 => n27147, B1 => n27141, B2 => 
                           n21951, ZN => n7346);
   U20239 : OAI22_X1 port map( A1 => n27429, A2 => n27147, B1 => n27141, B2 => 
                           n21950, ZN => n7347);
   U20240 : OAI22_X1 port map( A1 => n27432, A2 => n27147, B1 => n27141, B2 => 
                           n21949, ZN => n7348);
   U20241 : OAI22_X1 port map( A1 => n27435, A2 => n27147, B1 => n27141, B2 => 
                           n21948, ZN => n7349);
   U20242 : OAI22_X1 port map( A1 => n27438, A2 => n27147, B1 => n27141, B2 => 
                           n21947, ZN => n7350);
   U20243 : OAI22_X1 port map( A1 => n27441, A2 => n27147, B1 => n27141, B2 => 
                           n21946, ZN => n7351);
   U20244 : OAI22_X1 port map( A1 => n27444, A2 => n27147, B1 => n27141, B2 => 
                           n21945, ZN => n7352);
   U20245 : OAI22_X1 port map( A1 => n27447, A2 => n27147, B1 => n27141, B2 => 
                           n21944, ZN => n7353);
   U20246 : OAI22_X1 port map( A1 => n27450, A2 => n27147, B1 => n27141, B2 => 
                           n21943, ZN => n7354);
   U20247 : OAI22_X1 port map( A1 => n27453, A2 => n27147, B1 => n27141, B2 => 
                           n21942, ZN => n7355);
   U20248 : OAI22_X1 port map( A1 => n27456, A2 => n27147, B1 => n27141, B2 => 
                           n21941, ZN => n7356);
   U20249 : OAI22_X1 port map( A1 => n27459, A2 => n27148, B1 => n27141, B2 => 
                           n21940, ZN => n7357);
   U20250 : OAI22_X1 port map( A1 => n27319, A2 => n27072, B1 => n27066, B2 => 
                           n21747, ZN => n6926);
   U20251 : OAI22_X1 port map( A1 => n27322, A2 => n27072, B1 => n27066, B2 => 
                           n21746, ZN => n6927);
   U20252 : OAI22_X1 port map( A1 => n27325, A2 => n27072, B1 => n27066, B2 => 
                           n21745, ZN => n6928);
   U20253 : OAI22_X1 port map( A1 => n27328, A2 => n27072, B1 => n27066, B2 => 
                           n21744, ZN => n6929);
   U20254 : OAI22_X1 port map( A1 => n27331, A2 => n27072, B1 => n27066, B2 => 
                           n21743, ZN => n6930);
   U20255 : OAI22_X1 port map( A1 => n27334, A2 => n27072, B1 => n27066, B2 => 
                           n21742, ZN => n6931);
   U20256 : OAI22_X1 port map( A1 => n27337, A2 => n27072, B1 => n27066, B2 => 
                           n21741, ZN => n6932);
   U20257 : OAI22_X1 port map( A1 => n27340, A2 => n27072, B1 => n27066, B2 => 
                           n21740, ZN => n6933);
   U20258 : OAI22_X1 port map( A1 => n27343, A2 => n27072, B1 => n27066, B2 => 
                           n21739, ZN => n6934);
   U20259 : OAI22_X1 port map( A1 => n27346, A2 => n27072, B1 => n27066, B2 => 
                           n21738, ZN => n6935);
   U20260 : OAI22_X1 port map( A1 => n27349, A2 => n27072, B1 => n27066, B2 => 
                           n21737, ZN => n6936);
   U20261 : OAI22_X1 port map( A1 => n27352, A2 => n27073, B1 => n27066, B2 => 
                           n21736, ZN => n6937);
   U20262 : OAI22_X1 port map( A1 => n27355, A2 => n27073, B1 => n27067, B2 => 
                           n21735, ZN => n6938);
   U20263 : OAI22_X1 port map( A1 => n27358, A2 => n27073, B1 => n27067, B2 => 
                           n21734, ZN => n6939);
   U20264 : OAI22_X1 port map( A1 => n27361, A2 => n27073, B1 => n27067, B2 => 
                           n21733, ZN => n6940);
   U20265 : OAI22_X1 port map( A1 => n27364, A2 => n27073, B1 => n27067, B2 => 
                           n21732, ZN => n6941);
   U20266 : OAI22_X1 port map( A1 => n27367, A2 => n27073, B1 => n27067, B2 => 
                           n21731, ZN => n6942);
   U20267 : OAI22_X1 port map( A1 => n27370, A2 => n27073, B1 => n27067, B2 => 
                           n21730, ZN => n6943);
   U20268 : OAI22_X1 port map( A1 => n27373, A2 => n27073, B1 => n27067, B2 => 
                           n21729, ZN => n6944);
   U20269 : OAI22_X1 port map( A1 => n27376, A2 => n27073, B1 => n27067, B2 => 
                           n21728, ZN => n6945);
   U20270 : OAI22_X1 port map( A1 => n27379, A2 => n27073, B1 => n27067, B2 => 
                           n21727, ZN => n6946);
   U20271 : OAI22_X1 port map( A1 => n27382, A2 => n27073, B1 => n27067, B2 => 
                           n21726, ZN => n6947);
   U20272 : OAI22_X1 port map( A1 => n27385, A2 => n27073, B1 => n27067, B2 => 
                           n21725, ZN => n6948);
   U20273 : OAI22_X1 port map( A1 => n27388, A2 => n27074, B1 => n27067, B2 => 
                           n21724, ZN => n6949);
   U20274 : OAI22_X1 port map( A1 => n27391, A2 => n27074, B1 => n27068, B2 => 
                           n21723, ZN => n6950);
   U20275 : OAI22_X1 port map( A1 => n27394, A2 => n27074, B1 => n27068, B2 => 
                           n21722, ZN => n6951);
   U20276 : OAI22_X1 port map( A1 => n27397, A2 => n27074, B1 => n27068, B2 => 
                           n21721, ZN => n6952);
   U20277 : OAI22_X1 port map( A1 => n27400, A2 => n27074, B1 => n27068, B2 => 
                           n21720, ZN => n6953);
   U20278 : OAI22_X1 port map( A1 => n27403, A2 => n27074, B1 => n27068, B2 => 
                           n21719, ZN => n6954);
   U20279 : OAI22_X1 port map( A1 => n27406, A2 => n27074, B1 => n27068, B2 => 
                           n21718, ZN => n6955);
   U20280 : OAI22_X1 port map( A1 => n27409, A2 => n27074, B1 => n27068, B2 => 
                           n21717, ZN => n6956);
   U20281 : OAI22_X1 port map( A1 => n27412, A2 => n27074, B1 => n27068, B2 => 
                           n21716, ZN => n6957);
   U20282 : OAI22_X1 port map( A1 => n27415, A2 => n27074, B1 => n27068, B2 => 
                           n21715, ZN => n6958);
   U20283 : OAI22_X1 port map( A1 => n27418, A2 => n27074, B1 => n27068, B2 => 
                           n21714, ZN => n6959);
   U20284 : OAI22_X1 port map( A1 => n27421, A2 => n27074, B1 => n27068, B2 => 
                           n21713, ZN => n6960);
   U20285 : OAI22_X1 port map( A1 => n27424, A2 => n27075, B1 => n27068, B2 => 
                           n21712, ZN => n6961);
   U20286 : OAI22_X1 port map( A1 => n27427, A2 => n27075, B1 => n27069, B2 => 
                           n21711, ZN => n6962);
   U20287 : OAI22_X1 port map( A1 => n27430, A2 => n27075, B1 => n27069, B2 => 
                           n21710, ZN => n6963);
   U20288 : OAI22_X1 port map( A1 => n27433, A2 => n27075, B1 => n27069, B2 => 
                           n21709, ZN => n6964);
   U20289 : OAI22_X1 port map( A1 => n27436, A2 => n27075, B1 => n27069, B2 => 
                           n21708, ZN => n6965);
   U20290 : OAI22_X1 port map( A1 => n27439, A2 => n27075, B1 => n27069, B2 => 
                           n21707, ZN => n6966);
   U20291 : OAI22_X1 port map( A1 => n27442, A2 => n27075, B1 => n27069, B2 => 
                           n21706, ZN => n6967);
   U20292 : OAI22_X1 port map( A1 => n27445, A2 => n27075, B1 => n27069, B2 => 
                           n21705, ZN => n6968);
   U20293 : OAI22_X1 port map( A1 => n27448, A2 => n27075, B1 => n27069, B2 => 
                           n21704, ZN => n6969);
   U20294 : OAI22_X1 port map( A1 => n27451, A2 => n27075, B1 => n27069, B2 => 
                           n21703, ZN => n6970);
   U20295 : OAI22_X1 port map( A1 => n27454, A2 => n27075, B1 => n27069, B2 => 
                           n21702, ZN => n6971);
   U20296 : OAI22_X1 port map( A1 => n27457, A2 => n27075, B1 => n27069, B2 => 
                           n21701, ZN => n6972);
   U20297 : OAI22_X1 port map( A1 => n27460, A2 => n27076, B1 => n27069, B2 => 
                           n21700, ZN => n6973);
   U20298 : OAI22_X1 port map( A1 => n27320, A2 => n26964, B1 => n26958, B2 => 
                           n21627, ZN => n6350);
   U20299 : OAI22_X1 port map( A1 => n27323, A2 => n26964, B1 => n26958, B2 => 
                           n21626, ZN => n6351);
   U20300 : OAI22_X1 port map( A1 => n27326, A2 => n26964, B1 => n26958, B2 => 
                           n21625, ZN => n6352);
   U20301 : OAI22_X1 port map( A1 => n27329, A2 => n26964, B1 => n26958, B2 => 
                           n21624, ZN => n6353);
   U20302 : OAI22_X1 port map( A1 => n27332, A2 => n26964, B1 => n26958, B2 => 
                           n21623, ZN => n6354);
   U20303 : OAI22_X1 port map( A1 => n27335, A2 => n26964, B1 => n26958, B2 => 
                           n21622, ZN => n6355);
   U20304 : OAI22_X1 port map( A1 => n27338, A2 => n26964, B1 => n26958, B2 => 
                           n21621, ZN => n6356);
   U20305 : OAI22_X1 port map( A1 => n27341, A2 => n26964, B1 => n26958, B2 => 
                           n21620, ZN => n6357);
   U20306 : OAI22_X1 port map( A1 => n27344, A2 => n26964, B1 => n26958, B2 => 
                           n21619, ZN => n6358);
   U20307 : OAI22_X1 port map( A1 => n27347, A2 => n26964, B1 => n26958, B2 => 
                           n21618, ZN => n6359);
   U20308 : OAI22_X1 port map( A1 => n27350, A2 => n26964, B1 => n26958, B2 => 
                           n21617, ZN => n6360);
   U20309 : OAI22_X1 port map( A1 => n27353, A2 => n26965, B1 => n26958, B2 => 
                           n21616, ZN => n6361);
   U20310 : OAI22_X1 port map( A1 => n27356, A2 => n26965, B1 => n26959, B2 => 
                           n21615, ZN => n6362);
   U20311 : OAI22_X1 port map( A1 => n27359, A2 => n26965, B1 => n26959, B2 => 
                           n21614, ZN => n6363);
   U20312 : OAI22_X1 port map( A1 => n27362, A2 => n26965, B1 => n26959, B2 => 
                           n21613, ZN => n6364);
   U20313 : OAI22_X1 port map( A1 => n27365, A2 => n26965, B1 => n26959, B2 => 
                           n21612, ZN => n6365);
   U20314 : OAI22_X1 port map( A1 => n27368, A2 => n26965, B1 => n26959, B2 => 
                           n21611, ZN => n6366);
   U20315 : OAI22_X1 port map( A1 => n27371, A2 => n26965, B1 => n26959, B2 => 
                           n21610, ZN => n6367);
   U20316 : OAI22_X1 port map( A1 => n27374, A2 => n26965, B1 => n26959, B2 => 
                           n21609, ZN => n6368);
   U20317 : OAI22_X1 port map( A1 => n27377, A2 => n26965, B1 => n26959, B2 => 
                           n21608, ZN => n6369);
   U20318 : OAI22_X1 port map( A1 => n27380, A2 => n26965, B1 => n26959, B2 => 
                           n21607, ZN => n6370);
   U20319 : OAI22_X1 port map( A1 => n27383, A2 => n26965, B1 => n26959, B2 => 
                           n21606, ZN => n6371);
   U20320 : OAI22_X1 port map( A1 => n27386, A2 => n26965, B1 => n26959, B2 => 
                           n21605, ZN => n6372);
   U20321 : OAI22_X1 port map( A1 => n27389, A2 => n26966, B1 => n26959, B2 => 
                           n21604, ZN => n6373);
   U20322 : OAI22_X1 port map( A1 => n27392, A2 => n26966, B1 => n26960, B2 => 
                           n21603, ZN => n6374);
   U20323 : OAI22_X1 port map( A1 => n27395, A2 => n26966, B1 => n26960, B2 => 
                           n21602, ZN => n6375);
   U20324 : OAI22_X1 port map( A1 => n27398, A2 => n26966, B1 => n26960, B2 => 
                           n21601, ZN => n6376);
   U20325 : OAI22_X1 port map( A1 => n27401, A2 => n26966, B1 => n26960, B2 => 
                           n21600, ZN => n6377);
   U20326 : OAI22_X1 port map( A1 => n27404, A2 => n26966, B1 => n26960, B2 => 
                           n21599, ZN => n6378);
   U20327 : OAI22_X1 port map( A1 => n27407, A2 => n26966, B1 => n26960, B2 => 
                           n21598, ZN => n6379);
   U20328 : OAI22_X1 port map( A1 => n27410, A2 => n26966, B1 => n26960, B2 => 
                           n21597, ZN => n6380);
   U20329 : OAI22_X1 port map( A1 => n27413, A2 => n26966, B1 => n26960, B2 => 
                           n21596, ZN => n6381);
   U20330 : OAI22_X1 port map( A1 => n27416, A2 => n26966, B1 => n26960, B2 => 
                           n21595, ZN => n6382);
   U20331 : OAI22_X1 port map( A1 => n27419, A2 => n26966, B1 => n26960, B2 => 
                           n21594, ZN => n6383);
   U20332 : OAI22_X1 port map( A1 => n27422, A2 => n26966, B1 => n26960, B2 => 
                           n21593, ZN => n6384);
   U20333 : OAI22_X1 port map( A1 => n27425, A2 => n26967, B1 => n26960, B2 => 
                           n21592, ZN => n6385);
   U20334 : OAI22_X1 port map( A1 => n27428, A2 => n26967, B1 => n26961, B2 => 
                           n21591, ZN => n6386);
   U20335 : OAI22_X1 port map( A1 => n27431, A2 => n26967, B1 => n26961, B2 => 
                           n21590, ZN => n6387);
   U20336 : OAI22_X1 port map( A1 => n27434, A2 => n26967, B1 => n26961, B2 => 
                           n21589, ZN => n6388);
   U20337 : OAI22_X1 port map( A1 => n27437, A2 => n26967, B1 => n26961, B2 => 
                           n21588, ZN => n6389);
   U20338 : OAI22_X1 port map( A1 => n27440, A2 => n26967, B1 => n26961, B2 => 
                           n21587, ZN => n6390);
   U20339 : OAI22_X1 port map( A1 => n27443, A2 => n26967, B1 => n26961, B2 => 
                           n21586, ZN => n6391);
   U20340 : OAI22_X1 port map( A1 => n27446, A2 => n26967, B1 => n26961, B2 => 
                           n21585, ZN => n6392);
   U20341 : OAI22_X1 port map( A1 => n27449, A2 => n26967, B1 => n26961, B2 => 
                           n21584, ZN => n6393);
   U20342 : OAI22_X1 port map( A1 => n27452, A2 => n26967, B1 => n26961, B2 => 
                           n21583, ZN => n6394);
   U20343 : OAI22_X1 port map( A1 => n27455, A2 => n26967, B1 => n26961, B2 => 
                           n21582, ZN => n6395);
   U20344 : OAI22_X1 port map( A1 => n27458, A2 => n26967, B1 => n26961, B2 => 
                           n21581, ZN => n6396);
   U20345 : OAI22_X1 port map( A1 => n27461, A2 => n26968, B1 => n26961, B2 => 
                           n21580, ZN => n6397);
   U20346 : OAI22_X1 port map( A1 => n27318, A2 => n27216, B1 => n27210, B2 => 
                           n21567, ZN => n7694);
   U20347 : OAI22_X1 port map( A1 => n27321, A2 => n27216, B1 => n27210, B2 => 
                           n21566, ZN => n7695);
   U20348 : OAI22_X1 port map( A1 => n27324, A2 => n27216, B1 => n27210, B2 => 
                           n21565, ZN => n7696);
   U20349 : OAI22_X1 port map( A1 => n27327, A2 => n27216, B1 => n27210, B2 => 
                           n21564, ZN => n7697);
   U20350 : OAI22_X1 port map( A1 => n27330, A2 => n27216, B1 => n27210, B2 => 
                           n21563, ZN => n7698);
   U20351 : OAI22_X1 port map( A1 => n27333, A2 => n27216, B1 => n27210, B2 => 
                           n21562, ZN => n7699);
   U20352 : OAI22_X1 port map( A1 => n27336, A2 => n27216, B1 => n27210, B2 => 
                           n21561, ZN => n7700);
   U20353 : OAI22_X1 port map( A1 => n27339, A2 => n27216, B1 => n27210, B2 => 
                           n21560, ZN => n7701);
   U20354 : OAI22_X1 port map( A1 => n27342, A2 => n27216, B1 => n27210, B2 => 
                           n21559, ZN => n7702);
   U20355 : OAI22_X1 port map( A1 => n27345, A2 => n27216, B1 => n27210, B2 => 
                           n21558, ZN => n7703);
   U20356 : OAI22_X1 port map( A1 => n27348, A2 => n27216, B1 => n27210, B2 => 
                           n21557, ZN => n7704);
   U20357 : OAI22_X1 port map( A1 => n27351, A2 => n27217, B1 => n27210, B2 => 
                           n21556, ZN => n7705);
   U20358 : OAI22_X1 port map( A1 => n27354, A2 => n27217, B1 => n27211, B2 => 
                           n21555, ZN => n7706);
   U20359 : OAI22_X1 port map( A1 => n27357, A2 => n27217, B1 => n27211, B2 => 
                           n21554, ZN => n7707);
   U20360 : OAI22_X1 port map( A1 => n27360, A2 => n27217, B1 => n27211, B2 => 
                           n21553, ZN => n7708);
   U20361 : OAI22_X1 port map( A1 => n27363, A2 => n27217, B1 => n27211, B2 => 
                           n21552, ZN => n7709);
   U20362 : OAI22_X1 port map( A1 => n27366, A2 => n27217, B1 => n27211, B2 => 
                           n21551, ZN => n7710);
   U20363 : OAI22_X1 port map( A1 => n27369, A2 => n27217, B1 => n27211, B2 => 
                           n21550, ZN => n7711);
   U20364 : OAI22_X1 port map( A1 => n27372, A2 => n27217, B1 => n27211, B2 => 
                           n21549, ZN => n7712);
   U20365 : OAI22_X1 port map( A1 => n27375, A2 => n27217, B1 => n27211, B2 => 
                           n21548, ZN => n7713);
   U20366 : OAI22_X1 port map( A1 => n27378, A2 => n27217, B1 => n27211, B2 => 
                           n21547, ZN => n7714);
   U20367 : OAI22_X1 port map( A1 => n27381, A2 => n27217, B1 => n27211, B2 => 
                           n21546, ZN => n7715);
   U20368 : OAI22_X1 port map( A1 => n27384, A2 => n27217, B1 => n27211, B2 => 
                           n21545, ZN => n7716);
   U20369 : OAI22_X1 port map( A1 => n27387, A2 => n27218, B1 => n27211, B2 => 
                           n21544, ZN => n7717);
   U20370 : OAI22_X1 port map( A1 => n27390, A2 => n27218, B1 => n27212, B2 => 
                           n21543, ZN => n7718);
   U20371 : OAI22_X1 port map( A1 => n27393, A2 => n27218, B1 => n27212, B2 => 
                           n21542, ZN => n7719);
   U20372 : OAI22_X1 port map( A1 => n27396, A2 => n27218, B1 => n27212, B2 => 
                           n21541, ZN => n7720);
   U20373 : OAI22_X1 port map( A1 => n27399, A2 => n27218, B1 => n27212, B2 => 
                           n21540, ZN => n7721);
   U20374 : OAI22_X1 port map( A1 => n27402, A2 => n27218, B1 => n27212, B2 => 
                           n21539, ZN => n7722);
   U20375 : OAI22_X1 port map( A1 => n27405, A2 => n27218, B1 => n27212, B2 => 
                           n21538, ZN => n7723);
   U20376 : OAI22_X1 port map( A1 => n27408, A2 => n27218, B1 => n27212, B2 => 
                           n21537, ZN => n7724);
   U20377 : OAI22_X1 port map( A1 => n27411, A2 => n27218, B1 => n27212, B2 => 
                           n21536, ZN => n7725);
   U20378 : OAI22_X1 port map( A1 => n27414, A2 => n27218, B1 => n27212, B2 => 
                           n21535, ZN => n7726);
   U20379 : OAI22_X1 port map( A1 => n27417, A2 => n27218, B1 => n27212, B2 => 
                           n21534, ZN => n7727);
   U20380 : OAI22_X1 port map( A1 => n27420, A2 => n27218, B1 => n27212, B2 => 
                           n21533, ZN => n7728);
   U20381 : OAI22_X1 port map( A1 => n27423, A2 => n27219, B1 => n27212, B2 => 
                           n21532, ZN => n7729);
   U20382 : OAI22_X1 port map( A1 => n27426, A2 => n27219, B1 => n27213, B2 => 
                           n21531, ZN => n7730);
   U20383 : OAI22_X1 port map( A1 => n27429, A2 => n27219, B1 => n27213, B2 => 
                           n21530, ZN => n7731);
   U20384 : OAI22_X1 port map( A1 => n27432, A2 => n27219, B1 => n27213, B2 => 
                           n21529, ZN => n7732);
   U20385 : OAI22_X1 port map( A1 => n27435, A2 => n27219, B1 => n27213, B2 => 
                           n21528, ZN => n7733);
   U20386 : OAI22_X1 port map( A1 => n27438, A2 => n27219, B1 => n27213, B2 => 
                           n21527, ZN => n7734);
   U20387 : OAI22_X1 port map( A1 => n27441, A2 => n27219, B1 => n27213, B2 => 
                           n21526, ZN => n7735);
   U20388 : OAI22_X1 port map( A1 => n27444, A2 => n27219, B1 => n27213, B2 => 
                           n21525, ZN => n7736);
   U20389 : OAI22_X1 port map( A1 => n27447, A2 => n27219, B1 => n27213, B2 => 
                           n21524, ZN => n7737);
   U20390 : OAI22_X1 port map( A1 => n27450, A2 => n27219, B1 => n27213, B2 => 
                           n21523, ZN => n7738);
   U20391 : OAI22_X1 port map( A1 => n27453, A2 => n27219, B1 => n27213, B2 => 
                           n21522, ZN => n7739);
   U20392 : OAI22_X1 port map( A1 => n27456, A2 => n27219, B1 => n27213, B2 => 
                           n21521, ZN => n7740);
   U20393 : OAI22_X1 port map( A1 => n27459, A2 => n27220, B1 => n27213, B2 => 
                           n21520, ZN => n7741);
   U20394 : OAI22_X1 port map( A1 => n27318, A2 => n27240, B1 => n27234, B2 => 
                           n21407, ZN => n7822);
   U20395 : OAI22_X1 port map( A1 => n27321, A2 => n27240, B1 => n27234, B2 => 
                           n21406, ZN => n7823);
   U20396 : OAI22_X1 port map( A1 => n27324, A2 => n27240, B1 => n27234, B2 => 
                           n21405, ZN => n7824);
   U20397 : OAI22_X1 port map( A1 => n27327, A2 => n27240, B1 => n27234, B2 => 
                           n21404, ZN => n7825);
   U20398 : OAI22_X1 port map( A1 => n27330, A2 => n27240, B1 => n27234, B2 => 
                           n21403, ZN => n7826);
   U20399 : OAI22_X1 port map( A1 => n27333, A2 => n27240, B1 => n27234, B2 => 
                           n21402, ZN => n7827);
   U20400 : OAI22_X1 port map( A1 => n27336, A2 => n27240, B1 => n27234, B2 => 
                           n21401, ZN => n7828);
   U20401 : OAI22_X1 port map( A1 => n27339, A2 => n27240, B1 => n27234, B2 => 
                           n21400, ZN => n7829);
   U20402 : OAI22_X1 port map( A1 => n27342, A2 => n27240, B1 => n27234, B2 => 
                           n21399, ZN => n7830);
   U20403 : OAI22_X1 port map( A1 => n27345, A2 => n27240, B1 => n27234, B2 => 
                           n21398, ZN => n7831);
   U20404 : OAI22_X1 port map( A1 => n27348, A2 => n27240, B1 => n27234, B2 => 
                           n21397, ZN => n7832);
   U20405 : OAI22_X1 port map( A1 => n27351, A2 => n27241, B1 => n27234, B2 => 
                           n21396, ZN => n7833);
   U20406 : OAI22_X1 port map( A1 => n27354, A2 => n27241, B1 => n27235, B2 => 
                           n21395, ZN => n7834);
   U20407 : OAI22_X1 port map( A1 => n27357, A2 => n27241, B1 => n27235, B2 => 
                           n21394, ZN => n7835);
   U20408 : OAI22_X1 port map( A1 => n27360, A2 => n27241, B1 => n27235, B2 => 
                           n21393, ZN => n7836);
   U20409 : OAI22_X1 port map( A1 => n27363, A2 => n27241, B1 => n27235, B2 => 
                           n21392, ZN => n7837);
   U20410 : OAI22_X1 port map( A1 => n27366, A2 => n27241, B1 => n27235, B2 => 
                           n21391, ZN => n7838);
   U20411 : OAI22_X1 port map( A1 => n27369, A2 => n27241, B1 => n27235, B2 => 
                           n21390, ZN => n7839);
   U20412 : OAI22_X1 port map( A1 => n27372, A2 => n27241, B1 => n27235, B2 => 
                           n21389, ZN => n7840);
   U20413 : OAI22_X1 port map( A1 => n27375, A2 => n27241, B1 => n27235, B2 => 
                           n21388, ZN => n7841);
   U20414 : OAI22_X1 port map( A1 => n27378, A2 => n27241, B1 => n27235, B2 => 
                           n21387, ZN => n7842);
   U20415 : OAI22_X1 port map( A1 => n27381, A2 => n27241, B1 => n27235, B2 => 
                           n21386, ZN => n7843);
   U20416 : OAI22_X1 port map( A1 => n27384, A2 => n27241, B1 => n27235, B2 => 
                           n21385, ZN => n7844);
   U20417 : OAI22_X1 port map( A1 => n27387, A2 => n27242, B1 => n27235, B2 => 
                           n21384, ZN => n7845);
   U20418 : OAI22_X1 port map( A1 => n27390, A2 => n27242, B1 => n27236, B2 => 
                           n21383, ZN => n7846);
   U20419 : OAI22_X1 port map( A1 => n27393, A2 => n27242, B1 => n27236, B2 => 
                           n21382, ZN => n7847);
   U20420 : OAI22_X1 port map( A1 => n27396, A2 => n27242, B1 => n27236, B2 => 
                           n21381, ZN => n7848);
   U20421 : OAI22_X1 port map( A1 => n27399, A2 => n27242, B1 => n27236, B2 => 
                           n21380, ZN => n7849);
   U20422 : OAI22_X1 port map( A1 => n27402, A2 => n27242, B1 => n27236, B2 => 
                           n21379, ZN => n7850);
   U20423 : OAI22_X1 port map( A1 => n27405, A2 => n27242, B1 => n27236, B2 => 
                           n21378, ZN => n7851);
   U20424 : OAI22_X1 port map( A1 => n27408, A2 => n27242, B1 => n27236, B2 => 
                           n21377, ZN => n7852);
   U20425 : OAI22_X1 port map( A1 => n27411, A2 => n27242, B1 => n27236, B2 => 
                           n21376, ZN => n7853);
   U20426 : OAI22_X1 port map( A1 => n27414, A2 => n27242, B1 => n27236, B2 => 
                           n21375, ZN => n7854);
   U20427 : OAI22_X1 port map( A1 => n27417, A2 => n27242, B1 => n27236, B2 => 
                           n21374, ZN => n7855);
   U20428 : OAI22_X1 port map( A1 => n27420, A2 => n27242, B1 => n27236, B2 => 
                           n21373, ZN => n7856);
   U20429 : OAI22_X1 port map( A1 => n27423, A2 => n27243, B1 => n27236, B2 => 
                           n21372, ZN => n7857);
   U20430 : OAI22_X1 port map( A1 => n27426, A2 => n27243, B1 => n27237, B2 => 
                           n21371, ZN => n7858);
   U20431 : OAI22_X1 port map( A1 => n27429, A2 => n27243, B1 => n27237, B2 => 
                           n21370, ZN => n7859);
   U20432 : OAI22_X1 port map( A1 => n27432, A2 => n27243, B1 => n27237, B2 => 
                           n21369, ZN => n7860);
   U20433 : OAI22_X1 port map( A1 => n27435, A2 => n27243, B1 => n27237, B2 => 
                           n21368, ZN => n7861);
   U20434 : OAI22_X1 port map( A1 => n27438, A2 => n27243, B1 => n27237, B2 => 
                           n21367, ZN => n7862);
   U20435 : OAI22_X1 port map( A1 => n27441, A2 => n27243, B1 => n27237, B2 => 
                           n21366, ZN => n7863);
   U20436 : OAI22_X1 port map( A1 => n27444, A2 => n27243, B1 => n27237, B2 => 
                           n21365, ZN => n7864);
   U20437 : OAI22_X1 port map( A1 => n27447, A2 => n27243, B1 => n27237, B2 => 
                           n21364, ZN => n7865);
   U20438 : OAI22_X1 port map( A1 => n27450, A2 => n27243, B1 => n27237, B2 => 
                           n21363, ZN => n7866);
   U20439 : OAI22_X1 port map( A1 => n27453, A2 => n27243, B1 => n27237, B2 => 
                           n21362, ZN => n7867);
   U20440 : OAI22_X1 port map( A1 => n27456, A2 => n27243, B1 => n27237, B2 => 
                           n21361, ZN => n7868);
   U20441 : OAI22_X1 port map( A1 => n27459, A2 => n27244, B1 => n27237, B2 => 
                           n21360, ZN => n7869);
   U20442 : OAI22_X1 port map( A1 => n27319, A2 => n27000, B1 => n26994, B2 => 
                           n21347, ZN => n6542);
   U20443 : OAI22_X1 port map( A1 => n27322, A2 => n27000, B1 => n26994, B2 => 
                           n21346, ZN => n6543);
   U20444 : OAI22_X1 port map( A1 => n27325, A2 => n27000, B1 => n26994, B2 => 
                           n21345, ZN => n6544);
   U20445 : OAI22_X1 port map( A1 => n27328, A2 => n27000, B1 => n26994, B2 => 
                           n21344, ZN => n6545);
   U20446 : OAI22_X1 port map( A1 => n27331, A2 => n27000, B1 => n26994, B2 => 
                           n21343, ZN => n6546);
   U20447 : OAI22_X1 port map( A1 => n27334, A2 => n27000, B1 => n26994, B2 => 
                           n21342, ZN => n6547);
   U20448 : OAI22_X1 port map( A1 => n27337, A2 => n27000, B1 => n26994, B2 => 
                           n21341, ZN => n6548);
   U20449 : OAI22_X1 port map( A1 => n27340, A2 => n27000, B1 => n26994, B2 => 
                           n21340, ZN => n6549);
   U20450 : OAI22_X1 port map( A1 => n27343, A2 => n27000, B1 => n26994, B2 => 
                           n21339, ZN => n6550);
   U20451 : OAI22_X1 port map( A1 => n27346, A2 => n27000, B1 => n26994, B2 => 
                           n21338, ZN => n6551);
   U20452 : OAI22_X1 port map( A1 => n27349, A2 => n27000, B1 => n26994, B2 => 
                           n21337, ZN => n6552);
   U20453 : OAI22_X1 port map( A1 => n27352, A2 => n27001, B1 => n26994, B2 => 
                           n21336, ZN => n6553);
   U20454 : OAI22_X1 port map( A1 => n27355, A2 => n27001, B1 => n26995, B2 => 
                           n21335, ZN => n6554);
   U20455 : OAI22_X1 port map( A1 => n27358, A2 => n27001, B1 => n26995, B2 => 
                           n21334, ZN => n6555);
   U20456 : OAI22_X1 port map( A1 => n27361, A2 => n27001, B1 => n26995, B2 => 
                           n21333, ZN => n6556);
   U20457 : OAI22_X1 port map( A1 => n27364, A2 => n27001, B1 => n26995, B2 => 
                           n21332, ZN => n6557);
   U20458 : OAI22_X1 port map( A1 => n27367, A2 => n27001, B1 => n26995, B2 => 
                           n21331, ZN => n6558);
   U20459 : OAI22_X1 port map( A1 => n27370, A2 => n27001, B1 => n26995, B2 => 
                           n21330, ZN => n6559);
   U20460 : OAI22_X1 port map( A1 => n27373, A2 => n27001, B1 => n26995, B2 => 
                           n21329, ZN => n6560);
   U20461 : OAI22_X1 port map( A1 => n27376, A2 => n27001, B1 => n26995, B2 => 
                           n21328, ZN => n6561);
   U20462 : OAI22_X1 port map( A1 => n27379, A2 => n27001, B1 => n26995, B2 => 
                           n21327, ZN => n6562);
   U20463 : OAI22_X1 port map( A1 => n27382, A2 => n27001, B1 => n26995, B2 => 
                           n21326, ZN => n6563);
   U20464 : OAI22_X1 port map( A1 => n27385, A2 => n27001, B1 => n26995, B2 => 
                           n21325, ZN => n6564);
   U20465 : OAI22_X1 port map( A1 => n27388, A2 => n27002, B1 => n26995, B2 => 
                           n21324, ZN => n6565);
   U20466 : OAI22_X1 port map( A1 => n27391, A2 => n27002, B1 => n26996, B2 => 
                           n21323, ZN => n6566);
   U20467 : OAI22_X1 port map( A1 => n27394, A2 => n27002, B1 => n26996, B2 => 
                           n21322, ZN => n6567);
   U20468 : OAI22_X1 port map( A1 => n27397, A2 => n27002, B1 => n26996, B2 => 
                           n21321, ZN => n6568);
   U20469 : OAI22_X1 port map( A1 => n27400, A2 => n27002, B1 => n26996, B2 => 
                           n21320, ZN => n6569);
   U20470 : OAI22_X1 port map( A1 => n27403, A2 => n27002, B1 => n26996, B2 => 
                           n21319, ZN => n6570);
   U20471 : OAI22_X1 port map( A1 => n27406, A2 => n27002, B1 => n26996, B2 => 
                           n21318, ZN => n6571);
   U20472 : OAI22_X1 port map( A1 => n27409, A2 => n27002, B1 => n26996, B2 => 
                           n21317, ZN => n6572);
   U20473 : OAI22_X1 port map( A1 => n27412, A2 => n27002, B1 => n26996, B2 => 
                           n21316, ZN => n6573);
   U20474 : OAI22_X1 port map( A1 => n27415, A2 => n27002, B1 => n26996, B2 => 
                           n21315, ZN => n6574);
   U20475 : OAI22_X1 port map( A1 => n27418, A2 => n27002, B1 => n26996, B2 => 
                           n21314, ZN => n6575);
   U20476 : OAI22_X1 port map( A1 => n27421, A2 => n27002, B1 => n26996, B2 => 
                           n21313, ZN => n6576);
   U20477 : OAI22_X1 port map( A1 => n27424, A2 => n27003, B1 => n26996, B2 => 
                           n21312, ZN => n6577);
   U20478 : OAI22_X1 port map( A1 => n27427, A2 => n27003, B1 => n26997, B2 => 
                           n21311, ZN => n6578);
   U20479 : OAI22_X1 port map( A1 => n27430, A2 => n27003, B1 => n26997, B2 => 
                           n21310, ZN => n6579);
   U20480 : OAI22_X1 port map( A1 => n27433, A2 => n27003, B1 => n26997, B2 => 
                           n21309, ZN => n6580);
   U20481 : OAI22_X1 port map( A1 => n27436, A2 => n27003, B1 => n26997, B2 => 
                           n21308, ZN => n6581);
   U20482 : OAI22_X1 port map( A1 => n27439, A2 => n27003, B1 => n26997, B2 => 
                           n21307, ZN => n6582);
   U20483 : OAI22_X1 port map( A1 => n27442, A2 => n27003, B1 => n26997, B2 => 
                           n21306, ZN => n6583);
   U20484 : OAI22_X1 port map( A1 => n27445, A2 => n27003, B1 => n26997, B2 => 
                           n21305, ZN => n6584);
   U20485 : OAI22_X1 port map( A1 => n27448, A2 => n27003, B1 => n26997, B2 => 
                           n21304, ZN => n6585);
   U20486 : OAI22_X1 port map( A1 => n27451, A2 => n27003, B1 => n26997, B2 => 
                           n21303, ZN => n6586);
   U20487 : OAI22_X1 port map( A1 => n27454, A2 => n27003, B1 => n26997, B2 => 
                           n21302, ZN => n6587);
   U20488 : OAI22_X1 port map( A1 => n27457, A2 => n27003, B1 => n26997, B2 => 
                           n21301, ZN => n6588);
   U20489 : OAI22_X1 port map( A1 => n27460, A2 => n27004, B1 => n26997, B2 => 
                           n21300, ZN => n6589);
   U20490 : OAI22_X1 port map( A1 => n27319, A2 => n26976, B1 => n26970, B2 => 
                           n21227, ZN => n6414);
   U20491 : OAI22_X1 port map( A1 => n27322, A2 => n26976, B1 => n26970, B2 => 
                           n21226, ZN => n6415);
   U20492 : OAI22_X1 port map( A1 => n27325, A2 => n26976, B1 => n26970, B2 => 
                           n21225, ZN => n6416);
   U20493 : OAI22_X1 port map( A1 => n27328, A2 => n26976, B1 => n26970, B2 => 
                           n21224, ZN => n6417);
   U20494 : OAI22_X1 port map( A1 => n27331, A2 => n26976, B1 => n26970, B2 => 
                           n21223, ZN => n6418);
   U20495 : OAI22_X1 port map( A1 => n27334, A2 => n26976, B1 => n26970, B2 => 
                           n21222, ZN => n6419);
   U20496 : OAI22_X1 port map( A1 => n27337, A2 => n26976, B1 => n26970, B2 => 
                           n21221, ZN => n6420);
   U20497 : OAI22_X1 port map( A1 => n27340, A2 => n26976, B1 => n26970, B2 => 
                           n21220, ZN => n6421);
   U20498 : OAI22_X1 port map( A1 => n27343, A2 => n26976, B1 => n26970, B2 => 
                           n21219, ZN => n6422);
   U20499 : OAI22_X1 port map( A1 => n27346, A2 => n26976, B1 => n26970, B2 => 
                           n21218, ZN => n6423);
   U20500 : OAI22_X1 port map( A1 => n27349, A2 => n26976, B1 => n26970, B2 => 
                           n21217, ZN => n6424);
   U20501 : OAI22_X1 port map( A1 => n27352, A2 => n26977, B1 => n26970, B2 => 
                           n21216, ZN => n6425);
   U20502 : OAI22_X1 port map( A1 => n27355, A2 => n26977, B1 => n26971, B2 => 
                           n21215, ZN => n6426);
   U20503 : OAI22_X1 port map( A1 => n27358, A2 => n26977, B1 => n26971, B2 => 
                           n21214, ZN => n6427);
   U20504 : OAI22_X1 port map( A1 => n27361, A2 => n26977, B1 => n26971, B2 => 
                           n21213, ZN => n6428);
   U20505 : OAI22_X1 port map( A1 => n27364, A2 => n26977, B1 => n26971, B2 => 
                           n21212, ZN => n6429);
   U20506 : OAI22_X1 port map( A1 => n27367, A2 => n26977, B1 => n26971, B2 => 
                           n21211, ZN => n6430);
   U20507 : OAI22_X1 port map( A1 => n27370, A2 => n26977, B1 => n26971, B2 => 
                           n21210, ZN => n6431);
   U20508 : OAI22_X1 port map( A1 => n27373, A2 => n26977, B1 => n26971, B2 => 
                           n21209, ZN => n6432);
   U20509 : OAI22_X1 port map( A1 => n27376, A2 => n26977, B1 => n26971, B2 => 
                           n21208, ZN => n6433);
   U20510 : OAI22_X1 port map( A1 => n27379, A2 => n26977, B1 => n26971, B2 => 
                           n21207, ZN => n6434);
   U20511 : OAI22_X1 port map( A1 => n27382, A2 => n26977, B1 => n26971, B2 => 
                           n21206, ZN => n6435);
   U20512 : OAI22_X1 port map( A1 => n27385, A2 => n26977, B1 => n26971, B2 => 
                           n21205, ZN => n6436);
   U20513 : OAI22_X1 port map( A1 => n27388, A2 => n26978, B1 => n26971, B2 => 
                           n21204, ZN => n6437);
   U20514 : OAI22_X1 port map( A1 => n27391, A2 => n26978, B1 => n26972, B2 => 
                           n21203, ZN => n6438);
   U20515 : OAI22_X1 port map( A1 => n27394, A2 => n26978, B1 => n26972, B2 => 
                           n21202, ZN => n6439);
   U20516 : OAI22_X1 port map( A1 => n27397, A2 => n26978, B1 => n26972, B2 => 
                           n21201, ZN => n6440);
   U20517 : OAI22_X1 port map( A1 => n27400, A2 => n26978, B1 => n26972, B2 => 
                           n21200, ZN => n6441);
   U20518 : OAI22_X1 port map( A1 => n27403, A2 => n26978, B1 => n26972, B2 => 
                           n21199, ZN => n6442);
   U20519 : OAI22_X1 port map( A1 => n27406, A2 => n26978, B1 => n26972, B2 => 
                           n21198, ZN => n6443);
   U20520 : OAI22_X1 port map( A1 => n27409, A2 => n26978, B1 => n26972, B2 => 
                           n21197, ZN => n6444);
   U20521 : OAI22_X1 port map( A1 => n27412, A2 => n26978, B1 => n26972, B2 => 
                           n21196, ZN => n6445);
   U20522 : OAI22_X1 port map( A1 => n27415, A2 => n26978, B1 => n26972, B2 => 
                           n21195, ZN => n6446);
   U20523 : OAI22_X1 port map( A1 => n27418, A2 => n26978, B1 => n26972, B2 => 
                           n21194, ZN => n6447);
   U20524 : OAI22_X1 port map( A1 => n27421, A2 => n26978, B1 => n26972, B2 => 
                           n21193, ZN => n6448);
   U20525 : OAI22_X1 port map( A1 => n27424, A2 => n26979, B1 => n26972, B2 => 
                           n21192, ZN => n6449);
   U20526 : OAI22_X1 port map( A1 => n27427, A2 => n26979, B1 => n26973, B2 => 
                           n21191, ZN => n6450);
   U20527 : OAI22_X1 port map( A1 => n27430, A2 => n26979, B1 => n26973, B2 => 
                           n21190, ZN => n6451);
   U20528 : OAI22_X1 port map( A1 => n27433, A2 => n26979, B1 => n26973, B2 => 
                           n21189, ZN => n6452);
   U20529 : OAI22_X1 port map( A1 => n27436, A2 => n26979, B1 => n26973, B2 => 
                           n21188, ZN => n6453);
   U20530 : OAI22_X1 port map( A1 => n27439, A2 => n26979, B1 => n26973, B2 => 
                           n21187, ZN => n6454);
   U20531 : OAI22_X1 port map( A1 => n27442, A2 => n26979, B1 => n26973, B2 => 
                           n21186, ZN => n6455);
   U20532 : OAI22_X1 port map( A1 => n27445, A2 => n26979, B1 => n26973, B2 => 
                           n21185, ZN => n6456);
   U20533 : OAI22_X1 port map( A1 => n27448, A2 => n26979, B1 => n26973, B2 => 
                           n21184, ZN => n6457);
   U20534 : OAI22_X1 port map( A1 => n27451, A2 => n26979, B1 => n26973, B2 => 
                           n21183, ZN => n6458);
   U20535 : OAI22_X1 port map( A1 => n27454, A2 => n26979, B1 => n26973, B2 => 
                           n21182, ZN => n6459);
   U20536 : OAI22_X1 port map( A1 => n27457, A2 => n26979, B1 => n26973, B2 => 
                           n21181, ZN => n6460);
   U20537 : OAI22_X1 port map( A1 => n27460, A2 => n26980, B1 => n26973, B2 => 
                           n21180, ZN => n6461);
   U20538 : OAI22_X1 port map( A1 => n27319, A2 => n27108, B1 => n27102, B2 => 
                           n20822, ZN => n7118);
   U20539 : OAI22_X1 port map( A1 => n27322, A2 => n27108, B1 => n27102, B2 => 
                           n20821, ZN => n7119);
   U20540 : OAI22_X1 port map( A1 => n27325, A2 => n27108, B1 => n27102, B2 => 
                           n20820, ZN => n7120);
   U20541 : OAI22_X1 port map( A1 => n27328, A2 => n27108, B1 => n27102, B2 => 
                           n20819, ZN => n7121);
   U20542 : OAI22_X1 port map( A1 => n27331, A2 => n27108, B1 => n27102, B2 => 
                           n20818, ZN => n7122);
   U20543 : OAI22_X1 port map( A1 => n27334, A2 => n27108, B1 => n27102, B2 => 
                           n20817, ZN => n7123);
   U20544 : OAI22_X1 port map( A1 => n27337, A2 => n27108, B1 => n27102, B2 => 
                           n20816, ZN => n7124);
   U20545 : OAI22_X1 port map( A1 => n27340, A2 => n27108, B1 => n27102, B2 => 
                           n20815, ZN => n7125);
   U20546 : OAI22_X1 port map( A1 => n27343, A2 => n27108, B1 => n27102, B2 => 
                           n20814, ZN => n7126);
   U20547 : OAI22_X1 port map( A1 => n27346, A2 => n27108, B1 => n27102, B2 => 
                           n20813, ZN => n7127);
   U20548 : OAI22_X1 port map( A1 => n27349, A2 => n27108, B1 => n27102, B2 => 
                           n20812, ZN => n7128);
   U20549 : OAI22_X1 port map( A1 => n27352, A2 => n27109, B1 => n27102, B2 => 
                           n20811, ZN => n7129);
   U20550 : OAI22_X1 port map( A1 => n27355, A2 => n27109, B1 => n27103, B2 => 
                           n20810, ZN => n7130);
   U20551 : OAI22_X1 port map( A1 => n27358, A2 => n27109, B1 => n27103, B2 => 
                           n20809, ZN => n7131);
   U20552 : OAI22_X1 port map( A1 => n27361, A2 => n27109, B1 => n27103, B2 => 
                           n20808, ZN => n7132);
   U20553 : OAI22_X1 port map( A1 => n27364, A2 => n27109, B1 => n27103, B2 => 
                           n20807, ZN => n7133);
   U20554 : OAI22_X1 port map( A1 => n27367, A2 => n27109, B1 => n27103, B2 => 
                           n20806, ZN => n7134);
   U20555 : OAI22_X1 port map( A1 => n27370, A2 => n27109, B1 => n27103, B2 => 
                           n20805, ZN => n7135);
   U20556 : OAI22_X1 port map( A1 => n27373, A2 => n27109, B1 => n27103, B2 => 
                           n20804, ZN => n7136);
   U20557 : OAI22_X1 port map( A1 => n27376, A2 => n27109, B1 => n27103, B2 => 
                           n20803, ZN => n7137);
   U20558 : OAI22_X1 port map( A1 => n27379, A2 => n27109, B1 => n27103, B2 => 
                           n20802, ZN => n7138);
   U20559 : OAI22_X1 port map( A1 => n27382, A2 => n27109, B1 => n27103, B2 => 
                           n20801, ZN => n7139);
   U20560 : OAI22_X1 port map( A1 => n27385, A2 => n27109, B1 => n27103, B2 => 
                           n20800, ZN => n7140);
   U20561 : OAI22_X1 port map( A1 => n27388, A2 => n27110, B1 => n27103, B2 => 
                           n20799, ZN => n7141);
   U20562 : OAI22_X1 port map( A1 => n27391, A2 => n27110, B1 => n27104, B2 => 
                           n20798, ZN => n7142);
   U20563 : OAI22_X1 port map( A1 => n27394, A2 => n27110, B1 => n27104, B2 => 
                           n20797, ZN => n7143);
   U20564 : OAI22_X1 port map( A1 => n27397, A2 => n27110, B1 => n27104, B2 => 
                           n20796, ZN => n7144);
   U20565 : OAI22_X1 port map( A1 => n27400, A2 => n27110, B1 => n27104, B2 => 
                           n20795, ZN => n7145);
   U20566 : OAI22_X1 port map( A1 => n27403, A2 => n27110, B1 => n27104, B2 => 
                           n20794, ZN => n7146);
   U20567 : OAI22_X1 port map( A1 => n27406, A2 => n27110, B1 => n27104, B2 => 
                           n20793, ZN => n7147);
   U20568 : OAI22_X1 port map( A1 => n27409, A2 => n27110, B1 => n27104, B2 => 
                           n20792, ZN => n7148);
   U20569 : OAI22_X1 port map( A1 => n27412, A2 => n27110, B1 => n27104, B2 => 
                           n20791, ZN => n7149);
   U20570 : OAI22_X1 port map( A1 => n27415, A2 => n27110, B1 => n27104, B2 => 
                           n20790, ZN => n7150);
   U20571 : OAI22_X1 port map( A1 => n27418, A2 => n27110, B1 => n27104, B2 => 
                           n20789, ZN => n7151);
   U20572 : OAI22_X1 port map( A1 => n27421, A2 => n27110, B1 => n27104, B2 => 
                           n20788, ZN => n7152);
   U20573 : OAI22_X1 port map( A1 => n27424, A2 => n27111, B1 => n27104, B2 => 
                           n20787, ZN => n7153);
   U20574 : OAI22_X1 port map( A1 => n27427, A2 => n27111, B1 => n27105, B2 => 
                           n20786, ZN => n7154);
   U20575 : OAI22_X1 port map( A1 => n27430, A2 => n27111, B1 => n27105, B2 => 
                           n20785, ZN => n7155);
   U20576 : OAI22_X1 port map( A1 => n27433, A2 => n27111, B1 => n27105, B2 => 
                           n20784, ZN => n7156);
   U20577 : OAI22_X1 port map( A1 => n27436, A2 => n27111, B1 => n27105, B2 => 
                           n20783, ZN => n7157);
   U20578 : OAI22_X1 port map( A1 => n27439, A2 => n27111, B1 => n27105, B2 => 
                           n20782, ZN => n7158);
   U20579 : OAI22_X1 port map( A1 => n27442, A2 => n27111, B1 => n27105, B2 => 
                           n20781, ZN => n7159);
   U20580 : OAI22_X1 port map( A1 => n27445, A2 => n27111, B1 => n27105, B2 => 
                           n20780, ZN => n7160);
   U20581 : OAI22_X1 port map( A1 => n27448, A2 => n27111, B1 => n27105, B2 => 
                           n20779, ZN => n7161);
   U20582 : OAI22_X1 port map( A1 => n27451, A2 => n27111, B1 => n27105, B2 => 
                           n20778, ZN => n7162);
   U20583 : OAI22_X1 port map( A1 => n27454, A2 => n27111, B1 => n27105, B2 => 
                           n20777, ZN => n7163);
   U20584 : OAI22_X1 port map( A1 => n27457, A2 => n27111, B1 => n27105, B2 => 
                           n20776, ZN => n7164);
   U20585 : OAI22_X1 port map( A1 => n27460, A2 => n27112, B1 => n27105, B2 => 
                           n20775, ZN => n7165);
   U20586 : OAI22_X1 port map( A1 => n27318, A2 => n27132, B1 => n27126, B2 => 
                           n20759, ZN => n7246);
   U20587 : OAI22_X1 port map( A1 => n27321, A2 => n27132, B1 => n27126, B2 => 
                           n20758, ZN => n7247);
   U20588 : OAI22_X1 port map( A1 => n27324, A2 => n27132, B1 => n27126, B2 => 
                           n20757, ZN => n7248);
   U20589 : OAI22_X1 port map( A1 => n27327, A2 => n27132, B1 => n27126, B2 => 
                           n20756, ZN => n7249);
   U20590 : OAI22_X1 port map( A1 => n27330, A2 => n27132, B1 => n27126, B2 => 
                           n20755, ZN => n7250);
   U20591 : OAI22_X1 port map( A1 => n27333, A2 => n27132, B1 => n27126, B2 => 
                           n20754, ZN => n7251);
   U20592 : OAI22_X1 port map( A1 => n27336, A2 => n27132, B1 => n27126, B2 => 
                           n20753, ZN => n7252);
   U20593 : OAI22_X1 port map( A1 => n27339, A2 => n27132, B1 => n27126, B2 => 
                           n20752, ZN => n7253);
   U20594 : OAI22_X1 port map( A1 => n27342, A2 => n27132, B1 => n27126, B2 => 
                           n20751, ZN => n7254);
   U20595 : OAI22_X1 port map( A1 => n27345, A2 => n27132, B1 => n27126, B2 => 
                           n20750, ZN => n7255);
   U20596 : OAI22_X1 port map( A1 => n27348, A2 => n27132, B1 => n27126, B2 => 
                           n20749, ZN => n7256);
   U20597 : OAI22_X1 port map( A1 => n27351, A2 => n27133, B1 => n27126, B2 => 
                           n20748, ZN => n7257);
   U20598 : OAI22_X1 port map( A1 => n27354, A2 => n27133, B1 => n27127, B2 => 
                           n20747, ZN => n7258);
   U20599 : OAI22_X1 port map( A1 => n27357, A2 => n27133, B1 => n27127, B2 => 
                           n20746, ZN => n7259);
   U20600 : OAI22_X1 port map( A1 => n27360, A2 => n27133, B1 => n27127, B2 => 
                           n20745, ZN => n7260);
   U20601 : OAI22_X1 port map( A1 => n27363, A2 => n27133, B1 => n27127, B2 => 
                           n20744, ZN => n7261);
   U20602 : OAI22_X1 port map( A1 => n27366, A2 => n27133, B1 => n27127, B2 => 
                           n20743, ZN => n7262);
   U20603 : OAI22_X1 port map( A1 => n27369, A2 => n27133, B1 => n27127, B2 => 
                           n20742, ZN => n7263);
   U20604 : OAI22_X1 port map( A1 => n27372, A2 => n27133, B1 => n27127, B2 => 
                           n20741, ZN => n7264);
   U20605 : OAI22_X1 port map( A1 => n27375, A2 => n27133, B1 => n27127, B2 => 
                           n20740, ZN => n7265);
   U20606 : OAI22_X1 port map( A1 => n27378, A2 => n27133, B1 => n27127, B2 => 
                           n20739, ZN => n7266);
   U20607 : OAI22_X1 port map( A1 => n27381, A2 => n27133, B1 => n27127, B2 => 
                           n20738, ZN => n7267);
   U20608 : OAI22_X1 port map( A1 => n27384, A2 => n27133, B1 => n27127, B2 => 
                           n20737, ZN => n7268);
   U20609 : OAI22_X1 port map( A1 => n27387, A2 => n27134, B1 => n27127, B2 => 
                           n20736, ZN => n7269);
   U20610 : OAI22_X1 port map( A1 => n27390, A2 => n27134, B1 => n27128, B2 => 
                           n20735, ZN => n7270);
   U20611 : OAI22_X1 port map( A1 => n27393, A2 => n27134, B1 => n27128, B2 => 
                           n20734, ZN => n7271);
   U20612 : OAI22_X1 port map( A1 => n27396, A2 => n27134, B1 => n27128, B2 => 
                           n20733, ZN => n7272);
   U20613 : OAI22_X1 port map( A1 => n27399, A2 => n27134, B1 => n27128, B2 => 
                           n20732, ZN => n7273);
   U20614 : OAI22_X1 port map( A1 => n27402, A2 => n27134, B1 => n27128, B2 => 
                           n20731, ZN => n7274);
   U20615 : OAI22_X1 port map( A1 => n27405, A2 => n27134, B1 => n27128, B2 => 
                           n20730, ZN => n7275);
   U20616 : OAI22_X1 port map( A1 => n27408, A2 => n27134, B1 => n27128, B2 => 
                           n20729, ZN => n7276);
   U20617 : OAI22_X1 port map( A1 => n27411, A2 => n27134, B1 => n27128, B2 => 
                           n20728, ZN => n7277);
   U20618 : OAI22_X1 port map( A1 => n27414, A2 => n27134, B1 => n27128, B2 => 
                           n20727, ZN => n7278);
   U20619 : OAI22_X1 port map( A1 => n27417, A2 => n27134, B1 => n27128, B2 => 
                           n20726, ZN => n7279);
   U20620 : OAI22_X1 port map( A1 => n27420, A2 => n27134, B1 => n27128, B2 => 
                           n20725, ZN => n7280);
   U20621 : OAI22_X1 port map( A1 => n27423, A2 => n27135, B1 => n27128, B2 => 
                           n20724, ZN => n7281);
   U20622 : OAI22_X1 port map( A1 => n27426, A2 => n27135, B1 => n27129, B2 => 
                           n20723, ZN => n7282);
   U20623 : OAI22_X1 port map( A1 => n27429, A2 => n27135, B1 => n27129, B2 => 
                           n20722, ZN => n7283);
   U20624 : OAI22_X1 port map( A1 => n27432, A2 => n27135, B1 => n27129, B2 => 
                           n20721, ZN => n7284);
   U20625 : OAI22_X1 port map( A1 => n27435, A2 => n27135, B1 => n27129, B2 => 
                           n20720, ZN => n7285);
   U20626 : OAI22_X1 port map( A1 => n27438, A2 => n27135, B1 => n27129, B2 => 
                           n20719, ZN => n7286);
   U20627 : OAI22_X1 port map( A1 => n27441, A2 => n27135, B1 => n27129, B2 => 
                           n20718, ZN => n7287);
   U20628 : OAI22_X1 port map( A1 => n27444, A2 => n27135, B1 => n27129, B2 => 
                           n20717, ZN => n7288);
   U20629 : OAI22_X1 port map( A1 => n27447, A2 => n27135, B1 => n27129, B2 => 
                           n20716, ZN => n7289);
   U20630 : OAI22_X1 port map( A1 => n27450, A2 => n27135, B1 => n27129, B2 => 
                           n20715, ZN => n7290);
   U20631 : OAI22_X1 port map( A1 => n27453, A2 => n27135, B1 => n27129, B2 => 
                           n20714, ZN => n7291);
   U20632 : OAI22_X1 port map( A1 => n27456, A2 => n27135, B1 => n27129, B2 => 
                           n20713, ZN => n7292);
   U20633 : OAI22_X1 port map( A1 => n27459, A2 => n27136, B1 => n27129, B2 => 
                           n20712, ZN => n7293);
   U20634 : OAI22_X1 port map( A1 => n27462, A2 => n27172, B1 => n27166, B2 => 
                           n22511, ZN => n7486);
   U20635 : OAI22_X1 port map( A1 => n27465, A2 => n27172, B1 => n27166, B2 => 
                           n22510, ZN => n7487);
   U20636 : OAI22_X1 port map( A1 => n27468, A2 => n27172, B1 => n27166, B2 => 
                           n22509, ZN => n7488);
   U20637 : OAI22_X1 port map( A1 => n27471, A2 => n27172, B1 => n27166, B2 => 
                           n22508, ZN => n7489);
   U20638 : OAI22_X1 port map( A1 => n27463, A2 => n26992, B1 => n26986, B2 => 
                           n22503, ZN => n6526);
   U20639 : OAI22_X1 port map( A1 => n27466, A2 => n26992, B1 => n26986, B2 => 
                           n22502, ZN => n6527);
   U20640 : OAI22_X1 port map( A1 => n27469, A2 => n26992, B1 => n26986, B2 => 
                           n22501, ZN => n6528);
   U20641 : OAI22_X1 port map( A1 => n27472, A2 => n26992, B1 => n26986, B2 => 
                           n22500, ZN => n6529);
   U20642 : OAI22_X1 port map( A1 => n27462, A2 => n27184, B1 => n27178, B2 => 
                           n22259, ZN => n7550);
   U20643 : OAI22_X1 port map( A1 => n27465, A2 => n27184, B1 => n27178, B2 => 
                           n22258, ZN => n7551);
   U20644 : OAI22_X1 port map( A1 => n27468, A2 => n27184, B1 => n27178, B2 => 
                           n22257, ZN => n7552);
   U20645 : OAI22_X1 port map( A1 => n27471, A2 => n27184, B1 => n27178, B2 => 
                           n22256, ZN => n7553);
   U20646 : OAI22_X1 port map( A1 => n27463, A2 => n27052, B1 => n27046, B2 => 
                           n22251, ZN => n6846);
   U20647 : OAI22_X1 port map( A1 => n27466, A2 => n27052, B1 => n27046, B2 => 
                           n22250, ZN => n6847);
   U20648 : OAI22_X1 port map( A1 => n27469, A2 => n27052, B1 => n27046, B2 => 
                           n22249, ZN => n6848);
   U20649 : OAI22_X1 port map( A1 => n27472, A2 => n27052, B1 => n27046, B2 => 
                           n22248, ZN => n6849);
   U20650 : OAI22_X1 port map( A1 => n27462, A2 => n27196, B1 => n27190, B2 => 
                           n21511, ZN => n7614);
   U20651 : OAI22_X1 port map( A1 => n27465, A2 => n27196, B1 => n27190, B2 => 
                           n21510, ZN => n7615);
   U20652 : OAI22_X1 port map( A1 => n27468, A2 => n27196, B1 => n27190, B2 => 
                           n21509, ZN => n7616);
   U20653 : OAI22_X1 port map( A1 => n27471, A2 => n27196, B1 => n27190, B2 => 
                           n21508, ZN => n7617);
   U20654 : OAI22_X1 port map( A1 => n27462, A2 => n27148, B1 => n27142, B2 => 
                           n21507, ZN => n7358);
   U20655 : OAI22_X1 port map( A1 => n27465, A2 => n27148, B1 => n27142, B2 => 
                           n21506, ZN => n7359);
   U20656 : OAI22_X1 port map( A1 => n27468, A2 => n27148, B1 => n27142, B2 => 
                           n21505, ZN => n7360);
   U20657 : OAI22_X1 port map( A1 => n27471, A2 => n27148, B1 => n27142, B2 => 
                           n21504, ZN => n7361);
   U20658 : OAI22_X1 port map( A1 => n27463, A2 => n27076, B1 => n27070, B2 => 
                           n21491, ZN => n6974);
   U20659 : OAI22_X1 port map( A1 => n27466, A2 => n27076, B1 => n27070, B2 => 
                           n21490, ZN => n6975);
   U20660 : OAI22_X1 port map( A1 => n27469, A2 => n27076, B1 => n27070, B2 => 
                           n21489, ZN => n6976);
   U20661 : OAI22_X1 port map( A1 => n27472, A2 => n27076, B1 => n27070, B2 => 
                           n21488, ZN => n6977);
   U20662 : OAI22_X1 port map( A1 => n27464, A2 => n26968, B1 => n26962, B2 => 
                           n21483, ZN => n6398);
   U20663 : OAI22_X1 port map( A1 => n27467, A2 => n26968, B1 => n26962, B2 => 
                           n21482, ZN => n6399);
   U20664 : OAI22_X1 port map( A1 => n27470, A2 => n26968, B1 => n26962, B2 => 
                           n21481, ZN => n6400);
   U20665 : OAI22_X1 port map( A1 => n27473, A2 => n26968, B1 => n26962, B2 => 
                           n21480, ZN => n6401);
   U20666 : OAI22_X1 port map( A1 => n27462, A2 => n27220, B1 => n27214, B2 => 
                           n21179, ZN => n7742);
   U20667 : OAI22_X1 port map( A1 => n27465, A2 => n27220, B1 => n27214, B2 => 
                           n21178, ZN => n7743);
   U20668 : OAI22_X1 port map( A1 => n27468, A2 => n27220, B1 => n27214, B2 => 
                           n21177, ZN => n7744);
   U20669 : OAI22_X1 port map( A1 => n27471, A2 => n27220, B1 => n27214, B2 => 
                           n21176, ZN => n7745);
   U20670 : OAI22_X1 port map( A1 => n27462, A2 => n27244, B1 => n27238, B2 => 
                           n21171, ZN => n7870);
   U20671 : OAI22_X1 port map( A1 => n27465, A2 => n27244, B1 => n27238, B2 => 
                           n21170, ZN => n7871);
   U20672 : OAI22_X1 port map( A1 => n27468, A2 => n27244, B1 => n27238, B2 => 
                           n21169, ZN => n7872);
   U20673 : OAI22_X1 port map( A1 => n27471, A2 => n27244, B1 => n27238, B2 => 
                           n21168, ZN => n7873);
   U20674 : OAI22_X1 port map( A1 => n27463, A2 => n27004, B1 => n26998, B2 => 
                           n21167, ZN => n6590);
   U20675 : OAI22_X1 port map( A1 => n27466, A2 => n27004, B1 => n26998, B2 => 
                           n21166, ZN => n6591);
   U20676 : OAI22_X1 port map( A1 => n27469, A2 => n27004, B1 => n26998, B2 => 
                           n21165, ZN => n6592);
   U20677 : OAI22_X1 port map( A1 => n27472, A2 => n27004, B1 => n26998, B2 => 
                           n21164, ZN => n6593);
   U20678 : OAI22_X1 port map( A1 => n27463, A2 => n26980, B1 => n26974, B2 => 
                           n21159, ZN => n6462);
   U20679 : OAI22_X1 port map( A1 => n27466, A2 => n26980, B1 => n26974, B2 => 
                           n21158, ZN => n6463);
   U20680 : OAI22_X1 port map( A1 => n27469, A2 => n26980, B1 => n26974, B2 => 
                           n21157, ZN => n6464);
   U20681 : OAI22_X1 port map( A1 => n27472, A2 => n26980, B1 => n26974, B2 => 
                           n21156, ZN => n6465);
   U20682 : OAI22_X1 port map( A1 => n27472, A2 => n27112, B1 => n27106, B2 => 
                           n21155, ZN => n7169);
   U20683 : OAI22_X1 port map( A1 => n27463, A2 => n27112, B1 => n27106, B2 => 
                           n20774, ZN => n7166);
   U20684 : OAI22_X1 port map( A1 => n27466, A2 => n27112, B1 => n27106, B2 => 
                           n20773, ZN => n7167);
   U20685 : OAI22_X1 port map( A1 => n27469, A2 => n27112, B1 => n27106, B2 => 
                           n20772, ZN => n7168);
   U20686 : OAI22_X1 port map( A1 => n27462, A2 => n27136, B1 => n27130, B2 => 
                           n20711, ZN => n7294);
   U20687 : OAI22_X1 port map( A1 => n27465, A2 => n27136, B1 => n27130, B2 => 
                           n20710, ZN => n7295);
   U20688 : OAI22_X1 port map( A1 => n27468, A2 => n27136, B1 => n27130, B2 => 
                           n20709, ZN => n7296);
   U20689 : OAI22_X1 port map( A1 => n27471, A2 => n27136, B1 => n27130, B2 => 
                           n20708, ZN => n7297);
   U20690 : OAI22_X1 port map( A1 => n27282, A2 => n27167, B1 => n27161, B2 => 
                           n22691, ZN => n7426);
   U20691 : OAI22_X1 port map( A1 => n27285, A2 => n27167, B1 => n27161, B2 => 
                           n22690, ZN => n7427);
   U20692 : OAI22_X1 port map( A1 => n27288, A2 => n27167, B1 => n27161, B2 => 
                           n22689, ZN => n7428);
   U20693 : OAI22_X1 port map( A1 => n27291, A2 => n27167, B1 => n27161, B2 => 
                           n22688, ZN => n7429);
   U20694 : OAI22_X1 port map( A1 => n27294, A2 => n27167, B1 => n27161, B2 => 
                           n22687, ZN => n7430);
   U20695 : OAI22_X1 port map( A1 => n27297, A2 => n27167, B1 => n27161, B2 => 
                           n22686, ZN => n7431);
   U20696 : OAI22_X1 port map( A1 => n27300, A2 => n27167, B1 => n27161, B2 => 
                           n22685, ZN => n7432);
   U20697 : OAI22_X1 port map( A1 => n27303, A2 => n27167, B1 => n27161, B2 => 
                           n22684, ZN => n7433);
   U20698 : OAI22_X1 port map( A1 => n27306, A2 => n27167, B1 => n27161, B2 => 
                           n22683, ZN => n7434);
   U20699 : OAI22_X1 port map( A1 => n27309, A2 => n27167, B1 => n27161, B2 => 
                           n22682, ZN => n7435);
   U20700 : OAI22_X1 port map( A1 => n27312, A2 => n27167, B1 => n27161, B2 => 
                           n22681, ZN => n7436);
   U20701 : OAI22_X1 port map( A1 => n27315, A2 => n27168, B1 => n27161, B2 => 
                           n22680, ZN => n7437);
   U20702 : OAI22_X1 port map( A1 => n27283, A2 => n26987, B1 => n26981, B2 => 
                           n22571, ZN => n6466);
   U20703 : OAI22_X1 port map( A1 => n27286, A2 => n26987, B1 => n26981, B2 => 
                           n22570, ZN => n6467);
   U20704 : OAI22_X1 port map( A1 => n27289, A2 => n26987, B1 => n26981, B2 => 
                           n22569, ZN => n6468);
   U20705 : OAI22_X1 port map( A1 => n27292, A2 => n26987, B1 => n26981, B2 => 
                           n22568, ZN => n6469);
   U20706 : OAI22_X1 port map( A1 => n27295, A2 => n26987, B1 => n26981, B2 => 
                           n22567, ZN => n6470);
   U20707 : OAI22_X1 port map( A1 => n27298, A2 => n26987, B1 => n26981, B2 => 
                           n22566, ZN => n6471);
   U20708 : OAI22_X1 port map( A1 => n27301, A2 => n26987, B1 => n26981, B2 => 
                           n22565, ZN => n6472);
   U20709 : OAI22_X1 port map( A1 => n27304, A2 => n26987, B1 => n26981, B2 => 
                           n22564, ZN => n6473);
   U20710 : OAI22_X1 port map( A1 => n27307, A2 => n26987, B1 => n26981, B2 => 
                           n22563, ZN => n6474);
   U20711 : OAI22_X1 port map( A1 => n27310, A2 => n26987, B1 => n26981, B2 => 
                           n22562, ZN => n6475);
   U20712 : OAI22_X1 port map( A1 => n27313, A2 => n26987, B1 => n26981, B2 => 
                           n22561, ZN => n6476);
   U20713 : OAI22_X1 port map( A1 => n27316, A2 => n26988, B1 => n26981, B2 => 
                           n22560, ZN => n6477);
   U20714 : OAI22_X1 port map( A1 => n27282, A2 => n27179, B1 => n27173, B2 => 
                           n22499, ZN => n7490);
   U20715 : OAI22_X1 port map( A1 => n27285, A2 => n27179, B1 => n27173, B2 => 
                           n22498, ZN => n7491);
   U20716 : OAI22_X1 port map( A1 => n27288, A2 => n27179, B1 => n27173, B2 => 
                           n22497, ZN => n7492);
   U20717 : OAI22_X1 port map( A1 => n27291, A2 => n27179, B1 => n27173, B2 => 
                           n22496, ZN => n7493);
   U20718 : OAI22_X1 port map( A1 => n27294, A2 => n27179, B1 => n27173, B2 => 
                           n22495, ZN => n7494);
   U20719 : OAI22_X1 port map( A1 => n27297, A2 => n27179, B1 => n27173, B2 => 
                           n22494, ZN => n7495);
   U20720 : OAI22_X1 port map( A1 => n27300, A2 => n27179, B1 => n27173, B2 => 
                           n22493, ZN => n7496);
   U20721 : OAI22_X1 port map( A1 => n27303, A2 => n27179, B1 => n27173, B2 => 
                           n22492, ZN => n7497);
   U20722 : OAI22_X1 port map( A1 => n27306, A2 => n27179, B1 => n27173, B2 => 
                           n22491, ZN => n7498);
   U20723 : OAI22_X1 port map( A1 => n27309, A2 => n27179, B1 => n27173, B2 => 
                           n22490, ZN => n7499);
   U20724 : OAI22_X1 port map( A1 => n27312, A2 => n27179, B1 => n27173, B2 => 
                           n22489, ZN => n7500);
   U20725 : OAI22_X1 port map( A1 => n27315, A2 => n27180, B1 => n27173, B2 => 
                           n22488, ZN => n7501);
   U20726 : OAI22_X1 port map( A1 => n27283, A2 => n27047, B1 => n27041, B2 => 
                           n22379, ZN => n6786);
   U20727 : OAI22_X1 port map( A1 => n27286, A2 => n27047, B1 => n27041, B2 => 
                           n22378, ZN => n6787);
   U20728 : OAI22_X1 port map( A1 => n27289, A2 => n27047, B1 => n27041, B2 => 
                           n22377, ZN => n6788);
   U20729 : OAI22_X1 port map( A1 => n27292, A2 => n27047, B1 => n27041, B2 => 
                           n22376, ZN => n6789);
   U20730 : OAI22_X1 port map( A1 => n27295, A2 => n27047, B1 => n27041, B2 => 
                           n22375, ZN => n6790);
   U20731 : OAI22_X1 port map( A1 => n27298, A2 => n27047, B1 => n27041, B2 => 
                           n22374, ZN => n6791);
   U20732 : OAI22_X1 port map( A1 => n27301, A2 => n27047, B1 => n27041, B2 => 
                           n22373, ZN => n6792);
   U20733 : OAI22_X1 port map( A1 => n27304, A2 => n27047, B1 => n27041, B2 => 
                           n22372, ZN => n6793);
   U20734 : OAI22_X1 port map( A1 => n27307, A2 => n27047, B1 => n27041, B2 => 
                           n22371, ZN => n6794);
   U20735 : OAI22_X1 port map( A1 => n27310, A2 => n27047, B1 => n27041, B2 => 
                           n22370, ZN => n6795);
   U20736 : OAI22_X1 port map( A1 => n27313, A2 => n27047, B1 => n27041, B2 => 
                           n22369, ZN => n6796);
   U20737 : OAI22_X1 port map( A1 => n27316, A2 => n27048, B1 => n27041, B2 => 
                           n22368, ZN => n6797);
   U20738 : OAI22_X1 port map( A1 => n27282, A2 => n27191, B1 => n27185, B2 => 
                           n22059, ZN => n7554);
   U20739 : OAI22_X1 port map( A1 => n27285, A2 => n27191, B1 => n27185, B2 => 
                           n22058, ZN => n7555);
   U20740 : OAI22_X1 port map( A1 => n27288, A2 => n27191, B1 => n27185, B2 => 
                           n22057, ZN => n7556);
   U20741 : OAI22_X1 port map( A1 => n27291, A2 => n27191, B1 => n27185, B2 => 
                           n22056, ZN => n7557);
   U20742 : OAI22_X1 port map( A1 => n27294, A2 => n27191, B1 => n27185, B2 => 
                           n22055, ZN => n7558);
   U20743 : OAI22_X1 port map( A1 => n27297, A2 => n27191, B1 => n27185, B2 => 
                           n22054, ZN => n7559);
   U20744 : OAI22_X1 port map( A1 => n27300, A2 => n27191, B1 => n27185, B2 => 
                           n22053, ZN => n7560);
   U20745 : OAI22_X1 port map( A1 => n27303, A2 => n27191, B1 => n27185, B2 => 
                           n22052, ZN => n7561);
   U20746 : OAI22_X1 port map( A1 => n27306, A2 => n27191, B1 => n27185, B2 => 
                           n22051, ZN => n7562);
   U20747 : OAI22_X1 port map( A1 => n27309, A2 => n27191, B1 => n27185, B2 => 
                           n22050, ZN => n7563);
   U20748 : OAI22_X1 port map( A1 => n27312, A2 => n27191, B1 => n27185, B2 => 
                           n22049, ZN => n7564);
   U20749 : OAI22_X1 port map( A1 => n27315, A2 => n27192, B1 => n27185, B2 => 
                           n22048, ZN => n7565);
   U20750 : OAI22_X1 port map( A1 => n27282, A2 => n27143, B1 => n27137, B2 => 
                           n21999, ZN => n7298);
   U20751 : OAI22_X1 port map( A1 => n27285, A2 => n27143, B1 => n27137, B2 => 
                           n21998, ZN => n7299);
   U20752 : OAI22_X1 port map( A1 => n27288, A2 => n27143, B1 => n27137, B2 => 
                           n21997, ZN => n7300);
   U20753 : OAI22_X1 port map( A1 => n27291, A2 => n27143, B1 => n27137, B2 => 
                           n21996, ZN => n7301);
   U20754 : OAI22_X1 port map( A1 => n27294, A2 => n27143, B1 => n27137, B2 => 
                           n21995, ZN => n7302);
   U20755 : OAI22_X1 port map( A1 => n27297, A2 => n27143, B1 => n27137, B2 => 
                           n21994, ZN => n7303);
   U20756 : OAI22_X1 port map( A1 => n27300, A2 => n27143, B1 => n27137, B2 => 
                           n21993, ZN => n7304);
   U20757 : OAI22_X1 port map( A1 => n27303, A2 => n27143, B1 => n27137, B2 => 
                           n21992, ZN => n7305);
   U20758 : OAI22_X1 port map( A1 => n27306, A2 => n27143, B1 => n27137, B2 => 
                           n21991, ZN => n7306);
   U20759 : OAI22_X1 port map( A1 => n27309, A2 => n27143, B1 => n27137, B2 => 
                           n21990, ZN => n7307);
   U20760 : OAI22_X1 port map( A1 => n27312, A2 => n27143, B1 => n27137, B2 => 
                           n21989, ZN => n7308);
   U20761 : OAI22_X1 port map( A1 => n27315, A2 => n27144, B1 => n27137, B2 => 
                           n21988, ZN => n7309);
   U20762 : OAI22_X1 port map( A1 => n27283, A2 => n27071, B1 => n27065, B2 => 
                           n21759, ZN => n6914);
   U20763 : OAI22_X1 port map( A1 => n27286, A2 => n27071, B1 => n27065, B2 => 
                           n21758, ZN => n6915);
   U20764 : OAI22_X1 port map( A1 => n27289, A2 => n27071, B1 => n27065, B2 => 
                           n21757, ZN => n6916);
   U20765 : OAI22_X1 port map( A1 => n27292, A2 => n27071, B1 => n27065, B2 => 
                           n21756, ZN => n6917);
   U20766 : OAI22_X1 port map( A1 => n27295, A2 => n27071, B1 => n27065, B2 => 
                           n21755, ZN => n6918);
   U20767 : OAI22_X1 port map( A1 => n27298, A2 => n27071, B1 => n27065, B2 => 
                           n21754, ZN => n6919);
   U20768 : OAI22_X1 port map( A1 => n27301, A2 => n27071, B1 => n27065, B2 => 
                           n21753, ZN => n6920);
   U20769 : OAI22_X1 port map( A1 => n27304, A2 => n27071, B1 => n27065, B2 => 
                           n21752, ZN => n6921);
   U20770 : OAI22_X1 port map( A1 => n27307, A2 => n27071, B1 => n27065, B2 => 
                           n21751, ZN => n6922);
   U20771 : OAI22_X1 port map( A1 => n27310, A2 => n27071, B1 => n27065, B2 => 
                           n21750, ZN => n6923);
   U20772 : OAI22_X1 port map( A1 => n27313, A2 => n27071, B1 => n27065, B2 => 
                           n21749, ZN => n6924);
   U20773 : OAI22_X1 port map( A1 => n27316, A2 => n27072, B1 => n27065, B2 => 
                           n21748, ZN => n6925);
   U20774 : OAI22_X1 port map( A1 => n27284, A2 => n26963, B1 => n26957, B2 => 
                           n21639, ZN => n6338);
   U20775 : OAI22_X1 port map( A1 => n27287, A2 => n26963, B1 => n26957, B2 => 
                           n21638, ZN => n6339);
   U20776 : OAI22_X1 port map( A1 => n27290, A2 => n26963, B1 => n26957, B2 => 
                           n21637, ZN => n6340);
   U20777 : OAI22_X1 port map( A1 => n27293, A2 => n26963, B1 => n26957, B2 => 
                           n21636, ZN => n6341);
   U20778 : OAI22_X1 port map( A1 => n27296, A2 => n26963, B1 => n26957, B2 => 
                           n21635, ZN => n6342);
   U20779 : OAI22_X1 port map( A1 => n27299, A2 => n26963, B1 => n26957, B2 => 
                           n21634, ZN => n6343);
   U20780 : OAI22_X1 port map( A1 => n27302, A2 => n26963, B1 => n26957, B2 => 
                           n21633, ZN => n6344);
   U20781 : OAI22_X1 port map( A1 => n27305, A2 => n26963, B1 => n26957, B2 => 
                           n21632, ZN => n6345);
   U20782 : OAI22_X1 port map( A1 => n27308, A2 => n26963, B1 => n26957, B2 => 
                           n21631, ZN => n6346);
   U20783 : OAI22_X1 port map( A1 => n27311, A2 => n26963, B1 => n26957, B2 => 
                           n21630, ZN => n6347);
   U20784 : OAI22_X1 port map( A1 => n27314, A2 => n26963, B1 => n26957, B2 => 
                           n21629, ZN => n6348);
   U20785 : OAI22_X1 port map( A1 => n27317, A2 => n26964, B1 => n26957, B2 => 
                           n21628, ZN => n6349);
   U20786 : OAI22_X1 port map( A1 => n27282, A2 => n27215, B1 => n27209, B2 => 
                           n21579, ZN => n7682);
   U20787 : OAI22_X1 port map( A1 => n27285, A2 => n27215, B1 => n27209, B2 => 
                           n21578, ZN => n7683);
   U20788 : OAI22_X1 port map( A1 => n27288, A2 => n27215, B1 => n27209, B2 => 
                           n21577, ZN => n7684);
   U20789 : OAI22_X1 port map( A1 => n27291, A2 => n27215, B1 => n27209, B2 => 
                           n21576, ZN => n7685);
   U20790 : OAI22_X1 port map( A1 => n27294, A2 => n27215, B1 => n27209, B2 => 
                           n21575, ZN => n7686);
   U20791 : OAI22_X1 port map( A1 => n27297, A2 => n27215, B1 => n27209, B2 => 
                           n21574, ZN => n7687);
   U20792 : OAI22_X1 port map( A1 => n27300, A2 => n27215, B1 => n27209, B2 => 
                           n21573, ZN => n7688);
   U20793 : OAI22_X1 port map( A1 => n27303, A2 => n27215, B1 => n27209, B2 => 
                           n21572, ZN => n7689);
   U20794 : OAI22_X1 port map( A1 => n27306, A2 => n27215, B1 => n27209, B2 => 
                           n21571, ZN => n7690);
   U20795 : OAI22_X1 port map( A1 => n27309, A2 => n27215, B1 => n27209, B2 => 
                           n21570, ZN => n7691);
   U20796 : OAI22_X1 port map( A1 => n27312, A2 => n27215, B1 => n27209, B2 => 
                           n21569, ZN => n7692);
   U20797 : OAI22_X1 port map( A1 => n27315, A2 => n27216, B1 => n27209, B2 => 
                           n21568, ZN => n7693);
   U20798 : OAI22_X1 port map( A1 => n27282, A2 => n27239, B1 => n27233, B2 => 
                           n21419, ZN => n7810);
   U20799 : OAI22_X1 port map( A1 => n27285, A2 => n27239, B1 => n27233, B2 => 
                           n21418, ZN => n7811);
   U20800 : OAI22_X1 port map( A1 => n27288, A2 => n27239, B1 => n27233, B2 => 
                           n21417, ZN => n7812);
   U20801 : OAI22_X1 port map( A1 => n27291, A2 => n27239, B1 => n27233, B2 => 
                           n21416, ZN => n7813);
   U20802 : OAI22_X1 port map( A1 => n27294, A2 => n27239, B1 => n27233, B2 => 
                           n21415, ZN => n7814);
   U20803 : OAI22_X1 port map( A1 => n27297, A2 => n27239, B1 => n27233, B2 => 
                           n21414, ZN => n7815);
   U20804 : OAI22_X1 port map( A1 => n27300, A2 => n27239, B1 => n27233, B2 => 
                           n21413, ZN => n7816);
   U20805 : OAI22_X1 port map( A1 => n27303, A2 => n27239, B1 => n27233, B2 => 
                           n21412, ZN => n7817);
   U20806 : OAI22_X1 port map( A1 => n27306, A2 => n27239, B1 => n27233, B2 => 
                           n21411, ZN => n7818);
   U20807 : OAI22_X1 port map( A1 => n27309, A2 => n27239, B1 => n27233, B2 => 
                           n21410, ZN => n7819);
   U20808 : OAI22_X1 port map( A1 => n27312, A2 => n27239, B1 => n27233, B2 => 
                           n21409, ZN => n7820);
   U20809 : OAI22_X1 port map( A1 => n27315, A2 => n27240, B1 => n27233, B2 => 
                           n21408, ZN => n7821);
   U20810 : OAI22_X1 port map( A1 => n27283, A2 => n26999, B1 => n26993, B2 => 
                           n21359, ZN => n6530);
   U20811 : OAI22_X1 port map( A1 => n27286, A2 => n26999, B1 => n26993, B2 => 
                           n21358, ZN => n6531);
   U20812 : OAI22_X1 port map( A1 => n27289, A2 => n26999, B1 => n26993, B2 => 
                           n21357, ZN => n6532);
   U20813 : OAI22_X1 port map( A1 => n27292, A2 => n26999, B1 => n26993, B2 => 
                           n21356, ZN => n6533);
   U20814 : OAI22_X1 port map( A1 => n27295, A2 => n26999, B1 => n26993, B2 => 
                           n21355, ZN => n6534);
   U20815 : OAI22_X1 port map( A1 => n27298, A2 => n26999, B1 => n26993, B2 => 
                           n21354, ZN => n6535);
   U20816 : OAI22_X1 port map( A1 => n27301, A2 => n26999, B1 => n26993, B2 => 
                           n21353, ZN => n6536);
   U20817 : OAI22_X1 port map( A1 => n27304, A2 => n26999, B1 => n26993, B2 => 
                           n21352, ZN => n6537);
   U20818 : OAI22_X1 port map( A1 => n27307, A2 => n26999, B1 => n26993, B2 => 
                           n21351, ZN => n6538);
   U20819 : OAI22_X1 port map( A1 => n27310, A2 => n26999, B1 => n26993, B2 => 
                           n21350, ZN => n6539);
   U20820 : OAI22_X1 port map( A1 => n27313, A2 => n26999, B1 => n26993, B2 => 
                           n21349, ZN => n6540);
   U20821 : OAI22_X1 port map( A1 => n27316, A2 => n27000, B1 => n26993, B2 => 
                           n21348, ZN => n6541);
   U20822 : OAI22_X1 port map( A1 => n27283, A2 => n26975, B1 => n26969, B2 => 
                           n21239, ZN => n6402);
   U20823 : OAI22_X1 port map( A1 => n27286, A2 => n26975, B1 => n26969, B2 => 
                           n21238, ZN => n6403);
   U20824 : OAI22_X1 port map( A1 => n27289, A2 => n26975, B1 => n26969, B2 => 
                           n21237, ZN => n6404);
   U20825 : OAI22_X1 port map( A1 => n27292, A2 => n26975, B1 => n26969, B2 => 
                           n21236, ZN => n6405);
   U20826 : OAI22_X1 port map( A1 => n27295, A2 => n26975, B1 => n26969, B2 => 
                           n21235, ZN => n6406);
   U20827 : OAI22_X1 port map( A1 => n27298, A2 => n26975, B1 => n26969, B2 => 
                           n21234, ZN => n6407);
   U20828 : OAI22_X1 port map( A1 => n27301, A2 => n26975, B1 => n26969, B2 => 
                           n21233, ZN => n6408);
   U20829 : OAI22_X1 port map( A1 => n27304, A2 => n26975, B1 => n26969, B2 => 
                           n21232, ZN => n6409);
   U20830 : OAI22_X1 port map( A1 => n27307, A2 => n26975, B1 => n26969, B2 => 
                           n21231, ZN => n6410);
   U20831 : OAI22_X1 port map( A1 => n27310, A2 => n26975, B1 => n26969, B2 => 
                           n21230, ZN => n6411);
   U20832 : OAI22_X1 port map( A1 => n27313, A2 => n26975, B1 => n26969, B2 => 
                           n21229, ZN => n6412);
   U20833 : OAI22_X1 port map( A1 => n27316, A2 => n26976, B1 => n26969, B2 => 
                           n21228, ZN => n6413);
   U20834 : OAI22_X1 port map( A1 => n27283, A2 => n27107, B1 => n27101, B2 => 
                           n20834, ZN => n7106);
   U20835 : OAI22_X1 port map( A1 => n27286, A2 => n27107, B1 => n27101, B2 => 
                           n20833, ZN => n7107);
   U20836 : OAI22_X1 port map( A1 => n27289, A2 => n27107, B1 => n27101, B2 => 
                           n20832, ZN => n7108);
   U20837 : OAI22_X1 port map( A1 => n27292, A2 => n27107, B1 => n27101, B2 => 
                           n20831, ZN => n7109);
   U20838 : OAI22_X1 port map( A1 => n27295, A2 => n27107, B1 => n27101, B2 => 
                           n20830, ZN => n7110);
   U20839 : OAI22_X1 port map( A1 => n27298, A2 => n27107, B1 => n27101, B2 => 
                           n20829, ZN => n7111);
   U20840 : OAI22_X1 port map( A1 => n27301, A2 => n27107, B1 => n27101, B2 => 
                           n20828, ZN => n7112);
   U20841 : OAI22_X1 port map( A1 => n27304, A2 => n27107, B1 => n27101, B2 => 
                           n20827, ZN => n7113);
   U20842 : OAI22_X1 port map( A1 => n27307, A2 => n27107, B1 => n27101, B2 => 
                           n20826, ZN => n7114);
   U20843 : OAI22_X1 port map( A1 => n27310, A2 => n27107, B1 => n27101, B2 => 
                           n20825, ZN => n7115);
   U20844 : OAI22_X1 port map( A1 => n27313, A2 => n27107, B1 => n27101, B2 => 
                           n20824, ZN => n7116);
   U20845 : OAI22_X1 port map( A1 => n27316, A2 => n27108, B1 => n27101, B2 => 
                           n20823, ZN => n7117);
   U20846 : OAI22_X1 port map( A1 => n27282, A2 => n27131, B1 => n27125, B2 => 
                           n20771, ZN => n7234);
   U20847 : OAI22_X1 port map( A1 => n27285, A2 => n27131, B1 => n27125, B2 => 
                           n20770, ZN => n7235);
   U20848 : OAI22_X1 port map( A1 => n27288, A2 => n27131, B1 => n27125, B2 => 
                           n20769, ZN => n7236);
   U20849 : OAI22_X1 port map( A1 => n27291, A2 => n27131, B1 => n27125, B2 => 
                           n20768, ZN => n7237);
   U20850 : OAI22_X1 port map( A1 => n27294, A2 => n27131, B1 => n27125, B2 => 
                           n20767, ZN => n7238);
   U20851 : OAI22_X1 port map( A1 => n27297, A2 => n27131, B1 => n27125, B2 => 
                           n20766, ZN => n7239);
   U20852 : OAI22_X1 port map( A1 => n27300, A2 => n27131, B1 => n27125, B2 => 
                           n20765, ZN => n7240);
   U20853 : OAI22_X1 port map( A1 => n27303, A2 => n27131, B1 => n27125, B2 => 
                           n20764, ZN => n7241);
   U20854 : OAI22_X1 port map( A1 => n27306, A2 => n27131, B1 => n27125, B2 => 
                           n20763, ZN => n7242);
   U20855 : OAI22_X1 port map( A1 => n27309, A2 => n27131, B1 => n27125, B2 => 
                           n20762, ZN => n7243);
   U20856 : OAI22_X1 port map( A1 => n27312, A2 => n27131, B1 => n27125, B2 => 
                           n20761, ZN => n7244);
   U20857 : OAI22_X1 port map( A1 => n27315, A2 => n27132, B1 => n27125, B2 => 
                           n20760, ZN => n7245);
   U20858 : NAND2_X1 port map( A1 => n25136, A2 => n25137, ZN => n5763);
   U20859 : NOR4_X1 port map( A1 => n25156, A2 => n25157, A3 => n25158, A4 => 
                           n25159, ZN => n25136);
   U20860 : NOR4_X1 port map( A1 => n25138, A2 => n25139, A3 => n25140, A4 => 
                           n25141, ZN => n25137);
   U20861 : OAI221_X1 port map( B1 => n21579, B2 => n26495, C1 => n21419, C2 =>
                           n26489, A => n25162, ZN => n25157);
   U20862 : NAND2_X1 port map( A1 => n25118, A2 => n25119, ZN => n5765);
   U20863 : NOR4_X1 port map( A1 => n25128, A2 => n25129, A3 => n25130, A4 => 
                           n25131, ZN => n25118);
   U20864 : NOR4_X1 port map( A1 => n25120, A2 => n25121, A3 => n25122, A4 => 
                           n25123, ZN => n25119);
   U20865 : OAI221_X1 port map( B1 => n21578, B2 => n26495, C1 => n21418, C2 =>
                           n26489, A => n25134, ZN => n25129);
   U20866 : NAND2_X1 port map( A1 => n25100, A2 => n25101, ZN => n5767);
   U20867 : NOR4_X1 port map( A1 => n25110, A2 => n25111, A3 => n25112, A4 => 
                           n25113, ZN => n25100);
   U20868 : NOR4_X1 port map( A1 => n25102, A2 => n25103, A3 => n25104, A4 => 
                           n25105, ZN => n25101);
   U20869 : OAI221_X1 port map( B1 => n21577, B2 => n26495, C1 => n21417, C2 =>
                           n26489, A => n25116, ZN => n25111);
   U20870 : NAND2_X1 port map( A1 => n25082, A2 => n25083, ZN => n5769);
   U20871 : NOR4_X1 port map( A1 => n25092, A2 => n25093, A3 => n25094, A4 => 
                           n25095, ZN => n25082);
   U20872 : NOR4_X1 port map( A1 => n25084, A2 => n25085, A3 => n25086, A4 => 
                           n25087, ZN => n25083);
   U20873 : OAI221_X1 port map( B1 => n21576, B2 => n26495, C1 => n21416, C2 =>
                           n26489, A => n25098, ZN => n25093);
   U20874 : NAND2_X1 port map( A1 => n25064, A2 => n25065, ZN => n5771);
   U20875 : NOR4_X1 port map( A1 => n25074, A2 => n25075, A3 => n25076, A4 => 
                           n25077, ZN => n25064);
   U20876 : NOR4_X1 port map( A1 => n25066, A2 => n25067, A3 => n25068, A4 => 
                           n25069, ZN => n25065);
   U20877 : OAI221_X1 port map( B1 => n21575, B2 => n26495, C1 => n21415, C2 =>
                           n26489, A => n25080, ZN => n25075);
   U20878 : NAND2_X1 port map( A1 => n25046, A2 => n25047, ZN => n5773);
   U20879 : NOR4_X1 port map( A1 => n25056, A2 => n25057, A3 => n25058, A4 => 
                           n25059, ZN => n25046);
   U20880 : NOR4_X1 port map( A1 => n25048, A2 => n25049, A3 => n25050, A4 => 
                           n25051, ZN => n25047);
   U20881 : OAI221_X1 port map( B1 => n21574, B2 => n26495, C1 => n21414, C2 =>
                           n26489, A => n25062, ZN => n25057);
   U20882 : NAND2_X1 port map( A1 => n25028, A2 => n25029, ZN => n5775);
   U20883 : NOR4_X1 port map( A1 => n25038, A2 => n25039, A3 => n25040, A4 => 
                           n25041, ZN => n25028);
   U20884 : NOR4_X1 port map( A1 => n25030, A2 => n25031, A3 => n25032, A4 => 
                           n25033, ZN => n25029);
   U20885 : OAI221_X1 port map( B1 => n21573, B2 => n26495, C1 => n21413, C2 =>
                           n26489, A => n25044, ZN => n25039);
   U20886 : NAND2_X1 port map( A1 => n25010, A2 => n25011, ZN => n5777);
   U20887 : NOR4_X1 port map( A1 => n25020, A2 => n25021, A3 => n25022, A4 => 
                           n25023, ZN => n25010);
   U20888 : NOR4_X1 port map( A1 => n25012, A2 => n25013, A3 => n25014, A4 => 
                           n25015, ZN => n25011);
   U20889 : OAI221_X1 port map( B1 => n21572, B2 => n26495, C1 => n21412, C2 =>
                           n26489, A => n25026, ZN => n25021);
   U20890 : NAND2_X1 port map( A1 => n24992, A2 => n24993, ZN => n5779);
   U20891 : NOR4_X1 port map( A1 => n25002, A2 => n25003, A3 => n25004, A4 => 
                           n25005, ZN => n24992);
   U20892 : NOR4_X1 port map( A1 => n24994, A2 => n24995, A3 => n24996, A4 => 
                           n24997, ZN => n24993);
   U20893 : OAI221_X1 port map( B1 => n21571, B2 => n26495, C1 => n21411, C2 =>
                           n26489, A => n25008, ZN => n25003);
   U20894 : NAND2_X1 port map( A1 => n24974, A2 => n24975, ZN => n5781);
   U20895 : NOR4_X1 port map( A1 => n24984, A2 => n24985, A3 => n24986, A4 => 
                           n24987, ZN => n24974);
   U20896 : NOR4_X1 port map( A1 => n24976, A2 => n24977, A3 => n24978, A4 => 
                           n24979, ZN => n24975);
   U20897 : OAI221_X1 port map( B1 => n21570, B2 => n26495, C1 => n21410, C2 =>
                           n26489, A => n24990, ZN => n24985);
   U20898 : NAND2_X1 port map( A1 => n24956, A2 => n24957, ZN => n5783);
   U20899 : NOR4_X1 port map( A1 => n24966, A2 => n24967, A3 => n24968, A4 => 
                           n24969, ZN => n24956);
   U20900 : NOR4_X1 port map( A1 => n24958, A2 => n24959, A3 => n24960, A4 => 
                           n24961, ZN => n24957);
   U20901 : OAI221_X1 port map( B1 => n21569, B2 => n26495, C1 => n21409, C2 =>
                           n26489, A => n24972, ZN => n24967);
   U20902 : NAND2_X1 port map( A1 => n24938, A2 => n24939, ZN => n5785);
   U20903 : NOR4_X1 port map( A1 => n24948, A2 => n24949, A3 => n24950, A4 => 
                           n24951, ZN => n24938);
   U20904 : NOR4_X1 port map( A1 => n24940, A2 => n24941, A3 => n24942, A4 => 
                           n24943, ZN => n24939);
   U20905 : OAI221_X1 port map( B1 => n21568, B2 => n26495, C1 => n21408, C2 =>
                           n26489, A => n24954, ZN => n24949);
   U20906 : NAND2_X1 port map( A1 => n24920, A2 => n24921, ZN => n5787);
   U20907 : NOR4_X1 port map( A1 => n24930, A2 => n24931, A3 => n24932, A4 => 
                           n24933, ZN => n24920);
   U20908 : NOR4_X1 port map( A1 => n24922, A2 => n24923, A3 => n24924, A4 => 
                           n24925, ZN => n24921);
   U20909 : OAI221_X1 port map( B1 => n21567, B2 => n26496, C1 => n21407, C2 =>
                           n26490, A => n24936, ZN => n24931);
   U20910 : NAND2_X1 port map( A1 => n24902, A2 => n24903, ZN => n5789);
   U20911 : NOR4_X1 port map( A1 => n24912, A2 => n24913, A3 => n24914, A4 => 
                           n24915, ZN => n24902);
   U20912 : NOR4_X1 port map( A1 => n24904, A2 => n24905, A3 => n24906, A4 => 
                           n24907, ZN => n24903);
   U20913 : OAI221_X1 port map( B1 => n21566, B2 => n26496, C1 => n21406, C2 =>
                           n26490, A => n24918, ZN => n24913);
   U20914 : NAND2_X1 port map( A1 => n24884, A2 => n24885, ZN => n5791);
   U20915 : NOR4_X1 port map( A1 => n24894, A2 => n24895, A3 => n24896, A4 => 
                           n24897, ZN => n24884);
   U20916 : NOR4_X1 port map( A1 => n24886, A2 => n24887, A3 => n24888, A4 => 
                           n24889, ZN => n24885);
   U20917 : OAI221_X1 port map( B1 => n21565, B2 => n26496, C1 => n21405, C2 =>
                           n26490, A => n24900, ZN => n24895);
   U20918 : NAND2_X1 port map( A1 => n24866, A2 => n24867, ZN => n5793);
   U20919 : NOR4_X1 port map( A1 => n24876, A2 => n24877, A3 => n24878, A4 => 
                           n24879, ZN => n24866);
   U20920 : NOR4_X1 port map( A1 => n24868, A2 => n24869, A3 => n24870, A4 => 
                           n24871, ZN => n24867);
   U20921 : OAI221_X1 port map( B1 => n21564, B2 => n26496, C1 => n21404, C2 =>
                           n26490, A => n24882, ZN => n24877);
   U20922 : NAND2_X1 port map( A1 => n24848, A2 => n24849, ZN => n5795);
   U20923 : NOR4_X1 port map( A1 => n24858, A2 => n24859, A3 => n24860, A4 => 
                           n24861, ZN => n24848);
   U20924 : NOR4_X1 port map( A1 => n24850, A2 => n24851, A3 => n24852, A4 => 
                           n24853, ZN => n24849);
   U20925 : OAI221_X1 port map( B1 => n21563, B2 => n26496, C1 => n21403, C2 =>
                           n26490, A => n24864, ZN => n24859);
   U20926 : NAND2_X1 port map( A1 => n24830, A2 => n24831, ZN => n5797);
   U20927 : NOR4_X1 port map( A1 => n24840, A2 => n24841, A3 => n24842, A4 => 
                           n24843, ZN => n24830);
   U20928 : NOR4_X1 port map( A1 => n24832, A2 => n24833, A3 => n24834, A4 => 
                           n24835, ZN => n24831);
   U20929 : OAI221_X1 port map( B1 => n21562, B2 => n26496, C1 => n21402, C2 =>
                           n26490, A => n24846, ZN => n24841);
   U20930 : NAND2_X1 port map( A1 => n24812, A2 => n24813, ZN => n5799);
   U20931 : NOR4_X1 port map( A1 => n24822, A2 => n24823, A3 => n24824, A4 => 
                           n24825, ZN => n24812);
   U20932 : NOR4_X1 port map( A1 => n24814, A2 => n24815, A3 => n24816, A4 => 
                           n24817, ZN => n24813);
   U20933 : OAI221_X1 port map( B1 => n21561, B2 => n26496, C1 => n21401, C2 =>
                           n26490, A => n24828, ZN => n24823);
   U20934 : NAND2_X1 port map( A1 => n24794, A2 => n24795, ZN => n5801);
   U20935 : NOR4_X1 port map( A1 => n24804, A2 => n24805, A3 => n24806, A4 => 
                           n24807, ZN => n24794);
   U20936 : NOR4_X1 port map( A1 => n24796, A2 => n24797, A3 => n24798, A4 => 
                           n24799, ZN => n24795);
   U20937 : OAI221_X1 port map( B1 => n21560, B2 => n26496, C1 => n21400, C2 =>
                           n26490, A => n24810, ZN => n24805);
   U20938 : NAND2_X1 port map( A1 => n24776, A2 => n24777, ZN => n5803);
   U20939 : NOR4_X1 port map( A1 => n24786, A2 => n24787, A3 => n24788, A4 => 
                           n24789, ZN => n24776);
   U20940 : NOR4_X1 port map( A1 => n24778, A2 => n24779, A3 => n24780, A4 => 
                           n24781, ZN => n24777);
   U20941 : OAI221_X1 port map( B1 => n21559, B2 => n26496, C1 => n21399, C2 =>
                           n26490, A => n24792, ZN => n24787);
   U20942 : NAND2_X1 port map( A1 => n24758, A2 => n24759, ZN => n5805);
   U20943 : NOR4_X1 port map( A1 => n24768, A2 => n24769, A3 => n24770, A4 => 
                           n24771, ZN => n24758);
   U20944 : NOR4_X1 port map( A1 => n24760, A2 => n24761, A3 => n24762, A4 => 
                           n24763, ZN => n24759);
   U20945 : OAI221_X1 port map( B1 => n21558, B2 => n26496, C1 => n21398, C2 =>
                           n26490, A => n24774, ZN => n24769);
   U20946 : NAND2_X1 port map( A1 => n24740, A2 => n24741, ZN => n5807);
   U20947 : NOR4_X1 port map( A1 => n24750, A2 => n24751, A3 => n24752, A4 => 
                           n24753, ZN => n24740);
   U20948 : NOR4_X1 port map( A1 => n24742, A2 => n24743, A3 => n24744, A4 => 
                           n24745, ZN => n24741);
   U20949 : OAI221_X1 port map( B1 => n21557, B2 => n26496, C1 => n21397, C2 =>
                           n26490, A => n24756, ZN => n24751);
   U20950 : NAND2_X1 port map( A1 => n24722, A2 => n24723, ZN => n5809);
   U20951 : NOR4_X1 port map( A1 => n24732, A2 => n24733, A3 => n24734, A4 => 
                           n24735, ZN => n24722);
   U20952 : NOR4_X1 port map( A1 => n24724, A2 => n24725, A3 => n24726, A4 => 
                           n24727, ZN => n24723);
   U20953 : OAI221_X1 port map( B1 => n21556, B2 => n26496, C1 => n21396, C2 =>
                           n26490, A => n24738, ZN => n24733);
   U20954 : NAND2_X1 port map( A1 => n24704, A2 => n24705, ZN => n5811);
   U20955 : NOR4_X1 port map( A1 => n24714, A2 => n24715, A3 => n24716, A4 => 
                           n24717, ZN => n24704);
   U20956 : NOR4_X1 port map( A1 => n24706, A2 => n24707, A3 => n24708, A4 => 
                           n24709, ZN => n24705);
   U20957 : OAI221_X1 port map( B1 => n21555, B2 => n26497, C1 => n21395, C2 =>
                           n26491, A => n24720, ZN => n24715);
   U20958 : NAND2_X1 port map( A1 => n24686, A2 => n24687, ZN => n5813);
   U20959 : NOR4_X1 port map( A1 => n24696, A2 => n24697, A3 => n24698, A4 => 
                           n24699, ZN => n24686);
   U20960 : NOR4_X1 port map( A1 => n24688, A2 => n24689, A3 => n24690, A4 => 
                           n24691, ZN => n24687);
   U20961 : OAI221_X1 port map( B1 => n21554, B2 => n26497, C1 => n21394, C2 =>
                           n26491, A => n24702, ZN => n24697);
   U20962 : NAND2_X1 port map( A1 => n24668, A2 => n24669, ZN => n5815);
   U20963 : NOR4_X1 port map( A1 => n24678, A2 => n24679, A3 => n24680, A4 => 
                           n24681, ZN => n24668);
   U20964 : NOR4_X1 port map( A1 => n24670, A2 => n24671, A3 => n24672, A4 => 
                           n24673, ZN => n24669);
   U20965 : OAI221_X1 port map( B1 => n21553, B2 => n26497, C1 => n21393, C2 =>
                           n26491, A => n24684, ZN => n24679);
   U20966 : NAND2_X1 port map( A1 => n24650, A2 => n24651, ZN => n5817);
   U20967 : NOR4_X1 port map( A1 => n24660, A2 => n24661, A3 => n24662, A4 => 
                           n24663, ZN => n24650);
   U20968 : NOR4_X1 port map( A1 => n24652, A2 => n24653, A3 => n24654, A4 => 
                           n24655, ZN => n24651);
   U20969 : OAI221_X1 port map( B1 => n21552, B2 => n26497, C1 => n21392, C2 =>
                           n26491, A => n24666, ZN => n24661);
   U20970 : NAND2_X1 port map( A1 => n24632, A2 => n24633, ZN => n5819);
   U20971 : NOR4_X1 port map( A1 => n24642, A2 => n24643, A3 => n24644, A4 => 
                           n24645, ZN => n24632);
   U20972 : NOR4_X1 port map( A1 => n24634, A2 => n24635, A3 => n24636, A4 => 
                           n24637, ZN => n24633);
   U20973 : OAI221_X1 port map( B1 => n21551, B2 => n26497, C1 => n21391, C2 =>
                           n26491, A => n24648, ZN => n24643);
   U20974 : NAND2_X1 port map( A1 => n24614, A2 => n24615, ZN => n5821);
   U20975 : NOR4_X1 port map( A1 => n24624, A2 => n24625, A3 => n24626, A4 => 
                           n24627, ZN => n24614);
   U20976 : NOR4_X1 port map( A1 => n24616, A2 => n24617, A3 => n24618, A4 => 
                           n24619, ZN => n24615);
   U20977 : OAI221_X1 port map( B1 => n21550, B2 => n26497, C1 => n21390, C2 =>
                           n26491, A => n24630, ZN => n24625);
   U20978 : NAND2_X1 port map( A1 => n24596, A2 => n24597, ZN => n5823);
   U20979 : NOR4_X1 port map( A1 => n24606, A2 => n24607, A3 => n24608, A4 => 
                           n24609, ZN => n24596);
   U20980 : NOR4_X1 port map( A1 => n24598, A2 => n24599, A3 => n24600, A4 => 
                           n24601, ZN => n24597);
   U20981 : OAI221_X1 port map( B1 => n21549, B2 => n26497, C1 => n21389, C2 =>
                           n26491, A => n24612, ZN => n24607);
   U20982 : NAND2_X1 port map( A1 => n24578, A2 => n24579, ZN => n5825);
   U20983 : NOR4_X1 port map( A1 => n24588, A2 => n24589, A3 => n24590, A4 => 
                           n24591, ZN => n24578);
   U20984 : NOR4_X1 port map( A1 => n24580, A2 => n24581, A3 => n24582, A4 => 
                           n24583, ZN => n24579);
   U20985 : OAI221_X1 port map( B1 => n21548, B2 => n26497, C1 => n21388, C2 =>
                           n26491, A => n24594, ZN => n24589);
   U20986 : NAND2_X1 port map( A1 => n24560, A2 => n24561, ZN => n5827);
   U20987 : NOR4_X1 port map( A1 => n24570, A2 => n24571, A3 => n24572, A4 => 
                           n24573, ZN => n24560);
   U20988 : NOR4_X1 port map( A1 => n24562, A2 => n24563, A3 => n24564, A4 => 
                           n24565, ZN => n24561);
   U20989 : OAI221_X1 port map( B1 => n21547, B2 => n26497, C1 => n21387, C2 =>
                           n26491, A => n24576, ZN => n24571);
   U20990 : NAND2_X1 port map( A1 => n24542, A2 => n24543, ZN => n5829);
   U20991 : NOR4_X1 port map( A1 => n24552, A2 => n24553, A3 => n24554, A4 => 
                           n24555, ZN => n24542);
   U20992 : NOR4_X1 port map( A1 => n24544, A2 => n24545, A3 => n24546, A4 => 
                           n24547, ZN => n24543);
   U20993 : OAI221_X1 port map( B1 => n21546, B2 => n26497, C1 => n21386, C2 =>
                           n26491, A => n24558, ZN => n24553);
   U20994 : NAND2_X1 port map( A1 => n24524, A2 => n24525, ZN => n5831);
   U20995 : NOR4_X1 port map( A1 => n24534, A2 => n24535, A3 => n24536, A4 => 
                           n24537, ZN => n24524);
   U20996 : NOR4_X1 port map( A1 => n24526, A2 => n24527, A3 => n24528, A4 => 
                           n24529, ZN => n24525);
   U20997 : OAI221_X1 port map( B1 => n21545, B2 => n26497, C1 => n21385, C2 =>
                           n26491, A => n24540, ZN => n24535);
   U20998 : NAND2_X1 port map( A1 => n24506, A2 => n24507, ZN => n5833);
   U20999 : NOR4_X1 port map( A1 => n24516, A2 => n24517, A3 => n24518, A4 => 
                           n24519, ZN => n24506);
   U21000 : NOR4_X1 port map( A1 => n24508, A2 => n24509, A3 => n24510, A4 => 
                           n24511, ZN => n24507);
   U21001 : OAI221_X1 port map( B1 => n21544, B2 => n26497, C1 => n21384, C2 =>
                           n26491, A => n24522, ZN => n24517);
   U21002 : NAND2_X1 port map( A1 => n24488, A2 => n24489, ZN => n5835);
   U21003 : NOR4_X1 port map( A1 => n24498, A2 => n24499, A3 => n24500, A4 => 
                           n24501, ZN => n24488);
   U21004 : NOR4_X1 port map( A1 => n24490, A2 => n24491, A3 => n24492, A4 => 
                           n24493, ZN => n24489);
   U21005 : OAI221_X1 port map( B1 => n21543, B2 => n26498, C1 => n21383, C2 =>
                           n26492, A => n24504, ZN => n24499);
   U21006 : NAND2_X1 port map( A1 => n24470, A2 => n24471, ZN => n5837);
   U21007 : NOR4_X1 port map( A1 => n24480, A2 => n24481, A3 => n24482, A4 => 
                           n24483, ZN => n24470);
   U21008 : NOR4_X1 port map( A1 => n24472, A2 => n24473, A3 => n24474, A4 => 
                           n24475, ZN => n24471);
   U21009 : OAI221_X1 port map( B1 => n21542, B2 => n26498, C1 => n21382, C2 =>
                           n26492, A => n24486, ZN => n24481);
   U21010 : NAND2_X1 port map( A1 => n24452, A2 => n24453, ZN => n5839);
   U21011 : NOR4_X1 port map( A1 => n24462, A2 => n24463, A3 => n24464, A4 => 
                           n24465, ZN => n24452);
   U21012 : NOR4_X1 port map( A1 => n24454, A2 => n24455, A3 => n24456, A4 => 
                           n24457, ZN => n24453);
   U21013 : OAI221_X1 port map( B1 => n21541, B2 => n26498, C1 => n21381, C2 =>
                           n26492, A => n24468, ZN => n24463);
   U21014 : NAND2_X1 port map( A1 => n24434, A2 => n24435, ZN => n5841);
   U21015 : NOR4_X1 port map( A1 => n24444, A2 => n24445, A3 => n24446, A4 => 
                           n24447, ZN => n24434);
   U21016 : NOR4_X1 port map( A1 => n24436, A2 => n24437, A3 => n24438, A4 => 
                           n24439, ZN => n24435);
   U21017 : OAI221_X1 port map( B1 => n21540, B2 => n26498, C1 => n21380, C2 =>
                           n26492, A => n24450, ZN => n24445);
   U21018 : NAND2_X1 port map( A1 => n24416, A2 => n24417, ZN => n5843);
   U21019 : NOR4_X1 port map( A1 => n24426, A2 => n24427, A3 => n24428, A4 => 
                           n24429, ZN => n24416);
   U21020 : NOR4_X1 port map( A1 => n24418, A2 => n24419, A3 => n24420, A4 => 
                           n24421, ZN => n24417);
   U21021 : OAI221_X1 port map( B1 => n21539, B2 => n26498, C1 => n21379, C2 =>
                           n26492, A => n24432, ZN => n24427);
   U21022 : NAND2_X1 port map( A1 => n24398, A2 => n24399, ZN => n5845);
   U21023 : NOR4_X1 port map( A1 => n24408, A2 => n24409, A3 => n24410, A4 => 
                           n24411, ZN => n24398);
   U21024 : NOR4_X1 port map( A1 => n24400, A2 => n24401, A3 => n24402, A4 => 
                           n24403, ZN => n24399);
   U21025 : OAI221_X1 port map( B1 => n21538, B2 => n26498, C1 => n21378, C2 =>
                           n26492, A => n24414, ZN => n24409);
   U21026 : NAND2_X1 port map( A1 => n24380, A2 => n24381, ZN => n5847);
   U21027 : NOR4_X1 port map( A1 => n24390, A2 => n24391, A3 => n24392, A4 => 
                           n24393, ZN => n24380);
   U21028 : NOR4_X1 port map( A1 => n24382, A2 => n24383, A3 => n24384, A4 => 
                           n24385, ZN => n24381);
   U21029 : OAI221_X1 port map( B1 => n21537, B2 => n26498, C1 => n21377, C2 =>
                           n26492, A => n24396, ZN => n24391);
   U21030 : NAND2_X1 port map( A1 => n24362, A2 => n24363, ZN => n5849);
   U21031 : NOR4_X1 port map( A1 => n24372, A2 => n24373, A3 => n24374, A4 => 
                           n24375, ZN => n24362);
   U21032 : NOR4_X1 port map( A1 => n24364, A2 => n24365, A3 => n24366, A4 => 
                           n24367, ZN => n24363);
   U21033 : OAI221_X1 port map( B1 => n21536, B2 => n26498, C1 => n21376, C2 =>
                           n26492, A => n24378, ZN => n24373);
   U21034 : NAND2_X1 port map( A1 => n24344, A2 => n24345, ZN => n5851);
   U21035 : NOR4_X1 port map( A1 => n24354, A2 => n24355, A3 => n24356, A4 => 
                           n24357, ZN => n24344);
   U21036 : NOR4_X1 port map( A1 => n24346, A2 => n24347, A3 => n24348, A4 => 
                           n24349, ZN => n24345);
   U21037 : OAI221_X1 port map( B1 => n21535, B2 => n26498, C1 => n21375, C2 =>
                           n26492, A => n24360, ZN => n24355);
   U21038 : NAND2_X1 port map( A1 => n24326, A2 => n24327, ZN => n5853);
   U21039 : NOR4_X1 port map( A1 => n24336, A2 => n24337, A3 => n24338, A4 => 
                           n24339, ZN => n24326);
   U21040 : NOR4_X1 port map( A1 => n24328, A2 => n24329, A3 => n24330, A4 => 
                           n24331, ZN => n24327);
   U21041 : OAI221_X1 port map( B1 => n21534, B2 => n26498, C1 => n21374, C2 =>
                           n26492, A => n24342, ZN => n24337);
   U21042 : NAND2_X1 port map( A1 => n24308, A2 => n24309, ZN => n5855);
   U21043 : NOR4_X1 port map( A1 => n24318, A2 => n24319, A3 => n24320, A4 => 
                           n24321, ZN => n24308);
   U21044 : NOR4_X1 port map( A1 => n24310, A2 => n24311, A3 => n24312, A4 => 
                           n24313, ZN => n24309);
   U21045 : OAI221_X1 port map( B1 => n21533, B2 => n26498, C1 => n21373, C2 =>
                           n26492, A => n24324, ZN => n24319);
   U21046 : NAND2_X1 port map( A1 => n24290, A2 => n24291, ZN => n5857);
   U21047 : NOR4_X1 port map( A1 => n24300, A2 => n24301, A3 => n24302, A4 => 
                           n24303, ZN => n24290);
   U21048 : NOR4_X1 port map( A1 => n24292, A2 => n24293, A3 => n24294, A4 => 
                           n24295, ZN => n24291);
   U21049 : OAI221_X1 port map( B1 => n21532, B2 => n26498, C1 => n21372, C2 =>
                           n26492, A => n24306, ZN => n24301);
   U21050 : NAND2_X1 port map( A1 => n23937, A2 => n23938, ZN => n5891);
   U21051 : NOR4_X1 port map( A1 => n23957, A2 => n23958, A3 => n23959, A4 => 
                           n23960, ZN => n23937);
   U21052 : NOR4_X1 port map( A1 => n23939, A2 => n23940, A3 => n23941, A4 => 
                           n23942, ZN => n23938);
   U21053 : OAI221_X1 port map( B1 => n21579, B2 => n26720, C1 => n21419, C2 =>
                           n26714, A => n23963, ZN => n23958);
   U21054 : NAND2_X1 port map( A1 => n23919, A2 => n23920, ZN => n5893);
   U21055 : NOR4_X1 port map( A1 => n23929, A2 => n23930, A3 => n23931, A4 => 
                           n23932, ZN => n23919);
   U21056 : NOR4_X1 port map( A1 => n23921, A2 => n23922, A3 => n23923, A4 => 
                           n23924, ZN => n23920);
   U21057 : OAI221_X1 port map( B1 => n21578, B2 => n26720, C1 => n21418, C2 =>
                           n26714, A => n23935, ZN => n23930);
   U21058 : NAND2_X1 port map( A1 => n23901, A2 => n23902, ZN => n5895);
   U21059 : NOR4_X1 port map( A1 => n23911, A2 => n23912, A3 => n23913, A4 => 
                           n23914, ZN => n23901);
   U21060 : NOR4_X1 port map( A1 => n23903, A2 => n23904, A3 => n23905, A4 => 
                           n23906, ZN => n23902);
   U21061 : OAI221_X1 port map( B1 => n21577, B2 => n26720, C1 => n21417, C2 =>
                           n26714, A => n23917, ZN => n23912);
   U21062 : NAND2_X1 port map( A1 => n23883, A2 => n23884, ZN => n5897);
   U21063 : NOR4_X1 port map( A1 => n23893, A2 => n23894, A3 => n23895, A4 => 
                           n23896, ZN => n23883);
   U21064 : NOR4_X1 port map( A1 => n23885, A2 => n23886, A3 => n23887, A4 => 
                           n23888, ZN => n23884);
   U21065 : OAI221_X1 port map( B1 => n21576, B2 => n26720, C1 => n21416, C2 =>
                           n26714, A => n23899, ZN => n23894);
   U21066 : NAND2_X1 port map( A1 => n23865, A2 => n23866, ZN => n5899);
   U21067 : NOR4_X1 port map( A1 => n23875, A2 => n23876, A3 => n23877, A4 => 
                           n23878, ZN => n23865);
   U21068 : NOR4_X1 port map( A1 => n23867, A2 => n23868, A3 => n23869, A4 => 
                           n23870, ZN => n23866);
   U21069 : OAI221_X1 port map( B1 => n21575, B2 => n26720, C1 => n21415, C2 =>
                           n26714, A => n23881, ZN => n23876);
   U21070 : NAND2_X1 port map( A1 => n23847, A2 => n23848, ZN => n5901);
   U21071 : NOR4_X1 port map( A1 => n23857, A2 => n23858, A3 => n23859, A4 => 
                           n23860, ZN => n23847);
   U21072 : NOR4_X1 port map( A1 => n23849, A2 => n23850, A3 => n23851, A4 => 
                           n23852, ZN => n23848);
   U21073 : OAI221_X1 port map( B1 => n21574, B2 => n26720, C1 => n21414, C2 =>
                           n26714, A => n23863, ZN => n23858);
   U21074 : NAND2_X1 port map( A1 => n23829, A2 => n23830, ZN => n5903);
   U21075 : NOR4_X1 port map( A1 => n23839, A2 => n23840, A3 => n23841, A4 => 
                           n23842, ZN => n23829);
   U21076 : NOR4_X1 port map( A1 => n23831, A2 => n23832, A3 => n23833, A4 => 
                           n23834, ZN => n23830);
   U21077 : OAI221_X1 port map( B1 => n21573, B2 => n26720, C1 => n21413, C2 =>
                           n26714, A => n23845, ZN => n23840);
   U21078 : NAND2_X1 port map( A1 => n23811, A2 => n23812, ZN => n5905);
   U21079 : NOR4_X1 port map( A1 => n23821, A2 => n23822, A3 => n23823, A4 => 
                           n23824, ZN => n23811);
   U21080 : NOR4_X1 port map( A1 => n23813, A2 => n23814, A3 => n23815, A4 => 
                           n23816, ZN => n23812);
   U21081 : OAI221_X1 port map( B1 => n21572, B2 => n26720, C1 => n21412, C2 =>
                           n26714, A => n23827, ZN => n23822);
   U21082 : NAND2_X1 port map( A1 => n23793, A2 => n23794, ZN => n5907);
   U21083 : NOR4_X1 port map( A1 => n23803, A2 => n23804, A3 => n23805, A4 => 
                           n23806, ZN => n23793);
   U21084 : NOR4_X1 port map( A1 => n23795, A2 => n23796, A3 => n23797, A4 => 
                           n23798, ZN => n23794);
   U21085 : OAI221_X1 port map( B1 => n21571, B2 => n26720, C1 => n21411, C2 =>
                           n26714, A => n23809, ZN => n23804);
   U21086 : NAND2_X1 port map( A1 => n23775, A2 => n23776, ZN => n5909);
   U21087 : NOR4_X1 port map( A1 => n23785, A2 => n23786, A3 => n23787, A4 => 
                           n23788, ZN => n23775);
   U21088 : NOR4_X1 port map( A1 => n23777, A2 => n23778, A3 => n23779, A4 => 
                           n23780, ZN => n23776);
   U21089 : OAI221_X1 port map( B1 => n21570, B2 => n26720, C1 => n21410, C2 =>
                           n26714, A => n23791, ZN => n23786);
   U21090 : NAND2_X1 port map( A1 => n23757, A2 => n23758, ZN => n5911);
   U21091 : NOR4_X1 port map( A1 => n23767, A2 => n23768, A3 => n23769, A4 => 
                           n23770, ZN => n23757);
   U21092 : NOR4_X1 port map( A1 => n23759, A2 => n23760, A3 => n23761, A4 => 
                           n23762, ZN => n23758);
   U21093 : OAI221_X1 port map( B1 => n21569, B2 => n26720, C1 => n21409, C2 =>
                           n26714, A => n23773, ZN => n23768);
   U21094 : NAND2_X1 port map( A1 => n23739, A2 => n23740, ZN => n5913);
   U21095 : NOR4_X1 port map( A1 => n23749, A2 => n23750, A3 => n23751, A4 => 
                           n23752, ZN => n23739);
   U21096 : NOR4_X1 port map( A1 => n23741, A2 => n23742, A3 => n23743, A4 => 
                           n23744, ZN => n23740);
   U21097 : OAI221_X1 port map( B1 => n21568, B2 => n26720, C1 => n21408, C2 =>
                           n26714, A => n23755, ZN => n23750);
   U21098 : NAND2_X1 port map( A1 => n23721, A2 => n23722, ZN => n5915);
   U21099 : NOR4_X1 port map( A1 => n23731, A2 => n23732, A3 => n23733, A4 => 
                           n23734, ZN => n23721);
   U21100 : NOR4_X1 port map( A1 => n23723, A2 => n23724, A3 => n23725, A4 => 
                           n23726, ZN => n23722);
   U21101 : OAI221_X1 port map( B1 => n21567, B2 => n26721, C1 => n21407, C2 =>
                           n26715, A => n23737, ZN => n23732);
   U21102 : NAND2_X1 port map( A1 => n23703, A2 => n23704, ZN => n5917);
   U21103 : NOR4_X1 port map( A1 => n23713, A2 => n23714, A3 => n23715, A4 => 
                           n23716, ZN => n23703);
   U21104 : NOR4_X1 port map( A1 => n23705, A2 => n23706, A3 => n23707, A4 => 
                           n23708, ZN => n23704);
   U21105 : OAI221_X1 port map( B1 => n21566, B2 => n26721, C1 => n21406, C2 =>
                           n26715, A => n23719, ZN => n23714);
   U21106 : NAND2_X1 port map( A1 => n23685, A2 => n23686, ZN => n5919);
   U21107 : NOR4_X1 port map( A1 => n23695, A2 => n23696, A3 => n23697, A4 => 
                           n23698, ZN => n23685);
   U21108 : NOR4_X1 port map( A1 => n23687, A2 => n23688, A3 => n23689, A4 => 
                           n23690, ZN => n23686);
   U21109 : OAI221_X1 port map( B1 => n21565, B2 => n26721, C1 => n21405, C2 =>
                           n26715, A => n23701, ZN => n23696);
   U21110 : NAND2_X1 port map( A1 => n23667, A2 => n23668, ZN => n5921);
   U21111 : NOR4_X1 port map( A1 => n23677, A2 => n23678, A3 => n23679, A4 => 
                           n23680, ZN => n23667);
   U21112 : NOR4_X1 port map( A1 => n23669, A2 => n23670, A3 => n23671, A4 => 
                           n23672, ZN => n23668);
   U21113 : OAI221_X1 port map( B1 => n21564, B2 => n26721, C1 => n21404, C2 =>
                           n26715, A => n23683, ZN => n23678);
   U21114 : NAND2_X1 port map( A1 => n23649, A2 => n23650, ZN => n5923);
   U21115 : NOR4_X1 port map( A1 => n23659, A2 => n23660, A3 => n23661, A4 => 
                           n23662, ZN => n23649);
   U21116 : NOR4_X1 port map( A1 => n23651, A2 => n23652, A3 => n23653, A4 => 
                           n23654, ZN => n23650);
   U21117 : OAI221_X1 port map( B1 => n21563, B2 => n26721, C1 => n21403, C2 =>
                           n26715, A => n23665, ZN => n23660);
   U21118 : NAND2_X1 port map( A1 => n23631, A2 => n23632, ZN => n5925);
   U21119 : NOR4_X1 port map( A1 => n23641, A2 => n23642, A3 => n23643, A4 => 
                           n23644, ZN => n23631);
   U21120 : NOR4_X1 port map( A1 => n23633, A2 => n23634, A3 => n23635, A4 => 
                           n23636, ZN => n23632);
   U21121 : OAI221_X1 port map( B1 => n21562, B2 => n26721, C1 => n21402, C2 =>
                           n26715, A => n23647, ZN => n23642);
   U21122 : NAND2_X1 port map( A1 => n23613, A2 => n23614, ZN => n5927);
   U21123 : NOR4_X1 port map( A1 => n23623, A2 => n23624, A3 => n23625, A4 => 
                           n23626, ZN => n23613);
   U21124 : NOR4_X1 port map( A1 => n23615, A2 => n23616, A3 => n23617, A4 => 
                           n23618, ZN => n23614);
   U21125 : OAI221_X1 port map( B1 => n21561, B2 => n26721, C1 => n21401, C2 =>
                           n26715, A => n23629, ZN => n23624);
   U21126 : NAND2_X1 port map( A1 => n23595, A2 => n23596, ZN => n5929);
   U21127 : NOR4_X1 port map( A1 => n23605, A2 => n23606, A3 => n23607, A4 => 
                           n23608, ZN => n23595);
   U21128 : NOR4_X1 port map( A1 => n23597, A2 => n23598, A3 => n23599, A4 => 
                           n23600, ZN => n23596);
   U21129 : OAI221_X1 port map( B1 => n21560, B2 => n26721, C1 => n21400, C2 =>
                           n26715, A => n23611, ZN => n23606);
   U21130 : NAND2_X1 port map( A1 => n23577, A2 => n23578, ZN => n5931);
   U21131 : NOR4_X1 port map( A1 => n23587, A2 => n23588, A3 => n23589, A4 => 
                           n23590, ZN => n23577);
   U21132 : NOR4_X1 port map( A1 => n23579, A2 => n23580, A3 => n23581, A4 => 
                           n23582, ZN => n23578);
   U21133 : OAI221_X1 port map( B1 => n21559, B2 => n26721, C1 => n21399, C2 =>
                           n26715, A => n23593, ZN => n23588);
   U21134 : NAND2_X1 port map( A1 => n23559, A2 => n23560, ZN => n5933);
   U21135 : NOR4_X1 port map( A1 => n23569, A2 => n23570, A3 => n23571, A4 => 
                           n23572, ZN => n23559);
   U21136 : NOR4_X1 port map( A1 => n23561, A2 => n23562, A3 => n23563, A4 => 
                           n23564, ZN => n23560);
   U21137 : OAI221_X1 port map( B1 => n21558, B2 => n26721, C1 => n21398, C2 =>
                           n26715, A => n23575, ZN => n23570);
   U21138 : NAND2_X1 port map( A1 => n23541, A2 => n23542, ZN => n5935);
   U21139 : NOR4_X1 port map( A1 => n23551, A2 => n23552, A3 => n23553, A4 => 
                           n23554, ZN => n23541);
   U21140 : NOR4_X1 port map( A1 => n23543, A2 => n23544, A3 => n23545, A4 => 
                           n23546, ZN => n23542);
   U21141 : OAI221_X1 port map( B1 => n21557, B2 => n26721, C1 => n21397, C2 =>
                           n26715, A => n23557, ZN => n23552);
   U21142 : NAND2_X1 port map( A1 => n23523, A2 => n23524, ZN => n5937);
   U21143 : NOR4_X1 port map( A1 => n23533, A2 => n23534, A3 => n23535, A4 => 
                           n23536, ZN => n23523);
   U21144 : NOR4_X1 port map( A1 => n23525, A2 => n23526, A3 => n23527, A4 => 
                           n23528, ZN => n23524);
   U21145 : OAI221_X1 port map( B1 => n21556, B2 => n26721, C1 => n21396, C2 =>
                           n26715, A => n23539, ZN => n23534);
   U21146 : NAND2_X1 port map( A1 => n23505, A2 => n23506, ZN => n5939);
   U21147 : NOR4_X1 port map( A1 => n23515, A2 => n23516, A3 => n23517, A4 => 
                           n23518, ZN => n23505);
   U21148 : NOR4_X1 port map( A1 => n23507, A2 => n23508, A3 => n23509, A4 => 
                           n23510, ZN => n23506);
   U21149 : OAI221_X1 port map( B1 => n21555, B2 => n26722, C1 => n21395, C2 =>
                           n26716, A => n23521, ZN => n23516);
   U21150 : NAND2_X1 port map( A1 => n23487, A2 => n23488, ZN => n5941);
   U21151 : NOR4_X1 port map( A1 => n23497, A2 => n23498, A3 => n23499, A4 => 
                           n23500, ZN => n23487);
   U21152 : NOR4_X1 port map( A1 => n23489, A2 => n23490, A3 => n23491, A4 => 
                           n23492, ZN => n23488);
   U21153 : OAI221_X1 port map( B1 => n21554, B2 => n26722, C1 => n21394, C2 =>
                           n26716, A => n23503, ZN => n23498);
   U21154 : NAND2_X1 port map( A1 => n23469, A2 => n23470, ZN => n5943);
   U21155 : NOR4_X1 port map( A1 => n23479, A2 => n23480, A3 => n23481, A4 => 
                           n23482, ZN => n23469);
   U21156 : NOR4_X1 port map( A1 => n23471, A2 => n23472, A3 => n23473, A4 => 
                           n23474, ZN => n23470);
   U21157 : OAI221_X1 port map( B1 => n21553, B2 => n26722, C1 => n21393, C2 =>
                           n26716, A => n23485, ZN => n23480);
   U21158 : NAND2_X1 port map( A1 => n23451, A2 => n23452, ZN => n5945);
   U21159 : NOR4_X1 port map( A1 => n23461, A2 => n23462, A3 => n23463, A4 => 
                           n23464, ZN => n23451);
   U21160 : NOR4_X1 port map( A1 => n23453, A2 => n23454, A3 => n23455, A4 => 
                           n23456, ZN => n23452);
   U21161 : OAI221_X1 port map( B1 => n21552, B2 => n26722, C1 => n21392, C2 =>
                           n26716, A => n23467, ZN => n23462);
   U21162 : NAND2_X1 port map( A1 => n23433, A2 => n23434, ZN => n5947);
   U21163 : NOR4_X1 port map( A1 => n23443, A2 => n23444, A3 => n23445, A4 => 
                           n23446, ZN => n23433);
   U21164 : NOR4_X1 port map( A1 => n23435, A2 => n23436, A3 => n23437, A4 => 
                           n23438, ZN => n23434);
   U21165 : OAI221_X1 port map( B1 => n21551, B2 => n26722, C1 => n21391, C2 =>
                           n26716, A => n23449, ZN => n23444);
   U21166 : NAND2_X1 port map( A1 => n23415, A2 => n23416, ZN => n5949);
   U21167 : NOR4_X1 port map( A1 => n23425, A2 => n23426, A3 => n23427, A4 => 
                           n23428, ZN => n23415);
   U21168 : NOR4_X1 port map( A1 => n23417, A2 => n23418, A3 => n23419, A4 => 
                           n23420, ZN => n23416);
   U21169 : OAI221_X1 port map( B1 => n21550, B2 => n26722, C1 => n21390, C2 =>
                           n26716, A => n23431, ZN => n23426);
   U21170 : NAND2_X1 port map( A1 => n23397, A2 => n23398, ZN => n5951);
   U21171 : NOR4_X1 port map( A1 => n23407, A2 => n23408, A3 => n23409, A4 => 
                           n23410, ZN => n23397);
   U21172 : NOR4_X1 port map( A1 => n23399, A2 => n23400, A3 => n23401, A4 => 
                           n23402, ZN => n23398);
   U21173 : OAI221_X1 port map( B1 => n21549, B2 => n26722, C1 => n21389, C2 =>
                           n26716, A => n23413, ZN => n23408);
   U21174 : NAND2_X1 port map( A1 => n23379, A2 => n23380, ZN => n5953);
   U21175 : NOR4_X1 port map( A1 => n23389, A2 => n23390, A3 => n23391, A4 => 
                           n23392, ZN => n23379);
   U21176 : NOR4_X1 port map( A1 => n23381, A2 => n23382, A3 => n23383, A4 => 
                           n23384, ZN => n23380);
   U21177 : OAI221_X1 port map( B1 => n21548, B2 => n26722, C1 => n21388, C2 =>
                           n26716, A => n23395, ZN => n23390);
   U21178 : NAND2_X1 port map( A1 => n23361, A2 => n23362, ZN => n5955);
   U21179 : NOR4_X1 port map( A1 => n23371, A2 => n23372, A3 => n23373, A4 => 
                           n23374, ZN => n23361);
   U21180 : NOR4_X1 port map( A1 => n23363, A2 => n23364, A3 => n23365, A4 => 
                           n23366, ZN => n23362);
   U21181 : OAI221_X1 port map( B1 => n21547, B2 => n26722, C1 => n21387, C2 =>
                           n26716, A => n23377, ZN => n23372);
   U21182 : NAND2_X1 port map( A1 => n23343, A2 => n23344, ZN => n5957);
   U21183 : NOR4_X1 port map( A1 => n23353, A2 => n23354, A3 => n23355, A4 => 
                           n23356, ZN => n23343);
   U21184 : NOR4_X1 port map( A1 => n23345, A2 => n23346, A3 => n23347, A4 => 
                           n23348, ZN => n23344);
   U21185 : OAI221_X1 port map( B1 => n21546, B2 => n26722, C1 => n21386, C2 =>
                           n26716, A => n23359, ZN => n23354);
   U21186 : NAND2_X1 port map( A1 => n23325, A2 => n23326, ZN => n5959);
   U21187 : NOR4_X1 port map( A1 => n23335, A2 => n23336, A3 => n23337, A4 => 
                           n23338, ZN => n23325);
   U21188 : NOR4_X1 port map( A1 => n23327, A2 => n23328, A3 => n23329, A4 => 
                           n23330, ZN => n23326);
   U21189 : OAI221_X1 port map( B1 => n21545, B2 => n26722, C1 => n21385, C2 =>
                           n26716, A => n23341, ZN => n23336);
   U21190 : NAND2_X1 port map( A1 => n23307, A2 => n23308, ZN => n5961);
   U21191 : NOR4_X1 port map( A1 => n23317, A2 => n23318, A3 => n23319, A4 => 
                           n23320, ZN => n23307);
   U21192 : NOR4_X1 port map( A1 => n23309, A2 => n23310, A3 => n23311, A4 => 
                           n23312, ZN => n23308);
   U21193 : OAI221_X1 port map( B1 => n21544, B2 => n26722, C1 => n21384, C2 =>
                           n26716, A => n23323, ZN => n23318);
   U21194 : NAND2_X1 port map( A1 => n23289, A2 => n23290, ZN => n5963);
   U21195 : NOR4_X1 port map( A1 => n23299, A2 => n23300, A3 => n23301, A4 => 
                           n23302, ZN => n23289);
   U21196 : NOR4_X1 port map( A1 => n23291, A2 => n23292, A3 => n23293, A4 => 
                           n23294, ZN => n23290);
   U21197 : OAI221_X1 port map( B1 => n21543, B2 => n26723, C1 => n21383, C2 =>
                           n26717, A => n23305, ZN => n23300);
   U21198 : NAND2_X1 port map( A1 => n23271, A2 => n23272, ZN => n5965);
   U21199 : NOR4_X1 port map( A1 => n23281, A2 => n23282, A3 => n23283, A4 => 
                           n23284, ZN => n23271);
   U21200 : NOR4_X1 port map( A1 => n23273, A2 => n23274, A3 => n23275, A4 => 
                           n23276, ZN => n23272);
   U21201 : OAI221_X1 port map( B1 => n21542, B2 => n26723, C1 => n21382, C2 =>
                           n26717, A => n23287, ZN => n23282);
   U21202 : NAND2_X1 port map( A1 => n23253, A2 => n23254, ZN => n5967);
   U21203 : NOR4_X1 port map( A1 => n23263, A2 => n23264, A3 => n23265, A4 => 
                           n23266, ZN => n23253);
   U21204 : NOR4_X1 port map( A1 => n23255, A2 => n23256, A3 => n23257, A4 => 
                           n23258, ZN => n23254);
   U21205 : OAI221_X1 port map( B1 => n21541, B2 => n26723, C1 => n21381, C2 =>
                           n26717, A => n23269, ZN => n23264);
   U21206 : NAND2_X1 port map( A1 => n23235, A2 => n23236, ZN => n5969);
   U21207 : NOR4_X1 port map( A1 => n23245, A2 => n23246, A3 => n23247, A4 => 
                           n23248, ZN => n23235);
   U21208 : NOR4_X1 port map( A1 => n23237, A2 => n23238, A3 => n23239, A4 => 
                           n23240, ZN => n23236);
   U21209 : OAI221_X1 port map( B1 => n21540, B2 => n26723, C1 => n21380, C2 =>
                           n26717, A => n23251, ZN => n23246);
   U21210 : NAND2_X1 port map( A1 => n23217, A2 => n23218, ZN => n5971);
   U21211 : NOR4_X1 port map( A1 => n23227, A2 => n23228, A3 => n23229, A4 => 
                           n23230, ZN => n23217);
   U21212 : NOR4_X1 port map( A1 => n23219, A2 => n23220, A3 => n23221, A4 => 
                           n23222, ZN => n23218);
   U21213 : OAI221_X1 port map( B1 => n21539, B2 => n26723, C1 => n21379, C2 =>
                           n26717, A => n23233, ZN => n23228);
   U21214 : NAND2_X1 port map( A1 => n23199, A2 => n23200, ZN => n5973);
   U21215 : NOR4_X1 port map( A1 => n23209, A2 => n23210, A3 => n23211, A4 => 
                           n23212, ZN => n23199);
   U21216 : NOR4_X1 port map( A1 => n23201, A2 => n23202, A3 => n23203, A4 => 
                           n23204, ZN => n23200);
   U21217 : OAI221_X1 port map( B1 => n21538, B2 => n26723, C1 => n21378, C2 =>
                           n26717, A => n23215, ZN => n23210);
   U21218 : NAND2_X1 port map( A1 => n23181, A2 => n23182, ZN => n5975);
   U21219 : NOR4_X1 port map( A1 => n23191, A2 => n23192, A3 => n23193, A4 => 
                           n23194, ZN => n23181);
   U21220 : NOR4_X1 port map( A1 => n23183, A2 => n23184, A3 => n23185, A4 => 
                           n23186, ZN => n23182);
   U21221 : OAI221_X1 port map( B1 => n21537, B2 => n26723, C1 => n21377, C2 =>
                           n26717, A => n23197, ZN => n23192);
   U21222 : NAND2_X1 port map( A1 => n23163, A2 => n23164, ZN => n5977);
   U21223 : NOR4_X1 port map( A1 => n23173, A2 => n23174, A3 => n23175, A4 => 
                           n23176, ZN => n23163);
   U21224 : NOR4_X1 port map( A1 => n23165, A2 => n23166, A3 => n23167, A4 => 
                           n23168, ZN => n23164);
   U21225 : OAI221_X1 port map( B1 => n21536, B2 => n26723, C1 => n21376, C2 =>
                           n26717, A => n23179, ZN => n23174);
   U21226 : NAND2_X1 port map( A1 => n23145, A2 => n23146, ZN => n5979);
   U21227 : NOR4_X1 port map( A1 => n23155, A2 => n23156, A3 => n23157, A4 => 
                           n23158, ZN => n23145);
   U21228 : NOR4_X1 port map( A1 => n23147, A2 => n23148, A3 => n23149, A4 => 
                           n23150, ZN => n23146);
   U21229 : OAI221_X1 port map( B1 => n21535, B2 => n26723, C1 => n21375, C2 =>
                           n26717, A => n23161, ZN => n23156);
   U21230 : NAND2_X1 port map( A1 => n23127, A2 => n23128, ZN => n5981);
   U21231 : NOR4_X1 port map( A1 => n23137, A2 => n23138, A3 => n23139, A4 => 
                           n23140, ZN => n23127);
   U21232 : NOR4_X1 port map( A1 => n23129, A2 => n23130, A3 => n23131, A4 => 
                           n23132, ZN => n23128);
   U21233 : OAI221_X1 port map( B1 => n21534, B2 => n26723, C1 => n21374, C2 =>
                           n26717, A => n23143, ZN => n23138);
   U21234 : NAND2_X1 port map( A1 => n23109, A2 => n23110, ZN => n5983);
   U21235 : NOR4_X1 port map( A1 => n23119, A2 => n23120, A3 => n23121, A4 => 
                           n23122, ZN => n23109);
   U21236 : NOR4_X1 port map( A1 => n23111, A2 => n23112, A3 => n23113, A4 => 
                           n23114, ZN => n23110);
   U21237 : OAI221_X1 port map( B1 => n21533, B2 => n26723, C1 => n21373, C2 =>
                           n26717, A => n23125, ZN => n23120);
   U21238 : NAND2_X1 port map( A1 => n23091, A2 => n23092, ZN => n5985);
   U21239 : NOR4_X1 port map( A1 => n23101, A2 => n23102, A3 => n23103, A4 => 
                           n23104, ZN => n23091);
   U21240 : NOR4_X1 port map( A1 => n23093, A2 => n23094, A3 => n23095, A4 => 
                           n23096, ZN => n23092);
   U21241 : OAI221_X1 port map( B1 => n21532, B2 => n26723, C1 => n21372, C2 =>
                           n26717, A => n23107, ZN => n23102);
   U21242 : NAND2_X1 port map( A1 => n23968, A2 => n23969, ZN => n5889);
   U21243 : NOR4_X1 port map( A1 => n23995, A2 => n23996, A3 => n23997, A4 => 
                           n23998, ZN => n23968);
   U21244 : NOR4_X1 port map( A1 => n23970, A2 => n23971, A3 => n23972, A4 => 
                           n23973, ZN => n23969);
   U21245 : OAI221_X1 port map( B1 => n21176, B2 => n26500, C1 => n21168, C2 =>
                           n26494, A => n24011, ZN => n23996);
   U21246 : NAND2_X1 port map( A1 => n24056, A2 => n24057, ZN => n5883);
   U21247 : NOR4_X1 port map( A1 => n24066, A2 => n24067, A3 => n24068, A4 => 
                           n24069, ZN => n24056);
   U21248 : NOR4_X1 port map( A1 => n24058, A2 => n24059, A3 => n24060, A4 => 
                           n24061, ZN => n24057);
   U21249 : OAI221_X1 port map( B1 => n21179, B2 => n26500, C1 => n21171, C2 =>
                           n26494, A => n24072, ZN => n24067);
   U21250 : NAND2_X1 port map( A1 => n24038, A2 => n24039, ZN => n5885);
   U21251 : NOR4_X1 port map( A1 => n24048, A2 => n24049, A3 => n24050, A4 => 
                           n24051, ZN => n24038);
   U21252 : NOR4_X1 port map( A1 => n24040, A2 => n24041, A3 => n24042, A4 => 
                           n24043, ZN => n24039);
   U21253 : OAI221_X1 port map( B1 => n21178, B2 => n26500, C1 => n21170, C2 =>
                           n26494, A => n24054, ZN => n24049);
   U21254 : NAND2_X1 port map( A1 => n24020, A2 => n24021, ZN => n5887);
   U21255 : NOR4_X1 port map( A1 => n24030, A2 => n24031, A3 => n24032, A4 => 
                           n24033, ZN => n24020);
   U21256 : NOR4_X1 port map( A1 => n24022, A2 => n24023, A3 => n24024, A4 => 
                           n24025, ZN => n24021);
   U21257 : OAI221_X1 port map( B1 => n21177, B2 => n26500, C1 => n21169, C2 =>
                           n26494, A => n24036, ZN => n24031);
   U21258 : NAND2_X1 port map( A1 => n22857, A2 => n22858, ZN => n6011);
   U21259 : NOR4_X1 port map( A1 => n22867, A2 => n22868, A3 => n22869, A4 => 
                           n22870, ZN => n22857);
   U21260 : NOR4_X1 port map( A1 => n22859, A2 => n22860, A3 => n22861, A4 => 
                           n22862, ZN => n22858);
   U21261 : OAI221_X1 port map( B1 => n21179, B2 => n26725, C1 => n21171, C2 =>
                           n26719, A => n22873, ZN => n22868);
   U21262 : NAND2_X1 port map( A1 => n22839, A2 => n22840, ZN => n6013);
   U21263 : NOR4_X1 port map( A1 => n22849, A2 => n22850, A3 => n22851, A4 => 
                           n22852, ZN => n22839);
   U21264 : NOR4_X1 port map( A1 => n22841, A2 => n22842, A3 => n22843, A4 => 
                           n22844, ZN => n22840);
   U21265 : OAI221_X1 port map( B1 => n21178, B2 => n26725, C1 => n21170, C2 =>
                           n26719, A => n22855, ZN => n22850);
   U21266 : NAND2_X1 port map( A1 => n22821, A2 => n22822, ZN => n6015);
   U21267 : NOR4_X1 port map( A1 => n22831, A2 => n22832, A3 => n22833, A4 => 
                           n22834, ZN => n22821);
   U21268 : NOR4_X1 port map( A1 => n22823, A2 => n22824, A3 => n22825, A4 => 
                           n22826, ZN => n22822);
   U21269 : OAI221_X1 port map( B1 => n21177, B2 => n26725, C1 => n21169, C2 =>
                           n26719, A => n22837, ZN => n22832);
   U21270 : NAND2_X1 port map( A1 => n22769, A2 => n22770, ZN => n6017);
   U21271 : NOR4_X1 port map( A1 => n22796, A2 => n22797, A3 => n22798, A4 => 
                           n22799, ZN => n22769);
   U21272 : NOR4_X1 port map( A1 => n22771, A2 => n22772, A3 => n22773, A4 => 
                           n22774, ZN => n22770);
   U21273 : OAI221_X1 port map( B1 => n21176, B2 => n26725, C1 => n21168, C2 =>
                           n26719, A => n22812, ZN => n22797);
   U21274 : NAND2_X1 port map( A1 => n24272, A2 => n24273, ZN => n5859);
   U21275 : NOR4_X1 port map( A1 => n24282, A2 => n24283, A3 => n24284, A4 => 
                           n24285, ZN => n24272);
   U21276 : NOR4_X1 port map( A1 => n24274, A2 => n24275, A3 => n24276, A4 => 
                           n24277, ZN => n24273);
   U21277 : OAI221_X1 port map( B1 => n21531, B2 => n26499, C1 => n21371, C2 =>
                           n26493, A => n24288, ZN => n24283);
   U21278 : NAND2_X1 port map( A1 => n24254, A2 => n24255, ZN => n5861);
   U21279 : NOR4_X1 port map( A1 => n24264, A2 => n24265, A3 => n24266, A4 => 
                           n24267, ZN => n24254);
   U21280 : NOR4_X1 port map( A1 => n24256, A2 => n24257, A3 => n24258, A4 => 
                           n24259, ZN => n24255);
   U21281 : OAI221_X1 port map( B1 => n21530, B2 => n26499, C1 => n21370, C2 =>
                           n26493, A => n24270, ZN => n24265);
   U21282 : NAND2_X1 port map( A1 => n24236, A2 => n24237, ZN => n5863);
   U21283 : NOR4_X1 port map( A1 => n24246, A2 => n24247, A3 => n24248, A4 => 
                           n24249, ZN => n24236);
   U21284 : NOR4_X1 port map( A1 => n24238, A2 => n24239, A3 => n24240, A4 => 
                           n24241, ZN => n24237);
   U21285 : OAI221_X1 port map( B1 => n21529, B2 => n26499, C1 => n21369, C2 =>
                           n26493, A => n24252, ZN => n24247);
   U21286 : NAND2_X1 port map( A1 => n24218, A2 => n24219, ZN => n5865);
   U21287 : NOR4_X1 port map( A1 => n24228, A2 => n24229, A3 => n24230, A4 => 
                           n24231, ZN => n24218);
   U21288 : NOR4_X1 port map( A1 => n24220, A2 => n24221, A3 => n24222, A4 => 
                           n24223, ZN => n24219);
   U21289 : OAI221_X1 port map( B1 => n21528, B2 => n26499, C1 => n21368, C2 =>
                           n26493, A => n24234, ZN => n24229);
   U21290 : NAND2_X1 port map( A1 => n24200, A2 => n24201, ZN => n5867);
   U21291 : NOR4_X1 port map( A1 => n24210, A2 => n24211, A3 => n24212, A4 => 
                           n24213, ZN => n24200);
   U21292 : NOR4_X1 port map( A1 => n24202, A2 => n24203, A3 => n24204, A4 => 
                           n24205, ZN => n24201);
   U21293 : OAI221_X1 port map( B1 => n21527, B2 => n26499, C1 => n21367, C2 =>
                           n26493, A => n24216, ZN => n24211);
   U21294 : NAND2_X1 port map( A1 => n24182, A2 => n24183, ZN => n5869);
   U21295 : NOR4_X1 port map( A1 => n24192, A2 => n24193, A3 => n24194, A4 => 
                           n24195, ZN => n24182);
   U21296 : NOR4_X1 port map( A1 => n24184, A2 => n24185, A3 => n24186, A4 => 
                           n24187, ZN => n24183);
   U21297 : OAI221_X1 port map( B1 => n21526, B2 => n26499, C1 => n21366, C2 =>
                           n26493, A => n24198, ZN => n24193);
   U21298 : NAND2_X1 port map( A1 => n24164, A2 => n24165, ZN => n5871);
   U21299 : NOR4_X1 port map( A1 => n24174, A2 => n24175, A3 => n24176, A4 => 
                           n24177, ZN => n24164);
   U21300 : NOR4_X1 port map( A1 => n24166, A2 => n24167, A3 => n24168, A4 => 
                           n24169, ZN => n24165);
   U21301 : OAI221_X1 port map( B1 => n21525, B2 => n26499, C1 => n21365, C2 =>
                           n26493, A => n24180, ZN => n24175);
   U21302 : NAND2_X1 port map( A1 => n24146, A2 => n24147, ZN => n5873);
   U21303 : NOR4_X1 port map( A1 => n24156, A2 => n24157, A3 => n24158, A4 => 
                           n24159, ZN => n24146);
   U21304 : NOR4_X1 port map( A1 => n24148, A2 => n24149, A3 => n24150, A4 => 
                           n24151, ZN => n24147);
   U21305 : OAI221_X1 port map( B1 => n21524, B2 => n26499, C1 => n21364, C2 =>
                           n26493, A => n24162, ZN => n24157);
   U21306 : NAND2_X1 port map( A1 => n24128, A2 => n24129, ZN => n5875);
   U21307 : NOR4_X1 port map( A1 => n24138, A2 => n24139, A3 => n24140, A4 => 
                           n24141, ZN => n24128);
   U21308 : NOR4_X1 port map( A1 => n24130, A2 => n24131, A3 => n24132, A4 => 
                           n24133, ZN => n24129);
   U21309 : OAI221_X1 port map( B1 => n21523, B2 => n26499, C1 => n21363, C2 =>
                           n26493, A => n24144, ZN => n24139);
   U21310 : NAND2_X1 port map( A1 => n24110, A2 => n24111, ZN => n5877);
   U21311 : NOR4_X1 port map( A1 => n24120, A2 => n24121, A3 => n24122, A4 => 
                           n24123, ZN => n24110);
   U21312 : NOR4_X1 port map( A1 => n24112, A2 => n24113, A3 => n24114, A4 => 
                           n24115, ZN => n24111);
   U21313 : OAI221_X1 port map( B1 => n21522, B2 => n26499, C1 => n21362, C2 =>
                           n26493, A => n24126, ZN => n24121);
   U21314 : NAND2_X1 port map( A1 => n24092, A2 => n24093, ZN => n5879);
   U21315 : NOR4_X1 port map( A1 => n24102, A2 => n24103, A3 => n24104, A4 => 
                           n24105, ZN => n24092);
   U21316 : NOR4_X1 port map( A1 => n24094, A2 => n24095, A3 => n24096, A4 => 
                           n24097, ZN => n24093);
   U21317 : OAI221_X1 port map( B1 => n21521, B2 => n26499, C1 => n21361, C2 =>
                           n26493, A => n24108, ZN => n24103);
   U21318 : NAND2_X1 port map( A1 => n24074, A2 => n24075, ZN => n5881);
   U21319 : NOR4_X1 port map( A1 => n24084, A2 => n24085, A3 => n24086, A4 => 
                           n24087, ZN => n24074);
   U21320 : NOR4_X1 port map( A1 => n24076, A2 => n24077, A3 => n24078, A4 => 
                           n24079, ZN => n24075);
   U21321 : OAI221_X1 port map( B1 => n21520, B2 => n26499, C1 => n21360, C2 =>
                           n26493, A => n24090, ZN => n24085);
   U21322 : NAND2_X1 port map( A1 => n23073, A2 => n23074, ZN => n5987);
   U21323 : NOR4_X1 port map( A1 => n23083, A2 => n23084, A3 => n23085, A4 => 
                           n23086, ZN => n23073);
   U21324 : NOR4_X1 port map( A1 => n23075, A2 => n23076, A3 => n23077, A4 => 
                           n23078, ZN => n23074);
   U21325 : OAI221_X1 port map( B1 => n21531, B2 => n26724, C1 => n21371, C2 =>
                           n26718, A => n23089, ZN => n23084);
   U21326 : NAND2_X1 port map( A1 => n23055, A2 => n23056, ZN => n5989);
   U21327 : NOR4_X1 port map( A1 => n23065, A2 => n23066, A3 => n23067, A4 => 
                           n23068, ZN => n23055);
   U21328 : NOR4_X1 port map( A1 => n23057, A2 => n23058, A3 => n23059, A4 => 
                           n23060, ZN => n23056);
   U21329 : OAI221_X1 port map( B1 => n21530, B2 => n26724, C1 => n21370, C2 =>
                           n26718, A => n23071, ZN => n23066);
   U21330 : NAND2_X1 port map( A1 => n23037, A2 => n23038, ZN => n5991);
   U21331 : NOR4_X1 port map( A1 => n23047, A2 => n23048, A3 => n23049, A4 => 
                           n23050, ZN => n23037);
   U21332 : NOR4_X1 port map( A1 => n23039, A2 => n23040, A3 => n23041, A4 => 
                           n23042, ZN => n23038);
   U21333 : OAI221_X1 port map( B1 => n21529, B2 => n26724, C1 => n21369, C2 =>
                           n26718, A => n23053, ZN => n23048);
   U21334 : NAND2_X1 port map( A1 => n23019, A2 => n23020, ZN => n5993);
   U21335 : NOR4_X1 port map( A1 => n23029, A2 => n23030, A3 => n23031, A4 => 
                           n23032, ZN => n23019);
   U21336 : NOR4_X1 port map( A1 => n23021, A2 => n23022, A3 => n23023, A4 => 
                           n23024, ZN => n23020);
   U21337 : OAI221_X1 port map( B1 => n21528, B2 => n26724, C1 => n21368, C2 =>
                           n26718, A => n23035, ZN => n23030);
   U21338 : NAND2_X1 port map( A1 => n23001, A2 => n23002, ZN => n5995);
   U21339 : NOR4_X1 port map( A1 => n23011, A2 => n23012, A3 => n23013, A4 => 
                           n23014, ZN => n23001);
   U21340 : NOR4_X1 port map( A1 => n23003, A2 => n23004, A3 => n23005, A4 => 
                           n23006, ZN => n23002);
   U21341 : OAI221_X1 port map( B1 => n21527, B2 => n26724, C1 => n21367, C2 =>
                           n26718, A => n23017, ZN => n23012);
   U21342 : NAND2_X1 port map( A1 => n22983, A2 => n22984, ZN => n5997);
   U21343 : NOR4_X1 port map( A1 => n22993, A2 => n22994, A3 => n22995, A4 => 
                           n22996, ZN => n22983);
   U21344 : NOR4_X1 port map( A1 => n22985, A2 => n22986, A3 => n22987, A4 => 
                           n22988, ZN => n22984);
   U21345 : OAI221_X1 port map( B1 => n21526, B2 => n26724, C1 => n21366, C2 =>
                           n26718, A => n22999, ZN => n22994);
   U21346 : NAND2_X1 port map( A1 => n22965, A2 => n22966, ZN => n5999);
   U21347 : NOR4_X1 port map( A1 => n22975, A2 => n22976, A3 => n22977, A4 => 
                           n22978, ZN => n22965);
   U21348 : NOR4_X1 port map( A1 => n22967, A2 => n22968, A3 => n22969, A4 => 
                           n22970, ZN => n22966);
   U21349 : OAI221_X1 port map( B1 => n21525, B2 => n26724, C1 => n21365, C2 =>
                           n26718, A => n22981, ZN => n22976);
   U21350 : NAND2_X1 port map( A1 => n22947, A2 => n22948, ZN => n6001);
   U21351 : NOR4_X1 port map( A1 => n22957, A2 => n22958, A3 => n22959, A4 => 
                           n22960, ZN => n22947);
   U21352 : NOR4_X1 port map( A1 => n22949, A2 => n22950, A3 => n22951, A4 => 
                           n22952, ZN => n22948);
   U21353 : OAI221_X1 port map( B1 => n21524, B2 => n26724, C1 => n21364, C2 =>
                           n26718, A => n22963, ZN => n22958);
   U21354 : NAND2_X1 port map( A1 => n22929, A2 => n22930, ZN => n6003);
   U21355 : NOR4_X1 port map( A1 => n22939, A2 => n22940, A3 => n22941, A4 => 
                           n22942, ZN => n22929);
   U21356 : NOR4_X1 port map( A1 => n22931, A2 => n22932, A3 => n22933, A4 => 
                           n22934, ZN => n22930);
   U21357 : OAI221_X1 port map( B1 => n21523, B2 => n26724, C1 => n21363, C2 =>
                           n26718, A => n22945, ZN => n22940);
   U21358 : NAND2_X1 port map( A1 => n22911, A2 => n22912, ZN => n6005);
   U21359 : NOR4_X1 port map( A1 => n22921, A2 => n22922, A3 => n22923, A4 => 
                           n22924, ZN => n22911);
   U21360 : NOR4_X1 port map( A1 => n22913, A2 => n22914, A3 => n22915, A4 => 
                           n22916, ZN => n22912);
   U21361 : OAI221_X1 port map( B1 => n21522, B2 => n26724, C1 => n21362, C2 =>
                           n26718, A => n22927, ZN => n22922);
   U21362 : NAND2_X1 port map( A1 => n22893, A2 => n22894, ZN => n6007);
   U21363 : NOR4_X1 port map( A1 => n22903, A2 => n22904, A3 => n22905, A4 => 
                           n22906, ZN => n22893);
   U21364 : NOR4_X1 port map( A1 => n22895, A2 => n22896, A3 => n22897, A4 => 
                           n22898, ZN => n22894);
   U21365 : OAI221_X1 port map( B1 => n21521, B2 => n26724, C1 => n21361, C2 =>
                           n26718, A => n22909, ZN => n22904);
   U21366 : NAND2_X1 port map( A1 => n22875, A2 => n22876, ZN => n6009);
   U21367 : NOR4_X1 port map( A1 => n22885, A2 => n22886, A3 => n22887, A4 => 
                           n22888, ZN => n22875);
   U21368 : NOR4_X1 port map( A1 => n22877, A2 => n22878, A3 => n22879, A4 => 
                           n22880, ZN => n22876);
   U21369 : OAI221_X1 port map( B1 => n21520, B2 => n26724, C1 => n21360, C2 =>
                           n26718, A => n22891, ZN => n22886);
   U21370 : BUF_X1 port map( A => n24010, Z => n26489);
   U21371 : BUF_X1 port map( A => n24010, Z => n26490);
   U21372 : BUF_X1 port map( A => n24010, Z => n26491);
   U21373 : BUF_X1 port map( A => n24010, Z => n26492);
   U21374 : BUF_X1 port map( A => n22811, Z => n26714);
   U21375 : BUF_X1 port map( A => n22811, Z => n26715);
   U21376 : BUF_X1 port map( A => n22811, Z => n26716);
   U21377 : BUF_X1 port map( A => n22811, Z => n26717);
   U21378 : INV_X1 port map( A => n27487, ZN => n27477);
   U21379 : INV_X1 port map( A => n27487, ZN => n27478);
   U21380 : INV_X1 port map( A => n27487, ZN => n27479);
   U21381 : INV_X1 port map( A => n27487, ZN => n27480);
   U21382 : INV_X1 port map( A => n27487, ZN => n27481);
   U21383 : INV_X1 port map( A => n27487, ZN => n27483);
   U21384 : INV_X1 port map( A => n27487, ZN => n27482);
   U21385 : INV_X1 port map( A => n27487, ZN => n27485);
   U21386 : INV_X1 port map( A => n27487, ZN => n27486);
   U21387 : INV_X1 port map( A => n27487, ZN => n27484);
   U21388 : BUF_X1 port map( A => n24014, Z => n26471);
   U21389 : BUF_X1 port map( A => n24009, Z => n26495);
   U21390 : BUF_X1 port map( A => n24014, Z => n26472);
   U21391 : BUF_X1 port map( A => n24009, Z => n26496);
   U21392 : BUF_X1 port map( A => n24014, Z => n26473);
   U21393 : BUF_X1 port map( A => n24009, Z => n26497);
   U21394 : BUF_X1 port map( A => n24014, Z => n26474);
   U21395 : BUF_X1 port map( A => n24009, Z => n26498);
   U21396 : BUF_X1 port map( A => n22815, Z => n26696);
   U21397 : BUF_X1 port map( A => n22810, Z => n26720);
   U21398 : BUF_X1 port map( A => n22815, Z => n26697);
   U21399 : BUF_X1 port map( A => n22810, Z => n26721);
   U21400 : BUF_X1 port map( A => n22815, Z => n26698);
   U21401 : BUF_X1 port map( A => n22810, Z => n26722);
   U21402 : BUF_X1 port map( A => n22815, Z => n26699);
   U21403 : BUF_X1 port map( A => n22810, Z => n26723);
   U21404 : NOR3_X1 port map( A1 => n20640, A2 => n20643, A3 => n20639, ZN => 
                           n25143);
   U21405 : NOR3_X1 port map( A1 => n20635, A2 => n20638, A3 => n20634, ZN => 
                           n23944);
   U21406 : AND3_X1 port map( A1 => n20631, A2 => n20630, A3 => n22717, ZN => 
                           n22695);
   U21407 : NAND2_X1 port map( A1 => n22704, A2 => n22695, ZN => n22702);
   U21408 : NAND2_X1 port map( A1 => n22698, A2 => n22695, ZN => n22696);
   U21409 : NAND2_X1 port map( A1 => n22701, A2 => n22695, ZN => n22699);
   U21410 : AND3_X1 port map( A1 => n20642, A2 => n20641, A3 => n25164, ZN => 
                           n25151);
   U21411 : AND3_X1 port map( A1 => n20637, A2 => n20636, A3 => n23965, ZN => 
                           n23952);
   U21412 : BUF_X1 port map( A => n20707, Z => n27282);
   U21413 : BUF_X1 port map( A => n20706, Z => n27285);
   U21414 : BUF_X1 port map( A => n20705, Z => n27288);
   U21415 : BUF_X1 port map( A => n20704, Z => n27291);
   U21416 : BUF_X1 port map( A => n20703, Z => n27294);
   U21417 : BUF_X1 port map( A => n20702, Z => n27297);
   U21418 : BUF_X1 port map( A => n20701, Z => n27300);
   U21419 : BUF_X1 port map( A => n20700, Z => n27303);
   U21420 : BUF_X1 port map( A => n20699, Z => n27306);
   U21421 : BUF_X1 port map( A => n20698, Z => n27309);
   U21422 : BUF_X1 port map( A => n20697, Z => n27312);
   U21423 : BUF_X1 port map( A => n20696, Z => n27315);
   U21424 : BUF_X1 port map( A => n20695, Z => n27318);
   U21425 : BUF_X1 port map( A => n20694, Z => n27321);
   U21426 : BUF_X1 port map( A => n20693, Z => n27324);
   U21427 : BUF_X1 port map( A => n20692, Z => n27327);
   U21428 : BUF_X1 port map( A => n20691, Z => n27330);
   U21429 : BUF_X1 port map( A => n20690, Z => n27333);
   U21430 : BUF_X1 port map( A => n20689, Z => n27336);
   U21431 : BUF_X1 port map( A => n20688, Z => n27339);
   U21432 : BUF_X1 port map( A => n20687, Z => n27342);
   U21433 : BUF_X1 port map( A => n20686, Z => n27345);
   U21434 : BUF_X1 port map( A => n20685, Z => n27348);
   U21435 : BUF_X1 port map( A => n20684, Z => n27351);
   U21436 : BUF_X1 port map( A => n20683, Z => n27354);
   U21437 : BUF_X1 port map( A => n20682, Z => n27357);
   U21438 : BUF_X1 port map( A => n20681, Z => n27360);
   U21439 : BUF_X1 port map( A => n20680, Z => n27363);
   U21440 : BUF_X1 port map( A => n20679, Z => n27366);
   U21441 : BUF_X1 port map( A => n20678, Z => n27369);
   U21442 : BUF_X1 port map( A => n20677, Z => n27372);
   U21443 : BUF_X1 port map( A => n20676, Z => n27375);
   U21444 : BUF_X1 port map( A => n20675, Z => n27378);
   U21445 : BUF_X1 port map( A => n20674, Z => n27381);
   U21446 : BUF_X1 port map( A => n20673, Z => n27384);
   U21447 : BUF_X1 port map( A => n20672, Z => n27387);
   U21448 : BUF_X1 port map( A => n20671, Z => n27390);
   U21449 : BUF_X1 port map( A => n20670, Z => n27393);
   U21450 : BUF_X1 port map( A => n20669, Z => n27396);
   U21451 : BUF_X1 port map( A => n20668, Z => n27399);
   U21452 : BUF_X1 port map( A => n20667, Z => n27402);
   U21453 : BUF_X1 port map( A => n20666, Z => n27405);
   U21454 : BUF_X1 port map( A => n20665, Z => n27408);
   U21455 : BUF_X1 port map( A => n20664, Z => n27411);
   U21456 : BUF_X1 port map( A => n20663, Z => n27414);
   U21457 : BUF_X1 port map( A => n20662, Z => n27417);
   U21458 : BUF_X1 port map( A => n20661, Z => n27420);
   U21459 : BUF_X1 port map( A => n20660, Z => n27423);
   U21460 : BUF_X1 port map( A => n20659, Z => n27426);
   U21461 : BUF_X1 port map( A => n20658, Z => n27429);
   U21462 : BUF_X1 port map( A => n20657, Z => n27432);
   U21463 : BUF_X1 port map( A => n20656, Z => n27435);
   U21464 : BUF_X1 port map( A => n20655, Z => n27438);
   U21465 : BUF_X1 port map( A => n20654, Z => n27441);
   U21466 : BUF_X1 port map( A => n20653, Z => n27444);
   U21467 : BUF_X1 port map( A => n20652, Z => n27447);
   U21468 : BUF_X1 port map( A => n20651, Z => n27450);
   U21469 : BUF_X1 port map( A => n20650, Z => n27453);
   U21470 : BUF_X1 port map( A => n20649, Z => n27456);
   U21471 : BUF_X1 port map( A => n20648, Z => n27459);
   U21472 : BUF_X1 port map( A => n20647, Z => n27462);
   U21473 : BUF_X1 port map( A => n20646, Z => n27465);
   U21474 : BUF_X1 port map( A => n20645, Z => n27468);
   U21475 : BUF_X1 port map( A => n20644, Z => n27471);
   U21476 : BUF_X1 port map( A => n20644, Z => n27472);
   U21477 : BUF_X1 port map( A => n20707, Z => n27283);
   U21478 : BUF_X1 port map( A => n20706, Z => n27286);
   U21479 : BUF_X1 port map( A => n20705, Z => n27289);
   U21480 : BUF_X1 port map( A => n20704, Z => n27292);
   U21481 : BUF_X1 port map( A => n20703, Z => n27295);
   U21482 : BUF_X1 port map( A => n20702, Z => n27298);
   U21483 : BUF_X1 port map( A => n20701, Z => n27301);
   U21484 : BUF_X1 port map( A => n20700, Z => n27304);
   U21485 : BUF_X1 port map( A => n20699, Z => n27307);
   U21486 : BUF_X1 port map( A => n20698, Z => n27310);
   U21487 : BUF_X1 port map( A => n20697, Z => n27313);
   U21488 : BUF_X1 port map( A => n20696, Z => n27316);
   U21489 : BUF_X1 port map( A => n20695, Z => n27319);
   U21490 : BUF_X1 port map( A => n20694, Z => n27322);
   U21491 : BUF_X1 port map( A => n20693, Z => n27325);
   U21492 : BUF_X1 port map( A => n20692, Z => n27328);
   U21493 : BUF_X1 port map( A => n20691, Z => n27331);
   U21494 : BUF_X1 port map( A => n20690, Z => n27334);
   U21495 : BUF_X1 port map( A => n20689, Z => n27337);
   U21496 : BUF_X1 port map( A => n20688, Z => n27340);
   U21497 : BUF_X1 port map( A => n20687, Z => n27343);
   U21498 : BUF_X1 port map( A => n20686, Z => n27346);
   U21499 : BUF_X1 port map( A => n20685, Z => n27349);
   U21500 : BUF_X1 port map( A => n20684, Z => n27352);
   U21501 : BUF_X1 port map( A => n20683, Z => n27355);
   U21502 : BUF_X1 port map( A => n20682, Z => n27358);
   U21503 : BUF_X1 port map( A => n20681, Z => n27361);
   U21504 : BUF_X1 port map( A => n20680, Z => n27364);
   U21505 : BUF_X1 port map( A => n20679, Z => n27367);
   U21506 : BUF_X1 port map( A => n20678, Z => n27370);
   U21507 : BUF_X1 port map( A => n20677, Z => n27373);
   U21508 : BUF_X1 port map( A => n20676, Z => n27376);
   U21509 : BUF_X1 port map( A => n20675, Z => n27379);
   U21510 : BUF_X1 port map( A => n20674, Z => n27382);
   U21511 : BUF_X1 port map( A => n20673, Z => n27385);
   U21512 : BUF_X1 port map( A => n20672, Z => n27388);
   U21513 : BUF_X1 port map( A => n20671, Z => n27391);
   U21514 : BUF_X1 port map( A => n20670, Z => n27394);
   U21515 : BUF_X1 port map( A => n20669, Z => n27397);
   U21516 : BUF_X1 port map( A => n20668, Z => n27400);
   U21517 : BUF_X1 port map( A => n20667, Z => n27403);
   U21518 : BUF_X1 port map( A => n20666, Z => n27406);
   U21519 : BUF_X1 port map( A => n20665, Z => n27409);
   U21520 : BUF_X1 port map( A => n20664, Z => n27412);
   U21521 : BUF_X1 port map( A => n20663, Z => n27415);
   U21522 : BUF_X1 port map( A => n20662, Z => n27418);
   U21523 : BUF_X1 port map( A => n20661, Z => n27421);
   U21524 : BUF_X1 port map( A => n20660, Z => n27424);
   U21525 : BUF_X1 port map( A => n20659, Z => n27427);
   U21526 : BUF_X1 port map( A => n20658, Z => n27430);
   U21527 : BUF_X1 port map( A => n20657, Z => n27433);
   U21528 : BUF_X1 port map( A => n20656, Z => n27436);
   U21529 : BUF_X1 port map( A => n20655, Z => n27439);
   U21530 : BUF_X1 port map( A => n20654, Z => n27442);
   U21531 : BUF_X1 port map( A => n20653, Z => n27445);
   U21532 : BUF_X1 port map( A => n20652, Z => n27448);
   U21533 : BUF_X1 port map( A => n20651, Z => n27451);
   U21534 : BUF_X1 port map( A => n20650, Z => n27454);
   U21535 : BUF_X1 port map( A => n20649, Z => n27457);
   U21536 : BUF_X1 port map( A => n20648, Z => n27460);
   U21537 : BUF_X1 port map( A => n20647, Z => n27463);
   U21538 : BUF_X1 port map( A => n20646, Z => n27466);
   U21539 : BUF_X1 port map( A => n20645, Z => n27469);
   U21540 : NAND2_X1 port map( A1 => n25153, A2 => n25148, ZN => n23985);
   U21541 : NAND2_X1 port map( A1 => n25153, A2 => n25151, ZN => n24005);
   U21542 : NAND2_X1 port map( A1 => n23954, A2 => n23949, ZN => n22786);
   U21543 : NAND2_X1 port map( A1 => n23954, A2 => n23952, ZN => n22806);
   U21544 : NAND2_X1 port map( A1 => n22716, A2 => n22695, ZN => n22714);
   U21545 : NAND2_X1 port map( A1 => n22707, A2 => n22695, ZN => n22705);
   U21546 : NAND2_X1 port map( A1 => n22713, A2 => n22695, ZN => n22711);
   U21547 : NAND2_X1 port map( A1 => n22710, A2 => n22695, ZN => n22708);
   U21548 : NAND2_X1 port map( A1 => n25144, A2 => n25147, ZN => n23990);
   U21549 : NAND2_X1 port map( A1 => n25144, A2 => n25155, ZN => n24000);
   U21550 : NAND2_X1 port map( A1 => n23945, A2 => n23948, ZN => n22791);
   U21551 : NAND2_X1 port map( A1 => n23945, A2 => n23956, ZN => n22801);
   U21552 : NAND2_X1 port map( A1 => n22720, A2 => n22698, ZN => n22721);
   U21553 : NAND2_X1 port map( A1 => n22754, A2 => n22704, ZN => n22759);
   U21554 : NAND2_X1 port map( A1 => n22754, A2 => n22694, ZN => n22752);
   U21555 : NAND2_X1 port map( A1 => n22720, A2 => n22694, ZN => n22718);
   U21556 : NAND2_X1 port map( A1 => n22720, A2 => n22701, ZN => n22723);
   U21557 : NAND2_X1 port map( A1 => n22737, A2 => n22704, ZN => n22742);
   U21558 : NAND2_X1 port map( A1 => n22754, A2 => n22710, ZN => n22763);
   U21559 : NAND2_X1 port map( A1 => n22754, A2 => n22707, ZN => n22761);
   U21560 : NAND2_X1 port map( A1 => n22720, A2 => n22704, ZN => n22725);
   U21561 : NAND2_X1 port map( A1 => n22737, A2 => n22713, ZN => n22748);
   U21562 : NAND2_X1 port map( A1 => n22737, A2 => n22698, ZN => n22738);
   U21563 : NAND2_X1 port map( A1 => n22737, A2 => n22701, ZN => n22740);
   U21564 : NAND2_X1 port map( A1 => n22754, A2 => n22701, ZN => n22757);
   U21565 : NAND2_X1 port map( A1 => n22737, A2 => n22716, ZN => n22750);
   U21566 : NAND2_X1 port map( A1 => n22737, A2 => n22694, ZN => n22735);
   U21567 : NAND2_X1 port map( A1 => n22754, A2 => n22698, ZN => n22755);
   U21568 : NAND2_X1 port map( A1 => n22720, A2 => n22710, ZN => n22729);
   U21569 : NAND2_X1 port map( A1 => n22720, A2 => n22716, ZN => n22733);
   U21570 : NAND2_X1 port map( A1 => n22737, A2 => n22707, ZN => n22744);
   U21571 : NAND2_X1 port map( A1 => n22737, A2 => n22710, ZN => n22746);
   U21572 : NAND2_X1 port map( A1 => n22754, A2 => n22716, ZN => n22767);
   U21573 : NAND2_X1 port map( A1 => n22754, A2 => n22713, ZN => n22765);
   U21574 : NAND2_X1 port map( A1 => n22720, A2 => n22713, ZN => n22731);
   U21575 : NAND2_X1 port map( A1 => n22720, A2 => n22707, ZN => n22727);
   U21576 : NAND2_X1 port map( A1 => n25146, A2 => n25144, ZN => n23975);
   U21577 : NAND2_X1 port map( A1 => n23947, A2 => n23945, ZN => n22776);
   U21578 : BUF_X1 port map( A => n24010, Z => n26493);
   U21579 : BUF_X1 port map( A => n22811, Z => n26718);
   U21580 : BUF_X1 port map( A => n24015, Z => n26465);
   U21581 : BUF_X1 port map( A => n24015, Z => n26466);
   U21582 : BUF_X1 port map( A => n24015, Z => n26467);
   U21583 : BUF_X1 port map( A => n24015, Z => n26468);
   U21584 : BUF_X1 port map( A => n24015, Z => n26469);
   U21585 : BUF_X1 port map( A => n22816, Z => n26690);
   U21586 : BUF_X1 port map( A => n22816, Z => n26691);
   U21587 : BUF_X1 port map( A => n22816, Z => n26692);
   U21588 : BUF_X1 port map( A => n22816, Z => n26693);
   U21589 : BUF_X1 port map( A => n22816, Z => n26694);
   U21590 : BUF_X1 port map( A => n24014, Z => n26475);
   U21591 : BUF_X1 port map( A => n24009, Z => n26499);
   U21592 : BUF_X1 port map( A => n22815, Z => n26700);
   U21593 : BUF_X1 port map( A => n22810, Z => n26724);
   U21594 : BUF_X1 port map( A => n20626, Z => n27474);
   U21595 : BUF_X1 port map( A => n20626, Z => n27475);
   U21596 : BUF_X1 port map( A => n20707, Z => n27284);
   U21597 : BUF_X1 port map( A => n20706, Z => n27287);
   U21598 : BUF_X1 port map( A => n20705, Z => n27290);
   U21599 : BUF_X1 port map( A => n20704, Z => n27293);
   U21600 : BUF_X1 port map( A => n20703, Z => n27296);
   U21601 : BUF_X1 port map( A => n20702, Z => n27299);
   U21602 : BUF_X1 port map( A => n20701, Z => n27302);
   U21603 : BUF_X1 port map( A => n20700, Z => n27305);
   U21604 : BUF_X1 port map( A => n20699, Z => n27308);
   U21605 : BUF_X1 port map( A => n20698, Z => n27311);
   U21606 : BUF_X1 port map( A => n20697, Z => n27314);
   U21607 : BUF_X1 port map( A => n20696, Z => n27317);
   U21608 : BUF_X1 port map( A => n20695, Z => n27320);
   U21609 : BUF_X1 port map( A => n20694, Z => n27323);
   U21610 : BUF_X1 port map( A => n20693, Z => n27326);
   U21611 : BUF_X1 port map( A => n20692, Z => n27329);
   U21612 : BUF_X1 port map( A => n20691, Z => n27332);
   U21613 : BUF_X1 port map( A => n20690, Z => n27335);
   U21614 : BUF_X1 port map( A => n20689, Z => n27338);
   U21615 : BUF_X1 port map( A => n20688, Z => n27341);
   U21616 : BUF_X1 port map( A => n20687, Z => n27344);
   U21617 : BUF_X1 port map( A => n20686, Z => n27347);
   U21618 : BUF_X1 port map( A => n20685, Z => n27350);
   U21619 : BUF_X1 port map( A => n20684, Z => n27353);
   U21620 : BUF_X1 port map( A => n20683, Z => n27356);
   U21621 : BUF_X1 port map( A => n20682, Z => n27359);
   U21622 : BUF_X1 port map( A => n20681, Z => n27362);
   U21623 : BUF_X1 port map( A => n20680, Z => n27365);
   U21624 : BUF_X1 port map( A => n20679, Z => n27368);
   U21625 : BUF_X1 port map( A => n20678, Z => n27371);
   U21626 : BUF_X1 port map( A => n20677, Z => n27374);
   U21627 : BUF_X1 port map( A => n20676, Z => n27377);
   U21628 : BUF_X1 port map( A => n20675, Z => n27380);
   U21629 : BUF_X1 port map( A => n20674, Z => n27383);
   U21630 : BUF_X1 port map( A => n20673, Z => n27386);
   U21631 : BUF_X1 port map( A => n20672, Z => n27389);
   U21632 : BUF_X1 port map( A => n20671, Z => n27392);
   U21633 : BUF_X1 port map( A => n20670, Z => n27395);
   U21634 : BUF_X1 port map( A => n20669, Z => n27398);
   U21635 : BUF_X1 port map( A => n20668, Z => n27401);
   U21636 : BUF_X1 port map( A => n20667, Z => n27404);
   U21637 : BUF_X1 port map( A => n20666, Z => n27407);
   U21638 : BUF_X1 port map( A => n20665, Z => n27410);
   U21639 : BUF_X1 port map( A => n20664, Z => n27413);
   U21640 : BUF_X1 port map( A => n20663, Z => n27416);
   U21641 : BUF_X1 port map( A => n20662, Z => n27419);
   U21642 : BUF_X1 port map( A => n20661, Z => n27422);
   U21643 : BUF_X1 port map( A => n20660, Z => n27425);
   U21644 : BUF_X1 port map( A => n20659, Z => n27428);
   U21645 : BUF_X1 port map( A => n20658, Z => n27431);
   U21646 : BUF_X1 port map( A => n20657, Z => n27434);
   U21647 : BUF_X1 port map( A => n20656, Z => n27437);
   U21648 : BUF_X1 port map( A => n20655, Z => n27440);
   U21649 : BUF_X1 port map( A => n20654, Z => n27443);
   U21650 : BUF_X1 port map( A => n20653, Z => n27446);
   U21651 : BUF_X1 port map( A => n20652, Z => n27449);
   U21652 : BUF_X1 port map( A => n20651, Z => n27452);
   U21653 : BUF_X1 port map( A => n20650, Z => n27455);
   U21654 : BUF_X1 port map( A => n20649, Z => n27458);
   U21655 : BUF_X1 port map( A => n20648, Z => n27461);
   U21656 : BUF_X1 port map( A => n20647, Z => n27464);
   U21657 : BUF_X1 port map( A => n20646, Z => n27467);
   U21658 : BUF_X1 port map( A => n20645, Z => n27470);
   U21659 : BUF_X1 port map( A => n20644, Z => n27473);
   U21660 : BUF_X1 port map( A => n20626, Z => n27476);
   U21661 : NAND2_X1 port map( A1 => n25147, A2 => n25151, ZN => n23989);
   U21662 : NAND2_X1 port map( A1 => n25147, A2 => n25148, ZN => n23974);
   U21663 : NAND2_X1 port map( A1 => n23948, A2 => n23952, ZN => n22790);
   U21664 : NAND2_X1 port map( A1 => n23948, A2 => n23949, ZN => n22775);
   U21665 : NAND2_X1 port map( A1 => n25153, A2 => n25145, ZN => n23999);
   U21666 : NAND2_X1 port map( A1 => n23954, A2 => n23946, ZN => n22800);
   U21667 : NAND2_X1 port map( A1 => n25146, A2 => n25151, ZN => n23979);
   U21668 : NAND2_X1 port map( A1 => n23947, A2 => n23952, ZN => n22780);
   U21669 : NAND2_X1 port map( A1 => n25150, A2 => n25145, ZN => n23984);
   U21670 : NAND2_X1 port map( A1 => n23951, A2 => n23946, ZN => n22785);
   U21671 : NAND2_X1 port map( A1 => n25151, A2 => n25155, ZN => n24004);
   U21672 : NAND2_X1 port map( A1 => n23952, A2 => n23956, ZN => n22805);
   U21673 : NAND2_X1 port map( A1 => n22694, A2 => n22695, ZN => n22692);
   U21674 : AND3_X1 port map( A1 => n20642, A2 => n20641, A3 => n25165, ZN => 
                           n24012);
   U21675 : AND3_X1 port map( A1 => n20637, A2 => n20636, A3 => n23966, ZN => 
                           n22813);
   U21676 : AND2_X1 port map( A1 => n25147, A2 => n25145, ZN => n23988);
   U21677 : AND2_X1 port map( A1 => n23948, A2 => n23946, ZN => n22789);
   U21678 : AND2_X1 port map( A1 => n25153, A2 => n25144, ZN => n24002);
   U21679 : AND2_X1 port map( A1 => n23954, A2 => n23945, ZN => n22803);
   U21680 : AND2_X1 port map( A1 => n25155, A2 => n25148, ZN => n23993);
   U21681 : AND2_X1 port map( A1 => n23956, A2 => n23949, ZN => n22794);
   U21682 : AND2_X1 port map( A1 => n25146, A2 => n25145, ZN => n23983);
   U21683 : AND2_X1 port map( A1 => n25146, A2 => n25148, ZN => n24008);
   U21684 : AND2_X1 port map( A1 => n23947, A2 => n23946, ZN => n22784);
   U21685 : AND2_X1 port map( A1 => n23947, A2 => n23949, ZN => n22809);
   U21686 : AND2_X1 port map( A1 => n25150, A2 => n25148, ZN => n23982);
   U21687 : AND2_X1 port map( A1 => n23951, A2 => n23949, ZN => n22783);
   U21688 : AND2_X1 port map( A1 => n25143, A2 => n25145, ZN => n23977);
   U21689 : AND2_X1 port map( A1 => n25143, A2 => n25144, ZN => n23978);
   U21690 : AND2_X1 port map( A1 => n25143, A2 => n25148, ZN => n24007);
   U21691 : AND2_X1 port map( A1 => n23944, A2 => n23946, ZN => n22778);
   U21692 : AND2_X1 port map( A1 => n23944, A2 => n23945, ZN => n22779);
   U21693 : AND2_X1 port map( A1 => n23944, A2 => n23949, ZN => n22808);
   U21694 : AND2_X1 port map( A1 => n25145, A2 => n25155, ZN => n23994);
   U21695 : AND2_X1 port map( A1 => n23946, A2 => n23956, ZN => n22795);
   U21696 : AND2_X1 port map( A1 => n25163, A2 => n25148, ZN => n24017);
   U21697 : AND2_X1 port map( A1 => n25163, A2 => n25145, ZN => n24018);
   U21698 : AND2_X1 port map( A1 => n25163, A2 => n25151, ZN => n24019);
   U21699 : AND2_X1 port map( A1 => n25163, A2 => n25144, ZN => n24013);
   U21700 : AND2_X1 port map( A1 => n23964, A2 => n23949, ZN => n22818);
   U21701 : AND2_X1 port map( A1 => n23964, A2 => n23946, ZN => n22819);
   U21702 : AND2_X1 port map( A1 => n23964, A2 => n23952, ZN => n22820);
   U21703 : AND2_X1 port map( A1 => n23964, A2 => n23945, ZN => n22814);
   U21704 : AND2_X1 port map( A1 => n25151, A2 => n25150, ZN => n23992);
   U21705 : AND2_X1 port map( A1 => n25144, A2 => n25150, ZN => n23987);
   U21706 : AND2_X1 port map( A1 => n23952, A2 => n23951, ZN => n22793);
   U21707 : AND2_X1 port map( A1 => n23945, A2 => n23951, ZN => n22788);
   U21708 : BUF_X1 port map( A => n24003, Z => n26531);
   U21709 : BUF_X1 port map( A => n24003, Z => n26532);
   U21710 : BUF_X1 port map( A => n22804, Z => n26756);
   U21711 : BUF_X1 port map( A => n22804, Z => n26757);
   U21712 : OAI221_X1 port map( B1 => n21347, B2 => n26667, C1 => n21627, C2 =>
                           n26661, A => n24926, ZN => n24925);
   U21713 : AOI22_X1 port map( A1 => n26655, A2 => n9402, B1 => n26649, B2 => 
                           n19234, ZN => n24926);
   U21714 : OAI221_X1 port map( B1 => n20759, B2 => n26565, C1 => n21987, C2 =>
                           n26559, A => n24934, ZN => n24933);
   U21715 : AOI22_X1 port map( A1 => n26553, A2 => n19249, B1 => n26549, B2 => 
                           n4328, ZN => n24934);
   U21716 : OAI221_X1 port map( B1 => n21346, B2 => n26667, C1 => n21626, C2 =>
                           n26661, A => n24908, ZN => n24907);
   U21717 : AOI22_X1 port map( A1 => n26655, A2 => n9399, B1 => n26649, B2 => 
                           n19217, ZN => n24908);
   U21718 : OAI221_X1 port map( B1 => n20758, B2 => n26565, C1 => n21986, C2 =>
                           n26559, A => n24916, ZN => n24915);
   U21719 : AOI22_X1 port map( A1 => n26553, A2 => n19232, B1 => n26548, B2 => 
                           n4326, ZN => n24916);
   U21720 : OAI221_X1 port map( B1 => n21345, B2 => n26667, C1 => n21625, C2 =>
                           n26661, A => n24890, ZN => n24889);
   U21721 : AOI22_X1 port map( A1 => n26655, A2 => n9396, B1 => n26649, B2 => 
                           n19200, ZN => n24890);
   U21722 : OAI221_X1 port map( B1 => n20757, B2 => n26565, C1 => n21985, C2 =>
                           n26559, A => n24898, ZN => n24897);
   U21723 : AOI22_X1 port map( A1 => n26553, A2 => n19215, B1 => n26548, B2 => 
                           n4324, ZN => n24898);
   U21724 : OAI221_X1 port map( B1 => n21344, B2 => n26667, C1 => n21624, C2 =>
                           n26661, A => n24872, ZN => n24871);
   U21725 : AOI22_X1 port map( A1 => n26655, A2 => n9393, B1 => n26649, B2 => 
                           n19183, ZN => n24872);
   U21726 : OAI221_X1 port map( B1 => n20756, B2 => n26565, C1 => n21984, C2 =>
                           n26559, A => n24880, ZN => n24879);
   U21727 : AOI22_X1 port map( A1 => n26553, A2 => n19198, B1 => n26548, B2 => 
                           n4322, ZN => n24880);
   U21728 : OAI221_X1 port map( B1 => n21343, B2 => n26667, C1 => n21623, C2 =>
                           n26661, A => n24854, ZN => n24853);
   U21729 : AOI22_X1 port map( A1 => n26655, A2 => n9390, B1 => n26649, B2 => 
                           n19166, ZN => n24854);
   U21730 : OAI221_X1 port map( B1 => n20755, B2 => n26565, C1 => n21983, C2 =>
                           n26559, A => n24862, ZN => n24861);
   U21731 : AOI22_X1 port map( A1 => n26553, A2 => n19181, B1 => n26548, B2 => 
                           n4320, ZN => n24862);
   U21732 : OAI221_X1 port map( B1 => n21342, B2 => n26667, C1 => n21622, C2 =>
                           n26661, A => n24836, ZN => n24835);
   U21733 : AOI22_X1 port map( A1 => n26655, A2 => n9387, B1 => n26649, B2 => 
                           n19149, ZN => n24836);
   U21734 : OAI221_X1 port map( B1 => n20754, B2 => n26565, C1 => n21982, C2 =>
                           n26559, A => n24844, ZN => n24843);
   U21735 : AOI22_X1 port map( A1 => n26553, A2 => n19164, B1 => n26547, B2 => 
                           n4318, ZN => n24844);
   U21736 : OAI221_X1 port map( B1 => n21341, B2 => n26667, C1 => n21621, C2 =>
                           n26661, A => n24818, ZN => n24817);
   U21737 : AOI22_X1 port map( A1 => n26655, A2 => n9384, B1 => n26649, B2 => 
                           n19132, ZN => n24818);
   U21738 : OAI221_X1 port map( B1 => n20753, B2 => n26565, C1 => n21981, C2 =>
                           n26559, A => n24826, ZN => n24825);
   U21739 : AOI22_X1 port map( A1 => n26553, A2 => n19147, B1 => n26547, B2 => 
                           n4316, ZN => n24826);
   U21740 : OAI221_X1 port map( B1 => n21340, B2 => n26667, C1 => n21620, C2 =>
                           n26661, A => n24800, ZN => n24799);
   U21741 : AOI22_X1 port map( A1 => n26655, A2 => n9381, B1 => n26649, B2 => 
                           n19115, ZN => n24800);
   U21742 : OAI221_X1 port map( B1 => n20752, B2 => n26565, C1 => n21980, C2 =>
                           n26559, A => n24808, ZN => n24807);
   U21743 : AOI22_X1 port map( A1 => n26553, A2 => n19130, B1 => n26547, B2 => 
                           n4314, ZN => n24808);
   U21744 : OAI221_X1 port map( B1 => n21339, B2 => n26667, C1 => n21619, C2 =>
                           n26661, A => n24782, ZN => n24781);
   U21745 : AOI22_X1 port map( A1 => n26655, A2 => n9378, B1 => n26649, B2 => 
                           n19098, ZN => n24782);
   U21746 : OAI221_X1 port map( B1 => n20751, B2 => n26565, C1 => n21979, C2 =>
                           n26559, A => n24790, ZN => n24789);
   U21747 : AOI22_X1 port map( A1 => n26553, A2 => n19113, B1 => n26547, B2 => 
                           n4312, ZN => n24790);
   U21748 : OAI221_X1 port map( B1 => n21338, B2 => n26667, C1 => n21618, C2 =>
                           n26661, A => n24764, ZN => n24763);
   U21749 : AOI22_X1 port map( A1 => n26655, A2 => n9375, B1 => n26649, B2 => 
                           n19081, ZN => n24764);
   U21750 : OAI221_X1 port map( B1 => n20750, B2 => n26565, C1 => n21978, C2 =>
                           n26559, A => n24772, ZN => n24771);
   U21751 : AOI22_X1 port map( A1 => n26553, A2 => n19096, B1 => n26546, B2 => 
                           n4310, ZN => n24772);
   U21752 : OAI221_X1 port map( B1 => n21337, B2 => n26667, C1 => n21617, C2 =>
                           n26661, A => n24746, ZN => n24745);
   U21753 : AOI22_X1 port map( A1 => n26655, A2 => n9372, B1 => n26649, B2 => 
                           n19064, ZN => n24746);
   U21754 : OAI221_X1 port map( B1 => n20749, B2 => n26565, C1 => n21977, C2 =>
                           n26559, A => n24754, ZN => n24753);
   U21755 : AOI22_X1 port map( A1 => n26553, A2 => n19079, B1 => n26546, B2 => 
                           n4308, ZN => n24754);
   U21756 : OAI221_X1 port map( B1 => n21336, B2 => n26667, C1 => n21616, C2 =>
                           n26661, A => n24728, ZN => n24727);
   U21757 : AOI22_X1 port map( A1 => n26655, A2 => n9369, B1 => n26649, B2 => 
                           n19047, ZN => n24728);
   U21758 : OAI221_X1 port map( B1 => n20748, B2 => n26565, C1 => n21976, C2 =>
                           n26559, A => n24736, ZN => n24735);
   U21759 : AOI22_X1 port map( A1 => n26553, A2 => n19062, B1 => n26546, B2 => 
                           n4306, ZN => n24736);
   U21760 : OAI221_X1 port map( B1 => n21335, B2 => n26668, C1 => n21615, C2 =>
                           n26662, A => n24710, ZN => n24709);
   U21761 : AOI22_X1 port map( A1 => n26656, A2 => n9366, B1 => n26650, B2 => 
                           n19030, ZN => n24710);
   U21762 : OAI221_X1 port map( B1 => n20747, B2 => n26566, C1 => n21975, C2 =>
                           n26560, A => n24718, ZN => n24717);
   U21763 : AOI22_X1 port map( A1 => n26554, A2 => n19045, B1 => n26546, B2 => 
                           n4304, ZN => n24718);
   U21764 : OAI221_X1 port map( B1 => n21334, B2 => n26668, C1 => n21614, C2 =>
                           n26662, A => n24692, ZN => n24691);
   U21765 : AOI22_X1 port map( A1 => n26656, A2 => n9363, B1 => n26650, B2 => 
                           n19013, ZN => n24692);
   U21766 : OAI221_X1 port map( B1 => n20746, B2 => n26566, C1 => n21974, C2 =>
                           n26560, A => n24700, ZN => n24699);
   U21767 : AOI22_X1 port map( A1 => n26554, A2 => n19028, B1 => n26545, B2 => 
                           n4302, ZN => n24700);
   U21768 : OAI221_X1 port map( B1 => n21333, B2 => n26668, C1 => n21613, C2 =>
                           n26662, A => n24674, ZN => n24673);
   U21769 : AOI22_X1 port map( A1 => n26656, A2 => n9360, B1 => n26650, B2 => 
                           n18996, ZN => n24674);
   U21770 : OAI221_X1 port map( B1 => n20745, B2 => n26566, C1 => n21973, C2 =>
                           n26560, A => n24682, ZN => n24681);
   U21771 : AOI22_X1 port map( A1 => n26554, A2 => n19011, B1 => n26545, B2 => 
                           n4300, ZN => n24682);
   U21772 : OAI221_X1 port map( B1 => n21332, B2 => n26668, C1 => n21612, C2 =>
                           n26662, A => n24656, ZN => n24655);
   U21773 : AOI22_X1 port map( A1 => n26656, A2 => n9357, B1 => n26650, B2 => 
                           n18979, ZN => n24656);
   U21774 : OAI221_X1 port map( B1 => n20744, B2 => n26566, C1 => n21972, C2 =>
                           n26560, A => n24664, ZN => n24663);
   U21775 : AOI22_X1 port map( A1 => n26554, A2 => n18994, B1 => n26545, B2 => 
                           n4298, ZN => n24664);
   U21776 : OAI221_X1 port map( B1 => n21331, B2 => n26668, C1 => n21611, C2 =>
                           n26662, A => n24638, ZN => n24637);
   U21777 : AOI22_X1 port map( A1 => n26656, A2 => n9354, B1 => n26650, B2 => 
                           n18962, ZN => n24638);
   U21778 : OAI221_X1 port map( B1 => n20743, B2 => n26566, C1 => n21971, C2 =>
                           n26560, A => n24646, ZN => n24645);
   U21779 : AOI22_X1 port map( A1 => n26554, A2 => n18977, B1 => n26545, B2 => 
                           n4296, ZN => n24646);
   U21780 : OAI221_X1 port map( B1 => n21330, B2 => n26668, C1 => n21610, C2 =>
                           n26662, A => n24620, ZN => n24619);
   U21781 : AOI22_X1 port map( A1 => n26656, A2 => n9351, B1 => n26650, B2 => 
                           n18945, ZN => n24620);
   U21782 : OAI221_X1 port map( B1 => n20742, B2 => n26566, C1 => n21970, C2 =>
                           n26560, A => n24628, ZN => n24627);
   U21783 : AOI22_X1 port map( A1 => n26554, A2 => n18960, B1 => n26544, B2 => 
                           n4294, ZN => n24628);
   U21784 : OAI221_X1 port map( B1 => n21329, B2 => n26668, C1 => n21609, C2 =>
                           n26662, A => n24602, ZN => n24601);
   U21785 : AOI22_X1 port map( A1 => n26656, A2 => n9348, B1 => n26650, B2 => 
                           n18928, ZN => n24602);
   U21786 : OAI221_X1 port map( B1 => n20741, B2 => n26566, C1 => n21969, C2 =>
                           n26560, A => n24610, ZN => n24609);
   U21787 : AOI22_X1 port map( A1 => n26554, A2 => n18943, B1 => n26544, B2 => 
                           n4292, ZN => n24610);
   U21788 : OAI221_X1 port map( B1 => n21328, B2 => n26668, C1 => n21608, C2 =>
                           n26662, A => n24584, ZN => n24583);
   U21789 : AOI22_X1 port map( A1 => n26656, A2 => n9345, B1 => n26650, B2 => 
                           n18911, ZN => n24584);
   U21790 : OAI221_X1 port map( B1 => n20740, B2 => n26566, C1 => n21968, C2 =>
                           n26560, A => n24592, ZN => n24591);
   U21791 : AOI22_X1 port map( A1 => n26554, A2 => n18926, B1 => n26544, B2 => 
                           n4290, ZN => n24592);
   U21792 : OAI221_X1 port map( B1 => n21327, B2 => n26668, C1 => n21607, C2 =>
                           n26662, A => n24566, ZN => n24565);
   U21793 : AOI22_X1 port map( A1 => n26656, A2 => n9342, B1 => n26650, B2 => 
                           n18894, ZN => n24566);
   U21794 : OAI221_X1 port map( B1 => n20739, B2 => n26566, C1 => n21967, C2 =>
                           n26560, A => n24574, ZN => n24573);
   U21795 : AOI22_X1 port map( A1 => n26554, A2 => n18909, B1 => n26543, B2 => 
                           n4288, ZN => n24574);
   U21796 : OAI221_X1 port map( B1 => n21326, B2 => n26668, C1 => n21606, C2 =>
                           n26662, A => n24548, ZN => n24547);
   U21797 : AOI22_X1 port map( A1 => n26656, A2 => n9339, B1 => n26650, B2 => 
                           n18877, ZN => n24548);
   U21798 : OAI221_X1 port map( B1 => n20738, B2 => n26566, C1 => n21966, C2 =>
                           n26560, A => n24556, ZN => n24555);
   U21799 : AOI22_X1 port map( A1 => n26554, A2 => n18892, B1 => n26543, B2 => 
                           n4286, ZN => n24556);
   U21800 : OAI221_X1 port map( B1 => n21325, B2 => n26668, C1 => n21605, C2 =>
                           n26662, A => n24530, ZN => n24529);
   U21801 : AOI22_X1 port map( A1 => n26656, A2 => n9336, B1 => n26650, B2 => 
                           n18860, ZN => n24530);
   U21802 : OAI221_X1 port map( B1 => n20737, B2 => n26566, C1 => n21965, C2 =>
                           n26560, A => n24538, ZN => n24537);
   U21803 : AOI22_X1 port map( A1 => n26554, A2 => n18875, B1 => n26543, B2 => 
                           n4284, ZN => n24538);
   U21804 : OAI221_X1 port map( B1 => n21324, B2 => n26668, C1 => n21604, C2 =>
                           n26662, A => n24512, ZN => n24511);
   U21805 : AOI22_X1 port map( A1 => n26656, A2 => n9333, B1 => n26650, B2 => 
                           n18843, ZN => n24512);
   U21806 : OAI221_X1 port map( B1 => n20736, B2 => n26566, C1 => n21964, C2 =>
                           n26560, A => n24520, ZN => n24519);
   U21807 : AOI22_X1 port map( A1 => n26554, A2 => n18858, B1 => n26543, B2 => 
                           n4282, ZN => n24520);
   U21808 : OAI221_X1 port map( B1 => n21323, B2 => n26669, C1 => n21603, C2 =>
                           n26663, A => n24494, ZN => n24493);
   U21809 : AOI22_X1 port map( A1 => n26657, A2 => n9330, B1 => n26651, B2 => 
                           n18826, ZN => n24494);
   U21810 : OAI221_X1 port map( B1 => n20735, B2 => n26567, C1 => n21963, C2 =>
                           n26561, A => n24502, ZN => n24501);
   U21811 : AOI22_X1 port map( A1 => n26555, A2 => n18841, B1 => n26542, B2 => 
                           n4280, ZN => n24502);
   U21812 : OAI221_X1 port map( B1 => n21322, B2 => n26669, C1 => n21602, C2 =>
                           n26663, A => n24476, ZN => n24475);
   U21813 : AOI22_X1 port map( A1 => n26657, A2 => n9327, B1 => n26651, B2 => 
                           n18809, ZN => n24476);
   U21814 : OAI221_X1 port map( B1 => n20734, B2 => n26567, C1 => n21962, C2 =>
                           n26561, A => n24484, ZN => n24483);
   U21815 : AOI22_X1 port map( A1 => n26555, A2 => n18824, B1 => n26542, B2 => 
                           n4278, ZN => n24484);
   U21816 : OAI221_X1 port map( B1 => n21321, B2 => n26669, C1 => n21601, C2 =>
                           n26663, A => n24458, ZN => n24457);
   U21817 : AOI22_X1 port map( A1 => n26657, A2 => n9324, B1 => n26651, B2 => 
                           n18792, ZN => n24458);
   U21818 : OAI221_X1 port map( B1 => n20733, B2 => n26567, C1 => n21961, C2 =>
                           n26561, A => n24466, ZN => n24465);
   U21819 : AOI22_X1 port map( A1 => n26555, A2 => n18807, B1 => n26542, B2 => 
                           n4276, ZN => n24466);
   U21820 : OAI221_X1 port map( B1 => n21320, B2 => n26669, C1 => n21600, C2 =>
                           n26663, A => n24440, ZN => n24439);
   U21821 : AOI22_X1 port map( A1 => n26657, A2 => n9321, B1 => n26651, B2 => 
                           n18775, ZN => n24440);
   U21822 : OAI221_X1 port map( B1 => n20732, B2 => n26567, C1 => n21960, C2 =>
                           n26561, A => n24448, ZN => n24447);
   U21823 : AOI22_X1 port map( A1 => n26555, A2 => n18790, B1 => n26542, B2 => 
                           n4274, ZN => n24448);
   U21824 : OAI221_X1 port map( B1 => n21319, B2 => n26669, C1 => n21599, C2 =>
                           n26663, A => n24422, ZN => n24421);
   U21825 : AOI22_X1 port map( A1 => n26657, A2 => n9318, B1 => n26651, B2 => 
                           n18758, ZN => n24422);
   U21826 : OAI221_X1 port map( B1 => n20731, B2 => n26567, C1 => n21959, C2 =>
                           n26561, A => n24430, ZN => n24429);
   U21827 : AOI22_X1 port map( A1 => n26555, A2 => n18773, B1 => n26541, B2 => 
                           n4272, ZN => n24430);
   U21828 : OAI221_X1 port map( B1 => n21318, B2 => n26669, C1 => n21598, C2 =>
                           n26663, A => n24404, ZN => n24403);
   U21829 : AOI22_X1 port map( A1 => n26657, A2 => n9315, B1 => n26651, B2 => 
                           n18741, ZN => n24404);
   U21830 : OAI221_X1 port map( B1 => n20730, B2 => n26567, C1 => n21958, C2 =>
                           n26561, A => n24412, ZN => n24411);
   U21831 : AOI22_X1 port map( A1 => n26555, A2 => n18756, B1 => n26541, B2 => 
                           n4270, ZN => n24412);
   U21832 : OAI221_X1 port map( B1 => n21317, B2 => n26669, C1 => n21597, C2 =>
                           n26663, A => n24386, ZN => n24385);
   U21833 : AOI22_X1 port map( A1 => n26657, A2 => n9312, B1 => n26651, B2 => 
                           n18724, ZN => n24386);
   U21834 : OAI221_X1 port map( B1 => n20729, B2 => n26567, C1 => n21957, C2 =>
                           n26561, A => n24394, ZN => n24393);
   U21835 : AOI22_X1 port map( A1 => n26555, A2 => n18739, B1 => n26541, B2 => 
                           n4268, ZN => n24394);
   U21836 : OAI221_X1 port map( B1 => n21316, B2 => n26669, C1 => n21596, C2 =>
                           n26663, A => n24368, ZN => n24367);
   U21837 : AOI22_X1 port map( A1 => n26657, A2 => n9309, B1 => n26651, B2 => 
                           n18707, ZN => n24368);
   U21838 : OAI221_X1 port map( B1 => n20728, B2 => n26567, C1 => n21956, C2 =>
                           n26561, A => n24376, ZN => n24375);
   U21839 : AOI22_X1 port map( A1 => n26555, A2 => n18722, B1 => n26541, B2 => 
                           n4266, ZN => n24376);
   U21840 : OAI221_X1 port map( B1 => n21315, B2 => n26669, C1 => n21595, C2 =>
                           n26663, A => n24350, ZN => n24349);
   U21841 : AOI22_X1 port map( A1 => n26657, A2 => n9306, B1 => n26651, B2 => 
                           n18690, ZN => n24350);
   U21842 : OAI221_X1 port map( B1 => n20727, B2 => n26567, C1 => n21955, C2 =>
                           n26561, A => n24358, ZN => n24357);
   U21843 : AOI22_X1 port map( A1 => n26555, A2 => n18705, B1 => n26540, B2 => 
                           n4264, ZN => n24358);
   U21844 : OAI221_X1 port map( B1 => n21314, B2 => n26669, C1 => n21594, C2 =>
                           n26663, A => n24332, ZN => n24331);
   U21845 : AOI22_X1 port map( A1 => n26657, A2 => n9303, B1 => n26651, B2 => 
                           n18673, ZN => n24332);
   U21846 : OAI221_X1 port map( B1 => n20726, B2 => n26567, C1 => n21954, C2 =>
                           n26561, A => n24340, ZN => n24339);
   U21847 : AOI22_X1 port map( A1 => n26555, A2 => n18688, B1 => n26540, B2 => 
                           n4262, ZN => n24340);
   U21848 : OAI221_X1 port map( B1 => n21313, B2 => n26669, C1 => n21593, C2 =>
                           n26663, A => n24314, ZN => n24313);
   U21849 : AOI22_X1 port map( A1 => n26657, A2 => n9300, B1 => n26651, B2 => 
                           n18656, ZN => n24314);
   U21850 : OAI221_X1 port map( B1 => n20725, B2 => n26567, C1 => n21953, C2 =>
                           n26561, A => n24322, ZN => n24321);
   U21851 : AOI22_X1 port map( A1 => n26555, A2 => n18671, B1 => n26540, B2 => 
                           n4260, ZN => n24322);
   U21852 : OAI221_X1 port map( B1 => n21312, B2 => n26669, C1 => n21592, C2 =>
                           n26663, A => n24296, ZN => n24295);
   U21853 : AOI22_X1 port map( A1 => n26657, A2 => n9297, B1 => n26651, B2 => 
                           n18639, ZN => n24296);
   U21854 : OAI221_X1 port map( B1 => n20724, B2 => n26567, C1 => n21952, C2 =>
                           n26561, A => n24304, ZN => n24303);
   U21855 : AOI22_X1 port map( A1 => n26555, A2 => n18654, B1 => n26540, B2 => 
                           n4258, ZN => n24304);
   U21856 : OAI221_X1 port map( B1 => n21311, B2 => n26670, C1 => n21591, C2 =>
                           n26664, A => n24278, ZN => n24277);
   U21857 : AOI22_X1 port map( A1 => n26658, A2 => n9294, B1 => n26652, B2 => 
                           n18622, ZN => n24278);
   U21858 : OAI221_X1 port map( B1 => n20723, B2 => n26568, C1 => n21951, C2 =>
                           n26562, A => n24286, ZN => n24285);
   U21859 : AOI22_X1 port map( A1 => n26556, A2 => n18637, B1 => n26539, B2 => 
                           n4256, ZN => n24286);
   U21860 : OAI221_X1 port map( B1 => n21310, B2 => n26670, C1 => n21590, C2 =>
                           n26664, A => n24260, ZN => n24259);
   U21861 : AOI22_X1 port map( A1 => n26658, A2 => n9291, B1 => n26652, B2 => 
                           n18605, ZN => n24260);
   U21862 : OAI221_X1 port map( B1 => n20722, B2 => n26568, C1 => n21950, C2 =>
                           n26562, A => n24268, ZN => n24267);
   U21863 : AOI22_X1 port map( A1 => n26556, A2 => n18620, B1 => n26539, B2 => 
                           n4254, ZN => n24268);
   U21864 : OAI221_X1 port map( B1 => n21309, B2 => n26670, C1 => n21589, C2 =>
                           n26664, A => n24242, ZN => n24241);
   U21865 : AOI22_X1 port map( A1 => n26658, A2 => n9288, B1 => n26652, B2 => 
                           n18588, ZN => n24242);
   U21866 : OAI221_X1 port map( B1 => n20721, B2 => n26568, C1 => n21949, C2 =>
                           n26562, A => n24250, ZN => n24249);
   U21867 : AOI22_X1 port map( A1 => n26556, A2 => n18603, B1 => n26539, B2 => 
                           n4252, ZN => n24250);
   U21868 : OAI221_X1 port map( B1 => n21308, B2 => n26670, C1 => n21588, C2 =>
                           n26664, A => n24224, ZN => n24223);
   U21869 : AOI22_X1 port map( A1 => n26658, A2 => n9285, B1 => n26652, B2 => 
                           n18571, ZN => n24224);
   U21870 : OAI221_X1 port map( B1 => n20720, B2 => n26568, C1 => n21948, C2 =>
                           n26562, A => n24232, ZN => n24231);
   U21871 : AOI22_X1 port map( A1 => n26556, A2 => n18586, B1 => n26539, B2 => 
                           n4250, ZN => n24232);
   U21872 : OAI221_X1 port map( B1 => n21307, B2 => n26670, C1 => n21587, C2 =>
                           n26664, A => n24206, ZN => n24205);
   U21873 : AOI22_X1 port map( A1 => n26658, A2 => n9282, B1 => n26652, B2 => 
                           n18554, ZN => n24206);
   U21874 : OAI221_X1 port map( B1 => n20719, B2 => n26568, C1 => n21947, C2 =>
                           n26562, A => n24214, ZN => n24213);
   U21875 : AOI22_X1 port map( A1 => n26556, A2 => n18569, B1 => n26538, B2 => 
                           n4248, ZN => n24214);
   U21876 : OAI221_X1 port map( B1 => n21306, B2 => n26670, C1 => n21586, C2 =>
                           n26664, A => n24188, ZN => n24187);
   U21877 : AOI22_X1 port map( A1 => n26658, A2 => n9279, B1 => n26652, B2 => 
                           n18537, ZN => n24188);
   U21878 : OAI221_X1 port map( B1 => n20718, B2 => n26568, C1 => n21946, C2 =>
                           n26562, A => n24196, ZN => n24195);
   U21879 : AOI22_X1 port map( A1 => n26556, A2 => n18552, B1 => n26538, B2 => 
                           n4246, ZN => n24196);
   U21880 : OAI221_X1 port map( B1 => n21305, B2 => n26670, C1 => n21585, C2 =>
                           n26664, A => n24170, ZN => n24169);
   U21881 : AOI22_X1 port map( A1 => n26658, A2 => n9276, B1 => n26652, B2 => 
                           n18520, ZN => n24170);
   U21882 : OAI221_X1 port map( B1 => n20717, B2 => n26568, C1 => n21945, C2 =>
                           n26562, A => n24178, ZN => n24177);
   U21883 : AOI22_X1 port map( A1 => n26556, A2 => n18535, B1 => n26538, B2 => 
                           n4244, ZN => n24178);
   U21884 : OAI221_X1 port map( B1 => n21304, B2 => n26670, C1 => n21584, C2 =>
                           n26664, A => n24152, ZN => n24151);
   U21885 : AOI22_X1 port map( A1 => n26658, A2 => n9273, B1 => n26652, B2 => 
                           n18503, ZN => n24152);
   U21886 : OAI221_X1 port map( B1 => n20716, B2 => n26568, C1 => n21944, C2 =>
                           n26562, A => n24160, ZN => n24159);
   U21887 : AOI22_X1 port map( A1 => n26556, A2 => n18518, B1 => n26538, B2 => 
                           n4242, ZN => n24160);
   U21888 : OAI221_X1 port map( B1 => n21303, B2 => n26670, C1 => n21583, C2 =>
                           n26664, A => n24134, ZN => n24133);
   U21889 : AOI22_X1 port map( A1 => n26658, A2 => n9270, B1 => n26652, B2 => 
                           n18486, ZN => n24134);
   U21890 : OAI221_X1 port map( B1 => n20715, B2 => n26568, C1 => n21943, C2 =>
                           n26562, A => n24142, ZN => n24141);
   U21891 : AOI22_X1 port map( A1 => n26556, A2 => n18501, B1 => n26537, B2 => 
                           n4240, ZN => n24142);
   U21892 : OAI221_X1 port map( B1 => n21302, B2 => n26670, C1 => n21582, C2 =>
                           n26664, A => n24116, ZN => n24115);
   U21893 : AOI22_X1 port map( A1 => n26658, A2 => n9267, B1 => n26652, B2 => 
                           n18469, ZN => n24116);
   U21894 : OAI221_X1 port map( B1 => n20714, B2 => n26568, C1 => n21942, C2 =>
                           n26562, A => n24124, ZN => n24123);
   U21895 : AOI22_X1 port map( A1 => n26556, A2 => n18484, B1 => n26537, B2 => 
                           n4238, ZN => n24124);
   U21896 : OAI221_X1 port map( B1 => n21301, B2 => n26670, C1 => n21581, C2 =>
                           n26664, A => n24098, ZN => n24097);
   U21897 : AOI22_X1 port map( A1 => n26658, A2 => n9264, B1 => n26652, B2 => 
                           n18452, ZN => n24098);
   U21898 : OAI221_X1 port map( B1 => n20713, B2 => n26568, C1 => n21941, C2 =>
                           n26562, A => n24106, ZN => n24105);
   U21899 : AOI22_X1 port map( A1 => n26556, A2 => n18467, B1 => n26537, B2 => 
                           n4236, ZN => n24106);
   U21900 : OAI221_X1 port map( B1 => n21300, B2 => n26670, C1 => n21580, C2 =>
                           n26664, A => n24080, ZN => n24079);
   U21901 : AOI22_X1 port map( A1 => n26658, A2 => n9261, B1 => n26652, B2 => 
                           n18435, ZN => n24080);
   U21902 : OAI221_X1 port map( B1 => n20712, B2 => n26568, C1 => n21940, C2 =>
                           n26562, A => n24088, ZN => n24087);
   U21903 : AOI22_X1 port map( A1 => n26556, A2 => n18450, B1 => n26537, B2 => 
                           n4234, ZN => n24088);
   U21904 : OAI221_X1 port map( B1 => n21347, B2 => n26892, C1 => n21627, C2 =>
                           n26886, A => n23727, ZN => n23726);
   U21905 : AOI22_X1 port map( A1 => n26880, A2 => n9402, B1 => n26874, B2 => 
                           n19234, ZN => n23727);
   U21906 : OAI221_X1 port map( B1 => n20759, B2 => n26790, C1 => n21987, C2 =>
                           n26784, A => n23735, ZN => n23734);
   U21907 : AOI22_X1 port map( A1 => n26778, A2 => n19249, B1 => n26774, B2 => 
                           n4200, ZN => n23735);
   U21908 : OAI221_X1 port map( B1 => n21346, B2 => n26892, C1 => n21626, C2 =>
                           n26886, A => n23709, ZN => n23708);
   U21909 : AOI22_X1 port map( A1 => n26880, A2 => n9399, B1 => n26874, B2 => 
                           n19217, ZN => n23709);
   U21910 : OAI221_X1 port map( B1 => n20758, B2 => n26790, C1 => n21986, C2 =>
                           n26784, A => n23717, ZN => n23716);
   U21911 : AOI22_X1 port map( A1 => n26778, A2 => n19232, B1 => n26773, B2 => 
                           n4198, ZN => n23717);
   U21912 : OAI221_X1 port map( B1 => n21345, B2 => n26892, C1 => n21625, C2 =>
                           n26886, A => n23691, ZN => n23690);
   U21913 : AOI22_X1 port map( A1 => n26880, A2 => n9396, B1 => n26874, B2 => 
                           n19200, ZN => n23691);
   U21914 : OAI221_X1 port map( B1 => n20757, B2 => n26790, C1 => n21985, C2 =>
                           n26784, A => n23699, ZN => n23698);
   U21915 : AOI22_X1 port map( A1 => n26778, A2 => n19215, B1 => n26773, B2 => 
                           n4196, ZN => n23699);
   U21916 : OAI221_X1 port map( B1 => n21344, B2 => n26892, C1 => n21624, C2 =>
                           n26886, A => n23673, ZN => n23672);
   U21917 : AOI22_X1 port map( A1 => n26880, A2 => n9393, B1 => n26874, B2 => 
                           n19183, ZN => n23673);
   U21918 : OAI221_X1 port map( B1 => n20756, B2 => n26790, C1 => n21984, C2 =>
                           n26784, A => n23681, ZN => n23680);
   U21919 : AOI22_X1 port map( A1 => n26778, A2 => n19198, B1 => n26773, B2 => 
                           n4194, ZN => n23681);
   U21920 : OAI221_X1 port map( B1 => n21343, B2 => n26892, C1 => n21623, C2 =>
                           n26886, A => n23655, ZN => n23654);
   U21921 : AOI22_X1 port map( A1 => n26880, A2 => n9390, B1 => n26874, B2 => 
                           n19166, ZN => n23655);
   U21922 : OAI221_X1 port map( B1 => n20755, B2 => n26790, C1 => n21983, C2 =>
                           n26784, A => n23663, ZN => n23662);
   U21923 : AOI22_X1 port map( A1 => n26778, A2 => n19181, B1 => n26773, B2 => 
                           n4192, ZN => n23663);
   U21924 : OAI221_X1 port map( B1 => n21342, B2 => n26892, C1 => n21622, C2 =>
                           n26886, A => n23637, ZN => n23636);
   U21925 : AOI22_X1 port map( A1 => n26880, A2 => n9387, B1 => n26874, B2 => 
                           n19149, ZN => n23637);
   U21926 : OAI221_X1 port map( B1 => n20754, B2 => n26790, C1 => n21982, C2 =>
                           n26784, A => n23645, ZN => n23644);
   U21927 : AOI22_X1 port map( A1 => n26778, A2 => n19164, B1 => n26772, B2 => 
                           n4190, ZN => n23645);
   U21928 : OAI221_X1 port map( B1 => n21341, B2 => n26892, C1 => n21621, C2 =>
                           n26886, A => n23619, ZN => n23618);
   U21929 : AOI22_X1 port map( A1 => n26880, A2 => n9384, B1 => n26874, B2 => 
                           n19132, ZN => n23619);
   U21930 : OAI221_X1 port map( B1 => n20753, B2 => n26790, C1 => n21981, C2 =>
                           n26784, A => n23627, ZN => n23626);
   U21931 : AOI22_X1 port map( A1 => n26778, A2 => n19147, B1 => n26772, B2 => 
                           n4188, ZN => n23627);
   U21932 : OAI221_X1 port map( B1 => n21340, B2 => n26892, C1 => n21620, C2 =>
                           n26886, A => n23601, ZN => n23600);
   U21933 : AOI22_X1 port map( A1 => n26880, A2 => n9381, B1 => n26874, B2 => 
                           n19115, ZN => n23601);
   U21934 : OAI221_X1 port map( B1 => n20752, B2 => n26790, C1 => n21980, C2 =>
                           n26784, A => n23609, ZN => n23608);
   U21935 : AOI22_X1 port map( A1 => n26778, A2 => n19130, B1 => n26772, B2 => 
                           n4186, ZN => n23609);
   U21936 : OAI221_X1 port map( B1 => n21339, B2 => n26892, C1 => n21619, C2 =>
                           n26886, A => n23583, ZN => n23582);
   U21937 : AOI22_X1 port map( A1 => n26880, A2 => n9378, B1 => n26874, B2 => 
                           n19098, ZN => n23583);
   U21938 : OAI221_X1 port map( B1 => n20751, B2 => n26790, C1 => n21979, C2 =>
                           n26784, A => n23591, ZN => n23590);
   U21939 : AOI22_X1 port map( A1 => n26778, A2 => n19113, B1 => n26772, B2 => 
                           n4184, ZN => n23591);
   U21940 : OAI221_X1 port map( B1 => n21338, B2 => n26892, C1 => n21618, C2 =>
                           n26886, A => n23565, ZN => n23564);
   U21941 : AOI22_X1 port map( A1 => n26880, A2 => n9375, B1 => n26874, B2 => 
                           n19081, ZN => n23565);
   U21942 : OAI221_X1 port map( B1 => n20750, B2 => n26790, C1 => n21978, C2 =>
                           n26784, A => n23573, ZN => n23572);
   U21943 : AOI22_X1 port map( A1 => n26778, A2 => n19096, B1 => n26771, B2 => 
                           n4182, ZN => n23573);
   U21944 : OAI221_X1 port map( B1 => n21337, B2 => n26892, C1 => n21617, C2 =>
                           n26886, A => n23547, ZN => n23546);
   U21945 : AOI22_X1 port map( A1 => n26880, A2 => n9372, B1 => n26874, B2 => 
                           n19064, ZN => n23547);
   U21946 : OAI221_X1 port map( B1 => n20749, B2 => n26790, C1 => n21977, C2 =>
                           n26784, A => n23555, ZN => n23554);
   U21947 : AOI22_X1 port map( A1 => n26778, A2 => n19079, B1 => n26771, B2 => 
                           n4180, ZN => n23555);
   U21948 : OAI221_X1 port map( B1 => n21336, B2 => n26892, C1 => n21616, C2 =>
                           n26886, A => n23529, ZN => n23528);
   U21949 : AOI22_X1 port map( A1 => n26880, A2 => n9369, B1 => n26874, B2 => 
                           n19047, ZN => n23529);
   U21950 : OAI221_X1 port map( B1 => n20748, B2 => n26790, C1 => n21976, C2 =>
                           n26784, A => n23537, ZN => n23536);
   U21951 : AOI22_X1 port map( A1 => n26778, A2 => n19062, B1 => n26771, B2 => 
                           n4178, ZN => n23537);
   U21952 : OAI221_X1 port map( B1 => n21335, B2 => n26893, C1 => n21615, C2 =>
                           n26887, A => n23511, ZN => n23510);
   U21953 : AOI22_X1 port map( A1 => n26881, A2 => n9366, B1 => n26875, B2 => 
                           n19030, ZN => n23511);
   U21954 : OAI221_X1 port map( B1 => n20747, B2 => n26791, C1 => n21975, C2 =>
                           n26785, A => n23519, ZN => n23518);
   U21955 : AOI22_X1 port map( A1 => n26779, A2 => n19045, B1 => n26771, B2 => 
                           n4176, ZN => n23519);
   U21956 : OAI221_X1 port map( B1 => n21334, B2 => n26893, C1 => n21614, C2 =>
                           n26887, A => n23493, ZN => n23492);
   U21957 : AOI22_X1 port map( A1 => n26881, A2 => n9363, B1 => n26875, B2 => 
                           n19013, ZN => n23493);
   U21958 : OAI221_X1 port map( B1 => n20746, B2 => n26791, C1 => n21974, C2 =>
                           n26785, A => n23501, ZN => n23500);
   U21959 : AOI22_X1 port map( A1 => n26779, A2 => n19028, B1 => n26770, B2 => 
                           n4174, ZN => n23501);
   U21960 : OAI221_X1 port map( B1 => n21333, B2 => n26893, C1 => n21613, C2 =>
                           n26887, A => n23475, ZN => n23474);
   U21961 : AOI22_X1 port map( A1 => n26881, A2 => n9360, B1 => n26875, B2 => 
                           n18996, ZN => n23475);
   U21962 : OAI221_X1 port map( B1 => n20745, B2 => n26791, C1 => n21973, C2 =>
                           n26785, A => n23483, ZN => n23482);
   U21963 : AOI22_X1 port map( A1 => n26779, A2 => n19011, B1 => n26770, B2 => 
                           n4172, ZN => n23483);
   U21964 : OAI221_X1 port map( B1 => n21332, B2 => n26893, C1 => n21612, C2 =>
                           n26887, A => n23457, ZN => n23456);
   U21965 : AOI22_X1 port map( A1 => n26881, A2 => n9357, B1 => n26875, B2 => 
                           n18979, ZN => n23457);
   U21966 : OAI221_X1 port map( B1 => n20744, B2 => n26791, C1 => n21972, C2 =>
                           n26785, A => n23465, ZN => n23464);
   U21967 : AOI22_X1 port map( A1 => n26779, A2 => n18994, B1 => n26770, B2 => 
                           n4170, ZN => n23465);
   U21968 : OAI221_X1 port map( B1 => n21331, B2 => n26893, C1 => n21611, C2 =>
                           n26887, A => n23439, ZN => n23438);
   U21969 : AOI22_X1 port map( A1 => n26881, A2 => n9354, B1 => n26875, B2 => 
                           n18962, ZN => n23439);
   U21970 : OAI221_X1 port map( B1 => n20743, B2 => n26791, C1 => n21971, C2 =>
                           n26785, A => n23447, ZN => n23446);
   U21971 : AOI22_X1 port map( A1 => n26779, A2 => n18977, B1 => n26770, B2 => 
                           n4168, ZN => n23447);
   U21972 : OAI221_X1 port map( B1 => n21330, B2 => n26893, C1 => n21610, C2 =>
                           n26887, A => n23421, ZN => n23420);
   U21973 : AOI22_X1 port map( A1 => n26881, A2 => n9351, B1 => n26875, B2 => 
                           n18945, ZN => n23421);
   U21974 : OAI221_X1 port map( B1 => n20742, B2 => n26791, C1 => n21970, C2 =>
                           n26785, A => n23429, ZN => n23428);
   U21975 : AOI22_X1 port map( A1 => n26779, A2 => n18960, B1 => n26769, B2 => 
                           n4166, ZN => n23429);
   U21976 : OAI221_X1 port map( B1 => n21329, B2 => n26893, C1 => n21609, C2 =>
                           n26887, A => n23403, ZN => n23402);
   U21977 : AOI22_X1 port map( A1 => n26881, A2 => n9348, B1 => n26875, B2 => 
                           n18928, ZN => n23403);
   U21978 : OAI221_X1 port map( B1 => n20741, B2 => n26791, C1 => n21969, C2 =>
                           n26785, A => n23411, ZN => n23410);
   U21979 : AOI22_X1 port map( A1 => n26779, A2 => n18943, B1 => n26769, B2 => 
                           n4164, ZN => n23411);
   U21980 : OAI221_X1 port map( B1 => n21328, B2 => n26893, C1 => n21608, C2 =>
                           n26887, A => n23385, ZN => n23384);
   U21981 : AOI22_X1 port map( A1 => n26881, A2 => n9345, B1 => n26875, B2 => 
                           n18911, ZN => n23385);
   U21982 : OAI221_X1 port map( B1 => n20740, B2 => n26791, C1 => n21968, C2 =>
                           n26785, A => n23393, ZN => n23392);
   U21983 : AOI22_X1 port map( A1 => n26779, A2 => n18926, B1 => n26769, B2 => 
                           n4162, ZN => n23393);
   U21984 : OAI221_X1 port map( B1 => n21327, B2 => n26893, C1 => n21607, C2 =>
                           n26887, A => n23367, ZN => n23366);
   U21985 : AOI22_X1 port map( A1 => n26881, A2 => n9342, B1 => n26875, B2 => 
                           n18894, ZN => n23367);
   U21986 : OAI221_X1 port map( B1 => n20739, B2 => n26791, C1 => n21967, C2 =>
                           n26785, A => n23375, ZN => n23374);
   U21987 : AOI22_X1 port map( A1 => n26779, A2 => n18909, B1 => n26768, B2 => 
                           n4160, ZN => n23375);
   U21988 : OAI221_X1 port map( B1 => n21326, B2 => n26893, C1 => n21606, C2 =>
                           n26887, A => n23349, ZN => n23348);
   U21989 : AOI22_X1 port map( A1 => n26881, A2 => n9339, B1 => n26875, B2 => 
                           n18877, ZN => n23349);
   U21990 : OAI221_X1 port map( B1 => n20738, B2 => n26791, C1 => n21966, C2 =>
                           n26785, A => n23357, ZN => n23356);
   U21991 : AOI22_X1 port map( A1 => n26779, A2 => n18892, B1 => n26768, B2 => 
                           n4158, ZN => n23357);
   U21992 : OAI221_X1 port map( B1 => n21325, B2 => n26893, C1 => n21605, C2 =>
                           n26887, A => n23331, ZN => n23330);
   U21993 : AOI22_X1 port map( A1 => n26881, A2 => n9336, B1 => n26875, B2 => 
                           n18860, ZN => n23331);
   U21994 : OAI221_X1 port map( B1 => n20737, B2 => n26791, C1 => n21965, C2 =>
                           n26785, A => n23339, ZN => n23338);
   U21995 : AOI22_X1 port map( A1 => n26779, A2 => n18875, B1 => n26768, B2 => 
                           n4156, ZN => n23339);
   U21996 : OAI221_X1 port map( B1 => n21324, B2 => n26893, C1 => n21604, C2 =>
                           n26887, A => n23313, ZN => n23312);
   U21997 : AOI22_X1 port map( A1 => n26881, A2 => n9333, B1 => n26875, B2 => 
                           n18843, ZN => n23313);
   U21998 : OAI221_X1 port map( B1 => n20736, B2 => n26791, C1 => n21964, C2 =>
                           n26785, A => n23321, ZN => n23320);
   U21999 : AOI22_X1 port map( A1 => n26779, A2 => n18858, B1 => n26768, B2 => 
                           n4154, ZN => n23321);
   U22000 : OAI221_X1 port map( B1 => n21323, B2 => n26894, C1 => n21603, C2 =>
                           n26888, A => n23295, ZN => n23294);
   U22001 : AOI22_X1 port map( A1 => n26882, A2 => n9330, B1 => n26876, B2 => 
                           n18826, ZN => n23295);
   U22002 : OAI221_X1 port map( B1 => n20735, B2 => n26792, C1 => n21963, C2 =>
                           n26786, A => n23303, ZN => n23302);
   U22003 : AOI22_X1 port map( A1 => n26780, A2 => n18841, B1 => n26767, B2 => 
                           n4152, ZN => n23303);
   U22004 : OAI221_X1 port map( B1 => n21322, B2 => n26894, C1 => n21602, C2 =>
                           n26888, A => n23277, ZN => n23276);
   U22005 : AOI22_X1 port map( A1 => n26882, A2 => n9327, B1 => n26876, B2 => 
                           n18809, ZN => n23277);
   U22006 : OAI221_X1 port map( B1 => n20734, B2 => n26792, C1 => n21962, C2 =>
                           n26786, A => n23285, ZN => n23284);
   U22007 : AOI22_X1 port map( A1 => n26780, A2 => n18824, B1 => n26767, B2 => 
                           n4150, ZN => n23285);
   U22008 : OAI221_X1 port map( B1 => n21321, B2 => n26894, C1 => n21601, C2 =>
                           n26888, A => n23259, ZN => n23258);
   U22009 : AOI22_X1 port map( A1 => n26882, A2 => n9324, B1 => n26876, B2 => 
                           n18792, ZN => n23259);
   U22010 : OAI221_X1 port map( B1 => n20733, B2 => n26792, C1 => n21961, C2 =>
                           n26786, A => n23267, ZN => n23266);
   U22011 : AOI22_X1 port map( A1 => n26780, A2 => n18807, B1 => n26767, B2 => 
                           n4148, ZN => n23267);
   U22012 : OAI221_X1 port map( B1 => n21320, B2 => n26894, C1 => n21600, C2 =>
                           n26888, A => n23241, ZN => n23240);
   U22013 : AOI22_X1 port map( A1 => n26882, A2 => n9321, B1 => n26876, B2 => 
                           n18775, ZN => n23241);
   U22014 : OAI221_X1 port map( B1 => n20732, B2 => n26792, C1 => n21960, C2 =>
                           n26786, A => n23249, ZN => n23248);
   U22015 : AOI22_X1 port map( A1 => n26780, A2 => n18790, B1 => n26767, B2 => 
                           n4146, ZN => n23249);
   U22016 : OAI221_X1 port map( B1 => n21319, B2 => n26894, C1 => n21599, C2 =>
                           n26888, A => n23223, ZN => n23222);
   U22017 : AOI22_X1 port map( A1 => n26882, A2 => n9318, B1 => n26876, B2 => 
                           n18758, ZN => n23223);
   U22018 : OAI221_X1 port map( B1 => n20731, B2 => n26792, C1 => n21959, C2 =>
                           n26786, A => n23231, ZN => n23230);
   U22019 : AOI22_X1 port map( A1 => n26780, A2 => n18773, B1 => n26766, B2 => 
                           n4144, ZN => n23231);
   U22020 : OAI221_X1 port map( B1 => n21318, B2 => n26894, C1 => n21598, C2 =>
                           n26888, A => n23205, ZN => n23204);
   U22021 : AOI22_X1 port map( A1 => n26882, A2 => n9315, B1 => n26876, B2 => 
                           n18741, ZN => n23205);
   U22022 : OAI221_X1 port map( B1 => n20730, B2 => n26792, C1 => n21958, C2 =>
                           n26786, A => n23213, ZN => n23212);
   U22023 : AOI22_X1 port map( A1 => n26780, A2 => n18756, B1 => n26766, B2 => 
                           n4142, ZN => n23213);
   U22024 : OAI221_X1 port map( B1 => n21317, B2 => n26894, C1 => n21597, C2 =>
                           n26888, A => n23187, ZN => n23186);
   U22025 : AOI22_X1 port map( A1 => n26882, A2 => n9312, B1 => n26876, B2 => 
                           n18724, ZN => n23187);
   U22026 : OAI221_X1 port map( B1 => n20729, B2 => n26792, C1 => n21957, C2 =>
                           n26786, A => n23195, ZN => n23194);
   U22027 : AOI22_X1 port map( A1 => n26780, A2 => n18739, B1 => n26766, B2 => 
                           n4140, ZN => n23195);
   U22028 : OAI221_X1 port map( B1 => n21316, B2 => n26894, C1 => n21596, C2 =>
                           n26888, A => n23169, ZN => n23168);
   U22029 : AOI22_X1 port map( A1 => n26882, A2 => n9309, B1 => n26876, B2 => 
                           n18707, ZN => n23169);
   U22030 : OAI221_X1 port map( B1 => n20728, B2 => n26792, C1 => n21956, C2 =>
                           n26786, A => n23177, ZN => n23176);
   U22031 : AOI22_X1 port map( A1 => n26780, A2 => n18722, B1 => n26766, B2 => 
                           n4138, ZN => n23177);
   U22032 : OAI221_X1 port map( B1 => n21315, B2 => n26894, C1 => n21595, C2 =>
                           n26888, A => n23151, ZN => n23150);
   U22033 : AOI22_X1 port map( A1 => n26882, A2 => n9306, B1 => n26876, B2 => 
                           n18690, ZN => n23151);
   U22034 : OAI221_X1 port map( B1 => n20727, B2 => n26792, C1 => n21955, C2 =>
                           n26786, A => n23159, ZN => n23158);
   U22035 : AOI22_X1 port map( A1 => n26780, A2 => n18705, B1 => n26765, B2 => 
                           n4136, ZN => n23159);
   U22036 : OAI221_X1 port map( B1 => n21314, B2 => n26894, C1 => n21594, C2 =>
                           n26888, A => n23133, ZN => n23132);
   U22037 : AOI22_X1 port map( A1 => n26882, A2 => n9303, B1 => n26876, B2 => 
                           n18673, ZN => n23133);
   U22038 : OAI221_X1 port map( B1 => n20726, B2 => n26792, C1 => n21954, C2 =>
                           n26786, A => n23141, ZN => n23140);
   U22039 : AOI22_X1 port map( A1 => n26780, A2 => n18688, B1 => n26765, B2 => 
                           n4134, ZN => n23141);
   U22040 : OAI221_X1 port map( B1 => n21313, B2 => n26894, C1 => n21593, C2 =>
                           n26888, A => n23115, ZN => n23114);
   U22041 : AOI22_X1 port map( A1 => n26882, A2 => n9300, B1 => n26876, B2 => 
                           n18656, ZN => n23115);
   U22042 : OAI221_X1 port map( B1 => n20725, B2 => n26792, C1 => n21953, C2 =>
                           n26786, A => n23123, ZN => n23122);
   U22043 : AOI22_X1 port map( A1 => n26780, A2 => n18671, B1 => n26765, B2 => 
                           n4132, ZN => n23123);
   U22044 : OAI221_X1 port map( B1 => n21312, B2 => n26894, C1 => n21592, C2 =>
                           n26888, A => n23097, ZN => n23096);
   U22045 : AOI22_X1 port map( A1 => n26882, A2 => n9297, B1 => n26876, B2 => 
                           n18639, ZN => n23097);
   U22046 : OAI221_X1 port map( B1 => n20724, B2 => n26792, C1 => n21952, C2 =>
                           n26786, A => n23105, ZN => n23104);
   U22047 : AOI22_X1 port map( A1 => n26780, A2 => n18654, B1 => n26765, B2 => 
                           n4130, ZN => n23105);
   U22048 : OAI221_X1 port map( B1 => n21311, B2 => n26895, C1 => n21591, C2 =>
                           n26889, A => n23079, ZN => n23078);
   U22049 : AOI22_X1 port map( A1 => n26883, A2 => n9294, B1 => n26877, B2 => 
                           n18622, ZN => n23079);
   U22050 : OAI221_X1 port map( B1 => n20723, B2 => n26793, C1 => n21951, C2 =>
                           n26787, A => n23087, ZN => n23086);
   U22051 : AOI22_X1 port map( A1 => n26781, A2 => n18637, B1 => n26764, B2 => 
                           n4128, ZN => n23087);
   U22052 : OAI221_X1 port map( B1 => n21310, B2 => n26895, C1 => n21590, C2 =>
                           n26889, A => n23061, ZN => n23060);
   U22053 : AOI22_X1 port map( A1 => n26883, A2 => n9291, B1 => n26877, B2 => 
                           n18605, ZN => n23061);
   U22054 : OAI221_X1 port map( B1 => n20722, B2 => n26793, C1 => n21950, C2 =>
                           n26787, A => n23069, ZN => n23068);
   U22055 : AOI22_X1 port map( A1 => n26781, A2 => n18620, B1 => n26764, B2 => 
                           n4126, ZN => n23069);
   U22056 : OAI221_X1 port map( B1 => n21309, B2 => n26895, C1 => n21589, C2 =>
                           n26889, A => n23043, ZN => n23042);
   U22057 : AOI22_X1 port map( A1 => n26883, A2 => n9288, B1 => n26877, B2 => 
                           n18588, ZN => n23043);
   U22058 : OAI221_X1 port map( B1 => n20721, B2 => n26793, C1 => n21949, C2 =>
                           n26787, A => n23051, ZN => n23050);
   U22059 : AOI22_X1 port map( A1 => n26781, A2 => n18603, B1 => n26764, B2 => 
                           n4124, ZN => n23051);
   U22060 : OAI221_X1 port map( B1 => n21308, B2 => n26895, C1 => n21588, C2 =>
                           n26889, A => n23025, ZN => n23024);
   U22061 : AOI22_X1 port map( A1 => n26883, A2 => n9285, B1 => n26877, B2 => 
                           n18571, ZN => n23025);
   U22062 : OAI221_X1 port map( B1 => n20720, B2 => n26793, C1 => n21948, C2 =>
                           n26787, A => n23033, ZN => n23032);
   U22063 : AOI22_X1 port map( A1 => n26781, A2 => n18586, B1 => n26764, B2 => 
                           n4122, ZN => n23033);
   U22064 : OAI221_X1 port map( B1 => n21307, B2 => n26895, C1 => n21587, C2 =>
                           n26889, A => n23007, ZN => n23006);
   U22065 : AOI22_X1 port map( A1 => n26883, A2 => n9282, B1 => n26877, B2 => 
                           n18554, ZN => n23007);
   U22066 : OAI221_X1 port map( B1 => n20719, B2 => n26793, C1 => n21947, C2 =>
                           n26787, A => n23015, ZN => n23014);
   U22067 : AOI22_X1 port map( A1 => n26781, A2 => n18569, B1 => n26763, B2 => 
                           n4120, ZN => n23015);
   U22068 : OAI221_X1 port map( B1 => n21306, B2 => n26895, C1 => n21586, C2 =>
                           n26889, A => n22989, ZN => n22988);
   U22069 : AOI22_X1 port map( A1 => n26883, A2 => n9279, B1 => n26877, B2 => 
                           n18537, ZN => n22989);
   U22070 : OAI221_X1 port map( B1 => n20718, B2 => n26793, C1 => n21946, C2 =>
                           n26787, A => n22997, ZN => n22996);
   U22071 : AOI22_X1 port map( A1 => n26781, A2 => n18552, B1 => n26763, B2 => 
                           n4118, ZN => n22997);
   U22072 : OAI221_X1 port map( B1 => n21305, B2 => n26895, C1 => n21585, C2 =>
                           n26889, A => n22971, ZN => n22970);
   U22073 : AOI22_X1 port map( A1 => n26883, A2 => n9276, B1 => n26877, B2 => 
                           n18520, ZN => n22971);
   U22074 : OAI221_X1 port map( B1 => n20717, B2 => n26793, C1 => n21945, C2 =>
                           n26787, A => n22979, ZN => n22978);
   U22075 : AOI22_X1 port map( A1 => n26781, A2 => n18535, B1 => n26763, B2 => 
                           n4116, ZN => n22979);
   U22076 : OAI221_X1 port map( B1 => n21304, B2 => n26895, C1 => n21584, C2 =>
                           n26889, A => n22953, ZN => n22952);
   U22077 : AOI22_X1 port map( A1 => n26883, A2 => n9273, B1 => n26877, B2 => 
                           n18503, ZN => n22953);
   U22078 : OAI221_X1 port map( B1 => n20716, B2 => n26793, C1 => n21944, C2 =>
                           n26787, A => n22961, ZN => n22960);
   U22079 : AOI22_X1 port map( A1 => n26781, A2 => n18518, B1 => n26763, B2 => 
                           n4114, ZN => n22961);
   U22080 : OAI221_X1 port map( B1 => n21303, B2 => n26895, C1 => n21583, C2 =>
                           n26889, A => n22935, ZN => n22934);
   U22081 : AOI22_X1 port map( A1 => n26883, A2 => n9270, B1 => n26877, B2 => 
                           n18486, ZN => n22935);
   U22082 : OAI221_X1 port map( B1 => n20715, B2 => n26793, C1 => n21943, C2 =>
                           n26787, A => n22943, ZN => n22942);
   U22083 : AOI22_X1 port map( A1 => n26781, A2 => n18501, B1 => n26762, B2 => 
                           n4112, ZN => n22943);
   U22084 : OAI221_X1 port map( B1 => n21302, B2 => n26895, C1 => n21582, C2 =>
                           n26889, A => n22917, ZN => n22916);
   U22085 : AOI22_X1 port map( A1 => n26883, A2 => n9267, B1 => n26877, B2 => 
                           n18469, ZN => n22917);
   U22086 : OAI221_X1 port map( B1 => n20714, B2 => n26793, C1 => n21942, C2 =>
                           n26787, A => n22925, ZN => n22924);
   U22087 : AOI22_X1 port map( A1 => n26781, A2 => n18484, B1 => n26762, B2 => 
                           n4110, ZN => n22925);
   U22088 : OAI221_X1 port map( B1 => n21301, B2 => n26895, C1 => n21581, C2 =>
                           n26889, A => n22899, ZN => n22898);
   U22089 : AOI22_X1 port map( A1 => n26883, A2 => n9264, B1 => n26877, B2 => 
                           n18452, ZN => n22899);
   U22090 : OAI221_X1 port map( B1 => n20713, B2 => n26793, C1 => n21941, C2 =>
                           n26787, A => n22907, ZN => n22906);
   U22091 : AOI22_X1 port map( A1 => n26781, A2 => n18467, B1 => n26762, B2 => 
                           n4108, ZN => n22907);
   U22092 : OAI221_X1 port map( B1 => n21300, B2 => n26895, C1 => n21580, C2 =>
                           n26889, A => n22881, ZN => n22880);
   U22093 : AOI22_X1 port map( A1 => n26883, A2 => n9261, B1 => n26877, B2 => 
                           n18435, ZN => n22881);
   U22094 : OAI221_X1 port map( B1 => n20712, B2 => n26793, C1 => n21940, C2 =>
                           n26787, A => n22889, ZN => n22888);
   U22095 : AOI22_X1 port map( A1 => n26781, A2 => n18450, B1 => n26762, B2 => 
                           n4106, ZN => n22889);
   U22096 : OAI221_X1 port map( B1 => n21164, B2 => n26671, C1 => n21480, C2 =>
                           n26665, A => n23976, ZN => n23973);
   U22097 : AOI22_X1 port map( A1 => n26659, A2 => n9249, B1 => n26653, B2 => 
                           n18367, ZN => n23976);
   U22098 : OAI221_X1 port map( B1 => n20708, B2 => n26569, C1 => n21504, C2 =>
                           n26563, A => n24001, ZN => n23998);
   U22099 : AOI22_X1 port map( A1 => n26557, A2 => n18382, B1 => n26544, B2 => 
                           n4226, ZN => n24001);
   U22100 : OAI221_X1 port map( B1 => n21167, B2 => n26671, C1 => n21483, C2 =>
                           n26665, A => n24062, ZN => n24061);
   U22101 : AOI22_X1 port map( A1 => n26659, A2 => n9258, B1 => n26653, B2 => 
                           n18418, ZN => n24062);
   U22102 : OAI221_X1 port map( B1 => n20711, B2 => n26569, C1 => n21507, C2 =>
                           n26563, A => n24070, ZN => n24069);
   U22103 : AOI22_X1 port map( A1 => n26557, A2 => n18433, B1 => n26536, B2 => 
                           n4232, ZN => n24070);
   U22104 : OAI221_X1 port map( B1 => n21166, B2 => n26671, C1 => n21482, C2 =>
                           n26665, A => n24044, ZN => n24043);
   U22105 : AOI22_X1 port map( A1 => n26659, A2 => n9255, B1 => n26653, B2 => 
                           n18401, ZN => n24044);
   U22106 : OAI221_X1 port map( B1 => n20710, B2 => n26569, C1 => n21506, C2 =>
                           n26563, A => n24052, ZN => n24051);
   U22107 : AOI22_X1 port map( A1 => n26557, A2 => n18416, B1 => n26536, B2 => 
                           n4230, ZN => n24052);
   U22108 : OAI221_X1 port map( B1 => n21165, B2 => n26671, C1 => n21481, C2 =>
                           n26665, A => n24026, ZN => n24025);
   U22109 : AOI22_X1 port map( A1 => n26659, A2 => n9252, B1 => n26653, B2 => 
                           n18384, ZN => n24026);
   U22110 : OAI221_X1 port map( B1 => n20709, B2 => n26569, C1 => n21505, C2 =>
                           n26563, A => n24034, ZN => n24033);
   U22111 : AOI22_X1 port map( A1 => n26557, A2 => n18399, B1 => n26536, B2 => 
                           n4228, ZN => n24034);
   U22112 : OAI221_X1 port map( B1 => n21167, B2 => n26896, C1 => n21483, C2 =>
                           n26890, A => n22863, ZN => n22862);
   U22113 : AOI22_X1 port map( A1 => n26884, A2 => n9258, B1 => n26878, B2 => 
                           n18418, ZN => n22863);
   U22114 : OAI221_X1 port map( B1 => n20711, B2 => n26794, C1 => n21507, C2 =>
                           n26788, A => n22871, ZN => n22870);
   U22115 : AOI22_X1 port map( A1 => n26782, A2 => n18433, B1 => n26761, B2 => 
                           n4104, ZN => n22871);
   U22116 : OAI221_X1 port map( B1 => n21166, B2 => n26896, C1 => n21482, C2 =>
                           n26890, A => n22845, ZN => n22844);
   U22117 : AOI22_X1 port map( A1 => n26884, A2 => n9255, B1 => n26878, B2 => 
                           n18401, ZN => n22845);
   U22118 : OAI221_X1 port map( B1 => n20710, B2 => n26794, C1 => n21506, C2 =>
                           n26788, A => n22853, ZN => n22852);
   U22119 : AOI22_X1 port map( A1 => n26782, A2 => n18416, B1 => n26761, B2 => 
                           n4102, ZN => n22853);
   U22120 : OAI221_X1 port map( B1 => n21165, B2 => n26896, C1 => n21481, C2 =>
                           n26890, A => n22827, ZN => n22826);
   U22121 : AOI22_X1 port map( A1 => n26884, A2 => n9252, B1 => n26878, B2 => 
                           n18384, ZN => n22827);
   U22122 : OAI221_X1 port map( B1 => n20709, B2 => n26794, C1 => n21505, C2 =>
                           n26788, A => n22835, ZN => n22834);
   U22123 : AOI22_X1 port map( A1 => n26782, A2 => n18399, B1 => n26761, B2 => 
                           n4100, ZN => n22835);
   U22124 : OAI221_X1 port map( B1 => n21164, B2 => n26896, C1 => n21480, C2 =>
                           n26890, A => n22777, ZN => n22774);
   U22125 : AOI22_X1 port map( A1 => n26884, A2 => n9249, B1 => n26878, B2 => 
                           n18367, ZN => n22777);
   U22126 : OAI221_X1 port map( B1 => n20708, B2 => n26794, C1 => n21504, C2 =>
                           n26788, A => n22802, ZN => n22799);
   U22127 : AOI22_X1 port map( A1 => n26782, A2 => n18382, B1 => n26769, B2 => 
                           n4098, ZN => n22802);
   U22128 : OAI221_X1 port map( B1 => n21359, B2 => n26666, C1 => n21639, C2 =>
                           n26660, A => n25142, ZN => n25141);
   U22129 : AOI22_X1 port map( A1 => n26654, A2 => n9438, B1 => n26648, B2 => 
                           n19438, ZN => n25142);
   U22130 : OAI221_X1 port map( B1 => n20771, B2 => n26564, C1 => n21999, C2 =>
                           n26558, A => n25160, ZN => n25159);
   U22131 : AOI22_X1 port map( A1 => n26552, A2 => n19453, B1 => n26530, B2 => 
                           n4352, ZN => n25160);
   U22132 : OAI221_X1 port map( B1 => n21358, B2 => n26666, C1 => n21638, C2 =>
                           n26660, A => n25124, ZN => n25123);
   U22133 : AOI22_X1 port map( A1 => n26654, A2 => n9435, B1 => n26648, B2 => 
                           n19421, ZN => n25124);
   U22134 : OAI221_X1 port map( B1 => n20770, B2 => n26564, C1 => n21998, C2 =>
                           n26558, A => n25132, ZN => n25131);
   U22135 : AOI22_X1 port map( A1 => n26552, A2 => n19436, B1 => n26551, B2 => 
                           n4350, ZN => n25132);
   U22136 : OAI221_X1 port map( B1 => n21357, B2 => n26666, C1 => n21637, C2 =>
                           n26660, A => n25106, ZN => n25105);
   U22137 : AOI22_X1 port map( A1 => n26654, A2 => n9432, B1 => n26648, B2 => 
                           n19404, ZN => n25106);
   U22138 : OAI221_X1 port map( B1 => n20769, B2 => n26564, C1 => n21997, C2 =>
                           n26558, A => n25114, ZN => n25113);
   U22139 : AOI22_X1 port map( A1 => n26552, A2 => n19419, B1 => n26551, B2 => 
                           n4348, ZN => n25114);
   U22140 : OAI221_X1 port map( B1 => n21356, B2 => n26666, C1 => n21636, C2 =>
                           n26660, A => n25088, ZN => n25087);
   U22141 : AOI22_X1 port map( A1 => n26654, A2 => n9429, B1 => n26648, B2 => 
                           n19387, ZN => n25088);
   U22142 : OAI221_X1 port map( B1 => n20768, B2 => n26564, C1 => n21996, C2 =>
                           n26558, A => n25096, ZN => n25095);
   U22143 : AOI22_X1 port map( A1 => n26552, A2 => n19402, B1 => n26551, B2 => 
                           n4346, ZN => n25096);
   U22144 : OAI221_X1 port map( B1 => n21355, B2 => n26666, C1 => n21635, C2 =>
                           n26660, A => n25070, ZN => n25069);
   U22145 : AOI22_X1 port map( A1 => n26654, A2 => n9426, B1 => n26648, B2 => 
                           n19370, ZN => n25070);
   U22146 : OAI221_X1 port map( B1 => n20767, B2 => n26564, C1 => n21995, C2 =>
                           n26558, A => n25078, ZN => n25077);
   U22147 : AOI22_X1 port map( A1 => n26552, A2 => n19385, B1 => n26551, B2 => 
                           n4344, ZN => n25078);
   U22148 : OAI221_X1 port map( B1 => n21354, B2 => n26666, C1 => n21634, C2 =>
                           n26660, A => n25052, ZN => n25051);
   U22149 : AOI22_X1 port map( A1 => n26654, A2 => n9423, B1 => n26648, B2 => 
                           n19353, ZN => n25052);
   U22150 : OAI221_X1 port map( B1 => n20766, B2 => n26564, C1 => n21994, C2 =>
                           n26558, A => n25060, ZN => n25059);
   U22151 : AOI22_X1 port map( A1 => n26552, A2 => n19368, B1 => n26550, B2 => 
                           n4342, ZN => n25060);
   U22152 : OAI221_X1 port map( B1 => n21353, B2 => n26666, C1 => n21633, C2 =>
                           n26660, A => n25034, ZN => n25033);
   U22153 : AOI22_X1 port map( A1 => n26654, A2 => n9420, B1 => n26648, B2 => 
                           n19336, ZN => n25034);
   U22154 : OAI221_X1 port map( B1 => n20765, B2 => n26564, C1 => n21993, C2 =>
                           n26558, A => n25042, ZN => n25041);
   U22155 : AOI22_X1 port map( A1 => n26552, A2 => n19351, B1 => n26550, B2 => 
                           n4340, ZN => n25042);
   U22156 : OAI221_X1 port map( B1 => n21352, B2 => n26666, C1 => n21632, C2 =>
                           n26660, A => n25016, ZN => n25015);
   U22157 : AOI22_X1 port map( A1 => n26654, A2 => n9417, B1 => n26648, B2 => 
                           n19319, ZN => n25016);
   U22158 : OAI221_X1 port map( B1 => n20764, B2 => n26564, C1 => n21992, C2 =>
                           n26558, A => n25024, ZN => n25023);
   U22159 : AOI22_X1 port map( A1 => n26552, A2 => n19334, B1 => n26550, B2 => 
                           n4338, ZN => n25024);
   U22160 : OAI221_X1 port map( B1 => n21351, B2 => n26666, C1 => n21631, C2 =>
                           n26660, A => n24998, ZN => n24997);
   U22161 : AOI22_X1 port map( A1 => n26654, A2 => n9414, B1 => n26648, B2 => 
                           n19302, ZN => n24998);
   U22162 : OAI221_X1 port map( B1 => n20763, B2 => n26564, C1 => n21991, C2 =>
                           n26558, A => n25006, ZN => n25005);
   U22163 : AOI22_X1 port map( A1 => n26552, A2 => n19317, B1 => n26550, B2 => 
                           n4336, ZN => n25006);
   U22164 : OAI221_X1 port map( B1 => n21350, B2 => n26666, C1 => n21630, C2 =>
                           n26660, A => n24980, ZN => n24979);
   U22165 : AOI22_X1 port map( A1 => n26654, A2 => n9411, B1 => n26648, B2 => 
                           n19285, ZN => n24980);
   U22166 : OAI221_X1 port map( B1 => n20762, B2 => n26564, C1 => n21990, C2 =>
                           n26558, A => n24988, ZN => n24987);
   U22167 : AOI22_X1 port map( A1 => n26552, A2 => n19300, B1 => n26549, B2 => 
                           n4334, ZN => n24988);
   U22168 : OAI221_X1 port map( B1 => n21349, B2 => n26666, C1 => n21629, C2 =>
                           n26660, A => n24962, ZN => n24961);
   U22169 : AOI22_X1 port map( A1 => n26654, A2 => n9408, B1 => n26648, B2 => 
                           n19268, ZN => n24962);
   U22170 : OAI221_X1 port map( B1 => n20761, B2 => n26564, C1 => n21989, C2 =>
                           n26558, A => n24970, ZN => n24969);
   U22171 : AOI22_X1 port map( A1 => n26552, A2 => n19283, B1 => n26549, B2 => 
                           n4332, ZN => n24970);
   U22172 : OAI221_X1 port map( B1 => n21348, B2 => n26666, C1 => n21628, C2 =>
                           n26660, A => n24944, ZN => n24943);
   U22173 : AOI22_X1 port map( A1 => n26654, A2 => n9405, B1 => n26648, B2 => 
                           n19251, ZN => n24944);
   U22174 : OAI221_X1 port map( B1 => n20760, B2 => n26564, C1 => n21988, C2 =>
                           n26558, A => n24952, ZN => n24951);
   U22175 : AOI22_X1 port map( A1 => n26552, A2 => n19266, B1 => n26549, B2 => 
                           n4330, ZN => n24952);
   U22176 : OAI221_X1 port map( B1 => n21359, B2 => n26891, C1 => n21639, C2 =>
                           n26885, A => n23943, ZN => n23942);
   U22177 : AOI22_X1 port map( A1 => n26879, A2 => n9438, B1 => n26873, B2 => 
                           n19438, ZN => n23943);
   U22178 : OAI221_X1 port map( B1 => n20771, B2 => n26789, C1 => n21999, C2 =>
                           n26783, A => n23961, ZN => n23960);
   U22179 : AOI22_X1 port map( A1 => n26777, A2 => n19453, B1 => n26755, B2 => 
                           n4224, ZN => n23961);
   U22180 : OAI221_X1 port map( B1 => n21358, B2 => n26891, C1 => n21638, C2 =>
                           n26885, A => n23925, ZN => n23924);
   U22181 : AOI22_X1 port map( A1 => n26879, A2 => n9435, B1 => n26873, B2 => 
                           n19421, ZN => n23925);
   U22182 : OAI221_X1 port map( B1 => n20770, B2 => n26789, C1 => n21998, C2 =>
                           n26783, A => n23933, ZN => n23932);
   U22183 : AOI22_X1 port map( A1 => n26777, A2 => n19436, B1 => n26776, B2 => 
                           n4222, ZN => n23933);
   U22184 : OAI221_X1 port map( B1 => n21357, B2 => n26891, C1 => n21637, C2 =>
                           n26885, A => n23907, ZN => n23906);
   U22185 : AOI22_X1 port map( A1 => n26879, A2 => n9432, B1 => n26873, B2 => 
                           n19404, ZN => n23907);
   U22186 : OAI221_X1 port map( B1 => n20769, B2 => n26789, C1 => n21997, C2 =>
                           n26783, A => n23915, ZN => n23914);
   U22187 : AOI22_X1 port map( A1 => n26777, A2 => n19419, B1 => n26776, B2 => 
                           n4220, ZN => n23915);
   U22188 : OAI221_X1 port map( B1 => n21356, B2 => n26891, C1 => n21636, C2 =>
                           n26885, A => n23889, ZN => n23888);
   U22189 : AOI22_X1 port map( A1 => n26879, A2 => n9429, B1 => n26873, B2 => 
                           n19387, ZN => n23889);
   U22190 : OAI221_X1 port map( B1 => n20768, B2 => n26789, C1 => n21996, C2 =>
                           n26783, A => n23897, ZN => n23896);
   U22191 : AOI22_X1 port map( A1 => n26777, A2 => n19402, B1 => n26776, B2 => 
                           n4218, ZN => n23897);
   U22192 : OAI221_X1 port map( B1 => n21355, B2 => n26891, C1 => n21635, C2 =>
                           n26885, A => n23871, ZN => n23870);
   U22193 : AOI22_X1 port map( A1 => n26879, A2 => n9426, B1 => n26873, B2 => 
                           n19370, ZN => n23871);
   U22194 : OAI221_X1 port map( B1 => n20767, B2 => n26789, C1 => n21995, C2 =>
                           n26783, A => n23879, ZN => n23878);
   U22195 : AOI22_X1 port map( A1 => n26777, A2 => n19385, B1 => n26776, B2 => 
                           n4216, ZN => n23879);
   U22196 : OAI221_X1 port map( B1 => n21354, B2 => n26891, C1 => n21634, C2 =>
                           n26885, A => n23853, ZN => n23852);
   U22197 : AOI22_X1 port map( A1 => n26879, A2 => n9423, B1 => n26873, B2 => 
                           n19353, ZN => n23853);
   U22198 : OAI221_X1 port map( B1 => n20766, B2 => n26789, C1 => n21994, C2 =>
                           n26783, A => n23861, ZN => n23860);
   U22199 : AOI22_X1 port map( A1 => n26777, A2 => n19368, B1 => n26775, B2 => 
                           n4214, ZN => n23861);
   U22200 : OAI221_X1 port map( B1 => n21353, B2 => n26891, C1 => n21633, C2 =>
                           n26885, A => n23835, ZN => n23834);
   U22201 : AOI22_X1 port map( A1 => n26879, A2 => n9420, B1 => n26873, B2 => 
                           n19336, ZN => n23835);
   U22202 : OAI221_X1 port map( B1 => n20765, B2 => n26789, C1 => n21993, C2 =>
                           n26783, A => n23843, ZN => n23842);
   U22203 : AOI22_X1 port map( A1 => n26777, A2 => n19351, B1 => n26775, B2 => 
                           n4212, ZN => n23843);
   U22204 : OAI221_X1 port map( B1 => n21352, B2 => n26891, C1 => n21632, C2 =>
                           n26885, A => n23817, ZN => n23816);
   U22205 : AOI22_X1 port map( A1 => n26879, A2 => n9417, B1 => n26873, B2 => 
                           n19319, ZN => n23817);
   U22206 : OAI221_X1 port map( B1 => n20764, B2 => n26789, C1 => n21992, C2 =>
                           n26783, A => n23825, ZN => n23824);
   U22207 : AOI22_X1 port map( A1 => n26777, A2 => n19334, B1 => n26775, B2 => 
                           n4210, ZN => n23825);
   U22208 : OAI221_X1 port map( B1 => n21351, B2 => n26891, C1 => n21631, C2 =>
                           n26885, A => n23799, ZN => n23798);
   U22209 : AOI22_X1 port map( A1 => n26879, A2 => n9414, B1 => n26873, B2 => 
                           n19302, ZN => n23799);
   U22210 : OAI221_X1 port map( B1 => n20763, B2 => n26789, C1 => n21991, C2 =>
                           n26783, A => n23807, ZN => n23806);
   U22211 : AOI22_X1 port map( A1 => n26777, A2 => n19317, B1 => n26775, B2 => 
                           n4208, ZN => n23807);
   U22212 : OAI221_X1 port map( B1 => n21350, B2 => n26891, C1 => n21630, C2 =>
                           n26885, A => n23781, ZN => n23780);
   U22213 : AOI22_X1 port map( A1 => n26879, A2 => n9411, B1 => n26873, B2 => 
                           n19285, ZN => n23781);
   U22214 : OAI221_X1 port map( B1 => n20762, B2 => n26789, C1 => n21990, C2 =>
                           n26783, A => n23789, ZN => n23788);
   U22215 : AOI22_X1 port map( A1 => n26777, A2 => n19300, B1 => n26774, B2 => 
                           n4206, ZN => n23789);
   U22216 : OAI221_X1 port map( B1 => n21349, B2 => n26891, C1 => n21629, C2 =>
                           n26885, A => n23763, ZN => n23762);
   U22217 : AOI22_X1 port map( A1 => n26879, A2 => n9408, B1 => n26873, B2 => 
                           n19268, ZN => n23763);
   U22218 : OAI221_X1 port map( B1 => n20761, B2 => n26789, C1 => n21989, C2 =>
                           n26783, A => n23771, ZN => n23770);
   U22219 : AOI22_X1 port map( A1 => n26777, A2 => n19283, B1 => n26774, B2 => 
                           n4204, ZN => n23771);
   U22220 : OAI221_X1 port map( B1 => n21348, B2 => n26891, C1 => n21628, C2 =>
                           n26885, A => n23745, ZN => n23744);
   U22221 : AOI22_X1 port map( A1 => n26879, A2 => n9405, B1 => n26873, B2 => 
                           n19251, ZN => n23745);
   U22222 : OAI221_X1 port map( B1 => n20760, B2 => n26789, C1 => n21988, C2 =>
                           n26783, A => n23753, ZN => n23752);
   U22223 : AOI22_X1 port map( A1 => n26777, A2 => n19266, B1 => n26774, B2 => 
                           n4202, ZN => n23753);
   U22224 : OAI221_X1 port map( B1 => n22559, B2 => n26643, C1 => n21227, C2 =>
                           n26637, A => n24927, ZN => n24924);
   U22225 : AOI22_X1 port map( A1 => n26631, A2 => n25760, B1 => n26625, B2 => 
                           n8603, ZN => n24927);
   U22226 : OAI221_X1 port map( B1 => n22679, B2 => n26520, C1 => n22487, C2 =>
                           n26514, A => n24935, ZN => n24932);
   U22227 : AOI22_X1 port map( A1 => n26508, A2 => n26219, B1 => n26502, B2 => 
                           n26339, ZN => n24935);
   U22228 : OAI221_X1 port map( B1 => n22558, B2 => n26643, C1 => n21226, C2 =>
                           n26637, A => n24909, ZN => n24906);
   U22229 : AOI22_X1 port map( A1 => n26631, A2 => n25765, B1 => n26625, B2 => 
                           n8600, ZN => n24909);
   U22230 : OAI221_X1 port map( B1 => n22678, B2 => n26520, C1 => n22486, C2 =>
                           n26514, A => n24917, ZN => n24914);
   U22231 : AOI22_X1 port map( A1 => n26508, A2 => n26220, B1 => n26502, B2 => 
                           n26340, ZN => n24917);
   U22232 : OAI221_X1 port map( B1 => n22557, B2 => n26643, C1 => n21225, C2 =>
                           n26637, A => n24891, ZN => n24888);
   U22233 : AOI22_X1 port map( A1 => n26631, A2 => n25770, B1 => n26625, B2 => 
                           n8597, ZN => n24891);
   U22234 : OAI221_X1 port map( B1 => n22677, B2 => n26520, C1 => n22485, C2 =>
                           n26514, A => n24899, ZN => n24896);
   U22235 : AOI22_X1 port map( A1 => n26508, A2 => n26221, B1 => n26502, B2 => 
                           n26341, ZN => n24899);
   U22236 : OAI221_X1 port map( B1 => n22556, B2 => n26643, C1 => n21224, C2 =>
                           n26637, A => n24873, ZN => n24870);
   U22237 : AOI22_X1 port map( A1 => n26631, A2 => n25775, B1 => n26625, B2 => 
                           n8594, ZN => n24873);
   U22238 : OAI221_X1 port map( B1 => n22676, B2 => n26520, C1 => n22484, C2 =>
                           n26514, A => n24881, ZN => n24878);
   U22239 : AOI22_X1 port map( A1 => n26508, A2 => n26222, B1 => n26502, B2 => 
                           n26342, ZN => n24881);
   U22240 : OAI221_X1 port map( B1 => n22555, B2 => n26643, C1 => n21223, C2 =>
                           n26637, A => n24855, ZN => n24852);
   U22241 : AOI22_X1 port map( A1 => n26631, A2 => n25780, B1 => n26625, B2 => 
                           n8591, ZN => n24855);
   U22242 : OAI221_X1 port map( B1 => n22675, B2 => n26520, C1 => n22483, C2 =>
                           n26514, A => n24863, ZN => n24860);
   U22243 : AOI22_X1 port map( A1 => n26508, A2 => n26223, B1 => n26502, B2 => 
                           n26343, ZN => n24863);
   U22244 : OAI221_X1 port map( B1 => n22554, B2 => n26643, C1 => n21222, C2 =>
                           n26637, A => n24837, ZN => n24834);
   U22245 : AOI22_X1 port map( A1 => n26631, A2 => n25785, B1 => n26625, B2 => 
                           n8588, ZN => n24837);
   U22246 : OAI221_X1 port map( B1 => n22674, B2 => n26520, C1 => n22482, C2 =>
                           n26514, A => n24845, ZN => n24842);
   U22247 : AOI22_X1 port map( A1 => n26508, A2 => n26224, B1 => n26502, B2 => 
                           n26344, ZN => n24845);
   U22248 : OAI221_X1 port map( B1 => n22553, B2 => n26643, C1 => n21221, C2 =>
                           n26637, A => n24819, ZN => n24816);
   U22249 : AOI22_X1 port map( A1 => n26631, A2 => n25790, B1 => n26625, B2 => 
                           n8585, ZN => n24819);
   U22250 : OAI221_X1 port map( B1 => n22673, B2 => n26520, C1 => n22481, C2 =>
                           n26514, A => n24827, ZN => n24824);
   U22251 : AOI22_X1 port map( A1 => n26508, A2 => n26225, B1 => n26502, B2 => 
                           n26345, ZN => n24827);
   U22252 : OAI221_X1 port map( B1 => n22552, B2 => n26643, C1 => n21220, C2 =>
                           n26637, A => n24801, ZN => n24798);
   U22253 : AOI22_X1 port map( A1 => n26631, A2 => n25795, B1 => n26625, B2 => 
                           n8582, ZN => n24801);
   U22254 : OAI221_X1 port map( B1 => n22672, B2 => n26520, C1 => n22480, C2 =>
                           n26514, A => n24809, ZN => n24806);
   U22255 : AOI22_X1 port map( A1 => n26508, A2 => n26226, B1 => n26502, B2 => 
                           n26346, ZN => n24809);
   U22256 : OAI221_X1 port map( B1 => n22551, B2 => n26643, C1 => n21219, C2 =>
                           n26637, A => n24783, ZN => n24780);
   U22257 : AOI22_X1 port map( A1 => n26631, A2 => n25800, B1 => n26625, B2 => 
                           n8579, ZN => n24783);
   U22258 : OAI221_X1 port map( B1 => n22671, B2 => n26520, C1 => n22479, C2 =>
                           n26514, A => n24791, ZN => n24788);
   U22259 : AOI22_X1 port map( A1 => n26508, A2 => n26227, B1 => n26502, B2 => 
                           n26347, ZN => n24791);
   U22260 : OAI221_X1 port map( B1 => n22550, B2 => n26643, C1 => n21218, C2 =>
                           n26637, A => n24765, ZN => n24762);
   U22261 : AOI22_X1 port map( A1 => n26631, A2 => n25805, B1 => n26625, B2 => 
                           n8576, ZN => n24765);
   U22262 : OAI221_X1 port map( B1 => n22670, B2 => n26520, C1 => n22478, C2 =>
                           n26514, A => n24773, ZN => n24770);
   U22263 : AOI22_X1 port map( A1 => n26508, A2 => n26228, B1 => n26502, B2 => 
                           n26348, ZN => n24773);
   U22264 : OAI221_X1 port map( B1 => n22549, B2 => n26643, C1 => n21217, C2 =>
                           n26637, A => n24747, ZN => n24744);
   U22265 : AOI22_X1 port map( A1 => n26631, A2 => n25810, B1 => n26625, B2 => 
                           n8573, ZN => n24747);
   U22266 : OAI221_X1 port map( B1 => n22669, B2 => n26520, C1 => n22477, C2 =>
                           n26514, A => n24755, ZN => n24752);
   U22267 : AOI22_X1 port map( A1 => n26508, A2 => n26229, B1 => n26502, B2 => 
                           n26349, ZN => n24755);
   U22268 : OAI221_X1 port map( B1 => n22548, B2 => n26643, C1 => n21216, C2 =>
                           n26637, A => n24729, ZN => n24726);
   U22269 : AOI22_X1 port map( A1 => n26631, A2 => n25815, B1 => n26625, B2 => 
                           n8570, ZN => n24729);
   U22270 : OAI221_X1 port map( B1 => n22668, B2 => n26520, C1 => n22476, C2 =>
                           n26514, A => n24737, ZN => n24734);
   U22271 : AOI22_X1 port map( A1 => n26508, A2 => n26230, B1 => n26502, B2 => 
                           n26350, ZN => n24737);
   U22272 : OAI221_X1 port map( B1 => n22547, B2 => n26644, C1 => n21215, C2 =>
                           n26638, A => n24711, ZN => n24708);
   U22273 : AOI22_X1 port map( A1 => n26632, A2 => n25820, B1 => n26626, B2 => 
                           n8567, ZN => n24711);
   U22274 : OAI221_X1 port map( B1 => n22667, B2 => n26521, C1 => n22475, C2 =>
                           n26515, A => n24719, ZN => n24716);
   U22275 : AOI22_X1 port map( A1 => n26509, A2 => n26231, B1 => n26503, B2 => 
                           n26351, ZN => n24719);
   U22276 : OAI221_X1 port map( B1 => n22546, B2 => n26644, C1 => n21214, C2 =>
                           n26638, A => n24693, ZN => n24690);
   U22277 : AOI22_X1 port map( A1 => n26632, A2 => n25825, B1 => n26626, B2 => 
                           n8564, ZN => n24693);
   U22278 : OAI221_X1 port map( B1 => n22666, B2 => n26521, C1 => n22474, C2 =>
                           n26515, A => n24701, ZN => n24698);
   U22279 : AOI22_X1 port map( A1 => n26509, A2 => n26232, B1 => n26503, B2 => 
                           n26352, ZN => n24701);
   U22280 : OAI221_X1 port map( B1 => n22545, B2 => n26644, C1 => n21213, C2 =>
                           n26638, A => n24675, ZN => n24672);
   U22281 : AOI22_X1 port map( A1 => n26632, A2 => n25830, B1 => n26626, B2 => 
                           n8561, ZN => n24675);
   U22282 : OAI221_X1 port map( B1 => n22665, B2 => n26521, C1 => n22473, C2 =>
                           n26515, A => n24683, ZN => n24680);
   U22283 : AOI22_X1 port map( A1 => n26509, A2 => n26233, B1 => n26503, B2 => 
                           n26353, ZN => n24683);
   U22284 : OAI221_X1 port map( B1 => n22544, B2 => n26644, C1 => n21212, C2 =>
                           n26638, A => n24657, ZN => n24654);
   U22285 : AOI22_X1 port map( A1 => n26632, A2 => n25835, B1 => n26626, B2 => 
                           n8558, ZN => n24657);
   U22286 : OAI221_X1 port map( B1 => n22664, B2 => n26521, C1 => n22472, C2 =>
                           n26515, A => n24665, ZN => n24662);
   U22287 : AOI22_X1 port map( A1 => n26509, A2 => n26234, B1 => n26503, B2 => 
                           n26354, ZN => n24665);
   U22288 : OAI221_X1 port map( B1 => n22543, B2 => n26644, C1 => n21211, C2 =>
                           n26638, A => n24639, ZN => n24636);
   U22289 : AOI22_X1 port map( A1 => n26632, A2 => n25840, B1 => n26626, B2 => 
                           n8555, ZN => n24639);
   U22290 : OAI221_X1 port map( B1 => n22663, B2 => n26521, C1 => n22471, C2 =>
                           n26515, A => n24647, ZN => n24644);
   U22291 : AOI22_X1 port map( A1 => n26509, A2 => n26235, B1 => n26503, B2 => 
                           n26355, ZN => n24647);
   U22292 : OAI221_X1 port map( B1 => n22542, B2 => n26644, C1 => n21210, C2 =>
                           n26638, A => n24621, ZN => n24618);
   U22293 : AOI22_X1 port map( A1 => n26632, A2 => n25845, B1 => n26626, B2 => 
                           n8552, ZN => n24621);
   U22294 : OAI221_X1 port map( B1 => n22662, B2 => n26521, C1 => n22470, C2 =>
                           n26515, A => n24629, ZN => n24626);
   U22295 : AOI22_X1 port map( A1 => n26509, A2 => n26236, B1 => n26503, B2 => 
                           n26356, ZN => n24629);
   U22296 : OAI221_X1 port map( B1 => n22541, B2 => n26644, C1 => n21209, C2 =>
                           n26638, A => n24603, ZN => n24600);
   U22297 : AOI22_X1 port map( A1 => n26632, A2 => n25850, B1 => n26626, B2 => 
                           n8549, ZN => n24603);
   U22298 : OAI221_X1 port map( B1 => n22661, B2 => n26521, C1 => n22469, C2 =>
                           n26515, A => n24611, ZN => n24608);
   U22299 : AOI22_X1 port map( A1 => n26509, A2 => n26237, B1 => n26503, B2 => 
                           n26357, ZN => n24611);
   U22300 : OAI221_X1 port map( B1 => n22540, B2 => n26644, C1 => n21208, C2 =>
                           n26638, A => n24585, ZN => n24582);
   U22301 : AOI22_X1 port map( A1 => n26632, A2 => n25855, B1 => n26626, B2 => 
                           n8546, ZN => n24585);
   U22302 : OAI221_X1 port map( B1 => n22660, B2 => n26521, C1 => n22468, C2 =>
                           n26515, A => n24593, ZN => n24590);
   U22303 : AOI22_X1 port map( A1 => n26509, A2 => n26238, B1 => n26503, B2 => 
                           n26358, ZN => n24593);
   U22304 : OAI221_X1 port map( B1 => n22539, B2 => n26644, C1 => n21207, C2 =>
                           n26638, A => n24567, ZN => n24564);
   U22305 : AOI22_X1 port map( A1 => n26632, A2 => n25860, B1 => n26626, B2 => 
                           n8543, ZN => n24567);
   U22306 : OAI221_X1 port map( B1 => n22659, B2 => n26521, C1 => n22467, C2 =>
                           n26515, A => n24575, ZN => n24572);
   U22307 : AOI22_X1 port map( A1 => n26509, A2 => n26239, B1 => n26503, B2 => 
                           n26359, ZN => n24575);
   U22308 : OAI221_X1 port map( B1 => n22538, B2 => n26644, C1 => n21206, C2 =>
                           n26638, A => n24549, ZN => n24546);
   U22309 : AOI22_X1 port map( A1 => n26632, A2 => n25865, B1 => n26626, B2 => 
                           n8540, ZN => n24549);
   U22310 : OAI221_X1 port map( B1 => n22658, B2 => n26521, C1 => n22466, C2 =>
                           n26515, A => n24557, ZN => n24554);
   U22311 : AOI22_X1 port map( A1 => n26509, A2 => n26240, B1 => n26503, B2 => 
                           n26360, ZN => n24557);
   U22312 : OAI221_X1 port map( B1 => n22537, B2 => n26644, C1 => n21205, C2 =>
                           n26638, A => n24531, ZN => n24528);
   U22313 : AOI22_X1 port map( A1 => n26632, A2 => n25870, B1 => n26626, B2 => 
                           n8537, ZN => n24531);
   U22314 : OAI221_X1 port map( B1 => n22657, B2 => n26521, C1 => n22465, C2 =>
                           n26515, A => n24539, ZN => n24536);
   U22315 : AOI22_X1 port map( A1 => n26509, A2 => n26241, B1 => n26503, B2 => 
                           n26361, ZN => n24539);
   U22316 : OAI221_X1 port map( B1 => n22536, B2 => n26644, C1 => n21204, C2 =>
                           n26638, A => n24513, ZN => n24510);
   U22317 : AOI22_X1 port map( A1 => n26632, A2 => n25875, B1 => n26626, B2 => 
                           n8534, ZN => n24513);
   U22318 : OAI221_X1 port map( B1 => n22656, B2 => n26521, C1 => n22464, C2 =>
                           n26515, A => n24521, ZN => n24518);
   U22319 : AOI22_X1 port map( A1 => n26509, A2 => n26242, B1 => n26503, B2 => 
                           n26362, ZN => n24521);
   U22320 : OAI221_X1 port map( B1 => n22535, B2 => n26645, C1 => n21203, C2 =>
                           n26639, A => n24495, ZN => n24492);
   U22321 : AOI22_X1 port map( A1 => n26633, A2 => n25880, B1 => n26627, B2 => 
                           n8531, ZN => n24495);
   U22322 : OAI221_X1 port map( B1 => n22655, B2 => n26522, C1 => n22463, C2 =>
                           n26516, A => n24503, ZN => n24500);
   U22323 : AOI22_X1 port map( A1 => n26510, A2 => n26243, B1 => n26504, B2 => 
                           n26363, ZN => n24503);
   U22324 : OAI221_X1 port map( B1 => n22534, B2 => n26645, C1 => n21202, C2 =>
                           n26639, A => n24477, ZN => n24474);
   U22325 : AOI22_X1 port map( A1 => n26633, A2 => n25885, B1 => n26627, B2 => 
                           n8528, ZN => n24477);
   U22326 : OAI221_X1 port map( B1 => n22654, B2 => n26522, C1 => n22462, C2 =>
                           n26516, A => n24485, ZN => n24482);
   U22327 : AOI22_X1 port map( A1 => n26510, A2 => n26244, B1 => n26504, B2 => 
                           n26364, ZN => n24485);
   U22328 : OAI221_X1 port map( B1 => n22533, B2 => n26645, C1 => n21201, C2 =>
                           n26639, A => n24459, ZN => n24456);
   U22329 : AOI22_X1 port map( A1 => n26633, A2 => n25890, B1 => n26627, B2 => 
                           n8525, ZN => n24459);
   U22330 : OAI221_X1 port map( B1 => n22653, B2 => n26522, C1 => n22461, C2 =>
                           n26516, A => n24467, ZN => n24464);
   U22331 : AOI22_X1 port map( A1 => n26510, A2 => n26245, B1 => n26504, B2 => 
                           n26365, ZN => n24467);
   U22332 : OAI221_X1 port map( B1 => n22532, B2 => n26645, C1 => n21200, C2 =>
                           n26639, A => n24441, ZN => n24438);
   U22333 : AOI22_X1 port map( A1 => n26633, A2 => n25895, B1 => n26627, B2 => 
                           n8522, ZN => n24441);
   U22334 : OAI221_X1 port map( B1 => n22652, B2 => n26522, C1 => n22460, C2 =>
                           n26516, A => n24449, ZN => n24446);
   U22335 : AOI22_X1 port map( A1 => n26510, A2 => n26246, B1 => n26504, B2 => 
                           n26366, ZN => n24449);
   U22336 : OAI221_X1 port map( B1 => n22531, B2 => n26645, C1 => n21199, C2 =>
                           n26639, A => n24423, ZN => n24420);
   U22337 : AOI22_X1 port map( A1 => n26633, A2 => n25900, B1 => n26627, B2 => 
                           n8519, ZN => n24423);
   U22338 : OAI221_X1 port map( B1 => n22651, B2 => n26522, C1 => n22459, C2 =>
                           n26516, A => n24431, ZN => n24428);
   U22339 : AOI22_X1 port map( A1 => n26510, A2 => n26247, B1 => n26504, B2 => 
                           n26367, ZN => n24431);
   U22340 : OAI221_X1 port map( B1 => n22530, B2 => n26645, C1 => n21198, C2 =>
                           n26639, A => n24405, ZN => n24402);
   U22341 : AOI22_X1 port map( A1 => n26633, A2 => n25905, B1 => n26627, B2 => 
                           n8516, ZN => n24405);
   U22342 : OAI221_X1 port map( B1 => n22650, B2 => n26522, C1 => n22458, C2 =>
                           n26516, A => n24413, ZN => n24410);
   U22343 : AOI22_X1 port map( A1 => n26510, A2 => n26248, B1 => n26504, B2 => 
                           n26368, ZN => n24413);
   U22344 : OAI221_X1 port map( B1 => n22529, B2 => n26645, C1 => n21197, C2 =>
                           n26639, A => n24387, ZN => n24384);
   U22345 : AOI22_X1 port map( A1 => n26633, A2 => n25910, B1 => n26627, B2 => 
                           n8513, ZN => n24387);
   U22346 : OAI221_X1 port map( B1 => n22649, B2 => n26522, C1 => n22457, C2 =>
                           n26516, A => n24395, ZN => n24392);
   U22347 : AOI22_X1 port map( A1 => n26510, A2 => n26249, B1 => n26504, B2 => 
                           n26369, ZN => n24395);
   U22348 : OAI221_X1 port map( B1 => n22528, B2 => n26645, C1 => n21196, C2 =>
                           n26639, A => n24369, ZN => n24366);
   U22349 : AOI22_X1 port map( A1 => n26633, A2 => n25915, B1 => n26627, B2 => 
                           n8510, ZN => n24369);
   U22350 : OAI221_X1 port map( B1 => n22648, B2 => n26522, C1 => n22456, C2 =>
                           n26516, A => n24377, ZN => n24374);
   U22351 : AOI22_X1 port map( A1 => n26510, A2 => n26250, B1 => n26504, B2 => 
                           n26370, ZN => n24377);
   U22352 : OAI221_X1 port map( B1 => n22527, B2 => n26645, C1 => n21195, C2 =>
                           n26639, A => n24351, ZN => n24348);
   U22353 : AOI22_X1 port map( A1 => n26633, A2 => n25920, B1 => n26627, B2 => 
                           n8507, ZN => n24351);
   U22354 : OAI221_X1 port map( B1 => n22647, B2 => n26522, C1 => n22455, C2 =>
                           n26516, A => n24359, ZN => n24356);
   U22355 : AOI22_X1 port map( A1 => n26510, A2 => n26251, B1 => n26504, B2 => 
                           n26371, ZN => n24359);
   U22356 : OAI221_X1 port map( B1 => n22526, B2 => n26645, C1 => n21194, C2 =>
                           n26639, A => n24333, ZN => n24330);
   U22357 : AOI22_X1 port map( A1 => n26633, A2 => n25925, B1 => n26627, B2 => 
                           n8504, ZN => n24333);
   U22358 : OAI221_X1 port map( B1 => n22646, B2 => n26522, C1 => n22454, C2 =>
                           n26516, A => n24341, ZN => n24338);
   U22359 : AOI22_X1 port map( A1 => n26510, A2 => n26252, B1 => n26504, B2 => 
                           n26372, ZN => n24341);
   U22360 : OAI221_X1 port map( B1 => n22525, B2 => n26645, C1 => n21193, C2 =>
                           n26639, A => n24315, ZN => n24312);
   U22361 : AOI22_X1 port map( A1 => n26633, A2 => n25930, B1 => n26627, B2 => 
                           n8501, ZN => n24315);
   U22362 : OAI221_X1 port map( B1 => n22645, B2 => n26522, C1 => n22453, C2 =>
                           n26516, A => n24323, ZN => n24320);
   U22363 : AOI22_X1 port map( A1 => n26510, A2 => n26253, B1 => n26504, B2 => 
                           n26373, ZN => n24323);
   U22364 : OAI221_X1 port map( B1 => n22524, B2 => n26645, C1 => n21192, C2 =>
                           n26639, A => n24297, ZN => n24294);
   U22365 : AOI22_X1 port map( A1 => n26633, A2 => n25935, B1 => n26627, B2 => 
                           n8498, ZN => n24297);
   U22366 : OAI221_X1 port map( B1 => n22644, B2 => n26522, C1 => n22452, C2 =>
                           n26516, A => n24305, ZN => n24302);
   U22367 : AOI22_X1 port map( A1 => n26510, A2 => n26254, B1 => n26504, B2 => 
                           n26374, ZN => n24305);
   U22368 : OAI221_X1 port map( B1 => n22523, B2 => n26646, C1 => n21191, C2 =>
                           n26640, A => n24279, ZN => n24276);
   U22369 : AOI22_X1 port map( A1 => n26634, A2 => n25940, B1 => n26628, B2 => 
                           n8495, ZN => n24279);
   U22370 : OAI221_X1 port map( B1 => n22643, B2 => n26523, C1 => n22451, C2 =>
                           n26517, A => n24287, ZN => n24284);
   U22371 : AOI22_X1 port map( A1 => n26511, A2 => n26255, B1 => n26505, B2 => 
                           n26375, ZN => n24287);
   U22372 : OAI221_X1 port map( B1 => n22522, B2 => n26646, C1 => n21190, C2 =>
                           n26640, A => n24261, ZN => n24258);
   U22373 : AOI22_X1 port map( A1 => n26634, A2 => n25945, B1 => n26628, B2 => 
                           n8492, ZN => n24261);
   U22374 : OAI221_X1 port map( B1 => n22642, B2 => n26523, C1 => n22450, C2 =>
                           n26517, A => n24269, ZN => n24266);
   U22375 : AOI22_X1 port map( A1 => n26511, A2 => n26256, B1 => n26505, B2 => 
                           n26376, ZN => n24269);
   U22376 : OAI221_X1 port map( B1 => n22521, B2 => n26646, C1 => n21189, C2 =>
                           n26640, A => n24243, ZN => n24240);
   U22377 : AOI22_X1 port map( A1 => n26634, A2 => n25950, B1 => n26628, B2 => 
                           n8489, ZN => n24243);
   U22378 : OAI221_X1 port map( B1 => n22641, B2 => n26523, C1 => n22449, C2 =>
                           n26517, A => n24251, ZN => n24248);
   U22379 : AOI22_X1 port map( A1 => n26511, A2 => n26257, B1 => n26505, B2 => 
                           n26377, ZN => n24251);
   U22380 : OAI221_X1 port map( B1 => n22520, B2 => n26646, C1 => n21188, C2 =>
                           n26640, A => n24225, ZN => n24222);
   U22381 : AOI22_X1 port map( A1 => n26634, A2 => n25955, B1 => n26628, B2 => 
                           n8486, ZN => n24225);
   U22382 : OAI221_X1 port map( B1 => n22640, B2 => n26523, C1 => n22448, C2 =>
                           n26517, A => n24233, ZN => n24230);
   U22383 : AOI22_X1 port map( A1 => n26511, A2 => n26258, B1 => n26505, B2 => 
                           n26378, ZN => n24233);
   U22384 : OAI221_X1 port map( B1 => n22519, B2 => n26646, C1 => n21187, C2 =>
                           n26640, A => n24207, ZN => n24204);
   U22385 : AOI22_X1 port map( A1 => n26634, A2 => n25960, B1 => n26628, B2 => 
                           n8483, ZN => n24207);
   U22386 : OAI221_X1 port map( B1 => n22639, B2 => n26523, C1 => n22447, C2 =>
                           n26517, A => n24215, ZN => n24212);
   U22387 : AOI22_X1 port map( A1 => n26511, A2 => n26259, B1 => n26505, B2 => 
                           n26379, ZN => n24215);
   U22388 : OAI221_X1 port map( B1 => n22518, B2 => n26646, C1 => n21186, C2 =>
                           n26640, A => n24189, ZN => n24186);
   U22389 : AOI22_X1 port map( A1 => n26634, A2 => n25965, B1 => n26628, B2 => 
                           n8480, ZN => n24189);
   U22390 : OAI221_X1 port map( B1 => n22638, B2 => n26523, C1 => n22446, C2 =>
                           n26517, A => n24197, ZN => n24194);
   U22391 : AOI22_X1 port map( A1 => n26511, A2 => n26260, B1 => n26505, B2 => 
                           n26380, ZN => n24197);
   U22392 : OAI221_X1 port map( B1 => n22517, B2 => n26646, C1 => n21185, C2 =>
                           n26640, A => n24171, ZN => n24168);
   U22393 : AOI22_X1 port map( A1 => n26634, A2 => n25970, B1 => n26628, B2 => 
                           n8477, ZN => n24171);
   U22394 : OAI221_X1 port map( B1 => n22637, B2 => n26523, C1 => n22445, C2 =>
                           n26517, A => n24179, ZN => n24176);
   U22395 : AOI22_X1 port map( A1 => n26511, A2 => n26261, B1 => n26505, B2 => 
                           n26381, ZN => n24179);
   U22396 : OAI221_X1 port map( B1 => n22516, B2 => n26646, C1 => n21184, C2 =>
                           n26640, A => n24153, ZN => n24150);
   U22397 : AOI22_X1 port map( A1 => n26634, A2 => n25975, B1 => n26628, B2 => 
                           n8474, ZN => n24153);
   U22398 : OAI221_X1 port map( B1 => n22636, B2 => n26523, C1 => n22444, C2 =>
                           n26517, A => n24161, ZN => n24158);
   U22399 : AOI22_X1 port map( A1 => n26511, A2 => n26262, B1 => n26505, B2 => 
                           n26382, ZN => n24161);
   U22400 : OAI221_X1 port map( B1 => n22515, B2 => n26646, C1 => n21183, C2 =>
                           n26640, A => n24135, ZN => n24132);
   U22401 : AOI22_X1 port map( A1 => n26634, A2 => n25980, B1 => n26628, B2 => 
                           n8471, ZN => n24135);
   U22402 : OAI221_X1 port map( B1 => n22635, B2 => n26523, C1 => n22443, C2 =>
                           n26517, A => n24143, ZN => n24140);
   U22403 : AOI22_X1 port map( A1 => n26511, A2 => n26263, B1 => n26505, B2 => 
                           n26383, ZN => n24143);
   U22404 : OAI221_X1 port map( B1 => n22514, B2 => n26646, C1 => n21182, C2 =>
                           n26640, A => n24117, ZN => n24114);
   U22405 : AOI22_X1 port map( A1 => n26634, A2 => n25985, B1 => n26628, B2 => 
                           n8468, ZN => n24117);
   U22406 : OAI221_X1 port map( B1 => n22634, B2 => n26523, C1 => n22442, C2 =>
                           n26517, A => n24125, ZN => n24122);
   U22407 : AOI22_X1 port map( A1 => n26511, A2 => n26264, B1 => n26505, B2 => 
                           n26384, ZN => n24125);
   U22408 : OAI221_X1 port map( B1 => n22513, B2 => n26646, C1 => n21181, C2 =>
                           n26640, A => n24099, ZN => n24096);
   U22409 : AOI22_X1 port map( A1 => n26634, A2 => n25990, B1 => n26628, B2 => 
                           n8465, ZN => n24099);
   U22410 : OAI221_X1 port map( B1 => n22633, B2 => n26523, C1 => n22441, C2 =>
                           n26517, A => n24107, ZN => n24104);
   U22411 : AOI22_X1 port map( A1 => n26511, A2 => n26265, B1 => n26505, B2 => 
                           n26385, ZN => n24107);
   U22412 : OAI221_X1 port map( B1 => n22512, B2 => n26646, C1 => n21180, C2 =>
                           n26640, A => n24081, ZN => n24078);
   U22413 : AOI22_X1 port map( A1 => n26634, A2 => n25995, B1 => n26628, B2 => 
                           n8462, ZN => n24081);
   U22414 : OAI221_X1 port map( B1 => n22632, B2 => n26523, C1 => n22440, C2 =>
                           n26517, A => n24089, ZN => n24086);
   U22415 : AOI22_X1 port map( A1 => n26511, A2 => n26266, B1 => n26505, B2 => 
                           n26386, ZN => n24089);
   U22416 : OAI221_X1 port map( B1 => n22559, B2 => n26868, C1 => n21227, C2 =>
                           n26862, A => n23728, ZN => n23725);
   U22417 : AOI22_X1 port map( A1 => n26856, A2 => n25760, B1 => n26850, B2 => 
                           n8603, ZN => n23728);
   U22418 : OAI221_X1 port map( B1 => n22679, B2 => n26745, C1 => n22487, C2 =>
                           n26739, A => n23736, ZN => n23733);
   U22419 : AOI22_X1 port map( A1 => n26733, A2 => n26219, B1 => n26727, B2 => 
                           n26339, ZN => n23736);
   U22420 : OAI221_X1 port map( B1 => n22558, B2 => n26868, C1 => n21226, C2 =>
                           n26862, A => n23710, ZN => n23707);
   U22421 : AOI22_X1 port map( A1 => n26856, A2 => n25765, B1 => n26850, B2 => 
                           n8600, ZN => n23710);
   U22422 : OAI221_X1 port map( B1 => n22678, B2 => n26745, C1 => n22486, C2 =>
                           n26739, A => n23718, ZN => n23715);
   U22423 : AOI22_X1 port map( A1 => n26733, A2 => n26220, B1 => n26727, B2 => 
                           n26340, ZN => n23718);
   U22424 : OAI221_X1 port map( B1 => n22557, B2 => n26868, C1 => n21225, C2 =>
                           n26862, A => n23692, ZN => n23689);
   U22425 : AOI22_X1 port map( A1 => n26856, A2 => n25770, B1 => n26850, B2 => 
                           n8597, ZN => n23692);
   U22426 : OAI221_X1 port map( B1 => n22677, B2 => n26745, C1 => n22485, C2 =>
                           n26739, A => n23700, ZN => n23697);
   U22427 : AOI22_X1 port map( A1 => n26733, A2 => n26221, B1 => n26727, B2 => 
                           n26341, ZN => n23700);
   U22428 : OAI221_X1 port map( B1 => n22556, B2 => n26868, C1 => n21224, C2 =>
                           n26862, A => n23674, ZN => n23671);
   U22429 : AOI22_X1 port map( A1 => n26856, A2 => n25775, B1 => n26850, B2 => 
                           n8594, ZN => n23674);
   U22430 : OAI221_X1 port map( B1 => n22676, B2 => n26745, C1 => n22484, C2 =>
                           n26739, A => n23682, ZN => n23679);
   U22431 : AOI22_X1 port map( A1 => n26733, A2 => n26222, B1 => n26727, B2 => 
                           n26342, ZN => n23682);
   U22432 : OAI221_X1 port map( B1 => n22555, B2 => n26868, C1 => n21223, C2 =>
                           n26862, A => n23656, ZN => n23653);
   U22433 : AOI22_X1 port map( A1 => n26856, A2 => n25780, B1 => n26850, B2 => 
                           n8591, ZN => n23656);
   U22434 : OAI221_X1 port map( B1 => n22675, B2 => n26745, C1 => n22483, C2 =>
                           n26739, A => n23664, ZN => n23661);
   U22435 : AOI22_X1 port map( A1 => n26733, A2 => n26223, B1 => n26727, B2 => 
                           n26343, ZN => n23664);
   U22436 : OAI221_X1 port map( B1 => n22554, B2 => n26868, C1 => n21222, C2 =>
                           n26862, A => n23638, ZN => n23635);
   U22437 : AOI22_X1 port map( A1 => n26856, A2 => n25785, B1 => n26850, B2 => 
                           n8588, ZN => n23638);
   U22438 : OAI221_X1 port map( B1 => n22674, B2 => n26745, C1 => n22482, C2 =>
                           n26739, A => n23646, ZN => n23643);
   U22439 : AOI22_X1 port map( A1 => n26733, A2 => n26224, B1 => n26727, B2 => 
                           n26344, ZN => n23646);
   U22440 : OAI221_X1 port map( B1 => n22553, B2 => n26868, C1 => n21221, C2 =>
                           n26862, A => n23620, ZN => n23617);
   U22441 : AOI22_X1 port map( A1 => n26856, A2 => n25790, B1 => n26850, B2 => 
                           n8585, ZN => n23620);
   U22442 : OAI221_X1 port map( B1 => n22673, B2 => n26745, C1 => n22481, C2 =>
                           n26739, A => n23628, ZN => n23625);
   U22443 : AOI22_X1 port map( A1 => n26733, A2 => n26225, B1 => n26727, B2 => 
                           n26345, ZN => n23628);
   U22444 : OAI221_X1 port map( B1 => n22552, B2 => n26868, C1 => n21220, C2 =>
                           n26862, A => n23602, ZN => n23599);
   U22445 : AOI22_X1 port map( A1 => n26856, A2 => n25795, B1 => n26850, B2 => 
                           n8582, ZN => n23602);
   U22446 : OAI221_X1 port map( B1 => n22672, B2 => n26745, C1 => n22480, C2 =>
                           n26739, A => n23610, ZN => n23607);
   U22447 : AOI22_X1 port map( A1 => n26733, A2 => n26226, B1 => n26727, B2 => 
                           n26346, ZN => n23610);
   U22448 : OAI221_X1 port map( B1 => n22551, B2 => n26868, C1 => n21219, C2 =>
                           n26862, A => n23584, ZN => n23581);
   U22449 : AOI22_X1 port map( A1 => n26856, A2 => n25800, B1 => n26850, B2 => 
                           n8579, ZN => n23584);
   U22450 : OAI221_X1 port map( B1 => n22671, B2 => n26745, C1 => n22479, C2 =>
                           n26739, A => n23592, ZN => n23589);
   U22451 : AOI22_X1 port map( A1 => n26733, A2 => n26227, B1 => n26727, B2 => 
                           n26347, ZN => n23592);
   U22452 : OAI221_X1 port map( B1 => n22550, B2 => n26868, C1 => n21218, C2 =>
                           n26862, A => n23566, ZN => n23563);
   U22453 : AOI22_X1 port map( A1 => n26856, A2 => n25805, B1 => n26850, B2 => 
                           n8576, ZN => n23566);
   U22454 : OAI221_X1 port map( B1 => n22670, B2 => n26745, C1 => n22478, C2 =>
                           n26739, A => n23574, ZN => n23571);
   U22455 : AOI22_X1 port map( A1 => n26733, A2 => n26228, B1 => n26727, B2 => 
                           n26348, ZN => n23574);
   U22456 : OAI221_X1 port map( B1 => n22549, B2 => n26868, C1 => n21217, C2 =>
                           n26862, A => n23548, ZN => n23545);
   U22457 : AOI22_X1 port map( A1 => n26856, A2 => n25810, B1 => n26850, B2 => 
                           n8573, ZN => n23548);
   U22458 : OAI221_X1 port map( B1 => n22669, B2 => n26745, C1 => n22477, C2 =>
                           n26739, A => n23556, ZN => n23553);
   U22459 : AOI22_X1 port map( A1 => n26733, A2 => n26229, B1 => n26727, B2 => 
                           n26349, ZN => n23556);
   U22460 : OAI221_X1 port map( B1 => n22548, B2 => n26868, C1 => n21216, C2 =>
                           n26862, A => n23530, ZN => n23527);
   U22461 : AOI22_X1 port map( A1 => n26856, A2 => n25815, B1 => n26850, B2 => 
                           n8570, ZN => n23530);
   U22462 : OAI221_X1 port map( B1 => n22668, B2 => n26745, C1 => n22476, C2 =>
                           n26739, A => n23538, ZN => n23535);
   U22463 : AOI22_X1 port map( A1 => n26733, A2 => n26230, B1 => n26727, B2 => 
                           n26350, ZN => n23538);
   U22464 : OAI221_X1 port map( B1 => n22547, B2 => n26869, C1 => n21215, C2 =>
                           n26863, A => n23512, ZN => n23509);
   U22465 : AOI22_X1 port map( A1 => n26857, A2 => n25820, B1 => n26851, B2 => 
                           n8567, ZN => n23512);
   U22466 : OAI221_X1 port map( B1 => n22667, B2 => n26746, C1 => n22475, C2 =>
                           n26740, A => n23520, ZN => n23517);
   U22467 : AOI22_X1 port map( A1 => n26734, A2 => n26231, B1 => n26728, B2 => 
                           n26351, ZN => n23520);
   U22468 : OAI221_X1 port map( B1 => n22546, B2 => n26869, C1 => n21214, C2 =>
                           n26863, A => n23494, ZN => n23491);
   U22469 : AOI22_X1 port map( A1 => n26857, A2 => n25825, B1 => n26851, B2 => 
                           n8564, ZN => n23494);
   U22470 : OAI221_X1 port map( B1 => n22666, B2 => n26746, C1 => n22474, C2 =>
                           n26740, A => n23502, ZN => n23499);
   U22471 : AOI22_X1 port map( A1 => n26734, A2 => n26232, B1 => n26728, B2 => 
                           n26352, ZN => n23502);
   U22472 : OAI221_X1 port map( B1 => n22545, B2 => n26869, C1 => n21213, C2 =>
                           n26863, A => n23476, ZN => n23473);
   U22473 : AOI22_X1 port map( A1 => n26857, A2 => n25830, B1 => n26851, B2 => 
                           n8561, ZN => n23476);
   U22474 : OAI221_X1 port map( B1 => n22665, B2 => n26746, C1 => n22473, C2 =>
                           n26740, A => n23484, ZN => n23481);
   U22475 : AOI22_X1 port map( A1 => n26734, A2 => n26233, B1 => n26728, B2 => 
                           n26353, ZN => n23484);
   U22476 : OAI221_X1 port map( B1 => n22544, B2 => n26869, C1 => n21212, C2 =>
                           n26863, A => n23458, ZN => n23455);
   U22477 : AOI22_X1 port map( A1 => n26857, A2 => n25835, B1 => n26851, B2 => 
                           n8558, ZN => n23458);
   U22478 : OAI221_X1 port map( B1 => n22664, B2 => n26746, C1 => n22472, C2 =>
                           n26740, A => n23466, ZN => n23463);
   U22479 : AOI22_X1 port map( A1 => n26734, A2 => n26234, B1 => n26728, B2 => 
                           n26354, ZN => n23466);
   U22480 : OAI221_X1 port map( B1 => n22543, B2 => n26869, C1 => n21211, C2 =>
                           n26863, A => n23440, ZN => n23437);
   U22481 : AOI22_X1 port map( A1 => n26857, A2 => n25840, B1 => n26851, B2 => 
                           n8555, ZN => n23440);
   U22482 : OAI221_X1 port map( B1 => n22663, B2 => n26746, C1 => n22471, C2 =>
                           n26740, A => n23448, ZN => n23445);
   U22483 : AOI22_X1 port map( A1 => n26734, A2 => n26235, B1 => n26728, B2 => 
                           n26355, ZN => n23448);
   U22484 : OAI221_X1 port map( B1 => n22542, B2 => n26869, C1 => n21210, C2 =>
                           n26863, A => n23422, ZN => n23419);
   U22485 : AOI22_X1 port map( A1 => n26857, A2 => n25845, B1 => n26851, B2 => 
                           n8552, ZN => n23422);
   U22486 : OAI221_X1 port map( B1 => n22662, B2 => n26746, C1 => n22470, C2 =>
                           n26740, A => n23430, ZN => n23427);
   U22487 : AOI22_X1 port map( A1 => n26734, A2 => n26236, B1 => n26728, B2 => 
                           n26356, ZN => n23430);
   U22488 : OAI221_X1 port map( B1 => n22541, B2 => n26869, C1 => n21209, C2 =>
                           n26863, A => n23404, ZN => n23401);
   U22489 : AOI22_X1 port map( A1 => n26857, A2 => n25850, B1 => n26851, B2 => 
                           n8549, ZN => n23404);
   U22490 : OAI221_X1 port map( B1 => n22661, B2 => n26746, C1 => n22469, C2 =>
                           n26740, A => n23412, ZN => n23409);
   U22491 : AOI22_X1 port map( A1 => n26734, A2 => n26237, B1 => n26728, B2 => 
                           n26357, ZN => n23412);
   U22492 : OAI221_X1 port map( B1 => n22540, B2 => n26869, C1 => n21208, C2 =>
                           n26863, A => n23386, ZN => n23383);
   U22493 : AOI22_X1 port map( A1 => n26857, A2 => n25855, B1 => n26851, B2 => 
                           n8546, ZN => n23386);
   U22494 : OAI221_X1 port map( B1 => n22660, B2 => n26746, C1 => n22468, C2 =>
                           n26740, A => n23394, ZN => n23391);
   U22495 : AOI22_X1 port map( A1 => n26734, A2 => n26238, B1 => n26728, B2 => 
                           n26358, ZN => n23394);
   U22496 : OAI221_X1 port map( B1 => n22539, B2 => n26869, C1 => n21207, C2 =>
                           n26863, A => n23368, ZN => n23365);
   U22497 : AOI22_X1 port map( A1 => n26857, A2 => n25860, B1 => n26851, B2 => 
                           n8543, ZN => n23368);
   U22498 : OAI221_X1 port map( B1 => n22659, B2 => n26746, C1 => n22467, C2 =>
                           n26740, A => n23376, ZN => n23373);
   U22499 : AOI22_X1 port map( A1 => n26734, A2 => n26239, B1 => n26728, B2 => 
                           n26359, ZN => n23376);
   U22500 : OAI221_X1 port map( B1 => n22538, B2 => n26869, C1 => n21206, C2 =>
                           n26863, A => n23350, ZN => n23347);
   U22501 : AOI22_X1 port map( A1 => n26857, A2 => n25865, B1 => n26851, B2 => 
                           n8540, ZN => n23350);
   U22502 : OAI221_X1 port map( B1 => n22658, B2 => n26746, C1 => n22466, C2 =>
                           n26740, A => n23358, ZN => n23355);
   U22503 : AOI22_X1 port map( A1 => n26734, A2 => n26240, B1 => n26728, B2 => 
                           n26360, ZN => n23358);
   U22504 : OAI221_X1 port map( B1 => n22537, B2 => n26869, C1 => n21205, C2 =>
                           n26863, A => n23332, ZN => n23329);
   U22505 : AOI22_X1 port map( A1 => n26857, A2 => n25870, B1 => n26851, B2 => 
                           n8537, ZN => n23332);
   U22506 : OAI221_X1 port map( B1 => n22657, B2 => n26746, C1 => n22465, C2 =>
                           n26740, A => n23340, ZN => n23337);
   U22507 : AOI22_X1 port map( A1 => n26734, A2 => n26241, B1 => n26728, B2 => 
                           n26361, ZN => n23340);
   U22508 : OAI221_X1 port map( B1 => n22536, B2 => n26869, C1 => n21204, C2 =>
                           n26863, A => n23314, ZN => n23311);
   U22509 : AOI22_X1 port map( A1 => n26857, A2 => n25875, B1 => n26851, B2 => 
                           n8534, ZN => n23314);
   U22510 : OAI221_X1 port map( B1 => n22656, B2 => n26746, C1 => n22464, C2 =>
                           n26740, A => n23322, ZN => n23319);
   U22511 : AOI22_X1 port map( A1 => n26734, A2 => n26242, B1 => n26728, B2 => 
                           n26362, ZN => n23322);
   U22512 : OAI221_X1 port map( B1 => n22535, B2 => n26870, C1 => n21203, C2 =>
                           n26864, A => n23296, ZN => n23293);
   U22513 : AOI22_X1 port map( A1 => n26858, A2 => n25880, B1 => n26852, B2 => 
                           n8531, ZN => n23296);
   U22514 : OAI221_X1 port map( B1 => n22655, B2 => n26747, C1 => n22463, C2 =>
                           n26741, A => n23304, ZN => n23301);
   U22515 : AOI22_X1 port map( A1 => n26735, A2 => n26243, B1 => n26729, B2 => 
                           n26363, ZN => n23304);
   U22516 : OAI221_X1 port map( B1 => n22534, B2 => n26870, C1 => n21202, C2 =>
                           n26864, A => n23278, ZN => n23275);
   U22517 : AOI22_X1 port map( A1 => n26858, A2 => n25885, B1 => n26852, B2 => 
                           n8528, ZN => n23278);
   U22518 : OAI221_X1 port map( B1 => n22654, B2 => n26747, C1 => n22462, C2 =>
                           n26741, A => n23286, ZN => n23283);
   U22519 : AOI22_X1 port map( A1 => n26735, A2 => n26244, B1 => n26729, B2 => 
                           n26364, ZN => n23286);
   U22520 : OAI221_X1 port map( B1 => n22533, B2 => n26870, C1 => n21201, C2 =>
                           n26864, A => n23260, ZN => n23257);
   U22521 : AOI22_X1 port map( A1 => n26858, A2 => n25890, B1 => n26852, B2 => 
                           n8525, ZN => n23260);
   U22522 : OAI221_X1 port map( B1 => n22653, B2 => n26747, C1 => n22461, C2 =>
                           n26741, A => n23268, ZN => n23265);
   U22523 : AOI22_X1 port map( A1 => n26735, A2 => n26245, B1 => n26729, B2 => 
                           n26365, ZN => n23268);
   U22524 : OAI221_X1 port map( B1 => n22532, B2 => n26870, C1 => n21200, C2 =>
                           n26864, A => n23242, ZN => n23239);
   U22525 : AOI22_X1 port map( A1 => n26858, A2 => n25895, B1 => n26852, B2 => 
                           n8522, ZN => n23242);
   U22526 : OAI221_X1 port map( B1 => n22652, B2 => n26747, C1 => n22460, C2 =>
                           n26741, A => n23250, ZN => n23247);
   U22527 : AOI22_X1 port map( A1 => n26735, A2 => n26246, B1 => n26729, B2 => 
                           n26366, ZN => n23250);
   U22528 : OAI221_X1 port map( B1 => n22531, B2 => n26870, C1 => n21199, C2 =>
                           n26864, A => n23224, ZN => n23221);
   U22529 : AOI22_X1 port map( A1 => n26858, A2 => n25900, B1 => n26852, B2 => 
                           n8519, ZN => n23224);
   U22530 : OAI221_X1 port map( B1 => n22651, B2 => n26747, C1 => n22459, C2 =>
                           n26741, A => n23232, ZN => n23229);
   U22531 : AOI22_X1 port map( A1 => n26735, A2 => n26247, B1 => n26729, B2 => 
                           n26367, ZN => n23232);
   U22532 : OAI221_X1 port map( B1 => n22530, B2 => n26870, C1 => n21198, C2 =>
                           n26864, A => n23206, ZN => n23203);
   U22533 : AOI22_X1 port map( A1 => n26858, A2 => n25905, B1 => n26852, B2 => 
                           n8516, ZN => n23206);
   U22534 : OAI221_X1 port map( B1 => n22650, B2 => n26747, C1 => n22458, C2 =>
                           n26741, A => n23214, ZN => n23211);
   U22535 : AOI22_X1 port map( A1 => n26735, A2 => n26248, B1 => n26729, B2 => 
                           n26368, ZN => n23214);
   U22536 : OAI221_X1 port map( B1 => n22529, B2 => n26870, C1 => n21197, C2 =>
                           n26864, A => n23188, ZN => n23185);
   U22537 : AOI22_X1 port map( A1 => n26858, A2 => n25910, B1 => n26852, B2 => 
                           n8513, ZN => n23188);
   U22538 : OAI221_X1 port map( B1 => n22649, B2 => n26747, C1 => n22457, C2 =>
                           n26741, A => n23196, ZN => n23193);
   U22539 : AOI22_X1 port map( A1 => n26735, A2 => n26249, B1 => n26729, B2 => 
                           n26369, ZN => n23196);
   U22540 : OAI221_X1 port map( B1 => n22528, B2 => n26870, C1 => n21196, C2 =>
                           n26864, A => n23170, ZN => n23167);
   U22541 : AOI22_X1 port map( A1 => n26858, A2 => n25915, B1 => n26852, B2 => 
                           n8510, ZN => n23170);
   U22542 : OAI221_X1 port map( B1 => n22648, B2 => n26747, C1 => n22456, C2 =>
                           n26741, A => n23178, ZN => n23175);
   U22543 : AOI22_X1 port map( A1 => n26735, A2 => n26250, B1 => n26729, B2 => 
                           n26370, ZN => n23178);
   U22544 : OAI221_X1 port map( B1 => n22527, B2 => n26870, C1 => n21195, C2 =>
                           n26864, A => n23152, ZN => n23149);
   U22545 : AOI22_X1 port map( A1 => n26858, A2 => n25920, B1 => n26852, B2 => 
                           n8507, ZN => n23152);
   U22546 : OAI221_X1 port map( B1 => n22647, B2 => n26747, C1 => n22455, C2 =>
                           n26741, A => n23160, ZN => n23157);
   U22547 : AOI22_X1 port map( A1 => n26735, A2 => n26251, B1 => n26729, B2 => 
                           n26371, ZN => n23160);
   U22548 : OAI221_X1 port map( B1 => n22526, B2 => n26870, C1 => n21194, C2 =>
                           n26864, A => n23134, ZN => n23131);
   U22549 : AOI22_X1 port map( A1 => n26858, A2 => n25925, B1 => n26852, B2 => 
                           n8504, ZN => n23134);
   U22550 : OAI221_X1 port map( B1 => n22646, B2 => n26747, C1 => n22454, C2 =>
                           n26741, A => n23142, ZN => n23139);
   U22551 : AOI22_X1 port map( A1 => n26735, A2 => n26252, B1 => n26729, B2 => 
                           n26372, ZN => n23142);
   U22552 : OAI221_X1 port map( B1 => n22525, B2 => n26870, C1 => n21193, C2 =>
                           n26864, A => n23116, ZN => n23113);
   U22553 : AOI22_X1 port map( A1 => n26858, A2 => n25930, B1 => n26852, B2 => 
                           n8501, ZN => n23116);
   U22554 : OAI221_X1 port map( B1 => n22645, B2 => n26747, C1 => n22453, C2 =>
                           n26741, A => n23124, ZN => n23121);
   U22555 : AOI22_X1 port map( A1 => n26735, A2 => n26253, B1 => n26729, B2 => 
                           n26373, ZN => n23124);
   U22556 : OAI221_X1 port map( B1 => n22524, B2 => n26870, C1 => n21192, C2 =>
                           n26864, A => n23098, ZN => n23095);
   U22557 : AOI22_X1 port map( A1 => n26858, A2 => n25935, B1 => n26852, B2 => 
                           n8498, ZN => n23098);
   U22558 : OAI221_X1 port map( B1 => n22644, B2 => n26747, C1 => n22452, C2 =>
                           n26741, A => n23106, ZN => n23103);
   U22559 : AOI22_X1 port map( A1 => n26735, A2 => n26254, B1 => n26729, B2 => 
                           n26374, ZN => n23106);
   U22560 : OAI221_X1 port map( B1 => n22523, B2 => n26871, C1 => n21191, C2 =>
                           n26865, A => n23080, ZN => n23077);
   U22561 : AOI22_X1 port map( A1 => n26859, A2 => n25940, B1 => n26853, B2 => 
                           n8495, ZN => n23080);
   U22562 : OAI221_X1 port map( B1 => n22643, B2 => n26748, C1 => n22451, C2 =>
                           n26742, A => n23088, ZN => n23085);
   U22563 : AOI22_X1 port map( A1 => n26736, A2 => n26255, B1 => n26730, B2 => 
                           n26375, ZN => n23088);
   U22564 : OAI221_X1 port map( B1 => n22522, B2 => n26871, C1 => n21190, C2 =>
                           n26865, A => n23062, ZN => n23059);
   U22565 : AOI22_X1 port map( A1 => n26859, A2 => n25945, B1 => n26853, B2 => 
                           n8492, ZN => n23062);
   U22566 : OAI221_X1 port map( B1 => n22642, B2 => n26748, C1 => n22450, C2 =>
                           n26742, A => n23070, ZN => n23067);
   U22567 : AOI22_X1 port map( A1 => n26736, A2 => n26256, B1 => n26730, B2 => 
                           n26376, ZN => n23070);
   U22568 : OAI221_X1 port map( B1 => n22521, B2 => n26871, C1 => n21189, C2 =>
                           n26865, A => n23044, ZN => n23041);
   U22569 : AOI22_X1 port map( A1 => n26859, A2 => n25950, B1 => n26853, B2 => 
                           n8489, ZN => n23044);
   U22570 : OAI221_X1 port map( B1 => n22641, B2 => n26748, C1 => n22449, C2 =>
                           n26742, A => n23052, ZN => n23049);
   U22571 : AOI22_X1 port map( A1 => n26736, A2 => n26257, B1 => n26730, B2 => 
                           n26377, ZN => n23052);
   U22572 : OAI221_X1 port map( B1 => n22520, B2 => n26871, C1 => n21188, C2 =>
                           n26865, A => n23026, ZN => n23023);
   U22573 : AOI22_X1 port map( A1 => n26859, A2 => n25955, B1 => n26853, B2 => 
                           n8486, ZN => n23026);
   U22574 : OAI221_X1 port map( B1 => n22640, B2 => n26748, C1 => n22448, C2 =>
                           n26742, A => n23034, ZN => n23031);
   U22575 : AOI22_X1 port map( A1 => n26736, A2 => n26258, B1 => n26730, B2 => 
                           n26378, ZN => n23034);
   U22576 : OAI221_X1 port map( B1 => n22519, B2 => n26871, C1 => n21187, C2 =>
                           n26865, A => n23008, ZN => n23005);
   U22577 : AOI22_X1 port map( A1 => n26859, A2 => n25960, B1 => n26853, B2 => 
                           n8483, ZN => n23008);
   U22578 : OAI221_X1 port map( B1 => n22639, B2 => n26748, C1 => n22447, C2 =>
                           n26742, A => n23016, ZN => n23013);
   U22579 : AOI22_X1 port map( A1 => n26736, A2 => n26259, B1 => n26730, B2 => 
                           n26379, ZN => n23016);
   U22580 : OAI221_X1 port map( B1 => n22518, B2 => n26871, C1 => n21186, C2 =>
                           n26865, A => n22990, ZN => n22987);
   U22581 : AOI22_X1 port map( A1 => n26859, A2 => n25965, B1 => n26853, B2 => 
                           n8480, ZN => n22990);
   U22582 : OAI221_X1 port map( B1 => n22638, B2 => n26748, C1 => n22446, C2 =>
                           n26742, A => n22998, ZN => n22995);
   U22583 : AOI22_X1 port map( A1 => n26736, A2 => n26260, B1 => n26730, B2 => 
                           n26380, ZN => n22998);
   U22584 : OAI221_X1 port map( B1 => n22517, B2 => n26871, C1 => n21185, C2 =>
                           n26865, A => n22972, ZN => n22969);
   U22585 : AOI22_X1 port map( A1 => n26859, A2 => n25970, B1 => n26853, B2 => 
                           n8477, ZN => n22972);
   U22586 : OAI221_X1 port map( B1 => n22637, B2 => n26748, C1 => n22445, C2 =>
                           n26742, A => n22980, ZN => n22977);
   U22587 : AOI22_X1 port map( A1 => n26736, A2 => n26261, B1 => n26730, B2 => 
                           n26381, ZN => n22980);
   U22588 : OAI221_X1 port map( B1 => n22516, B2 => n26871, C1 => n21184, C2 =>
                           n26865, A => n22954, ZN => n22951);
   U22589 : AOI22_X1 port map( A1 => n26859, A2 => n25975, B1 => n26853, B2 => 
                           n8474, ZN => n22954);
   U22590 : OAI221_X1 port map( B1 => n22636, B2 => n26748, C1 => n22444, C2 =>
                           n26742, A => n22962, ZN => n22959);
   U22591 : AOI22_X1 port map( A1 => n26736, A2 => n26262, B1 => n26730, B2 => 
                           n26382, ZN => n22962);
   U22592 : OAI221_X1 port map( B1 => n22515, B2 => n26871, C1 => n21183, C2 =>
                           n26865, A => n22936, ZN => n22933);
   U22593 : AOI22_X1 port map( A1 => n26859, A2 => n25980, B1 => n26853, B2 => 
                           n8471, ZN => n22936);
   U22594 : OAI221_X1 port map( B1 => n22635, B2 => n26748, C1 => n22443, C2 =>
                           n26742, A => n22944, ZN => n22941);
   U22595 : AOI22_X1 port map( A1 => n26736, A2 => n26263, B1 => n26730, B2 => 
                           n26383, ZN => n22944);
   U22596 : OAI221_X1 port map( B1 => n22514, B2 => n26871, C1 => n21182, C2 =>
                           n26865, A => n22918, ZN => n22915);
   U22597 : AOI22_X1 port map( A1 => n26859, A2 => n25985, B1 => n26853, B2 => 
                           n8468, ZN => n22918);
   U22598 : OAI221_X1 port map( B1 => n22634, B2 => n26748, C1 => n22442, C2 =>
                           n26742, A => n22926, ZN => n22923);
   U22599 : AOI22_X1 port map( A1 => n26736, A2 => n26264, B1 => n26730, B2 => 
                           n26384, ZN => n22926);
   U22600 : OAI221_X1 port map( B1 => n22513, B2 => n26871, C1 => n21181, C2 =>
                           n26865, A => n22900, ZN => n22897);
   U22601 : AOI22_X1 port map( A1 => n26859, A2 => n25990, B1 => n26853, B2 => 
                           n8465, ZN => n22900);
   U22602 : OAI221_X1 port map( B1 => n22633, B2 => n26748, C1 => n22441, C2 =>
                           n26742, A => n22908, ZN => n22905);
   U22603 : AOI22_X1 port map( A1 => n26736, A2 => n26265, B1 => n26730, B2 => 
                           n26385, ZN => n22908);
   U22604 : OAI221_X1 port map( B1 => n22512, B2 => n26871, C1 => n21180, C2 =>
                           n26865, A => n22882, ZN => n22879);
   U22605 : AOI22_X1 port map( A1 => n26859, A2 => n25995, B1 => n26853, B2 => 
                           n8462, ZN => n22882);
   U22606 : OAI221_X1 port map( B1 => n22632, B2 => n26748, C1 => n22440, C2 =>
                           n26742, A => n22890, ZN => n22887);
   U22607 : AOI22_X1 port map( A1 => n26736, A2 => n26266, B1 => n26730, B2 => 
                           n26386, ZN => n22890);
   U22608 : OAI221_X1 port map( B1 => n22500, B2 => n26647, C1 => n21156, C2 =>
                           n26641, A => n23981, ZN => n23972);
   U22609 : AOI22_X1 port map( A1 => n26635, A2 => n25695, B1 => n26629, B2 => 
                           n8450, ZN => n23981);
   U22610 : OAI221_X1 port map( B1 => n22508, B2 => n26524, C1 => n22256, C2 =>
                           n26518, A => n24006, ZN => n23997);
   U22611 : AOI22_X1 port map( A1 => n26512, A2 => n26194, B1 => n26506, B2 => 
                           n26198, ZN => n24006);
   U22612 : OAI221_X1 port map( B1 => n22503, B2 => n26647, C1 => n21159, C2 =>
                           n26641, A => n24063, ZN => n24060);
   U22613 : AOI22_X1 port map( A1 => n26635, A2 => n25680, B1 => n26629, B2 => 
                           n8459, ZN => n24063);
   U22614 : OAI221_X1 port map( B1 => n22511, B2 => n26524, C1 => n22259, C2 =>
                           n26518, A => n24071, ZN => n24068);
   U22615 : AOI22_X1 port map( A1 => n26512, A2 => n26191, B1 => n26506, B2 => 
                           n26195, ZN => n24071);
   U22616 : OAI221_X1 port map( B1 => n22502, B2 => n26647, C1 => n21158, C2 =>
                           n26641, A => n24045, ZN => n24042);
   U22617 : AOI22_X1 port map( A1 => n26635, A2 => n25685, B1 => n26629, B2 => 
                           n8456, ZN => n24045);
   U22618 : OAI221_X1 port map( B1 => n22510, B2 => n26524, C1 => n22258, C2 =>
                           n26518, A => n24053, ZN => n24050);
   U22619 : AOI22_X1 port map( A1 => n26512, A2 => n26192, B1 => n26506, B2 => 
                           n26196, ZN => n24053);
   U22620 : OAI221_X1 port map( B1 => n22501, B2 => n26647, C1 => n21157, C2 =>
                           n26641, A => n24027, ZN => n24024);
   U22621 : AOI22_X1 port map( A1 => n26635, A2 => n25690, B1 => n26629, B2 => 
                           n8453, ZN => n24027);
   U22622 : OAI221_X1 port map( B1 => n22509, B2 => n26524, C1 => n22257, C2 =>
                           n26518, A => n24035, ZN => n24032);
   U22623 : AOI22_X1 port map( A1 => n26512, A2 => n26193, B1 => n26506, B2 => 
                           n26197, ZN => n24035);
   U22624 : OAI221_X1 port map( B1 => n22503, B2 => n26872, C1 => n21159, C2 =>
                           n26866, A => n22864, ZN => n22861);
   U22625 : AOI22_X1 port map( A1 => n26860, A2 => n25680, B1 => n26854, B2 => 
                           n8459, ZN => n22864);
   U22626 : OAI221_X1 port map( B1 => n22511, B2 => n26749, C1 => n22259, C2 =>
                           n26743, A => n22872, ZN => n22869);
   U22627 : AOI22_X1 port map( A1 => n26737, A2 => n26191, B1 => n26731, B2 => 
                           n26195, ZN => n22872);
   U22628 : OAI221_X1 port map( B1 => n22502, B2 => n26872, C1 => n21158, C2 =>
                           n26866, A => n22846, ZN => n22843);
   U22629 : AOI22_X1 port map( A1 => n26860, A2 => n25685, B1 => n26854, B2 => 
                           n8456, ZN => n22846);
   U22630 : OAI221_X1 port map( B1 => n22510, B2 => n26749, C1 => n22258, C2 =>
                           n26743, A => n22854, ZN => n22851);
   U22631 : AOI22_X1 port map( A1 => n26737, A2 => n26192, B1 => n26731, B2 => 
                           n26196, ZN => n22854);
   U22632 : OAI221_X1 port map( B1 => n22501, B2 => n26872, C1 => n21157, C2 =>
                           n26866, A => n22828, ZN => n22825);
   U22633 : AOI22_X1 port map( A1 => n26860, A2 => n25690, B1 => n26854, B2 => 
                           n8453, ZN => n22828);
   U22634 : OAI221_X1 port map( B1 => n22509, B2 => n26749, C1 => n22257, C2 =>
                           n26743, A => n22836, ZN => n22833);
   U22635 : AOI22_X1 port map( A1 => n26737, A2 => n26193, B1 => n26731, B2 => 
                           n26197, ZN => n22836);
   U22636 : OAI221_X1 port map( B1 => n22500, B2 => n26872, C1 => n21156, C2 =>
                           n26866, A => n22782, ZN => n22773);
   U22637 : AOI22_X1 port map( A1 => n26860, A2 => n25695, B1 => n26854, B2 => 
                           n8450, ZN => n22782);
   U22638 : OAI221_X1 port map( B1 => n22508, B2 => n26749, C1 => n22256, C2 =>
                           n26743, A => n22807, ZN => n22798);
   U22639 : AOI22_X1 port map( A1 => n26737, A2 => n26194, B1 => n26731, B2 => 
                           n26198, ZN => n22807);
   U22640 : OAI221_X1 port map( B1 => n22571, B2 => n26642, C1 => n21239, C2 =>
                           n26636, A => n25149, ZN => n25140);
   U22641 : AOI22_X1 port map( A1 => n26630, A2 => n25700, B1 => n26624, B2 => 
                           n8639, ZN => n25149);
   U22642 : OAI221_X1 port map( B1 => n22691, B2 => n26519, C1 => n22499, C2 =>
                           n26513, A => n25161, ZN => n25158);
   U22643 : AOI22_X1 port map( A1 => n26507, A2 => n26207, B1 => n26501, B2 => 
                           n26327, ZN => n25161);
   U22644 : OAI221_X1 port map( B1 => n22570, B2 => n26642, C1 => n21238, C2 =>
                           n26636, A => n25125, ZN => n25122);
   U22645 : AOI22_X1 port map( A1 => n26630, A2 => n25705, B1 => n26624, B2 => 
                           n8636, ZN => n25125);
   U22646 : OAI221_X1 port map( B1 => n22690, B2 => n26519, C1 => n22498, C2 =>
                           n26513, A => n25133, ZN => n25130);
   U22647 : AOI22_X1 port map( A1 => n26507, A2 => n26208, B1 => n26501, B2 => 
                           n26328, ZN => n25133);
   U22648 : OAI221_X1 port map( B1 => n22569, B2 => n26642, C1 => n21237, C2 =>
                           n26636, A => n25107, ZN => n25104);
   U22649 : AOI22_X1 port map( A1 => n26630, A2 => n25710, B1 => n26624, B2 => 
                           n8633, ZN => n25107);
   U22650 : OAI221_X1 port map( B1 => n22689, B2 => n26519, C1 => n22497, C2 =>
                           n26513, A => n25115, ZN => n25112);
   U22651 : AOI22_X1 port map( A1 => n26507, A2 => n26209, B1 => n26501, B2 => 
                           n26329, ZN => n25115);
   U22652 : OAI221_X1 port map( B1 => n22568, B2 => n26642, C1 => n21236, C2 =>
                           n26636, A => n25089, ZN => n25086);
   U22653 : AOI22_X1 port map( A1 => n26630, A2 => n25715, B1 => n26624, B2 => 
                           n8630, ZN => n25089);
   U22654 : OAI221_X1 port map( B1 => n22688, B2 => n26519, C1 => n22496, C2 =>
                           n26513, A => n25097, ZN => n25094);
   U22655 : AOI22_X1 port map( A1 => n26507, A2 => n26210, B1 => n26501, B2 => 
                           n26330, ZN => n25097);
   U22656 : OAI221_X1 port map( B1 => n22567, B2 => n26642, C1 => n21235, C2 =>
                           n26636, A => n25071, ZN => n25068);
   U22657 : AOI22_X1 port map( A1 => n26630, A2 => n25720, B1 => n26624, B2 => 
                           n8627, ZN => n25071);
   U22658 : OAI221_X1 port map( B1 => n22687, B2 => n26519, C1 => n22495, C2 =>
                           n26513, A => n25079, ZN => n25076);
   U22659 : AOI22_X1 port map( A1 => n26507, A2 => n26211, B1 => n26501, B2 => 
                           n26331, ZN => n25079);
   U22660 : OAI221_X1 port map( B1 => n22566, B2 => n26642, C1 => n21234, C2 =>
                           n26636, A => n25053, ZN => n25050);
   U22661 : AOI22_X1 port map( A1 => n26630, A2 => n25725, B1 => n26624, B2 => 
                           n8624, ZN => n25053);
   U22662 : OAI221_X1 port map( B1 => n22686, B2 => n26519, C1 => n22494, C2 =>
                           n26513, A => n25061, ZN => n25058);
   U22663 : AOI22_X1 port map( A1 => n26507, A2 => n26212, B1 => n26501, B2 => 
                           n26332, ZN => n25061);
   U22664 : OAI221_X1 port map( B1 => n22565, B2 => n26642, C1 => n21233, C2 =>
                           n26636, A => n25035, ZN => n25032);
   U22665 : AOI22_X1 port map( A1 => n26630, A2 => n25730, B1 => n26624, B2 => 
                           n8621, ZN => n25035);
   U22666 : OAI221_X1 port map( B1 => n22685, B2 => n26519, C1 => n22493, C2 =>
                           n26513, A => n25043, ZN => n25040);
   U22667 : AOI22_X1 port map( A1 => n26507, A2 => n26213, B1 => n26501, B2 => 
                           n26333, ZN => n25043);
   U22668 : OAI221_X1 port map( B1 => n22564, B2 => n26642, C1 => n21232, C2 =>
                           n26636, A => n25017, ZN => n25014);
   U22669 : AOI22_X1 port map( A1 => n26630, A2 => n25735, B1 => n26624, B2 => 
                           n8618, ZN => n25017);
   U22670 : OAI221_X1 port map( B1 => n22684, B2 => n26519, C1 => n22492, C2 =>
                           n26513, A => n25025, ZN => n25022);
   U22671 : AOI22_X1 port map( A1 => n26507, A2 => n26214, B1 => n26501, B2 => 
                           n26334, ZN => n25025);
   U22672 : OAI221_X1 port map( B1 => n22563, B2 => n26642, C1 => n21231, C2 =>
                           n26636, A => n24999, ZN => n24996);
   U22673 : AOI22_X1 port map( A1 => n26630, A2 => n25740, B1 => n26624, B2 => 
                           n8615, ZN => n24999);
   U22674 : OAI221_X1 port map( B1 => n22683, B2 => n26519, C1 => n22491, C2 =>
                           n26513, A => n25007, ZN => n25004);
   U22675 : AOI22_X1 port map( A1 => n26507, A2 => n26215, B1 => n26501, B2 => 
                           n26335, ZN => n25007);
   U22676 : OAI221_X1 port map( B1 => n22562, B2 => n26642, C1 => n21230, C2 =>
                           n26636, A => n24981, ZN => n24978);
   U22677 : AOI22_X1 port map( A1 => n26630, A2 => n25745, B1 => n26624, B2 => 
                           n8612, ZN => n24981);
   U22678 : OAI221_X1 port map( B1 => n22682, B2 => n26519, C1 => n22490, C2 =>
                           n26513, A => n24989, ZN => n24986);
   U22679 : AOI22_X1 port map( A1 => n26507, A2 => n26216, B1 => n26501, B2 => 
                           n26336, ZN => n24989);
   U22680 : OAI221_X1 port map( B1 => n22561, B2 => n26642, C1 => n21229, C2 =>
                           n26636, A => n24963, ZN => n24960);
   U22681 : AOI22_X1 port map( A1 => n26630, A2 => n25750, B1 => n26624, B2 => 
                           n8609, ZN => n24963);
   U22682 : OAI221_X1 port map( B1 => n22681, B2 => n26519, C1 => n22489, C2 =>
                           n26513, A => n24971, ZN => n24968);
   U22683 : AOI22_X1 port map( A1 => n26507, A2 => n26217, B1 => n26501, B2 => 
                           n26337, ZN => n24971);
   U22684 : OAI221_X1 port map( B1 => n22560, B2 => n26642, C1 => n21228, C2 =>
                           n26636, A => n24945, ZN => n24942);
   U22685 : AOI22_X1 port map( A1 => n26630, A2 => n25755, B1 => n26624, B2 => 
                           n8606, ZN => n24945);
   U22686 : OAI221_X1 port map( B1 => n22680, B2 => n26519, C1 => n22488, C2 =>
                           n26513, A => n24953, ZN => n24950);
   U22687 : AOI22_X1 port map( A1 => n26507, A2 => n26218, B1 => n26501, B2 => 
                           n26338, ZN => n24953);
   U22688 : OAI221_X1 port map( B1 => n22571, B2 => n26867, C1 => n21239, C2 =>
                           n26861, A => n23950, ZN => n23941);
   U22689 : AOI22_X1 port map( A1 => n26855, A2 => n25700, B1 => n26849, B2 => 
                           n8639, ZN => n23950);
   U22690 : OAI221_X1 port map( B1 => n22691, B2 => n26744, C1 => n22499, C2 =>
                           n26738, A => n23962, ZN => n23959);
   U22691 : AOI22_X1 port map( A1 => n26732, A2 => n26207, B1 => n26726, B2 => 
                           n26327, ZN => n23962);
   U22692 : OAI221_X1 port map( B1 => n22570, B2 => n26867, C1 => n21238, C2 =>
                           n26861, A => n23926, ZN => n23923);
   U22693 : AOI22_X1 port map( A1 => n26855, A2 => n25705, B1 => n26849, B2 => 
                           n8636, ZN => n23926);
   U22694 : OAI221_X1 port map( B1 => n22690, B2 => n26744, C1 => n22498, C2 =>
                           n26738, A => n23934, ZN => n23931);
   U22695 : AOI22_X1 port map( A1 => n26732, A2 => n26208, B1 => n26726, B2 => 
                           n26328, ZN => n23934);
   U22696 : OAI221_X1 port map( B1 => n22569, B2 => n26867, C1 => n21237, C2 =>
                           n26861, A => n23908, ZN => n23905);
   U22697 : AOI22_X1 port map( A1 => n26855, A2 => n25710, B1 => n26849, B2 => 
                           n8633, ZN => n23908);
   U22698 : OAI221_X1 port map( B1 => n22689, B2 => n26744, C1 => n22497, C2 =>
                           n26738, A => n23916, ZN => n23913);
   U22699 : AOI22_X1 port map( A1 => n26732, A2 => n26209, B1 => n26726, B2 => 
                           n26329, ZN => n23916);
   U22700 : OAI221_X1 port map( B1 => n22568, B2 => n26867, C1 => n21236, C2 =>
                           n26861, A => n23890, ZN => n23887);
   U22701 : AOI22_X1 port map( A1 => n26855, A2 => n25715, B1 => n26849, B2 => 
                           n8630, ZN => n23890);
   U22702 : OAI221_X1 port map( B1 => n22688, B2 => n26744, C1 => n22496, C2 =>
                           n26738, A => n23898, ZN => n23895);
   U22703 : AOI22_X1 port map( A1 => n26732, A2 => n26210, B1 => n26726, B2 => 
                           n26330, ZN => n23898);
   U22704 : OAI221_X1 port map( B1 => n22567, B2 => n26867, C1 => n21235, C2 =>
                           n26861, A => n23872, ZN => n23869);
   U22705 : AOI22_X1 port map( A1 => n26855, A2 => n25720, B1 => n26849, B2 => 
                           n8627, ZN => n23872);
   U22706 : OAI221_X1 port map( B1 => n22687, B2 => n26744, C1 => n22495, C2 =>
                           n26738, A => n23880, ZN => n23877);
   U22707 : AOI22_X1 port map( A1 => n26732, A2 => n26211, B1 => n26726, B2 => 
                           n26331, ZN => n23880);
   U22708 : OAI221_X1 port map( B1 => n22566, B2 => n26867, C1 => n21234, C2 =>
                           n26861, A => n23854, ZN => n23851);
   U22709 : AOI22_X1 port map( A1 => n26855, A2 => n25725, B1 => n26849, B2 => 
                           n8624, ZN => n23854);
   U22710 : OAI221_X1 port map( B1 => n22686, B2 => n26744, C1 => n22494, C2 =>
                           n26738, A => n23862, ZN => n23859);
   U22711 : AOI22_X1 port map( A1 => n26732, A2 => n26212, B1 => n26726, B2 => 
                           n26332, ZN => n23862);
   U22712 : OAI221_X1 port map( B1 => n22565, B2 => n26867, C1 => n21233, C2 =>
                           n26861, A => n23836, ZN => n23833);
   U22713 : AOI22_X1 port map( A1 => n26855, A2 => n25730, B1 => n26849, B2 => 
                           n8621, ZN => n23836);
   U22714 : OAI221_X1 port map( B1 => n22685, B2 => n26744, C1 => n22493, C2 =>
                           n26738, A => n23844, ZN => n23841);
   U22715 : AOI22_X1 port map( A1 => n26732, A2 => n26213, B1 => n26726, B2 => 
                           n26333, ZN => n23844);
   U22716 : OAI221_X1 port map( B1 => n22564, B2 => n26867, C1 => n21232, C2 =>
                           n26861, A => n23818, ZN => n23815);
   U22717 : AOI22_X1 port map( A1 => n26855, A2 => n25735, B1 => n26849, B2 => 
                           n8618, ZN => n23818);
   U22718 : OAI221_X1 port map( B1 => n22684, B2 => n26744, C1 => n22492, C2 =>
                           n26738, A => n23826, ZN => n23823);
   U22719 : AOI22_X1 port map( A1 => n26732, A2 => n26214, B1 => n26726, B2 => 
                           n26334, ZN => n23826);
   U22720 : OAI221_X1 port map( B1 => n22563, B2 => n26867, C1 => n21231, C2 =>
                           n26861, A => n23800, ZN => n23797);
   U22721 : AOI22_X1 port map( A1 => n26855, A2 => n25740, B1 => n26849, B2 => 
                           n8615, ZN => n23800);
   U22722 : OAI221_X1 port map( B1 => n22683, B2 => n26744, C1 => n22491, C2 =>
                           n26738, A => n23808, ZN => n23805);
   U22723 : AOI22_X1 port map( A1 => n26732, A2 => n26215, B1 => n26726, B2 => 
                           n26335, ZN => n23808);
   U22724 : OAI221_X1 port map( B1 => n22562, B2 => n26867, C1 => n21230, C2 =>
                           n26861, A => n23782, ZN => n23779);
   U22725 : AOI22_X1 port map( A1 => n26855, A2 => n25745, B1 => n26849, B2 => 
                           n8612, ZN => n23782);
   U22726 : OAI221_X1 port map( B1 => n22682, B2 => n26744, C1 => n22490, C2 =>
                           n26738, A => n23790, ZN => n23787);
   U22727 : AOI22_X1 port map( A1 => n26732, A2 => n26216, B1 => n26726, B2 => 
                           n26336, ZN => n23790);
   U22728 : OAI221_X1 port map( B1 => n22561, B2 => n26867, C1 => n21229, C2 =>
                           n26861, A => n23764, ZN => n23761);
   U22729 : AOI22_X1 port map( A1 => n26855, A2 => n25750, B1 => n26849, B2 => 
                           n8609, ZN => n23764);
   U22730 : OAI221_X1 port map( B1 => n22681, B2 => n26744, C1 => n22489, C2 =>
                           n26738, A => n23772, ZN => n23769);
   U22731 : AOI22_X1 port map( A1 => n26732, A2 => n26217, B1 => n26726, B2 => 
                           n26337, ZN => n23772);
   U22732 : OAI221_X1 port map( B1 => n22560, B2 => n26867, C1 => n21228, C2 =>
                           n26861, A => n23746, ZN => n23743);
   U22733 : AOI22_X1 port map( A1 => n26855, A2 => n25755, B1 => n26849, B2 => 
                           n8606, ZN => n23746);
   U22734 : OAI221_X1 port map( B1 => n22680, B2 => n26744, C1 => n22488, C2 =>
                           n26738, A => n23754, ZN => n23751);
   U22735 : AOI22_X1 port map( A1 => n26732, A2 => n26218, B1 => n26726, B2 => 
                           n26338, ZN => n23754);
   U22736 : OAI221_X1 port map( B1 => n9620, B2 => n26619, C1 => n20822, C2 => 
                           n26613, A => n24928, ZN => n24923);
   U22737 : AOI22_X1 port map( A1 => n26607, A2 => n25761, B1 => n26601, B2 => 
                           n21022, ZN => n24928);
   U22738 : OAI221_X1 port map( B1 => n9619, B2 => n26619, C1 => n20821, C2 => 
                           n26613, A => n24910, ZN => n24905);
   U22739 : AOI22_X1 port map( A1 => n26607, A2 => n25766, B1 => n26601, B2 => 
                           n21021, ZN => n24910);
   U22740 : OAI221_X1 port map( B1 => n9618, B2 => n26619, C1 => n20820, C2 => 
                           n26613, A => n24892, ZN => n24887);
   U22741 : AOI22_X1 port map( A1 => n26607, A2 => n25771, B1 => n26601, B2 => 
                           n21020, ZN => n24892);
   U22742 : OAI221_X1 port map( B1 => n9617, B2 => n26619, C1 => n20819, C2 => 
                           n26613, A => n24874, ZN => n24869);
   U22743 : AOI22_X1 port map( A1 => n26607, A2 => n25776, B1 => n26601, B2 => 
                           n21019, ZN => n24874);
   U22744 : OAI221_X1 port map( B1 => n9616, B2 => n26619, C1 => n20818, C2 => 
                           n26613, A => n24856, ZN => n24851);
   U22745 : AOI22_X1 port map( A1 => n26607, A2 => n25781, B1 => n26601, B2 => 
                           n21018, ZN => n24856);
   U22746 : OAI221_X1 port map( B1 => n9615, B2 => n26619, C1 => n20817, C2 => 
                           n26613, A => n24838, ZN => n24833);
   U22747 : AOI22_X1 port map( A1 => n26607, A2 => n25786, B1 => n26601, B2 => 
                           n21017, ZN => n24838);
   U22748 : OAI221_X1 port map( B1 => n9614, B2 => n26619, C1 => n20816, C2 => 
                           n26613, A => n24820, ZN => n24815);
   U22749 : AOI22_X1 port map( A1 => n26607, A2 => n25791, B1 => n26601, B2 => 
                           n21016, ZN => n24820);
   U22750 : OAI221_X1 port map( B1 => n9613, B2 => n26619, C1 => n20815, C2 => 
                           n26613, A => n24802, ZN => n24797);
   U22751 : AOI22_X1 port map( A1 => n26607, A2 => n25796, B1 => n26601, B2 => 
                           n21015, ZN => n24802);
   U22752 : OAI221_X1 port map( B1 => n9612, B2 => n26619, C1 => n20814, C2 => 
                           n26613, A => n24784, ZN => n24779);
   U22753 : AOI22_X1 port map( A1 => n26607, A2 => n25801, B1 => n26601, B2 => 
                           n21014, ZN => n24784);
   U22754 : OAI221_X1 port map( B1 => n9611, B2 => n26619, C1 => n20813, C2 => 
                           n26613, A => n24766, ZN => n24761);
   U22755 : AOI22_X1 port map( A1 => n26607, A2 => n25806, B1 => n26601, B2 => 
                           n21013, ZN => n24766);
   U22756 : OAI221_X1 port map( B1 => n9610, B2 => n26619, C1 => n20812, C2 => 
                           n26613, A => n24748, ZN => n24743);
   U22757 : AOI22_X1 port map( A1 => n26607, A2 => n25811, B1 => n26601, B2 => 
                           n21012, ZN => n24748);
   U22758 : OAI221_X1 port map( B1 => n9609, B2 => n26619, C1 => n20811, C2 => 
                           n26613, A => n24730, ZN => n24725);
   U22759 : AOI22_X1 port map( A1 => n26607, A2 => n25816, B1 => n26601, B2 => 
                           n21011, ZN => n24730);
   U22760 : OAI221_X1 port map( B1 => n9608, B2 => n26620, C1 => n20810, C2 => 
                           n26614, A => n24712, ZN => n24707);
   U22761 : AOI22_X1 port map( A1 => n26608, A2 => n25821, B1 => n26602, B2 => 
                           n21010, ZN => n24712);
   U22762 : OAI221_X1 port map( B1 => n9607, B2 => n26620, C1 => n20809, C2 => 
                           n26614, A => n24694, ZN => n24689);
   U22763 : AOI22_X1 port map( A1 => n26608, A2 => n25826, B1 => n26602, B2 => 
                           n21009, ZN => n24694);
   U22764 : OAI221_X1 port map( B1 => n9606, B2 => n26620, C1 => n20808, C2 => 
                           n26614, A => n24676, ZN => n24671);
   U22765 : AOI22_X1 port map( A1 => n26608, A2 => n25831, B1 => n26602, B2 => 
                           n21008, ZN => n24676);
   U22766 : OAI221_X1 port map( B1 => n9605, B2 => n26620, C1 => n20807, C2 => 
                           n26614, A => n24658, ZN => n24653);
   U22767 : AOI22_X1 port map( A1 => n26608, A2 => n25836, B1 => n26602, B2 => 
                           n21007, ZN => n24658);
   U22768 : OAI221_X1 port map( B1 => n9604, B2 => n26620, C1 => n20806, C2 => 
                           n26614, A => n24640, ZN => n24635);
   U22769 : AOI22_X1 port map( A1 => n26608, A2 => n25841, B1 => n26602, B2 => 
                           n21006, ZN => n24640);
   U22770 : OAI221_X1 port map( B1 => n9603, B2 => n26620, C1 => n20805, C2 => 
                           n26614, A => n24622, ZN => n24617);
   U22771 : AOI22_X1 port map( A1 => n26608, A2 => n25846, B1 => n26602, B2 => 
                           n21005, ZN => n24622);
   U22772 : OAI221_X1 port map( B1 => n9602, B2 => n26620, C1 => n20804, C2 => 
                           n26614, A => n24604, ZN => n24599);
   U22773 : AOI22_X1 port map( A1 => n26608, A2 => n25851, B1 => n26602, B2 => 
                           n21004, ZN => n24604);
   U22774 : OAI221_X1 port map( B1 => n9601, B2 => n26620, C1 => n20803, C2 => 
                           n26614, A => n24586, ZN => n24581);
   U22775 : AOI22_X1 port map( A1 => n26608, A2 => n25856, B1 => n26602, B2 => 
                           n21003, ZN => n24586);
   U22776 : OAI221_X1 port map( B1 => n9600, B2 => n26620, C1 => n20802, C2 => 
                           n26614, A => n24568, ZN => n24563);
   U22777 : AOI22_X1 port map( A1 => n26608, A2 => n25861, B1 => n26602, B2 => 
                           n21002, ZN => n24568);
   U22778 : OAI221_X1 port map( B1 => n9599, B2 => n26620, C1 => n20801, C2 => 
                           n26614, A => n24550, ZN => n24545);
   U22779 : AOI22_X1 port map( A1 => n26608, A2 => n25866, B1 => n26602, B2 => 
                           n21001, ZN => n24550);
   U22780 : OAI221_X1 port map( B1 => n9598, B2 => n26620, C1 => n20800, C2 => 
                           n26614, A => n24532, ZN => n24527);
   U22781 : AOI22_X1 port map( A1 => n26608, A2 => n25871, B1 => n26602, B2 => 
                           n21000, ZN => n24532);
   U22782 : OAI221_X1 port map( B1 => n9597, B2 => n26620, C1 => n20799, C2 => 
                           n26614, A => n24514, ZN => n24509);
   U22783 : AOI22_X1 port map( A1 => n26608, A2 => n25876, B1 => n26602, B2 => 
                           n20999, ZN => n24514);
   U22784 : OAI221_X1 port map( B1 => n9596, B2 => n26621, C1 => n20798, C2 => 
                           n26615, A => n24496, ZN => n24491);
   U22785 : AOI22_X1 port map( A1 => n26609, A2 => n25881, B1 => n26603, B2 => 
                           n20998, ZN => n24496);
   U22786 : OAI221_X1 port map( B1 => n9595, B2 => n26621, C1 => n20797, C2 => 
                           n26615, A => n24478, ZN => n24473);
   U22787 : AOI22_X1 port map( A1 => n26609, A2 => n25886, B1 => n26603, B2 => 
                           n20997, ZN => n24478);
   U22788 : OAI221_X1 port map( B1 => n9594, B2 => n26621, C1 => n20796, C2 => 
                           n26615, A => n24460, ZN => n24455);
   U22789 : AOI22_X1 port map( A1 => n26609, A2 => n25891, B1 => n26603, B2 => 
                           n20996, ZN => n24460);
   U22790 : OAI221_X1 port map( B1 => n9593, B2 => n26621, C1 => n20795, C2 => 
                           n26615, A => n24442, ZN => n24437);
   U22791 : AOI22_X1 port map( A1 => n26609, A2 => n25896, B1 => n26603, B2 => 
                           n20995, ZN => n24442);
   U22792 : OAI221_X1 port map( B1 => n9592, B2 => n26621, C1 => n20794, C2 => 
                           n26615, A => n24424, ZN => n24419);
   U22793 : AOI22_X1 port map( A1 => n26609, A2 => n25901, B1 => n26603, B2 => 
                           n20994, ZN => n24424);
   U22794 : OAI221_X1 port map( B1 => n9591, B2 => n26621, C1 => n20793, C2 => 
                           n26615, A => n24406, ZN => n24401);
   U22795 : AOI22_X1 port map( A1 => n26609, A2 => n25906, B1 => n26603, B2 => 
                           n20993, ZN => n24406);
   U22796 : OAI221_X1 port map( B1 => n9590, B2 => n26621, C1 => n20792, C2 => 
                           n26615, A => n24388, ZN => n24383);
   U22797 : AOI22_X1 port map( A1 => n26609, A2 => n25911, B1 => n26603, B2 => 
                           n20992, ZN => n24388);
   U22798 : OAI221_X1 port map( B1 => n9589, B2 => n26621, C1 => n20791, C2 => 
                           n26615, A => n24370, ZN => n24365);
   U22799 : AOI22_X1 port map( A1 => n26609, A2 => n25916, B1 => n26603, B2 => 
                           n20991, ZN => n24370);
   U22800 : OAI221_X1 port map( B1 => n9588, B2 => n26621, C1 => n20790, C2 => 
                           n26615, A => n24352, ZN => n24347);
   U22801 : AOI22_X1 port map( A1 => n26609, A2 => n25921, B1 => n26603, B2 => 
                           n20990, ZN => n24352);
   U22802 : OAI221_X1 port map( B1 => n9587, B2 => n26621, C1 => n20789, C2 => 
                           n26615, A => n24334, ZN => n24329);
   U22803 : AOI22_X1 port map( A1 => n26609, A2 => n25926, B1 => n26603, B2 => 
                           n20989, ZN => n24334);
   U22804 : OAI221_X1 port map( B1 => n9586, B2 => n26621, C1 => n20788, C2 => 
                           n26615, A => n24316, ZN => n24311);
   U22805 : AOI22_X1 port map( A1 => n26609, A2 => n25931, B1 => n26603, B2 => 
                           n20988, ZN => n24316);
   U22806 : OAI221_X1 port map( B1 => n9585, B2 => n26621, C1 => n20787, C2 => 
                           n26615, A => n24298, ZN => n24293);
   U22807 : AOI22_X1 port map( A1 => n26609, A2 => n25936, B1 => n26603, B2 => 
                           n20987, ZN => n24298);
   U22808 : OAI221_X1 port map( B1 => n9620, B2 => n26844, C1 => n20822, C2 => 
                           n26838, A => n23729, ZN => n23724);
   U22809 : AOI22_X1 port map( A1 => n26832, A2 => n25761, B1 => n26826, B2 => 
                           n21022, ZN => n23729);
   U22810 : OAI221_X1 port map( B1 => n9619, B2 => n26844, C1 => n20821, C2 => 
                           n26838, A => n23711, ZN => n23706);
   U22811 : AOI22_X1 port map( A1 => n26832, A2 => n25766, B1 => n26826, B2 => 
                           n21021, ZN => n23711);
   U22812 : OAI221_X1 port map( B1 => n9618, B2 => n26844, C1 => n20820, C2 => 
                           n26838, A => n23693, ZN => n23688);
   U22813 : AOI22_X1 port map( A1 => n26832, A2 => n25771, B1 => n26826, B2 => 
                           n21020, ZN => n23693);
   U22814 : OAI221_X1 port map( B1 => n9617, B2 => n26844, C1 => n20819, C2 => 
                           n26838, A => n23675, ZN => n23670);
   U22815 : AOI22_X1 port map( A1 => n26832, A2 => n25776, B1 => n26826, B2 => 
                           n21019, ZN => n23675);
   U22816 : OAI221_X1 port map( B1 => n9616, B2 => n26844, C1 => n20818, C2 => 
                           n26838, A => n23657, ZN => n23652);
   U22817 : AOI22_X1 port map( A1 => n26832, A2 => n25781, B1 => n26826, B2 => 
                           n21018, ZN => n23657);
   U22818 : OAI221_X1 port map( B1 => n9615, B2 => n26844, C1 => n20817, C2 => 
                           n26838, A => n23639, ZN => n23634);
   U22819 : AOI22_X1 port map( A1 => n26832, A2 => n25786, B1 => n26826, B2 => 
                           n21017, ZN => n23639);
   U22820 : OAI221_X1 port map( B1 => n9614, B2 => n26844, C1 => n20816, C2 => 
                           n26838, A => n23621, ZN => n23616);
   U22821 : AOI22_X1 port map( A1 => n26832, A2 => n25791, B1 => n26826, B2 => 
                           n21016, ZN => n23621);
   U22822 : OAI221_X1 port map( B1 => n9613, B2 => n26844, C1 => n20815, C2 => 
                           n26838, A => n23603, ZN => n23598);
   U22823 : AOI22_X1 port map( A1 => n26832, A2 => n25796, B1 => n26826, B2 => 
                           n21015, ZN => n23603);
   U22824 : OAI221_X1 port map( B1 => n9612, B2 => n26844, C1 => n20814, C2 => 
                           n26838, A => n23585, ZN => n23580);
   U22825 : AOI22_X1 port map( A1 => n26832, A2 => n25801, B1 => n26826, B2 => 
                           n21014, ZN => n23585);
   U22826 : OAI221_X1 port map( B1 => n9611, B2 => n26844, C1 => n20813, C2 => 
                           n26838, A => n23567, ZN => n23562);
   U22827 : AOI22_X1 port map( A1 => n26832, A2 => n25806, B1 => n26826, B2 => 
                           n21013, ZN => n23567);
   U22828 : OAI221_X1 port map( B1 => n9610, B2 => n26844, C1 => n20812, C2 => 
                           n26838, A => n23549, ZN => n23544);
   U22829 : AOI22_X1 port map( A1 => n26832, A2 => n25811, B1 => n26826, B2 => 
                           n21012, ZN => n23549);
   U22830 : OAI221_X1 port map( B1 => n9609, B2 => n26844, C1 => n20811, C2 => 
                           n26838, A => n23531, ZN => n23526);
   U22831 : AOI22_X1 port map( A1 => n26832, A2 => n25816, B1 => n26826, B2 => 
                           n21011, ZN => n23531);
   U22832 : OAI221_X1 port map( B1 => n9608, B2 => n26845, C1 => n20810, C2 => 
                           n26839, A => n23513, ZN => n23508);
   U22833 : AOI22_X1 port map( A1 => n26833, A2 => n25821, B1 => n26827, B2 => 
                           n21010, ZN => n23513);
   U22834 : OAI221_X1 port map( B1 => n9607, B2 => n26845, C1 => n20809, C2 => 
                           n26839, A => n23495, ZN => n23490);
   U22835 : AOI22_X1 port map( A1 => n26833, A2 => n25826, B1 => n26827, B2 => 
                           n21009, ZN => n23495);
   U22836 : OAI221_X1 port map( B1 => n9606, B2 => n26845, C1 => n20808, C2 => 
                           n26839, A => n23477, ZN => n23472);
   U22837 : AOI22_X1 port map( A1 => n26833, A2 => n25831, B1 => n26827, B2 => 
                           n21008, ZN => n23477);
   U22838 : OAI221_X1 port map( B1 => n9605, B2 => n26845, C1 => n20807, C2 => 
                           n26839, A => n23459, ZN => n23454);
   U22839 : AOI22_X1 port map( A1 => n26833, A2 => n25836, B1 => n26827, B2 => 
                           n21007, ZN => n23459);
   U22840 : OAI221_X1 port map( B1 => n9604, B2 => n26845, C1 => n20806, C2 => 
                           n26839, A => n23441, ZN => n23436);
   U22841 : AOI22_X1 port map( A1 => n26833, A2 => n25841, B1 => n26827, B2 => 
                           n21006, ZN => n23441);
   U22842 : OAI221_X1 port map( B1 => n9603, B2 => n26845, C1 => n20805, C2 => 
                           n26839, A => n23423, ZN => n23418);
   U22843 : AOI22_X1 port map( A1 => n26833, A2 => n25846, B1 => n26827, B2 => 
                           n21005, ZN => n23423);
   U22844 : OAI221_X1 port map( B1 => n9602, B2 => n26845, C1 => n20804, C2 => 
                           n26839, A => n23405, ZN => n23400);
   U22845 : AOI22_X1 port map( A1 => n26833, A2 => n25851, B1 => n26827, B2 => 
                           n21004, ZN => n23405);
   U22846 : OAI221_X1 port map( B1 => n9601, B2 => n26845, C1 => n20803, C2 => 
                           n26839, A => n23387, ZN => n23382);
   U22847 : AOI22_X1 port map( A1 => n26833, A2 => n25856, B1 => n26827, B2 => 
                           n21003, ZN => n23387);
   U22848 : OAI221_X1 port map( B1 => n9600, B2 => n26845, C1 => n20802, C2 => 
                           n26839, A => n23369, ZN => n23364);
   U22849 : AOI22_X1 port map( A1 => n26833, A2 => n25861, B1 => n26827, B2 => 
                           n21002, ZN => n23369);
   U22850 : OAI221_X1 port map( B1 => n9599, B2 => n26845, C1 => n20801, C2 => 
                           n26839, A => n23351, ZN => n23346);
   U22851 : AOI22_X1 port map( A1 => n26833, A2 => n25866, B1 => n26827, B2 => 
                           n21001, ZN => n23351);
   U22852 : OAI221_X1 port map( B1 => n9598, B2 => n26845, C1 => n20800, C2 => 
                           n26839, A => n23333, ZN => n23328);
   U22853 : AOI22_X1 port map( A1 => n26833, A2 => n25871, B1 => n26827, B2 => 
                           n21000, ZN => n23333);
   U22854 : OAI221_X1 port map( B1 => n9597, B2 => n26845, C1 => n20799, C2 => 
                           n26839, A => n23315, ZN => n23310);
   U22855 : AOI22_X1 port map( A1 => n26833, A2 => n25876, B1 => n26827, B2 => 
                           n20999, ZN => n23315);
   U22856 : OAI221_X1 port map( B1 => n9596, B2 => n26846, C1 => n20798, C2 => 
                           n26840, A => n23297, ZN => n23292);
   U22857 : AOI22_X1 port map( A1 => n26834, A2 => n25881, B1 => n26828, B2 => 
                           n20998, ZN => n23297);
   U22858 : OAI221_X1 port map( B1 => n9595, B2 => n26846, C1 => n20797, C2 => 
                           n26840, A => n23279, ZN => n23274);
   U22859 : AOI22_X1 port map( A1 => n26834, A2 => n25886, B1 => n26828, B2 => 
                           n20997, ZN => n23279);
   U22860 : OAI221_X1 port map( B1 => n9594, B2 => n26846, C1 => n20796, C2 => 
                           n26840, A => n23261, ZN => n23256);
   U22861 : AOI22_X1 port map( A1 => n26834, A2 => n25891, B1 => n26828, B2 => 
                           n20996, ZN => n23261);
   U22862 : OAI221_X1 port map( B1 => n9593, B2 => n26846, C1 => n20795, C2 => 
                           n26840, A => n23243, ZN => n23238);
   U22863 : AOI22_X1 port map( A1 => n26834, A2 => n25896, B1 => n26828, B2 => 
                           n20995, ZN => n23243);
   U22864 : OAI221_X1 port map( B1 => n9592, B2 => n26846, C1 => n20794, C2 => 
                           n26840, A => n23225, ZN => n23220);
   U22865 : AOI22_X1 port map( A1 => n26834, A2 => n25901, B1 => n26828, B2 => 
                           n20994, ZN => n23225);
   U22866 : OAI221_X1 port map( B1 => n9591, B2 => n26846, C1 => n20793, C2 => 
                           n26840, A => n23207, ZN => n23202);
   U22867 : AOI22_X1 port map( A1 => n26834, A2 => n25906, B1 => n26828, B2 => 
                           n20993, ZN => n23207);
   U22868 : OAI221_X1 port map( B1 => n9590, B2 => n26846, C1 => n20792, C2 => 
                           n26840, A => n23189, ZN => n23184);
   U22869 : AOI22_X1 port map( A1 => n26834, A2 => n25911, B1 => n26828, B2 => 
                           n20992, ZN => n23189);
   U22870 : OAI221_X1 port map( B1 => n9589, B2 => n26846, C1 => n20791, C2 => 
                           n26840, A => n23171, ZN => n23166);
   U22871 : AOI22_X1 port map( A1 => n26834, A2 => n25916, B1 => n26828, B2 => 
                           n20991, ZN => n23171);
   U22872 : OAI221_X1 port map( B1 => n9588, B2 => n26846, C1 => n20790, C2 => 
                           n26840, A => n23153, ZN => n23148);
   U22873 : AOI22_X1 port map( A1 => n26834, A2 => n25921, B1 => n26828, B2 => 
                           n20990, ZN => n23153);
   U22874 : OAI221_X1 port map( B1 => n9587, B2 => n26846, C1 => n20789, C2 => 
                           n26840, A => n23135, ZN => n23130);
   U22875 : AOI22_X1 port map( A1 => n26834, A2 => n25926, B1 => n26828, B2 => 
                           n20989, ZN => n23135);
   U22876 : OAI221_X1 port map( B1 => n9586, B2 => n26846, C1 => n20788, C2 => 
                           n26840, A => n23117, ZN => n23112);
   U22877 : AOI22_X1 port map( A1 => n26834, A2 => n25931, B1 => n26828, B2 => 
                           n20988, ZN => n23117);
   U22878 : OAI221_X1 port map( B1 => n9585, B2 => n26846, C1 => n20787, C2 => 
                           n26840, A => n23099, ZN => n23094);
   U22879 : AOI22_X1 port map( A1 => n26834, A2 => n25936, B1 => n26828, B2 => 
                           n20987, ZN => n23099);
   U22880 : OAI221_X1 port map( B1 => n9569, B2 => n26623, C1 => n21155, C2 => 
                           n26617, A => n23986, ZN => n23971);
   U22881 : AOI22_X1 port map( A1 => n26611, A2 => n25696, B1 => n26605, B2 => 
                           n20963, ZN => n23986);
   U22882 : OAI221_X1 port map( B1 => n9572, B2 => n26623, C1 => n20774, C2 => 
                           n26617, A => n24064, ZN => n24059);
   U22883 : AOI22_X1 port map( A1 => n26611, A2 => n25681, B1 => n26605, B2 => 
                           n20966, ZN => n24064);
   U22884 : OAI221_X1 port map( B1 => n9571, B2 => n26623, C1 => n20773, C2 => 
                           n26617, A => n24046, ZN => n24041);
   U22885 : AOI22_X1 port map( A1 => n26611, A2 => n25686, B1 => n26605, B2 => 
                           n20965, ZN => n24046);
   U22886 : OAI221_X1 port map( B1 => n9570, B2 => n26623, C1 => n20772, C2 => 
                           n26617, A => n24028, ZN => n24023);
   U22887 : AOI22_X1 port map( A1 => n26611, A2 => n25691, B1 => n26605, B2 => 
                           n20964, ZN => n24028);
   U22888 : OAI221_X1 port map( B1 => n9572, B2 => n26848, C1 => n20774, C2 => 
                           n26842, A => n22865, ZN => n22860);
   U22889 : AOI22_X1 port map( A1 => n26836, A2 => n25681, B1 => n26830, B2 => 
                           n20966, ZN => n22865);
   U22890 : OAI221_X1 port map( B1 => n9571, B2 => n26848, C1 => n20773, C2 => 
                           n26842, A => n22847, ZN => n22842);
   U22891 : AOI22_X1 port map( A1 => n26836, A2 => n25686, B1 => n26830, B2 => 
                           n20965, ZN => n22847);
   U22892 : OAI221_X1 port map( B1 => n9570, B2 => n26848, C1 => n20772, C2 => 
                           n26842, A => n22829, ZN => n22824);
   U22893 : AOI22_X1 port map( A1 => n26836, A2 => n25691, B1 => n26830, B2 => 
                           n20964, ZN => n22829);
   U22894 : OAI221_X1 port map( B1 => n9569, B2 => n26848, C1 => n21155, C2 => 
                           n26842, A => n22787, ZN => n22772);
   U22895 : AOI22_X1 port map( A1 => n26836, A2 => n25696, B1 => n26830, B2 => 
                           n20963, ZN => n22787);
   U22896 : OAI221_X1 port map( B1 => n21747, B2 => n26595, C1 => n22367, C2 =>
                           n26589, A => n24929, ZN => n24922);
   U22897 : AOI222_X1 port map( A1 => n26583, A2 => n25762, B1 => n26577, B2 =>
                           n21082, C1 => n26571, C2 => n21142, ZN => n24929);
   U22898 : OAI221_X1 port map( B1 => n21746, B2 => n26595, C1 => n22366, C2 =>
                           n26589, A => n24911, ZN => n24904);
   U22899 : AOI222_X1 port map( A1 => n26583, A2 => n25767, B1 => n26577, B2 =>
                           n21081, C1 => n26571, C2 => n21141, ZN => n24911);
   U22900 : OAI221_X1 port map( B1 => n21745, B2 => n26595, C1 => n22365, C2 =>
                           n26589, A => n24893, ZN => n24886);
   U22901 : AOI222_X1 port map( A1 => n26583, A2 => n25772, B1 => n26577, B2 =>
                           n21080, C1 => n26571, C2 => n21140, ZN => n24893);
   U22902 : OAI221_X1 port map( B1 => n21744, B2 => n26595, C1 => n22364, C2 =>
                           n26589, A => n24875, ZN => n24868);
   U22903 : AOI222_X1 port map( A1 => n26583, A2 => n25777, B1 => n26577, B2 =>
                           n21079, C1 => n26571, C2 => n21139, ZN => n24875);
   U22904 : OAI221_X1 port map( B1 => n21743, B2 => n26595, C1 => n22363, C2 =>
                           n26589, A => n24857, ZN => n24850);
   U22905 : AOI222_X1 port map( A1 => n26583, A2 => n25782, B1 => n26577, B2 =>
                           n21078, C1 => n26571, C2 => n21138, ZN => n24857);
   U22906 : OAI221_X1 port map( B1 => n21742, B2 => n26595, C1 => n22362, C2 =>
                           n26589, A => n24839, ZN => n24832);
   U22907 : AOI222_X1 port map( A1 => n26583, A2 => n25787, B1 => n26577, B2 =>
                           n21077, C1 => n26571, C2 => n21137, ZN => n24839);
   U22908 : OAI221_X1 port map( B1 => n21741, B2 => n26595, C1 => n22361, C2 =>
                           n26589, A => n24821, ZN => n24814);
   U22909 : AOI222_X1 port map( A1 => n26583, A2 => n25792, B1 => n26577, B2 =>
                           n21076, C1 => n26571, C2 => n21136, ZN => n24821);
   U22910 : OAI221_X1 port map( B1 => n21740, B2 => n26595, C1 => n22360, C2 =>
                           n26589, A => n24803, ZN => n24796);
   U22911 : AOI222_X1 port map( A1 => n26583, A2 => n25797, B1 => n26577, B2 =>
                           n21075, C1 => n26571, C2 => n21135, ZN => n24803);
   U22912 : OAI221_X1 port map( B1 => n21739, B2 => n26595, C1 => n22359, C2 =>
                           n26589, A => n24785, ZN => n24778);
   U22913 : AOI222_X1 port map( A1 => n26583, A2 => n25802, B1 => n26577, B2 =>
                           n21074, C1 => n26571, C2 => n21134, ZN => n24785);
   U22914 : OAI221_X1 port map( B1 => n21738, B2 => n26595, C1 => n22358, C2 =>
                           n26589, A => n24767, ZN => n24760);
   U22915 : AOI222_X1 port map( A1 => n26583, A2 => n25807, B1 => n26577, B2 =>
                           n21073, C1 => n26571, C2 => n21133, ZN => n24767);
   U22916 : OAI221_X1 port map( B1 => n21737, B2 => n26595, C1 => n22357, C2 =>
                           n26589, A => n24749, ZN => n24742);
   U22917 : AOI222_X1 port map( A1 => n26583, A2 => n25812, B1 => n26577, B2 =>
                           n21072, C1 => n26571, C2 => n21132, ZN => n24749);
   U22918 : OAI221_X1 port map( B1 => n21736, B2 => n26595, C1 => n22356, C2 =>
                           n26589, A => n24731, ZN => n24724);
   U22919 : AOI222_X1 port map( A1 => n26583, A2 => n25817, B1 => n26577, B2 =>
                           n21071, C1 => n26571, C2 => n21131, ZN => n24731);
   U22920 : OAI221_X1 port map( B1 => n21735, B2 => n26596, C1 => n22355, C2 =>
                           n26590, A => n24713, ZN => n24706);
   U22921 : AOI222_X1 port map( A1 => n26584, A2 => n25822, B1 => n26578, B2 =>
                           n21070, C1 => n26572, C2 => n21130, ZN => n24713);
   U22922 : OAI221_X1 port map( B1 => n21734, B2 => n26596, C1 => n22354, C2 =>
                           n26590, A => n24695, ZN => n24688);
   U22923 : AOI222_X1 port map( A1 => n26584, A2 => n25827, B1 => n26578, B2 =>
                           n21069, C1 => n26572, C2 => n21129, ZN => n24695);
   U22924 : OAI221_X1 port map( B1 => n21733, B2 => n26596, C1 => n22353, C2 =>
                           n26590, A => n24677, ZN => n24670);
   U22925 : AOI222_X1 port map( A1 => n26584, A2 => n25832, B1 => n26578, B2 =>
                           n21068, C1 => n26572, C2 => n21128, ZN => n24677);
   U22926 : OAI221_X1 port map( B1 => n21732, B2 => n26596, C1 => n22352, C2 =>
                           n26590, A => n24659, ZN => n24652);
   U22927 : AOI222_X1 port map( A1 => n26584, A2 => n25837, B1 => n26578, B2 =>
                           n21067, C1 => n26572, C2 => n21127, ZN => n24659);
   U22928 : OAI221_X1 port map( B1 => n21731, B2 => n26596, C1 => n22351, C2 =>
                           n26590, A => n24641, ZN => n24634);
   U22929 : AOI222_X1 port map( A1 => n26584, A2 => n25842, B1 => n26578, B2 =>
                           n21066, C1 => n26572, C2 => n21126, ZN => n24641);
   U22930 : OAI221_X1 port map( B1 => n21730, B2 => n26596, C1 => n22350, C2 =>
                           n26590, A => n24623, ZN => n24616);
   U22931 : AOI222_X1 port map( A1 => n26584, A2 => n25847, B1 => n26578, B2 =>
                           n21065, C1 => n26572, C2 => n21125, ZN => n24623);
   U22932 : OAI221_X1 port map( B1 => n21729, B2 => n26596, C1 => n22349, C2 =>
                           n26590, A => n24605, ZN => n24598);
   U22933 : AOI222_X1 port map( A1 => n26584, A2 => n25852, B1 => n26578, B2 =>
                           n21064, C1 => n26572, C2 => n21124, ZN => n24605);
   U22934 : OAI221_X1 port map( B1 => n21728, B2 => n26596, C1 => n22348, C2 =>
                           n26590, A => n24587, ZN => n24580);
   U22935 : AOI222_X1 port map( A1 => n26584, A2 => n25857, B1 => n26578, B2 =>
                           n21063, C1 => n26572, C2 => n21123, ZN => n24587);
   U22936 : OAI221_X1 port map( B1 => n21727, B2 => n26596, C1 => n22347, C2 =>
                           n26590, A => n24569, ZN => n24562);
   U22937 : AOI222_X1 port map( A1 => n26584, A2 => n25862, B1 => n26578, B2 =>
                           n21062, C1 => n26572, C2 => n21122, ZN => n24569);
   U22938 : OAI221_X1 port map( B1 => n21726, B2 => n26596, C1 => n22346, C2 =>
                           n26590, A => n24551, ZN => n24544);
   U22939 : AOI222_X1 port map( A1 => n26584, A2 => n25867, B1 => n26578, B2 =>
                           n21061, C1 => n26572, C2 => n21121, ZN => n24551);
   U22940 : OAI221_X1 port map( B1 => n21725, B2 => n26596, C1 => n22345, C2 =>
                           n26590, A => n24533, ZN => n24526);
   U22941 : AOI222_X1 port map( A1 => n26584, A2 => n25872, B1 => n26578, B2 =>
                           n21060, C1 => n26572, C2 => n21120, ZN => n24533);
   U22942 : OAI221_X1 port map( B1 => n21724, B2 => n26596, C1 => n22344, C2 =>
                           n26590, A => n24515, ZN => n24508);
   U22943 : AOI222_X1 port map( A1 => n26584, A2 => n25877, B1 => n26578, B2 =>
                           n21059, C1 => n26572, C2 => n21119, ZN => n24515);
   U22944 : OAI221_X1 port map( B1 => n21723, B2 => n26597, C1 => n22343, C2 =>
                           n26591, A => n24497, ZN => n24490);
   U22945 : AOI222_X1 port map( A1 => n26585, A2 => n25882, B1 => n26579, B2 =>
                           n21058, C1 => n26573, C2 => n21118, ZN => n24497);
   U22946 : OAI221_X1 port map( B1 => n21722, B2 => n26597, C1 => n22342, C2 =>
                           n26591, A => n24479, ZN => n24472);
   U22947 : AOI222_X1 port map( A1 => n26585, A2 => n25887, B1 => n26579, B2 =>
                           n21057, C1 => n26573, C2 => n21117, ZN => n24479);
   U22948 : OAI221_X1 port map( B1 => n21721, B2 => n26597, C1 => n22341, C2 =>
                           n26591, A => n24461, ZN => n24454);
   U22949 : AOI222_X1 port map( A1 => n26585, A2 => n25892, B1 => n26579, B2 =>
                           n21056, C1 => n26573, C2 => n21116, ZN => n24461);
   U22950 : OAI221_X1 port map( B1 => n21720, B2 => n26597, C1 => n22340, C2 =>
                           n26591, A => n24443, ZN => n24436);
   U22951 : AOI222_X1 port map( A1 => n26585, A2 => n25897, B1 => n26579, B2 =>
                           n21055, C1 => n26573, C2 => n21115, ZN => n24443);
   U22952 : OAI221_X1 port map( B1 => n21719, B2 => n26597, C1 => n22339, C2 =>
                           n26591, A => n24425, ZN => n24418);
   U22953 : AOI222_X1 port map( A1 => n26585, A2 => n25902, B1 => n26579, B2 =>
                           n21054, C1 => n26573, C2 => n21114, ZN => n24425);
   U22954 : OAI221_X1 port map( B1 => n21718, B2 => n26597, C1 => n22338, C2 =>
                           n26591, A => n24407, ZN => n24400);
   U22955 : AOI222_X1 port map( A1 => n26585, A2 => n25907, B1 => n26579, B2 =>
                           n21053, C1 => n26573, C2 => n21113, ZN => n24407);
   U22956 : OAI221_X1 port map( B1 => n21717, B2 => n26597, C1 => n22337, C2 =>
                           n26591, A => n24389, ZN => n24382);
   U22957 : AOI222_X1 port map( A1 => n26585, A2 => n25912, B1 => n26579, B2 =>
                           n21052, C1 => n26573, C2 => n21112, ZN => n24389);
   U22958 : OAI221_X1 port map( B1 => n21716, B2 => n26597, C1 => n22336, C2 =>
                           n26591, A => n24371, ZN => n24364);
   U22959 : AOI222_X1 port map( A1 => n26585, A2 => n25917, B1 => n26579, B2 =>
                           n21051, C1 => n26573, C2 => n21111, ZN => n24371);
   U22960 : OAI221_X1 port map( B1 => n21715, B2 => n26597, C1 => n22335, C2 =>
                           n26591, A => n24353, ZN => n24346);
   U22961 : AOI222_X1 port map( A1 => n26585, A2 => n25922, B1 => n26579, B2 =>
                           n21050, C1 => n26573, C2 => n21110, ZN => n24353);
   U22962 : OAI221_X1 port map( B1 => n21714, B2 => n26597, C1 => n22334, C2 =>
                           n26591, A => n24335, ZN => n24328);
   U22963 : AOI222_X1 port map( A1 => n26585, A2 => n25927, B1 => n26579, B2 =>
                           n21049, C1 => n26573, C2 => n21109, ZN => n24335);
   U22964 : OAI221_X1 port map( B1 => n21713, B2 => n26597, C1 => n22333, C2 =>
                           n26591, A => n24317, ZN => n24310);
   U22965 : AOI222_X1 port map( A1 => n26585, A2 => n25932, B1 => n26579, B2 =>
                           n21048, C1 => n26573, C2 => n21108, ZN => n24317);
   U22966 : OAI221_X1 port map( B1 => n21712, B2 => n26597, C1 => n22332, C2 =>
                           n26591, A => n24299, ZN => n24292);
   U22967 : AOI222_X1 port map( A1 => n26585, A2 => n25937, B1 => n26579, B2 =>
                           n21047, C1 => n26573, C2 => n21107, ZN => n24299);
   U22968 : OAI221_X1 port map( B1 => n21711, B2 => n26598, C1 => n22331, C2 =>
                           n26592, A => n24281, ZN => n24274);
   U22969 : AOI222_X1 port map( A1 => n26586, A2 => n25942, B1 => n26580, B2 =>
                           n21046, C1 => n26574, C2 => n21106, ZN => n24281);
   U22970 : OAI221_X1 port map( B1 => n21710, B2 => n26598, C1 => n22330, C2 =>
                           n26592, A => n24263, ZN => n24256);
   U22971 : AOI222_X1 port map( A1 => n26586, A2 => n25947, B1 => n26580, B2 =>
                           n21045, C1 => n26574, C2 => n21105, ZN => n24263);
   U22972 : OAI221_X1 port map( B1 => n21709, B2 => n26598, C1 => n22329, C2 =>
                           n26592, A => n24245, ZN => n24238);
   U22973 : AOI222_X1 port map( A1 => n26586, A2 => n25952, B1 => n26580, B2 =>
                           n21044, C1 => n26574, C2 => n21104, ZN => n24245);
   U22974 : OAI221_X1 port map( B1 => n21708, B2 => n26598, C1 => n22328, C2 =>
                           n26592, A => n24227, ZN => n24220);
   U22975 : AOI222_X1 port map( A1 => n26586, A2 => n25957, B1 => n26580, B2 =>
                           n21043, C1 => n26574, C2 => n21103, ZN => n24227);
   U22976 : OAI221_X1 port map( B1 => n21707, B2 => n26598, C1 => n22327, C2 =>
                           n26592, A => n24209, ZN => n24202);
   U22977 : AOI222_X1 port map( A1 => n26586, A2 => n25962, B1 => n26580, B2 =>
                           n21042, C1 => n26574, C2 => n21102, ZN => n24209);
   U22978 : OAI221_X1 port map( B1 => n21706, B2 => n26598, C1 => n22326, C2 =>
                           n26592, A => n24191, ZN => n24184);
   U22979 : AOI222_X1 port map( A1 => n26586, A2 => n25967, B1 => n26580, B2 =>
                           n21041, C1 => n26574, C2 => n21101, ZN => n24191);
   U22980 : OAI221_X1 port map( B1 => n21705, B2 => n26598, C1 => n22325, C2 =>
                           n26592, A => n24173, ZN => n24166);
   U22981 : AOI222_X1 port map( A1 => n26586, A2 => n25972, B1 => n26580, B2 =>
                           n21040, C1 => n26574, C2 => n21100, ZN => n24173);
   U22982 : OAI221_X1 port map( B1 => n21704, B2 => n26598, C1 => n22324, C2 =>
                           n26592, A => n24155, ZN => n24148);
   U22983 : AOI222_X1 port map( A1 => n26586, A2 => n25977, B1 => n26580, B2 =>
                           n21039, C1 => n26574, C2 => n21099, ZN => n24155);
   U22984 : OAI221_X1 port map( B1 => n21703, B2 => n26598, C1 => n22323, C2 =>
                           n26592, A => n24137, ZN => n24130);
   U22985 : AOI222_X1 port map( A1 => n26586, A2 => n25982, B1 => n26580, B2 =>
                           n21038, C1 => n26574, C2 => n21098, ZN => n24137);
   U22986 : OAI221_X1 port map( B1 => n21702, B2 => n26598, C1 => n22322, C2 =>
                           n26592, A => n24119, ZN => n24112);
   U22987 : AOI222_X1 port map( A1 => n26586, A2 => n25987, B1 => n26580, B2 =>
                           n21037, C1 => n26574, C2 => n21097, ZN => n24119);
   U22988 : OAI221_X1 port map( B1 => n21701, B2 => n26598, C1 => n22321, C2 =>
                           n26592, A => n24101, ZN => n24094);
   U22989 : AOI222_X1 port map( A1 => n26586, A2 => n25992, B1 => n26580, B2 =>
                           n21036, C1 => n26574, C2 => n21096, ZN => n24101);
   U22990 : OAI221_X1 port map( B1 => n21700, B2 => n26598, C1 => n22320, C2 =>
                           n26592, A => n24083, ZN => n24076);
   U22991 : AOI222_X1 port map( A1 => n26586, A2 => n25997, B1 => n26580, B2 =>
                           n21035, C1 => n26574, C2 => n21095, ZN => n24083);
   U22992 : OAI221_X1 port map( B1 => n21747, B2 => n26820, C1 => n22367, C2 =>
                           n26814, A => n23730, ZN => n23723);
   U22993 : AOI222_X1 port map( A1 => n26808, A2 => n25762, B1 => n26802, B2 =>
                           n21082, C1 => n26796, C2 => n21142, ZN => n23730);
   U22994 : OAI221_X1 port map( B1 => n21746, B2 => n26820, C1 => n22366, C2 =>
                           n26814, A => n23712, ZN => n23705);
   U22995 : AOI222_X1 port map( A1 => n26808, A2 => n25767, B1 => n26802, B2 =>
                           n21081, C1 => n26796, C2 => n21141, ZN => n23712);
   U22996 : OAI221_X1 port map( B1 => n21745, B2 => n26820, C1 => n22365, C2 =>
                           n26814, A => n23694, ZN => n23687);
   U22997 : AOI222_X1 port map( A1 => n26808, A2 => n25772, B1 => n26802, B2 =>
                           n21080, C1 => n26796, C2 => n21140, ZN => n23694);
   U22998 : OAI221_X1 port map( B1 => n21744, B2 => n26820, C1 => n22364, C2 =>
                           n26814, A => n23676, ZN => n23669);
   U22999 : AOI222_X1 port map( A1 => n26808, A2 => n25777, B1 => n26802, B2 =>
                           n21079, C1 => n26796, C2 => n21139, ZN => n23676);
   U23000 : OAI221_X1 port map( B1 => n21743, B2 => n26820, C1 => n22363, C2 =>
                           n26814, A => n23658, ZN => n23651);
   U23001 : AOI222_X1 port map( A1 => n26808, A2 => n25782, B1 => n26802, B2 =>
                           n21078, C1 => n26796, C2 => n21138, ZN => n23658);
   U23002 : OAI221_X1 port map( B1 => n21742, B2 => n26820, C1 => n22362, C2 =>
                           n26814, A => n23640, ZN => n23633);
   U23003 : AOI222_X1 port map( A1 => n26808, A2 => n25787, B1 => n26802, B2 =>
                           n21077, C1 => n26796, C2 => n21137, ZN => n23640);
   U23004 : OAI221_X1 port map( B1 => n21741, B2 => n26820, C1 => n22361, C2 =>
                           n26814, A => n23622, ZN => n23615);
   U23005 : AOI222_X1 port map( A1 => n26808, A2 => n25792, B1 => n26802, B2 =>
                           n21076, C1 => n26796, C2 => n21136, ZN => n23622);
   U23006 : OAI221_X1 port map( B1 => n21740, B2 => n26820, C1 => n22360, C2 =>
                           n26814, A => n23604, ZN => n23597);
   U23007 : AOI222_X1 port map( A1 => n26808, A2 => n25797, B1 => n26802, B2 =>
                           n21075, C1 => n26796, C2 => n21135, ZN => n23604);
   U23008 : OAI221_X1 port map( B1 => n21739, B2 => n26820, C1 => n22359, C2 =>
                           n26814, A => n23586, ZN => n23579);
   U23009 : AOI222_X1 port map( A1 => n26808, A2 => n25802, B1 => n26802, B2 =>
                           n21074, C1 => n26796, C2 => n21134, ZN => n23586);
   U23010 : OAI221_X1 port map( B1 => n21738, B2 => n26820, C1 => n22358, C2 =>
                           n26814, A => n23568, ZN => n23561);
   U23011 : AOI222_X1 port map( A1 => n26808, A2 => n25807, B1 => n26802, B2 =>
                           n21073, C1 => n26796, C2 => n21133, ZN => n23568);
   U23012 : OAI221_X1 port map( B1 => n21737, B2 => n26820, C1 => n22357, C2 =>
                           n26814, A => n23550, ZN => n23543);
   U23013 : AOI222_X1 port map( A1 => n26808, A2 => n25812, B1 => n26802, B2 =>
                           n21072, C1 => n26796, C2 => n21132, ZN => n23550);
   U23014 : OAI221_X1 port map( B1 => n21736, B2 => n26820, C1 => n22356, C2 =>
                           n26814, A => n23532, ZN => n23525);
   U23015 : AOI222_X1 port map( A1 => n26808, A2 => n25817, B1 => n26802, B2 =>
                           n21071, C1 => n26796, C2 => n21131, ZN => n23532);
   U23016 : OAI221_X1 port map( B1 => n21735, B2 => n26821, C1 => n22355, C2 =>
                           n26815, A => n23514, ZN => n23507);
   U23017 : AOI222_X1 port map( A1 => n26809, A2 => n25822, B1 => n26803, B2 =>
                           n21070, C1 => n26797, C2 => n21130, ZN => n23514);
   U23018 : OAI221_X1 port map( B1 => n21734, B2 => n26821, C1 => n22354, C2 =>
                           n26815, A => n23496, ZN => n23489);
   U23019 : AOI222_X1 port map( A1 => n26809, A2 => n25827, B1 => n26803, B2 =>
                           n21069, C1 => n26797, C2 => n21129, ZN => n23496);
   U23020 : OAI221_X1 port map( B1 => n21733, B2 => n26821, C1 => n22353, C2 =>
                           n26815, A => n23478, ZN => n23471);
   U23021 : AOI222_X1 port map( A1 => n26809, A2 => n25832, B1 => n26803, B2 =>
                           n21068, C1 => n26797, C2 => n21128, ZN => n23478);
   U23022 : OAI221_X1 port map( B1 => n21732, B2 => n26821, C1 => n22352, C2 =>
                           n26815, A => n23460, ZN => n23453);
   U23023 : AOI222_X1 port map( A1 => n26809, A2 => n25837, B1 => n26803, B2 =>
                           n21067, C1 => n26797, C2 => n21127, ZN => n23460);
   U23024 : OAI221_X1 port map( B1 => n21731, B2 => n26821, C1 => n22351, C2 =>
                           n26815, A => n23442, ZN => n23435);
   U23025 : AOI222_X1 port map( A1 => n26809, A2 => n25842, B1 => n26803, B2 =>
                           n21066, C1 => n26797, C2 => n21126, ZN => n23442);
   U23026 : OAI221_X1 port map( B1 => n21730, B2 => n26821, C1 => n22350, C2 =>
                           n26815, A => n23424, ZN => n23417);
   U23027 : AOI222_X1 port map( A1 => n26809, A2 => n25847, B1 => n26803, B2 =>
                           n21065, C1 => n26797, C2 => n21125, ZN => n23424);
   U23028 : OAI221_X1 port map( B1 => n21729, B2 => n26821, C1 => n22349, C2 =>
                           n26815, A => n23406, ZN => n23399);
   U23029 : AOI222_X1 port map( A1 => n26809, A2 => n25852, B1 => n26803, B2 =>
                           n21064, C1 => n26797, C2 => n21124, ZN => n23406);
   U23030 : OAI221_X1 port map( B1 => n21728, B2 => n26821, C1 => n22348, C2 =>
                           n26815, A => n23388, ZN => n23381);
   U23031 : AOI222_X1 port map( A1 => n26809, A2 => n25857, B1 => n26803, B2 =>
                           n21063, C1 => n26797, C2 => n21123, ZN => n23388);
   U23032 : OAI221_X1 port map( B1 => n21727, B2 => n26821, C1 => n22347, C2 =>
                           n26815, A => n23370, ZN => n23363);
   U23033 : AOI222_X1 port map( A1 => n26809, A2 => n25862, B1 => n26803, B2 =>
                           n21062, C1 => n26797, C2 => n21122, ZN => n23370);
   U23034 : OAI221_X1 port map( B1 => n21726, B2 => n26821, C1 => n22346, C2 =>
                           n26815, A => n23352, ZN => n23345);
   U23035 : AOI222_X1 port map( A1 => n26809, A2 => n25867, B1 => n26803, B2 =>
                           n21061, C1 => n26797, C2 => n21121, ZN => n23352);
   U23036 : OAI221_X1 port map( B1 => n21725, B2 => n26821, C1 => n22345, C2 =>
                           n26815, A => n23334, ZN => n23327);
   U23037 : AOI222_X1 port map( A1 => n26809, A2 => n25872, B1 => n26803, B2 =>
                           n21060, C1 => n26797, C2 => n21120, ZN => n23334);
   U23038 : OAI221_X1 port map( B1 => n21724, B2 => n26821, C1 => n22344, C2 =>
                           n26815, A => n23316, ZN => n23309);
   U23039 : AOI222_X1 port map( A1 => n26809, A2 => n25877, B1 => n26803, B2 =>
                           n21059, C1 => n26797, C2 => n21119, ZN => n23316);
   U23040 : OAI221_X1 port map( B1 => n21723, B2 => n26822, C1 => n22343, C2 =>
                           n26816, A => n23298, ZN => n23291);
   U23041 : AOI222_X1 port map( A1 => n26810, A2 => n25882, B1 => n26804, B2 =>
                           n21058, C1 => n26798, C2 => n21118, ZN => n23298);
   U23042 : OAI221_X1 port map( B1 => n21722, B2 => n26822, C1 => n22342, C2 =>
                           n26816, A => n23280, ZN => n23273);
   U23043 : AOI222_X1 port map( A1 => n26810, A2 => n25887, B1 => n26804, B2 =>
                           n21057, C1 => n26798, C2 => n21117, ZN => n23280);
   U23044 : OAI221_X1 port map( B1 => n21721, B2 => n26822, C1 => n22341, C2 =>
                           n26816, A => n23262, ZN => n23255);
   U23045 : AOI222_X1 port map( A1 => n26810, A2 => n25892, B1 => n26804, B2 =>
                           n21056, C1 => n26798, C2 => n21116, ZN => n23262);
   U23046 : OAI221_X1 port map( B1 => n21720, B2 => n26822, C1 => n22340, C2 =>
                           n26816, A => n23244, ZN => n23237);
   U23047 : AOI222_X1 port map( A1 => n26810, A2 => n25897, B1 => n26804, B2 =>
                           n21055, C1 => n26798, C2 => n21115, ZN => n23244);
   U23048 : OAI221_X1 port map( B1 => n21719, B2 => n26822, C1 => n22339, C2 =>
                           n26816, A => n23226, ZN => n23219);
   U23049 : AOI222_X1 port map( A1 => n26810, A2 => n25902, B1 => n26804, B2 =>
                           n21054, C1 => n26798, C2 => n21114, ZN => n23226);
   U23050 : OAI221_X1 port map( B1 => n21718, B2 => n26822, C1 => n22338, C2 =>
                           n26816, A => n23208, ZN => n23201);
   U23051 : AOI222_X1 port map( A1 => n26810, A2 => n25907, B1 => n26804, B2 =>
                           n21053, C1 => n26798, C2 => n21113, ZN => n23208);
   U23052 : OAI221_X1 port map( B1 => n21717, B2 => n26822, C1 => n22337, C2 =>
                           n26816, A => n23190, ZN => n23183);
   U23053 : AOI222_X1 port map( A1 => n26810, A2 => n25912, B1 => n26804, B2 =>
                           n21052, C1 => n26798, C2 => n21112, ZN => n23190);
   U23054 : OAI221_X1 port map( B1 => n21716, B2 => n26822, C1 => n22336, C2 =>
                           n26816, A => n23172, ZN => n23165);
   U23055 : AOI222_X1 port map( A1 => n26810, A2 => n25917, B1 => n26804, B2 =>
                           n21051, C1 => n26798, C2 => n21111, ZN => n23172);
   U23056 : OAI221_X1 port map( B1 => n21715, B2 => n26822, C1 => n22335, C2 =>
                           n26816, A => n23154, ZN => n23147);
   U23057 : AOI222_X1 port map( A1 => n26810, A2 => n25922, B1 => n26804, B2 =>
                           n21050, C1 => n26798, C2 => n21110, ZN => n23154);
   U23058 : OAI221_X1 port map( B1 => n21714, B2 => n26822, C1 => n22334, C2 =>
                           n26816, A => n23136, ZN => n23129);
   U23059 : AOI222_X1 port map( A1 => n26810, A2 => n25927, B1 => n26804, B2 =>
                           n21049, C1 => n26798, C2 => n21109, ZN => n23136);
   U23060 : OAI221_X1 port map( B1 => n21713, B2 => n26822, C1 => n22333, C2 =>
                           n26816, A => n23118, ZN => n23111);
   U23061 : AOI222_X1 port map( A1 => n26810, A2 => n25932, B1 => n26804, B2 =>
                           n21048, C1 => n26798, C2 => n21108, ZN => n23118);
   U23062 : OAI221_X1 port map( B1 => n21712, B2 => n26822, C1 => n22332, C2 =>
                           n26816, A => n23100, ZN => n23093);
   U23063 : AOI222_X1 port map( A1 => n26810, A2 => n25937, B1 => n26804, B2 =>
                           n21047, C1 => n26798, C2 => n21107, ZN => n23100);
   U23064 : OAI221_X1 port map( B1 => n21711, B2 => n26823, C1 => n22331, C2 =>
                           n26817, A => n23082, ZN => n23075);
   U23065 : AOI222_X1 port map( A1 => n26811, A2 => n25942, B1 => n26805, B2 =>
                           n21046, C1 => n26799, C2 => n21106, ZN => n23082);
   U23066 : OAI221_X1 port map( B1 => n21710, B2 => n26823, C1 => n22330, C2 =>
                           n26817, A => n23064, ZN => n23057);
   U23067 : AOI222_X1 port map( A1 => n26811, A2 => n25947, B1 => n26805, B2 =>
                           n21045, C1 => n26799, C2 => n21105, ZN => n23064);
   U23068 : OAI221_X1 port map( B1 => n21709, B2 => n26823, C1 => n22329, C2 =>
                           n26817, A => n23046, ZN => n23039);
   U23069 : AOI222_X1 port map( A1 => n26811, A2 => n25952, B1 => n26805, B2 =>
                           n21044, C1 => n26799, C2 => n21104, ZN => n23046);
   U23070 : OAI221_X1 port map( B1 => n21708, B2 => n26823, C1 => n22328, C2 =>
                           n26817, A => n23028, ZN => n23021);
   U23071 : AOI222_X1 port map( A1 => n26811, A2 => n25957, B1 => n26805, B2 =>
                           n21043, C1 => n26799, C2 => n21103, ZN => n23028);
   U23072 : OAI221_X1 port map( B1 => n21707, B2 => n26823, C1 => n22327, C2 =>
                           n26817, A => n23010, ZN => n23003);
   U23073 : AOI222_X1 port map( A1 => n26811, A2 => n25962, B1 => n26805, B2 =>
                           n21042, C1 => n26799, C2 => n21102, ZN => n23010);
   U23074 : OAI221_X1 port map( B1 => n21706, B2 => n26823, C1 => n22326, C2 =>
                           n26817, A => n22992, ZN => n22985);
   U23075 : AOI222_X1 port map( A1 => n26811, A2 => n25967, B1 => n26805, B2 =>
                           n21041, C1 => n26799, C2 => n21101, ZN => n22992);
   U23076 : OAI221_X1 port map( B1 => n21705, B2 => n26823, C1 => n22325, C2 =>
                           n26817, A => n22974, ZN => n22967);
   U23077 : AOI222_X1 port map( A1 => n26811, A2 => n25972, B1 => n26805, B2 =>
                           n21040, C1 => n26799, C2 => n21100, ZN => n22974);
   U23078 : OAI221_X1 port map( B1 => n21704, B2 => n26823, C1 => n22324, C2 =>
                           n26817, A => n22956, ZN => n22949);
   U23079 : AOI222_X1 port map( A1 => n26811, A2 => n25977, B1 => n26805, B2 =>
                           n21039, C1 => n26799, C2 => n21099, ZN => n22956);
   U23080 : OAI221_X1 port map( B1 => n21703, B2 => n26823, C1 => n22323, C2 =>
                           n26817, A => n22938, ZN => n22931);
   U23081 : AOI222_X1 port map( A1 => n26811, A2 => n25982, B1 => n26805, B2 =>
                           n21038, C1 => n26799, C2 => n21098, ZN => n22938);
   U23082 : OAI221_X1 port map( B1 => n21702, B2 => n26823, C1 => n22322, C2 =>
                           n26817, A => n22920, ZN => n22913);
   U23083 : AOI222_X1 port map( A1 => n26811, A2 => n25987, B1 => n26805, B2 =>
                           n21037, C1 => n26799, C2 => n21097, ZN => n22920);
   U23084 : OAI221_X1 port map( B1 => n21701, B2 => n26823, C1 => n22321, C2 =>
                           n26817, A => n22902, ZN => n22895);
   U23085 : AOI222_X1 port map( A1 => n26811, A2 => n25992, B1 => n26805, B2 =>
                           n21036, C1 => n26799, C2 => n21096, ZN => n22902);
   U23086 : OAI221_X1 port map( B1 => n21700, B2 => n26823, C1 => n22320, C2 =>
                           n26817, A => n22884, ZN => n22877);
   U23087 : AOI222_X1 port map( A1 => n26811, A2 => n25997, B1 => n26805, B2 =>
                           n21035, C1 => n26799, C2 => n21095, ZN => n22884);
   U23088 : OAI221_X1 port map( B1 => n21508, B2 => n26476, C1 => n27473, C2 =>
                           n26470, A => n24016, ZN => n23995);
   U23089 : AOI222_X1 port map( A1 => n26464, A2 => n25558, B1 => n26458, B2 =>
                           n25574, C1 => n26452, C2 => n25582, ZN => n24016);
   U23090 : OAI221_X1 port map( B1 => n21511, B2 => n26476, C1 => n27464, C2 =>
                           n26470, A => n24073, ZN => n24066);
   U23091 : AOI222_X1 port map( A1 => n26464, A2 => n25555, B1 => n26458, B2 =>
                           n25571, C1 => n26452, C2 => n25579, ZN => n24073);
   U23092 : OAI221_X1 port map( B1 => n21510, B2 => n26476, C1 => n27467, C2 =>
                           n26470, A => n24055, ZN => n24048);
   U23093 : AOI222_X1 port map( A1 => n26464, A2 => n25556, B1 => n26458, B2 =>
                           n25572, C1 => n26452, C2 => n25580, ZN => n24055);
   U23094 : OAI221_X1 port map( B1 => n21509, B2 => n26476, C1 => n27470, C2 =>
                           n26470, A => n24037, ZN => n24030);
   U23095 : AOI222_X1 port map( A1 => n26464, A2 => n25557, B1 => n26458, B2 =>
                           n25573, C1 => n26452, C2 => n25581, ZN => n24037);
   U23096 : OAI221_X1 port map( B1 => n21511, B2 => n26701, C1 => n27464, C2 =>
                           n26695, A => n22874, ZN => n22867);
   U23097 : AOI222_X1 port map( A1 => n26689, A2 => n25555, B1 => n26683, B2 =>
                           n25571, C1 => n26677, C2 => n25579, ZN => n22874);
   U23098 : OAI221_X1 port map( B1 => n21510, B2 => n26701, C1 => n27467, C2 =>
                           n26695, A => n22856, ZN => n22849);
   U23099 : AOI222_X1 port map( A1 => n26689, A2 => n25556, B1 => n26683, B2 =>
                           n25572, C1 => n26677, C2 => n25580, ZN => n22856);
   U23100 : OAI221_X1 port map( B1 => n21509, B2 => n26701, C1 => n27470, C2 =>
                           n26695, A => n22838, ZN => n22831);
   U23101 : AOI222_X1 port map( A1 => n26689, A2 => n25557, B1 => n26683, B2 =>
                           n25573, C1 => n26677, C2 => n25581, ZN => n22838);
   U23102 : OAI221_X1 port map( B1 => n21508, B2 => n26701, C1 => n27473, C2 =>
                           n26695, A => n22817, ZN => n22796);
   U23103 : AOI222_X1 port map( A1 => n26689, A2 => n25558, B1 => n26683, B2 =>
                           n25574, C1 => n26677, C2 => n25582, ZN => n22817);
   U23104 : OAI221_X1 port map( B1 => n21488, B2 => n26599, C1 => n22248, C2 =>
                           n26593, A => n23991, ZN => n23970);
   U23105 : AOI222_X1 port map( A1 => n26587, A2 => n25697, B1 => n26581, B2 =>
                           n20967, C1 => n26575, C2 => n20971, ZN => n23991);
   U23106 : OAI221_X1 port map( B1 => n21491, B2 => n26599, C1 => n22251, C2 =>
                           n26593, A => n24065, ZN => n24058);
   U23107 : AOI222_X1 port map( A1 => n26587, A2 => n25682, B1 => n26581, B2 =>
                           n20970, C1 => n26575, C2 => n20974, ZN => n24065);
   U23108 : OAI221_X1 port map( B1 => n21490, B2 => n26599, C1 => n22250, C2 =>
                           n26593, A => n24047, ZN => n24040);
   U23109 : AOI222_X1 port map( A1 => n26587, A2 => n25687, B1 => n26581, B2 =>
                           n20969, C1 => n26575, C2 => n20973, ZN => n24047);
   U23110 : OAI221_X1 port map( B1 => n21489, B2 => n26599, C1 => n22249, C2 =>
                           n26593, A => n24029, ZN => n24022);
   U23111 : AOI222_X1 port map( A1 => n26587, A2 => n25692, B1 => n26581, B2 =>
                           n20968, C1 => n26575, C2 => n20972, ZN => n24029);
   U23112 : OAI221_X1 port map( B1 => n21491, B2 => n26824, C1 => n22251, C2 =>
                           n26818, A => n22866, ZN => n22859);
   U23113 : AOI222_X1 port map( A1 => n26812, A2 => n25682, B1 => n26806, B2 =>
                           n20970, C1 => n26800, C2 => n20974, ZN => n22866);
   U23114 : OAI221_X1 port map( B1 => n21490, B2 => n26824, C1 => n22250, C2 =>
                           n26818, A => n22848, ZN => n22841);
   U23115 : AOI222_X1 port map( A1 => n26812, A2 => n25687, B1 => n26806, B2 =>
                           n20969, C1 => n26800, C2 => n20973, ZN => n22848);
   U23116 : OAI221_X1 port map( B1 => n21489, B2 => n26824, C1 => n22249, C2 =>
                           n26818, A => n22830, ZN => n22823);
   U23117 : AOI222_X1 port map( A1 => n26812, A2 => n25692, B1 => n26806, B2 =>
                           n20968, C1 => n26800, C2 => n20972, ZN => n22830);
   U23118 : OAI221_X1 port map( B1 => n21488, B2 => n26824, C1 => n22248, C2 =>
                           n26818, A => n22792, ZN => n22771);
   U23119 : AOI222_X1 port map( A1 => n26812, A2 => n25697, B1 => n26806, B2 =>
                           n20967, C1 => n26800, C2 => n20971, ZN => n22792);
   U23120 : OAI221_X1 port map( B1 => n9632, B2 => n26618, C1 => n20834, C2 => 
                           n26612, A => n25152, ZN => n25139);
   U23121 : AOI22_X1 port map( A1 => n26606, A2 => n25701, B1 => n26600, B2 => 
                           n21034, ZN => n25152);
   U23122 : OAI221_X1 port map( B1 => n9631, B2 => n26618, C1 => n20833, C2 => 
                           n26612, A => n25126, ZN => n25121);
   U23123 : AOI22_X1 port map( A1 => n26606, A2 => n25706, B1 => n26600, B2 => 
                           n21033, ZN => n25126);
   U23124 : OAI221_X1 port map( B1 => n9630, B2 => n26618, C1 => n20832, C2 => 
                           n26612, A => n25108, ZN => n25103);
   U23125 : AOI22_X1 port map( A1 => n26606, A2 => n25711, B1 => n26600, B2 => 
                           n21032, ZN => n25108);
   U23126 : OAI221_X1 port map( B1 => n9629, B2 => n26618, C1 => n20831, C2 => 
                           n26612, A => n25090, ZN => n25085);
   U23127 : AOI22_X1 port map( A1 => n26606, A2 => n25716, B1 => n26600, B2 => 
                           n21031, ZN => n25090);
   U23128 : OAI221_X1 port map( B1 => n9628, B2 => n26618, C1 => n20830, C2 => 
                           n26612, A => n25072, ZN => n25067);
   U23129 : AOI22_X1 port map( A1 => n26606, A2 => n25721, B1 => n26600, B2 => 
                           n21030, ZN => n25072);
   U23130 : OAI221_X1 port map( B1 => n9627, B2 => n26618, C1 => n20829, C2 => 
                           n26612, A => n25054, ZN => n25049);
   U23131 : AOI22_X1 port map( A1 => n26606, A2 => n25726, B1 => n26600, B2 => 
                           n21029, ZN => n25054);
   U23132 : OAI221_X1 port map( B1 => n9626, B2 => n26618, C1 => n20828, C2 => 
                           n26612, A => n25036, ZN => n25031);
   U23133 : AOI22_X1 port map( A1 => n26606, A2 => n25731, B1 => n26600, B2 => 
                           n21028, ZN => n25036);
   U23134 : OAI221_X1 port map( B1 => n9625, B2 => n26618, C1 => n20827, C2 => 
                           n26612, A => n25018, ZN => n25013);
   U23135 : AOI22_X1 port map( A1 => n26606, A2 => n25736, B1 => n26600, B2 => 
                           n21027, ZN => n25018);
   U23136 : OAI221_X1 port map( B1 => n9624, B2 => n26618, C1 => n20826, C2 => 
                           n26612, A => n25000, ZN => n24995);
   U23137 : AOI22_X1 port map( A1 => n26606, A2 => n25741, B1 => n26600, B2 => 
                           n21026, ZN => n25000);
   U23138 : OAI221_X1 port map( B1 => n9623, B2 => n26618, C1 => n20825, C2 => 
                           n26612, A => n24982, ZN => n24977);
   U23139 : AOI22_X1 port map( A1 => n26606, A2 => n25746, B1 => n26600, B2 => 
                           n21025, ZN => n24982);
   U23140 : OAI221_X1 port map( B1 => n9622, B2 => n26618, C1 => n20824, C2 => 
                           n26612, A => n24964, ZN => n24959);
   U23141 : AOI22_X1 port map( A1 => n26606, A2 => n25751, B1 => n26600, B2 => 
                           n21024, ZN => n24964);
   U23142 : OAI221_X1 port map( B1 => n9621, B2 => n26618, C1 => n20823, C2 => 
                           n26612, A => n24946, ZN => n24941);
   U23143 : AOI22_X1 port map( A1 => n26606, A2 => n25756, B1 => n26600, B2 => 
                           n21023, ZN => n24946);
   U23144 : OAI221_X1 port map( B1 => n9632, B2 => n26843, C1 => n20834, C2 => 
                           n26837, A => n23953, ZN => n23940);
   U23145 : AOI22_X1 port map( A1 => n26831, A2 => n25701, B1 => n26825, B2 => 
                           n21034, ZN => n23953);
   U23146 : OAI221_X1 port map( B1 => n9631, B2 => n26843, C1 => n20833, C2 => 
                           n26837, A => n23927, ZN => n23922);
   U23147 : AOI22_X1 port map( A1 => n26831, A2 => n25706, B1 => n26825, B2 => 
                           n21033, ZN => n23927);
   U23148 : OAI221_X1 port map( B1 => n9630, B2 => n26843, C1 => n20832, C2 => 
                           n26837, A => n23909, ZN => n23904);
   U23149 : AOI22_X1 port map( A1 => n26831, A2 => n25711, B1 => n26825, B2 => 
                           n21032, ZN => n23909);
   U23150 : OAI221_X1 port map( B1 => n9629, B2 => n26843, C1 => n20831, C2 => 
                           n26837, A => n23891, ZN => n23886);
   U23151 : AOI22_X1 port map( A1 => n26831, A2 => n25716, B1 => n26825, B2 => 
                           n21031, ZN => n23891);
   U23152 : OAI221_X1 port map( B1 => n9628, B2 => n26843, C1 => n20830, C2 => 
                           n26837, A => n23873, ZN => n23868);
   U23153 : AOI22_X1 port map( A1 => n26831, A2 => n25721, B1 => n26825, B2 => 
                           n21030, ZN => n23873);
   U23154 : OAI221_X1 port map( B1 => n9627, B2 => n26843, C1 => n20829, C2 => 
                           n26837, A => n23855, ZN => n23850);
   U23155 : AOI22_X1 port map( A1 => n26831, A2 => n25726, B1 => n26825, B2 => 
                           n21029, ZN => n23855);
   U23156 : OAI221_X1 port map( B1 => n9626, B2 => n26843, C1 => n20828, C2 => 
                           n26837, A => n23837, ZN => n23832);
   U23157 : AOI22_X1 port map( A1 => n26831, A2 => n25731, B1 => n26825, B2 => 
                           n21028, ZN => n23837);
   U23158 : OAI221_X1 port map( B1 => n9625, B2 => n26843, C1 => n20827, C2 => 
                           n26837, A => n23819, ZN => n23814);
   U23159 : AOI22_X1 port map( A1 => n26831, A2 => n25736, B1 => n26825, B2 => 
                           n21027, ZN => n23819);
   U23160 : OAI221_X1 port map( B1 => n9624, B2 => n26843, C1 => n20826, C2 => 
                           n26837, A => n23801, ZN => n23796);
   U23161 : AOI22_X1 port map( A1 => n26831, A2 => n25741, B1 => n26825, B2 => 
                           n21026, ZN => n23801);
   U23162 : OAI221_X1 port map( B1 => n9623, B2 => n26843, C1 => n20825, C2 => 
                           n26837, A => n23783, ZN => n23778);
   U23163 : AOI22_X1 port map( A1 => n26831, A2 => n25746, B1 => n26825, B2 => 
                           n21025, ZN => n23783);
   U23164 : OAI221_X1 port map( B1 => n9622, B2 => n26843, C1 => n20824, C2 => 
                           n26837, A => n23765, ZN => n23760);
   U23165 : AOI22_X1 port map( A1 => n26831, A2 => n25751, B1 => n26825, B2 => 
                           n21024, ZN => n23765);
   U23166 : OAI221_X1 port map( B1 => n9621, B2 => n26843, C1 => n20823, C2 => 
                           n26837, A => n23747, ZN => n23742);
   U23167 : AOI22_X1 port map( A1 => n26831, A2 => n25756, B1 => n26825, B2 => 
                           n21023, ZN => n23747);
   U23168 : OAI221_X1 port map( B1 => n22059, B2 => n26471, C1 => n27284, C2 =>
                           n26465, A => n25166, ZN => n25156);
   U23169 : AOI222_X1 port map( A1 => n26459, A2 => n25595, B1 => n26453, B2 =>
                           n25619, C1 => n26447, C2 => n25667, ZN => n25166);
   U23170 : OAI221_X1 port map( B1 => n22058, B2 => n26471, C1 => n27287, C2 =>
                           n26465, A => n25135, ZN => n25128);
   U23171 : AOI222_X1 port map( A1 => n26459, A2 => n25596, B1 => n26453, B2 =>
                           n25620, C1 => n26447, C2 => n25668, ZN => n25135);
   U23172 : OAI221_X1 port map( B1 => n22057, B2 => n26471, C1 => n27290, C2 =>
                           n26465, A => n25117, ZN => n25110);
   U23173 : AOI222_X1 port map( A1 => n26459, A2 => n25597, B1 => n26453, B2 =>
                           n25621, C1 => n26447, C2 => n25669, ZN => n25117);
   U23174 : OAI221_X1 port map( B1 => n22056, B2 => n26471, C1 => n27293, C2 =>
                           n26465, A => n25099, ZN => n25092);
   U23175 : AOI222_X1 port map( A1 => n26459, A2 => n25598, B1 => n26453, B2 =>
                           n25622, C1 => n26447, C2 => n25670, ZN => n25099);
   U23176 : OAI221_X1 port map( B1 => n22055, B2 => n26471, C1 => n27296, C2 =>
                           n26465, A => n25081, ZN => n25074);
   U23177 : AOI222_X1 port map( A1 => n26459, A2 => n25599, B1 => n26453, B2 =>
                           n25623, C1 => n26447, C2 => n25671, ZN => n25081);
   U23178 : OAI221_X1 port map( B1 => n22054, B2 => n26471, C1 => n27299, C2 =>
                           n26465, A => n25063, ZN => n25056);
   U23179 : AOI222_X1 port map( A1 => n26459, A2 => n25600, B1 => n26453, B2 =>
                           n25624, C1 => n26447, C2 => n25672, ZN => n25063);
   U23180 : OAI221_X1 port map( B1 => n22053, B2 => n26471, C1 => n27302, C2 =>
                           n26465, A => n25045, ZN => n25038);
   U23181 : AOI222_X1 port map( A1 => n26459, A2 => n25601, B1 => n26453, B2 =>
                           n25625, C1 => n26447, C2 => n25673, ZN => n25045);
   U23182 : OAI221_X1 port map( B1 => n22052, B2 => n26471, C1 => n27305, C2 =>
                           n26465, A => n25027, ZN => n25020);
   U23183 : AOI222_X1 port map( A1 => n26459, A2 => n25602, B1 => n26453, B2 =>
                           n25626, C1 => n26447, C2 => n25674, ZN => n25027);
   U23184 : OAI221_X1 port map( B1 => n22051, B2 => n26471, C1 => n27308, C2 =>
                           n26465, A => n25009, ZN => n25002);
   U23185 : AOI222_X1 port map( A1 => n26459, A2 => n25603, B1 => n26453, B2 =>
                           n25627, C1 => n26447, C2 => n25675, ZN => n25009);
   U23186 : OAI221_X1 port map( B1 => n22050, B2 => n26471, C1 => n27311, C2 =>
                           n26465, A => n24991, ZN => n24984);
   U23187 : AOI222_X1 port map( A1 => n26459, A2 => n25604, B1 => n26453, B2 =>
                           n25628, C1 => n26447, C2 => n25676, ZN => n24991);
   U23188 : OAI221_X1 port map( B1 => n22049, B2 => n26471, C1 => n27314, C2 =>
                           n26465, A => n24973, ZN => n24966);
   U23189 : AOI222_X1 port map( A1 => n26459, A2 => n25605, B1 => n26453, B2 =>
                           n25629, C1 => n26447, C2 => n25677, ZN => n24973);
   U23190 : OAI221_X1 port map( B1 => n22048, B2 => n26471, C1 => n27317, C2 =>
                           n26465, A => n24955, ZN => n24948);
   U23191 : AOI222_X1 port map( A1 => n26459, A2 => n25606, B1 => n26453, B2 =>
                           n25630, C1 => n26447, C2 => n25678, ZN => n24955);
   U23192 : OAI221_X1 port map( B1 => n22047, B2 => n26472, C1 => n27320, C2 =>
                           n26466, A => n24937, ZN => n24930);
   U23193 : AOI222_X1 port map( A1 => n26460, A2 => n25215, B1 => n26454, B2 =>
                           n25407, C1 => n26448, C2 => n25503, ZN => n24937);
   U23194 : OAI221_X1 port map( B1 => n22046, B2 => n26472, C1 => n27323, C2 =>
                           n26466, A => n24919, ZN => n24912);
   U23195 : AOI222_X1 port map( A1 => n26460, A2 => n25216, B1 => n26454, B2 =>
                           n25408, C1 => n26448, C2 => n25504, ZN => n24919);
   U23196 : OAI221_X1 port map( B1 => n22045, B2 => n26472, C1 => n27326, C2 =>
                           n26466, A => n24901, ZN => n24894);
   U23197 : AOI222_X1 port map( A1 => n26460, A2 => n25217, B1 => n26454, B2 =>
                           n25409, C1 => n26448, C2 => n25505, ZN => n24901);
   U23198 : OAI221_X1 port map( B1 => n22044, B2 => n26472, C1 => n27329, C2 =>
                           n26466, A => n24883, ZN => n24876);
   U23199 : AOI222_X1 port map( A1 => n26460, A2 => n25218, B1 => n26454, B2 =>
                           n25410, C1 => n26448, C2 => n25506, ZN => n24883);
   U23200 : OAI221_X1 port map( B1 => n22043, B2 => n26472, C1 => n27332, C2 =>
                           n26466, A => n24865, ZN => n24858);
   U23201 : AOI222_X1 port map( A1 => n26460, A2 => n25219, B1 => n26454, B2 =>
                           n25411, C1 => n26448, C2 => n25507, ZN => n24865);
   U23202 : OAI221_X1 port map( B1 => n22042, B2 => n26472, C1 => n27335, C2 =>
                           n26466, A => n24847, ZN => n24840);
   U23203 : AOI222_X1 port map( A1 => n26460, A2 => n25220, B1 => n26454, B2 =>
                           n25412, C1 => n26448, C2 => n25508, ZN => n24847);
   U23204 : OAI221_X1 port map( B1 => n22041, B2 => n26472, C1 => n27338, C2 =>
                           n26466, A => n24829, ZN => n24822);
   U23205 : AOI222_X1 port map( A1 => n26460, A2 => n25221, B1 => n26454, B2 =>
                           n25413, C1 => n26448, C2 => n25509, ZN => n24829);
   U23206 : OAI221_X1 port map( B1 => n22040, B2 => n26472, C1 => n27341, C2 =>
                           n26466, A => n24811, ZN => n24804);
   U23207 : AOI222_X1 port map( A1 => n26460, A2 => n25222, B1 => n26454, B2 =>
                           n25414, C1 => n26448, C2 => n25510, ZN => n24811);
   U23208 : OAI221_X1 port map( B1 => n22039, B2 => n26472, C1 => n27344, C2 =>
                           n26466, A => n24793, ZN => n24786);
   U23209 : AOI222_X1 port map( A1 => n26460, A2 => n25223, B1 => n26454, B2 =>
                           n25415, C1 => n26448, C2 => n25511, ZN => n24793);
   U23210 : OAI221_X1 port map( B1 => n22038, B2 => n26472, C1 => n27347, C2 =>
                           n26466, A => n24775, ZN => n24768);
   U23211 : AOI222_X1 port map( A1 => n26460, A2 => n25224, B1 => n26454, B2 =>
                           n25416, C1 => n26448, C2 => n25512, ZN => n24775);
   U23212 : OAI221_X1 port map( B1 => n22037, B2 => n26472, C1 => n27350, C2 =>
                           n26466, A => n24757, ZN => n24750);
   U23213 : AOI222_X1 port map( A1 => n26460, A2 => n25225, B1 => n26454, B2 =>
                           n25417, C1 => n26448, C2 => n25513, ZN => n24757);
   U23214 : OAI221_X1 port map( B1 => n22036, B2 => n26472, C1 => n27353, C2 =>
                           n26466, A => n24739, ZN => n24732);
   U23215 : AOI222_X1 port map( A1 => n26460, A2 => n25226, B1 => n26454, B2 =>
                           n25418, C1 => n26448, C2 => n25514, ZN => n24739);
   U23216 : OAI221_X1 port map( B1 => n22035, B2 => n26473, C1 => n27356, C2 =>
                           n26467, A => n24721, ZN => n24714);
   U23217 : AOI222_X1 port map( A1 => n26461, A2 => n25227, B1 => n26455, B2 =>
                           n25419, C1 => n26449, C2 => n25515, ZN => n24721);
   U23218 : OAI221_X1 port map( B1 => n22034, B2 => n26473, C1 => n27359, C2 =>
                           n26467, A => n24703, ZN => n24696);
   U23219 : AOI222_X1 port map( A1 => n26461, A2 => n25228, B1 => n26455, B2 =>
                           n25420, C1 => n26449, C2 => n25516, ZN => n24703);
   U23220 : OAI221_X1 port map( B1 => n22033, B2 => n26473, C1 => n27362, C2 =>
                           n26467, A => n24685, ZN => n24678);
   U23221 : AOI222_X1 port map( A1 => n26461, A2 => n25229, B1 => n26455, B2 =>
                           n25421, C1 => n26449, C2 => n25517, ZN => n24685);
   U23222 : OAI221_X1 port map( B1 => n22032, B2 => n26473, C1 => n27365, C2 =>
                           n26467, A => n24667, ZN => n24660);
   U23223 : AOI222_X1 port map( A1 => n26461, A2 => n25230, B1 => n26455, B2 =>
                           n25422, C1 => n26449, C2 => n25518, ZN => n24667);
   U23224 : OAI221_X1 port map( B1 => n22031, B2 => n26473, C1 => n27368, C2 =>
                           n26467, A => n24649, ZN => n24642);
   U23225 : AOI222_X1 port map( A1 => n26461, A2 => n25231, B1 => n26455, B2 =>
                           n25423, C1 => n26449, C2 => n25519, ZN => n24649);
   U23226 : OAI221_X1 port map( B1 => n22030, B2 => n26473, C1 => n27371, C2 =>
                           n26467, A => n24631, ZN => n24624);
   U23227 : AOI222_X1 port map( A1 => n26461, A2 => n25232, B1 => n26455, B2 =>
                           n25424, C1 => n26449, C2 => n25520, ZN => n24631);
   U23228 : OAI221_X1 port map( B1 => n22029, B2 => n26473, C1 => n27374, C2 =>
                           n26467, A => n24613, ZN => n24606);
   U23229 : AOI222_X1 port map( A1 => n26461, A2 => n25233, B1 => n26455, B2 =>
                           n25425, C1 => n26449, C2 => n25521, ZN => n24613);
   U23230 : OAI221_X1 port map( B1 => n22028, B2 => n26473, C1 => n27377, C2 =>
                           n26467, A => n24595, ZN => n24588);
   U23231 : AOI222_X1 port map( A1 => n26461, A2 => n25234, B1 => n26455, B2 =>
                           n25426, C1 => n26449, C2 => n25522, ZN => n24595);
   U23232 : OAI221_X1 port map( B1 => n22027, B2 => n26473, C1 => n27380, C2 =>
                           n26467, A => n24577, ZN => n24570);
   U23233 : AOI222_X1 port map( A1 => n26461, A2 => n25235, B1 => n26455, B2 =>
                           n25427, C1 => n26449, C2 => n25523, ZN => n24577);
   U23234 : OAI221_X1 port map( B1 => n22026, B2 => n26473, C1 => n27383, C2 =>
                           n26467, A => n24559, ZN => n24552);
   U23235 : AOI222_X1 port map( A1 => n26461, A2 => n25236, B1 => n26455, B2 =>
                           n25428, C1 => n26449, C2 => n25524, ZN => n24559);
   U23236 : OAI221_X1 port map( B1 => n22025, B2 => n26473, C1 => n27386, C2 =>
                           n26467, A => n24541, ZN => n24534);
   U23237 : AOI222_X1 port map( A1 => n26461, A2 => n25237, B1 => n26455, B2 =>
                           n25429, C1 => n26449, C2 => n25525, ZN => n24541);
   U23238 : OAI221_X1 port map( B1 => n22024, B2 => n26473, C1 => n27389, C2 =>
                           n26467, A => n24523, ZN => n24516);
   U23239 : AOI222_X1 port map( A1 => n26461, A2 => n25238, B1 => n26455, B2 =>
                           n25430, C1 => n26449, C2 => n25526, ZN => n24523);
   U23240 : OAI221_X1 port map( B1 => n22023, B2 => n26474, C1 => n27392, C2 =>
                           n26468, A => n24505, ZN => n24498);
   U23241 : AOI222_X1 port map( A1 => n26462, A2 => n25239, B1 => n26456, B2 =>
                           n25431, C1 => n26450, C2 => n25527, ZN => n24505);
   U23242 : OAI221_X1 port map( B1 => n22022, B2 => n26474, C1 => n27395, C2 =>
                           n26468, A => n24487, ZN => n24480);
   U23243 : AOI222_X1 port map( A1 => n26462, A2 => n25240, B1 => n26456, B2 =>
                           n25432, C1 => n26450, C2 => n25528, ZN => n24487);
   U23244 : OAI221_X1 port map( B1 => n22021, B2 => n26474, C1 => n27398, C2 =>
                           n26468, A => n24469, ZN => n24462);
   U23245 : AOI222_X1 port map( A1 => n26462, A2 => n25241, B1 => n26456, B2 =>
                           n25433, C1 => n26450, C2 => n25529, ZN => n24469);
   U23246 : OAI221_X1 port map( B1 => n22020, B2 => n26474, C1 => n27401, C2 =>
                           n26468, A => n24451, ZN => n24444);
   U23247 : AOI222_X1 port map( A1 => n26462, A2 => n25242, B1 => n26456, B2 =>
                           n25434, C1 => n26450, C2 => n25530, ZN => n24451);
   U23248 : OAI221_X1 port map( B1 => n22019, B2 => n26474, C1 => n27404, C2 =>
                           n26468, A => n24433, ZN => n24426);
   U23249 : AOI222_X1 port map( A1 => n26462, A2 => n25243, B1 => n26456, B2 =>
                           n25435, C1 => n26450, C2 => n25531, ZN => n24433);
   U23250 : OAI221_X1 port map( B1 => n22018, B2 => n26474, C1 => n27407, C2 =>
                           n26468, A => n24415, ZN => n24408);
   U23251 : AOI222_X1 port map( A1 => n26462, A2 => n25244, B1 => n26456, B2 =>
                           n25436, C1 => n26450, C2 => n25532, ZN => n24415);
   U23252 : OAI221_X1 port map( B1 => n22017, B2 => n26474, C1 => n27410, C2 =>
                           n26468, A => n24397, ZN => n24390);
   U23253 : AOI222_X1 port map( A1 => n26462, A2 => n25245, B1 => n26456, B2 =>
                           n25437, C1 => n26450, C2 => n25533, ZN => n24397);
   U23254 : OAI221_X1 port map( B1 => n22016, B2 => n26474, C1 => n27413, C2 =>
                           n26468, A => n24379, ZN => n24372);
   U23255 : AOI222_X1 port map( A1 => n26462, A2 => n25246, B1 => n26456, B2 =>
                           n25438, C1 => n26450, C2 => n25534, ZN => n24379);
   U23256 : OAI221_X1 port map( B1 => n22015, B2 => n26474, C1 => n27416, C2 =>
                           n26468, A => n24361, ZN => n24354);
   U23257 : AOI222_X1 port map( A1 => n26462, A2 => n25247, B1 => n26456, B2 =>
                           n25439, C1 => n26450, C2 => n25535, ZN => n24361);
   U23258 : OAI221_X1 port map( B1 => n22014, B2 => n26474, C1 => n27419, C2 =>
                           n26468, A => n24343, ZN => n24336);
   U23259 : AOI222_X1 port map( A1 => n26462, A2 => n25248, B1 => n26456, B2 =>
                           n25440, C1 => n26450, C2 => n25536, ZN => n24343);
   U23260 : OAI221_X1 port map( B1 => n22013, B2 => n26474, C1 => n27422, C2 =>
                           n26468, A => n24325, ZN => n24318);
   U23261 : AOI222_X1 port map( A1 => n26462, A2 => n25249, B1 => n26456, B2 =>
                           n25441, C1 => n26450, C2 => n25537, ZN => n24325);
   U23262 : OAI221_X1 port map( B1 => n22012, B2 => n26474, C1 => n27425, C2 =>
                           n26468, A => n24307, ZN => n24300);
   U23263 : AOI222_X1 port map( A1 => n26462, A2 => n25250, B1 => n26456, B2 =>
                           n25442, C1 => n26450, C2 => n25538, ZN => n24307);
   U23264 : OAI221_X1 port map( B1 => n22059, B2 => n26696, C1 => n27284, C2 =>
                           n26690, A => n23967, ZN => n23957);
   U23265 : AOI222_X1 port map( A1 => n26684, A2 => n25595, B1 => n26678, B2 =>
                           n25619, C1 => n26672, C2 => n25667, ZN => n23967);
   U23266 : OAI221_X1 port map( B1 => n22058, B2 => n26696, C1 => n27287, C2 =>
                           n26690, A => n23936, ZN => n23929);
   U23267 : AOI222_X1 port map( A1 => n26684, A2 => n25596, B1 => n26678, B2 =>
                           n25620, C1 => n26672, C2 => n25668, ZN => n23936);
   U23268 : OAI221_X1 port map( B1 => n22057, B2 => n26696, C1 => n27290, C2 =>
                           n26690, A => n23918, ZN => n23911);
   U23269 : AOI222_X1 port map( A1 => n26684, A2 => n25597, B1 => n26678, B2 =>
                           n25621, C1 => n26672, C2 => n25669, ZN => n23918);
   U23270 : OAI221_X1 port map( B1 => n22056, B2 => n26696, C1 => n27293, C2 =>
                           n26690, A => n23900, ZN => n23893);
   U23271 : AOI222_X1 port map( A1 => n26684, A2 => n25598, B1 => n26678, B2 =>
                           n25622, C1 => n26672, C2 => n25670, ZN => n23900);
   U23272 : OAI221_X1 port map( B1 => n22055, B2 => n26696, C1 => n27296, C2 =>
                           n26690, A => n23882, ZN => n23875);
   U23273 : AOI222_X1 port map( A1 => n26684, A2 => n25599, B1 => n26678, B2 =>
                           n25623, C1 => n26672, C2 => n25671, ZN => n23882);
   U23274 : OAI221_X1 port map( B1 => n22054, B2 => n26696, C1 => n27299, C2 =>
                           n26690, A => n23864, ZN => n23857);
   U23275 : AOI222_X1 port map( A1 => n26684, A2 => n25600, B1 => n26678, B2 =>
                           n25624, C1 => n26672, C2 => n25672, ZN => n23864);
   U23276 : OAI221_X1 port map( B1 => n22053, B2 => n26696, C1 => n27302, C2 =>
                           n26690, A => n23846, ZN => n23839);
   U23277 : AOI222_X1 port map( A1 => n26684, A2 => n25601, B1 => n26678, B2 =>
                           n25625, C1 => n26672, C2 => n25673, ZN => n23846);
   U23278 : OAI221_X1 port map( B1 => n22052, B2 => n26696, C1 => n27305, C2 =>
                           n26690, A => n23828, ZN => n23821);
   U23279 : AOI222_X1 port map( A1 => n26684, A2 => n25602, B1 => n26678, B2 =>
                           n25626, C1 => n26672, C2 => n25674, ZN => n23828);
   U23280 : OAI221_X1 port map( B1 => n22051, B2 => n26696, C1 => n27308, C2 =>
                           n26690, A => n23810, ZN => n23803);
   U23281 : AOI222_X1 port map( A1 => n26684, A2 => n25603, B1 => n26678, B2 =>
                           n25627, C1 => n26672, C2 => n25675, ZN => n23810);
   U23282 : OAI221_X1 port map( B1 => n22050, B2 => n26696, C1 => n27311, C2 =>
                           n26690, A => n23792, ZN => n23785);
   U23283 : AOI222_X1 port map( A1 => n26684, A2 => n25604, B1 => n26678, B2 =>
                           n25628, C1 => n26672, C2 => n25676, ZN => n23792);
   U23284 : OAI221_X1 port map( B1 => n22049, B2 => n26696, C1 => n27314, C2 =>
                           n26690, A => n23774, ZN => n23767);
   U23285 : AOI222_X1 port map( A1 => n26684, A2 => n25605, B1 => n26678, B2 =>
                           n25629, C1 => n26672, C2 => n25677, ZN => n23774);
   U23286 : OAI221_X1 port map( B1 => n22048, B2 => n26696, C1 => n27317, C2 =>
                           n26690, A => n23756, ZN => n23749);
   U23287 : AOI222_X1 port map( A1 => n26684, A2 => n25606, B1 => n26678, B2 =>
                           n25630, C1 => n26672, C2 => n25678, ZN => n23756);
   U23288 : OAI221_X1 port map( B1 => n22047, B2 => n26697, C1 => n27320, C2 =>
                           n26691, A => n23738, ZN => n23731);
   U23289 : AOI222_X1 port map( A1 => n26685, A2 => n25215, B1 => n26679, B2 =>
                           n25407, C1 => n26673, C2 => n25503, ZN => n23738);
   U23290 : OAI221_X1 port map( B1 => n22046, B2 => n26697, C1 => n27323, C2 =>
                           n26691, A => n23720, ZN => n23713);
   U23291 : AOI222_X1 port map( A1 => n26685, A2 => n25216, B1 => n26679, B2 =>
                           n25408, C1 => n26673, C2 => n25504, ZN => n23720);
   U23292 : OAI221_X1 port map( B1 => n22045, B2 => n26697, C1 => n27326, C2 =>
                           n26691, A => n23702, ZN => n23695);
   U23293 : AOI222_X1 port map( A1 => n26685, A2 => n25217, B1 => n26679, B2 =>
                           n25409, C1 => n26673, C2 => n25505, ZN => n23702);
   U23294 : OAI221_X1 port map( B1 => n22044, B2 => n26697, C1 => n27329, C2 =>
                           n26691, A => n23684, ZN => n23677);
   U23295 : AOI222_X1 port map( A1 => n26685, A2 => n25218, B1 => n26679, B2 =>
                           n25410, C1 => n26673, C2 => n25506, ZN => n23684);
   U23296 : OAI221_X1 port map( B1 => n22043, B2 => n26697, C1 => n27332, C2 =>
                           n26691, A => n23666, ZN => n23659);
   U23297 : AOI222_X1 port map( A1 => n26685, A2 => n25219, B1 => n26679, B2 =>
                           n25411, C1 => n26673, C2 => n25507, ZN => n23666);
   U23298 : OAI221_X1 port map( B1 => n22042, B2 => n26697, C1 => n27335, C2 =>
                           n26691, A => n23648, ZN => n23641);
   U23299 : AOI222_X1 port map( A1 => n26685, A2 => n25220, B1 => n26679, B2 =>
                           n25412, C1 => n26673, C2 => n25508, ZN => n23648);
   U23300 : OAI221_X1 port map( B1 => n22041, B2 => n26697, C1 => n27338, C2 =>
                           n26691, A => n23630, ZN => n23623);
   U23301 : AOI222_X1 port map( A1 => n26685, A2 => n25221, B1 => n26679, B2 =>
                           n25413, C1 => n26673, C2 => n25509, ZN => n23630);
   U23302 : OAI221_X1 port map( B1 => n22040, B2 => n26697, C1 => n27341, C2 =>
                           n26691, A => n23612, ZN => n23605);
   U23303 : AOI222_X1 port map( A1 => n26685, A2 => n25222, B1 => n26679, B2 =>
                           n25414, C1 => n26673, C2 => n25510, ZN => n23612);
   U23304 : OAI221_X1 port map( B1 => n22039, B2 => n26697, C1 => n27344, C2 =>
                           n26691, A => n23594, ZN => n23587);
   U23305 : AOI222_X1 port map( A1 => n26685, A2 => n25223, B1 => n26679, B2 =>
                           n25415, C1 => n26673, C2 => n25511, ZN => n23594);
   U23306 : OAI221_X1 port map( B1 => n22038, B2 => n26697, C1 => n27347, C2 =>
                           n26691, A => n23576, ZN => n23569);
   U23307 : AOI222_X1 port map( A1 => n26685, A2 => n25224, B1 => n26679, B2 =>
                           n25416, C1 => n26673, C2 => n25512, ZN => n23576);
   U23308 : OAI221_X1 port map( B1 => n22037, B2 => n26697, C1 => n27350, C2 =>
                           n26691, A => n23558, ZN => n23551);
   U23309 : AOI222_X1 port map( A1 => n26685, A2 => n25225, B1 => n26679, B2 =>
                           n25417, C1 => n26673, C2 => n25513, ZN => n23558);
   U23310 : OAI221_X1 port map( B1 => n22036, B2 => n26697, C1 => n27353, C2 =>
                           n26691, A => n23540, ZN => n23533);
   U23311 : AOI222_X1 port map( A1 => n26685, A2 => n25226, B1 => n26679, B2 =>
                           n25418, C1 => n26673, C2 => n25514, ZN => n23540);
   U23312 : OAI221_X1 port map( B1 => n22035, B2 => n26698, C1 => n27356, C2 =>
                           n26692, A => n23522, ZN => n23515);
   U23313 : AOI222_X1 port map( A1 => n26686, A2 => n25227, B1 => n26680, B2 =>
                           n25419, C1 => n26674, C2 => n25515, ZN => n23522);
   U23314 : OAI221_X1 port map( B1 => n22034, B2 => n26698, C1 => n27359, C2 =>
                           n26692, A => n23504, ZN => n23497);
   U23315 : AOI222_X1 port map( A1 => n26686, A2 => n25228, B1 => n26680, B2 =>
                           n25420, C1 => n26674, C2 => n25516, ZN => n23504);
   U23316 : OAI221_X1 port map( B1 => n22033, B2 => n26698, C1 => n27362, C2 =>
                           n26692, A => n23486, ZN => n23479);
   U23317 : AOI222_X1 port map( A1 => n26686, A2 => n25229, B1 => n26680, B2 =>
                           n25421, C1 => n26674, C2 => n25517, ZN => n23486);
   U23318 : OAI221_X1 port map( B1 => n22032, B2 => n26698, C1 => n27365, C2 =>
                           n26692, A => n23468, ZN => n23461);
   U23319 : AOI222_X1 port map( A1 => n26686, A2 => n25230, B1 => n26680, B2 =>
                           n25422, C1 => n26674, C2 => n25518, ZN => n23468);
   U23320 : OAI221_X1 port map( B1 => n22031, B2 => n26698, C1 => n27368, C2 =>
                           n26692, A => n23450, ZN => n23443);
   U23321 : AOI222_X1 port map( A1 => n26686, A2 => n25231, B1 => n26680, B2 =>
                           n25423, C1 => n26674, C2 => n25519, ZN => n23450);
   U23322 : OAI221_X1 port map( B1 => n22030, B2 => n26698, C1 => n27371, C2 =>
                           n26692, A => n23432, ZN => n23425);
   U23323 : AOI222_X1 port map( A1 => n26686, A2 => n25232, B1 => n26680, B2 =>
                           n25424, C1 => n26674, C2 => n25520, ZN => n23432);
   U23324 : OAI221_X1 port map( B1 => n22029, B2 => n26698, C1 => n27374, C2 =>
                           n26692, A => n23414, ZN => n23407);
   U23325 : AOI222_X1 port map( A1 => n26686, A2 => n25233, B1 => n26680, B2 =>
                           n25425, C1 => n26674, C2 => n25521, ZN => n23414);
   U23326 : OAI221_X1 port map( B1 => n22028, B2 => n26698, C1 => n27377, C2 =>
                           n26692, A => n23396, ZN => n23389);
   U23327 : AOI222_X1 port map( A1 => n26686, A2 => n25234, B1 => n26680, B2 =>
                           n25426, C1 => n26674, C2 => n25522, ZN => n23396);
   U23328 : OAI221_X1 port map( B1 => n22027, B2 => n26698, C1 => n27380, C2 =>
                           n26692, A => n23378, ZN => n23371);
   U23329 : AOI222_X1 port map( A1 => n26686, A2 => n25235, B1 => n26680, B2 =>
                           n25427, C1 => n26674, C2 => n25523, ZN => n23378);
   U23330 : OAI221_X1 port map( B1 => n22026, B2 => n26698, C1 => n27383, C2 =>
                           n26692, A => n23360, ZN => n23353);
   U23331 : AOI222_X1 port map( A1 => n26686, A2 => n25236, B1 => n26680, B2 =>
                           n25428, C1 => n26674, C2 => n25524, ZN => n23360);
   U23332 : OAI221_X1 port map( B1 => n22025, B2 => n26698, C1 => n27386, C2 =>
                           n26692, A => n23342, ZN => n23335);
   U23333 : AOI222_X1 port map( A1 => n26686, A2 => n25237, B1 => n26680, B2 =>
                           n25429, C1 => n26674, C2 => n25525, ZN => n23342);
   U23334 : OAI221_X1 port map( B1 => n22024, B2 => n26698, C1 => n27389, C2 =>
                           n26692, A => n23324, ZN => n23317);
   U23335 : AOI222_X1 port map( A1 => n26686, A2 => n25238, B1 => n26680, B2 =>
                           n25430, C1 => n26674, C2 => n25526, ZN => n23324);
   U23336 : OAI221_X1 port map( B1 => n22023, B2 => n26699, C1 => n27392, C2 =>
                           n26693, A => n23306, ZN => n23299);
   U23337 : AOI222_X1 port map( A1 => n26687, A2 => n25239, B1 => n26681, B2 =>
                           n25431, C1 => n26675, C2 => n25527, ZN => n23306);
   U23338 : OAI221_X1 port map( B1 => n22022, B2 => n26699, C1 => n27395, C2 =>
                           n26693, A => n23288, ZN => n23281);
   U23339 : AOI222_X1 port map( A1 => n26687, A2 => n25240, B1 => n26681, B2 =>
                           n25432, C1 => n26675, C2 => n25528, ZN => n23288);
   U23340 : OAI221_X1 port map( B1 => n22021, B2 => n26699, C1 => n27398, C2 =>
                           n26693, A => n23270, ZN => n23263);
   U23341 : AOI222_X1 port map( A1 => n26687, A2 => n25241, B1 => n26681, B2 =>
                           n25433, C1 => n26675, C2 => n25529, ZN => n23270);
   U23342 : OAI221_X1 port map( B1 => n22020, B2 => n26699, C1 => n27401, C2 =>
                           n26693, A => n23252, ZN => n23245);
   U23343 : AOI222_X1 port map( A1 => n26687, A2 => n25242, B1 => n26681, B2 =>
                           n25434, C1 => n26675, C2 => n25530, ZN => n23252);
   U23344 : OAI221_X1 port map( B1 => n22019, B2 => n26699, C1 => n27404, C2 =>
                           n26693, A => n23234, ZN => n23227);
   U23345 : AOI222_X1 port map( A1 => n26687, A2 => n25243, B1 => n26681, B2 =>
                           n25435, C1 => n26675, C2 => n25531, ZN => n23234);
   U23346 : OAI221_X1 port map( B1 => n22018, B2 => n26699, C1 => n27407, C2 =>
                           n26693, A => n23216, ZN => n23209);
   U23347 : AOI222_X1 port map( A1 => n26687, A2 => n25244, B1 => n26681, B2 =>
                           n25436, C1 => n26675, C2 => n25532, ZN => n23216);
   U23348 : OAI221_X1 port map( B1 => n22017, B2 => n26699, C1 => n27410, C2 =>
                           n26693, A => n23198, ZN => n23191);
   U23349 : AOI222_X1 port map( A1 => n26687, A2 => n25245, B1 => n26681, B2 =>
                           n25437, C1 => n26675, C2 => n25533, ZN => n23198);
   U23350 : OAI221_X1 port map( B1 => n22016, B2 => n26699, C1 => n27413, C2 =>
                           n26693, A => n23180, ZN => n23173);
   U23351 : AOI222_X1 port map( A1 => n26687, A2 => n25246, B1 => n26681, B2 =>
                           n25438, C1 => n26675, C2 => n25534, ZN => n23180);
   U23352 : OAI221_X1 port map( B1 => n22015, B2 => n26699, C1 => n27416, C2 =>
                           n26693, A => n23162, ZN => n23155);
   U23353 : AOI222_X1 port map( A1 => n26687, A2 => n25247, B1 => n26681, B2 =>
                           n25439, C1 => n26675, C2 => n25535, ZN => n23162);
   U23354 : OAI221_X1 port map( B1 => n22014, B2 => n26699, C1 => n27419, C2 =>
                           n26693, A => n23144, ZN => n23137);
   U23355 : AOI222_X1 port map( A1 => n26687, A2 => n25248, B1 => n26681, B2 =>
                           n25440, C1 => n26675, C2 => n25536, ZN => n23144);
   U23356 : OAI221_X1 port map( B1 => n22013, B2 => n26699, C1 => n27422, C2 =>
                           n26693, A => n23126, ZN => n23119);
   U23357 : AOI222_X1 port map( A1 => n26687, A2 => n25249, B1 => n26681, B2 =>
                           n25441, C1 => n26675, C2 => n25537, ZN => n23126);
   U23358 : OAI221_X1 port map( B1 => n22012, B2 => n26699, C1 => n27425, C2 =>
                           n26693, A => n23108, ZN => n23101);
   U23359 : AOI222_X1 port map( A1 => n26687, A2 => n25250, B1 => n26681, B2 =>
                           n25442, C1 => n26675, C2 => n25538, ZN => n23108);
   U23360 : OAI221_X1 port map( B1 => n21759, B2 => n26594, C1 => n22379, C2 =>
                           n26588, A => n25154, ZN => n25138);
   U23361 : AOI222_X1 port map( A1 => n26582, A2 => n25702, B1 => n26576, B2 =>
                           n21094, C1 => n26570, C2 => n21154, ZN => n25154);
   U23362 : OAI221_X1 port map( B1 => n21758, B2 => n26594, C1 => n22378, C2 =>
                           n26588, A => n25127, ZN => n25120);
   U23363 : AOI222_X1 port map( A1 => n26582, A2 => n25707, B1 => n26576, B2 =>
                           n21093, C1 => n26570, C2 => n21153, ZN => n25127);
   U23364 : OAI221_X1 port map( B1 => n21757, B2 => n26594, C1 => n22377, C2 =>
                           n26588, A => n25109, ZN => n25102);
   U23365 : AOI222_X1 port map( A1 => n26582, A2 => n25712, B1 => n26576, B2 =>
                           n21092, C1 => n26570, C2 => n21152, ZN => n25109);
   U23366 : OAI221_X1 port map( B1 => n21756, B2 => n26594, C1 => n22376, C2 =>
                           n26588, A => n25091, ZN => n25084);
   U23367 : AOI222_X1 port map( A1 => n26582, A2 => n25717, B1 => n26576, B2 =>
                           n21091, C1 => n26570, C2 => n21151, ZN => n25091);
   U23368 : OAI221_X1 port map( B1 => n21755, B2 => n26594, C1 => n22375, C2 =>
                           n26588, A => n25073, ZN => n25066);
   U23369 : AOI222_X1 port map( A1 => n26582, A2 => n25722, B1 => n26576, B2 =>
                           n21090, C1 => n26570, C2 => n21150, ZN => n25073);
   U23370 : OAI221_X1 port map( B1 => n21754, B2 => n26594, C1 => n22374, C2 =>
                           n26588, A => n25055, ZN => n25048);
   U23371 : AOI222_X1 port map( A1 => n26582, A2 => n25727, B1 => n26576, B2 =>
                           n21089, C1 => n26570, C2 => n21149, ZN => n25055);
   U23372 : OAI221_X1 port map( B1 => n21753, B2 => n26594, C1 => n22373, C2 =>
                           n26588, A => n25037, ZN => n25030);
   U23373 : AOI222_X1 port map( A1 => n26582, A2 => n25732, B1 => n26576, B2 =>
                           n21088, C1 => n26570, C2 => n21148, ZN => n25037);
   U23374 : OAI221_X1 port map( B1 => n21752, B2 => n26594, C1 => n22372, C2 =>
                           n26588, A => n25019, ZN => n25012);
   U23375 : AOI222_X1 port map( A1 => n26582, A2 => n25737, B1 => n26576, B2 =>
                           n21087, C1 => n26570, C2 => n21147, ZN => n25019);
   U23376 : OAI221_X1 port map( B1 => n21751, B2 => n26594, C1 => n22371, C2 =>
                           n26588, A => n25001, ZN => n24994);
   U23377 : AOI222_X1 port map( A1 => n26582, A2 => n25742, B1 => n26576, B2 =>
                           n21086, C1 => n26570, C2 => n21146, ZN => n25001);
   U23378 : OAI221_X1 port map( B1 => n21750, B2 => n26594, C1 => n22370, C2 =>
                           n26588, A => n24983, ZN => n24976);
   U23379 : AOI222_X1 port map( A1 => n26582, A2 => n25747, B1 => n26576, B2 =>
                           n21085, C1 => n26570, C2 => n21145, ZN => n24983);
   U23380 : OAI221_X1 port map( B1 => n21749, B2 => n26594, C1 => n22369, C2 =>
                           n26588, A => n24965, ZN => n24958);
   U23381 : AOI222_X1 port map( A1 => n26582, A2 => n25752, B1 => n26576, B2 =>
                           n21084, C1 => n26570, C2 => n21144, ZN => n24965);
   U23382 : OAI221_X1 port map( B1 => n21748, B2 => n26594, C1 => n22368, C2 =>
                           n26588, A => n24947, ZN => n24940);
   U23383 : AOI222_X1 port map( A1 => n26582, A2 => n25757, B1 => n26576, B2 =>
                           n21083, C1 => n26570, C2 => n21143, ZN => n24947);
   U23384 : OAI221_X1 port map( B1 => n22011, B2 => n26475, C1 => n27428, C2 =>
                           n26469, A => n24289, ZN => n24282);
   U23385 : AOI222_X1 port map( A1 => n26463, A2 => n25251, B1 => n26457, B2 =>
                           n25443, C1 => n26451, C2 => n25539, ZN => n24289);
   U23386 : OAI221_X1 port map( B1 => n22010, B2 => n26475, C1 => n27431, C2 =>
                           n26469, A => n24271, ZN => n24264);
   U23387 : AOI222_X1 port map( A1 => n26463, A2 => n25252, B1 => n26457, B2 =>
                           n25444, C1 => n26451, C2 => n25540, ZN => n24271);
   U23388 : OAI221_X1 port map( B1 => n22009, B2 => n26475, C1 => n27434, C2 =>
                           n26469, A => n24253, ZN => n24246);
   U23389 : AOI222_X1 port map( A1 => n26463, A2 => n25253, B1 => n26457, B2 =>
                           n25445, C1 => n26451, C2 => n25541, ZN => n24253);
   U23390 : OAI221_X1 port map( B1 => n22008, B2 => n26475, C1 => n27437, C2 =>
                           n26469, A => n24235, ZN => n24228);
   U23391 : AOI222_X1 port map( A1 => n26463, A2 => n25254, B1 => n26457, B2 =>
                           n25446, C1 => n26451, C2 => n25542, ZN => n24235);
   U23392 : OAI221_X1 port map( B1 => n22007, B2 => n26475, C1 => n27440, C2 =>
                           n26469, A => n24217, ZN => n24210);
   U23393 : AOI222_X1 port map( A1 => n26463, A2 => n25255, B1 => n26457, B2 =>
                           n25447, C1 => n26451, C2 => n25543, ZN => n24217);
   U23394 : OAI221_X1 port map( B1 => n22006, B2 => n26475, C1 => n27443, C2 =>
                           n26469, A => n24199, ZN => n24192);
   U23395 : AOI222_X1 port map( A1 => n26463, A2 => n25256, B1 => n26457, B2 =>
                           n25448, C1 => n26451, C2 => n25544, ZN => n24199);
   U23396 : OAI221_X1 port map( B1 => n22005, B2 => n26475, C1 => n27446, C2 =>
                           n26469, A => n24181, ZN => n24174);
   U23397 : AOI222_X1 port map( A1 => n26463, A2 => n25257, B1 => n26457, B2 =>
                           n25449, C1 => n26451, C2 => n25545, ZN => n24181);
   U23398 : OAI221_X1 port map( B1 => n22004, B2 => n26475, C1 => n27449, C2 =>
                           n26469, A => n24163, ZN => n24156);
   U23399 : AOI222_X1 port map( A1 => n26463, A2 => n25258, B1 => n26457, B2 =>
                           n25450, C1 => n26451, C2 => n25546, ZN => n24163);
   U23400 : OAI221_X1 port map( B1 => n22003, B2 => n26475, C1 => n27452, C2 =>
                           n26469, A => n24145, ZN => n24138);
   U23401 : AOI222_X1 port map( A1 => n26463, A2 => n25259, B1 => n26457, B2 =>
                           n25451, C1 => n26451, C2 => n25547, ZN => n24145);
   U23402 : OAI221_X1 port map( B1 => n22002, B2 => n26475, C1 => n27455, C2 =>
                           n26469, A => n24127, ZN => n24120);
   U23403 : AOI222_X1 port map( A1 => n26463, A2 => n25260, B1 => n26457, B2 =>
                           n25452, C1 => n26451, C2 => n25548, ZN => n24127);
   U23404 : OAI221_X1 port map( B1 => n22001, B2 => n26475, C1 => n27458, C2 =>
                           n26469, A => n24109, ZN => n24102);
   U23405 : AOI222_X1 port map( A1 => n26463, A2 => n25261, B1 => n26457, B2 =>
                           n25453, C1 => n26451, C2 => n25549, ZN => n24109);
   U23406 : OAI221_X1 port map( B1 => n22000, B2 => n26475, C1 => n27461, C2 =>
                           n26469, A => n24091, ZN => n24084);
   U23407 : AOI222_X1 port map( A1 => n26463, A2 => n25262, B1 => n26457, B2 =>
                           n25454, C1 => n26451, C2 => n25550, ZN => n24091);
   U23408 : OAI221_X1 port map( B1 => n21759, B2 => n26819, C1 => n22379, C2 =>
                           n26813, A => n23955, ZN => n23939);
   U23409 : AOI222_X1 port map( A1 => n26807, A2 => n25702, B1 => n26801, B2 =>
                           n21094, C1 => n26795, C2 => n21154, ZN => n23955);
   U23410 : OAI221_X1 port map( B1 => n21758, B2 => n26819, C1 => n22378, C2 =>
                           n26813, A => n23928, ZN => n23921);
   U23411 : AOI222_X1 port map( A1 => n26807, A2 => n25707, B1 => n26801, B2 =>
                           n21093, C1 => n26795, C2 => n21153, ZN => n23928);
   U23412 : OAI221_X1 port map( B1 => n21757, B2 => n26819, C1 => n22377, C2 =>
                           n26813, A => n23910, ZN => n23903);
   U23413 : AOI222_X1 port map( A1 => n26807, A2 => n25712, B1 => n26801, B2 =>
                           n21092, C1 => n26795, C2 => n21152, ZN => n23910);
   U23414 : OAI221_X1 port map( B1 => n21756, B2 => n26819, C1 => n22376, C2 =>
                           n26813, A => n23892, ZN => n23885);
   U23415 : AOI222_X1 port map( A1 => n26807, A2 => n25717, B1 => n26801, B2 =>
                           n21091, C1 => n26795, C2 => n21151, ZN => n23892);
   U23416 : OAI221_X1 port map( B1 => n21755, B2 => n26819, C1 => n22375, C2 =>
                           n26813, A => n23874, ZN => n23867);
   U23417 : AOI222_X1 port map( A1 => n26807, A2 => n25722, B1 => n26801, B2 =>
                           n21090, C1 => n26795, C2 => n21150, ZN => n23874);
   U23418 : OAI221_X1 port map( B1 => n21754, B2 => n26819, C1 => n22374, C2 =>
                           n26813, A => n23856, ZN => n23849);
   U23419 : AOI222_X1 port map( A1 => n26807, A2 => n25727, B1 => n26801, B2 =>
                           n21089, C1 => n26795, C2 => n21149, ZN => n23856);
   U23420 : OAI221_X1 port map( B1 => n21753, B2 => n26819, C1 => n22373, C2 =>
                           n26813, A => n23838, ZN => n23831);
   U23421 : AOI222_X1 port map( A1 => n26807, A2 => n25732, B1 => n26801, B2 =>
                           n21088, C1 => n26795, C2 => n21148, ZN => n23838);
   U23422 : OAI221_X1 port map( B1 => n21752, B2 => n26819, C1 => n22372, C2 =>
                           n26813, A => n23820, ZN => n23813);
   U23423 : AOI222_X1 port map( A1 => n26807, A2 => n25737, B1 => n26801, B2 =>
                           n21087, C1 => n26795, C2 => n21147, ZN => n23820);
   U23424 : OAI221_X1 port map( B1 => n21751, B2 => n26819, C1 => n22371, C2 =>
                           n26813, A => n23802, ZN => n23795);
   U23425 : AOI222_X1 port map( A1 => n26807, A2 => n25742, B1 => n26801, B2 =>
                           n21086, C1 => n26795, C2 => n21146, ZN => n23802);
   U23426 : OAI221_X1 port map( B1 => n21750, B2 => n26819, C1 => n22370, C2 =>
                           n26813, A => n23784, ZN => n23777);
   U23427 : AOI222_X1 port map( A1 => n26807, A2 => n25747, B1 => n26801, B2 =>
                           n21085, C1 => n26795, C2 => n21145, ZN => n23784);
   U23428 : OAI221_X1 port map( B1 => n21749, B2 => n26819, C1 => n22369, C2 =>
                           n26813, A => n23766, ZN => n23759);
   U23429 : AOI222_X1 port map( A1 => n26807, A2 => n25752, B1 => n26801, B2 =>
                           n21084, C1 => n26795, C2 => n21144, ZN => n23766);
   U23430 : OAI221_X1 port map( B1 => n21748, B2 => n26819, C1 => n22368, C2 =>
                           n26813, A => n23748, ZN => n23741);
   U23431 : AOI222_X1 port map( A1 => n26807, A2 => n25757, B1 => n26801, B2 =>
                           n21083, C1 => n26795, C2 => n21143, ZN => n23748);
   U23432 : OAI221_X1 port map( B1 => n22011, B2 => n26700, C1 => n27428, C2 =>
                           n26694, A => n23090, ZN => n23083);
   U23433 : AOI222_X1 port map( A1 => n26688, A2 => n25251, B1 => n26682, B2 =>
                           n25443, C1 => n26676, C2 => n25539, ZN => n23090);
   U23434 : OAI221_X1 port map( B1 => n22010, B2 => n26700, C1 => n27431, C2 =>
                           n26694, A => n23072, ZN => n23065);
   U23435 : AOI222_X1 port map( A1 => n26688, A2 => n25252, B1 => n26682, B2 =>
                           n25444, C1 => n26676, C2 => n25540, ZN => n23072);
   U23436 : OAI221_X1 port map( B1 => n22009, B2 => n26700, C1 => n27434, C2 =>
                           n26694, A => n23054, ZN => n23047);
   U23437 : AOI222_X1 port map( A1 => n26688, A2 => n25253, B1 => n26682, B2 =>
                           n25445, C1 => n26676, C2 => n25541, ZN => n23054);
   U23438 : OAI221_X1 port map( B1 => n22008, B2 => n26700, C1 => n27437, C2 =>
                           n26694, A => n23036, ZN => n23029);
   U23439 : AOI222_X1 port map( A1 => n26688, A2 => n25254, B1 => n26682, B2 =>
                           n25446, C1 => n26676, C2 => n25542, ZN => n23036);
   U23440 : OAI221_X1 port map( B1 => n22007, B2 => n26700, C1 => n27440, C2 =>
                           n26694, A => n23018, ZN => n23011);
   U23441 : AOI222_X1 port map( A1 => n26688, A2 => n25255, B1 => n26682, B2 =>
                           n25447, C1 => n26676, C2 => n25543, ZN => n23018);
   U23442 : OAI221_X1 port map( B1 => n22006, B2 => n26700, C1 => n27443, C2 =>
                           n26694, A => n23000, ZN => n22993);
   U23443 : AOI222_X1 port map( A1 => n26688, A2 => n25256, B1 => n26682, B2 =>
                           n25448, C1 => n26676, C2 => n25544, ZN => n23000);
   U23444 : OAI221_X1 port map( B1 => n22005, B2 => n26700, C1 => n27446, C2 =>
                           n26694, A => n22982, ZN => n22975);
   U23445 : AOI222_X1 port map( A1 => n26688, A2 => n25257, B1 => n26682, B2 =>
                           n25449, C1 => n26676, C2 => n25545, ZN => n22982);
   U23446 : OAI221_X1 port map( B1 => n22004, B2 => n26700, C1 => n27449, C2 =>
                           n26694, A => n22964, ZN => n22957);
   U23447 : AOI222_X1 port map( A1 => n26688, A2 => n25258, B1 => n26682, B2 =>
                           n25450, C1 => n26676, C2 => n25546, ZN => n22964);
   U23448 : OAI221_X1 port map( B1 => n22003, B2 => n26700, C1 => n27452, C2 =>
                           n26694, A => n22946, ZN => n22939);
   U23449 : AOI222_X1 port map( A1 => n26688, A2 => n25259, B1 => n26682, B2 =>
                           n25451, C1 => n26676, C2 => n25547, ZN => n22946);
   U23450 : OAI221_X1 port map( B1 => n22002, B2 => n26700, C1 => n27455, C2 =>
                           n26694, A => n22928, ZN => n22921);
   U23451 : AOI222_X1 port map( A1 => n26688, A2 => n25260, B1 => n26682, B2 =>
                           n25452, C1 => n26676, C2 => n25548, ZN => n22928);
   U23452 : OAI221_X1 port map( B1 => n22001, B2 => n26700, C1 => n27458, C2 =>
                           n26694, A => n22910, ZN => n22903);
   U23453 : AOI222_X1 port map( A1 => n26688, A2 => n25261, B1 => n26682, B2 =>
                           n25453, C1 => n26676, C2 => n25549, ZN => n22910);
   U23454 : OAI221_X1 port map( B1 => n22000, B2 => n26700, C1 => n27461, C2 =>
                           n26694, A => n22892, ZN => n22885);
   U23455 : AOI222_X1 port map( A1 => n26688, A2 => n25262, B1 => n26682, B2 =>
                           n25454, C1 => n26676, C2 => n25550, ZN => n22892);
   U23456 : OAI22_X1 port map( A1 => n27320, A2 => n26952, B1 => n26946, B2 => 
                           n22619, ZN => n6286);
   U23457 : OAI22_X1 port map( A1 => n27323, A2 => n26952, B1 => n26946, B2 => 
                           n22618, ZN => n6287);
   U23458 : OAI22_X1 port map( A1 => n27326, A2 => n26952, B1 => n26946, B2 => 
                           n22617, ZN => n6288);
   U23459 : OAI22_X1 port map( A1 => n27329, A2 => n26952, B1 => n26946, B2 => 
                           n22616, ZN => n6289);
   U23460 : OAI22_X1 port map( A1 => n27332, A2 => n26952, B1 => n26946, B2 => 
                           n22615, ZN => n6290);
   U23461 : OAI22_X1 port map( A1 => n27335, A2 => n26952, B1 => n26946, B2 => 
                           n22614, ZN => n6291);
   U23462 : OAI22_X1 port map( A1 => n27338, A2 => n26952, B1 => n26946, B2 => 
                           n22613, ZN => n6292);
   U23463 : OAI22_X1 port map( A1 => n27341, A2 => n26952, B1 => n26946, B2 => 
                           n22612, ZN => n6293);
   U23464 : OAI22_X1 port map( A1 => n27344, A2 => n26952, B1 => n26946, B2 => 
                           n22611, ZN => n6294);
   U23465 : OAI22_X1 port map( A1 => n27347, A2 => n26952, B1 => n26946, B2 => 
                           n22610, ZN => n6295);
   U23466 : OAI22_X1 port map( A1 => n27350, A2 => n26952, B1 => n26946, B2 => 
                           n22609, ZN => n6296);
   U23467 : OAI22_X1 port map( A1 => n27353, A2 => n26953, B1 => n26946, B2 => 
                           n22608, ZN => n6297);
   U23468 : OAI22_X1 port map( A1 => n27356, A2 => n26953, B1 => n26947, B2 => 
                           n22607, ZN => n6298);
   U23469 : OAI22_X1 port map( A1 => n27359, A2 => n26953, B1 => n26947, B2 => 
                           n22606, ZN => n6299);
   U23470 : OAI22_X1 port map( A1 => n27362, A2 => n26953, B1 => n26947, B2 => 
                           n22605, ZN => n6300);
   U23471 : OAI22_X1 port map( A1 => n27365, A2 => n26953, B1 => n26947, B2 => 
                           n22604, ZN => n6301);
   U23472 : OAI22_X1 port map( A1 => n27368, A2 => n26953, B1 => n26947, B2 => 
                           n22603, ZN => n6302);
   U23473 : OAI22_X1 port map( A1 => n27371, A2 => n26953, B1 => n26947, B2 => 
                           n22602, ZN => n6303);
   U23474 : OAI22_X1 port map( A1 => n27374, A2 => n26953, B1 => n26947, B2 => 
                           n22601, ZN => n6304);
   U23475 : OAI22_X1 port map( A1 => n27377, A2 => n26953, B1 => n26947, B2 => 
                           n22600, ZN => n6305);
   U23476 : OAI22_X1 port map( A1 => n27380, A2 => n26953, B1 => n26947, B2 => 
                           n22599, ZN => n6306);
   U23477 : OAI22_X1 port map( A1 => n27383, A2 => n26953, B1 => n26947, B2 => 
                           n22598, ZN => n6307);
   U23478 : OAI22_X1 port map( A1 => n27386, A2 => n26953, B1 => n26947, B2 => 
                           n22597, ZN => n6308);
   U23479 : OAI22_X1 port map( A1 => n27389, A2 => n26954, B1 => n26947, B2 => 
                           n22596, ZN => n6309);
   U23480 : OAI22_X1 port map( A1 => n27392, A2 => n26954, B1 => n26948, B2 => 
                           n22595, ZN => n6310);
   U23481 : OAI22_X1 port map( A1 => n27395, A2 => n26954, B1 => n26948, B2 => 
                           n22594, ZN => n6311);
   U23482 : OAI22_X1 port map( A1 => n27398, A2 => n26954, B1 => n26948, B2 => 
                           n22593, ZN => n6312);
   U23483 : OAI22_X1 port map( A1 => n27401, A2 => n26954, B1 => n26948, B2 => 
                           n22592, ZN => n6313);
   U23484 : OAI22_X1 port map( A1 => n27404, A2 => n26954, B1 => n26948, B2 => 
                           n22591, ZN => n6314);
   U23485 : OAI22_X1 port map( A1 => n27407, A2 => n26954, B1 => n26948, B2 => 
                           n22590, ZN => n6315);
   U23486 : OAI22_X1 port map( A1 => n27410, A2 => n26954, B1 => n26948, B2 => 
                           n22589, ZN => n6316);
   U23487 : OAI22_X1 port map( A1 => n27413, A2 => n26954, B1 => n26948, B2 => 
                           n22588, ZN => n6317);
   U23488 : OAI22_X1 port map( A1 => n27416, A2 => n26954, B1 => n26948, B2 => 
                           n22587, ZN => n6318);
   U23489 : OAI22_X1 port map( A1 => n27419, A2 => n26954, B1 => n26948, B2 => 
                           n22586, ZN => n6319);
   U23490 : OAI22_X1 port map( A1 => n27422, A2 => n26954, B1 => n26948, B2 => 
                           n22585, ZN => n6320);
   U23491 : OAI22_X1 port map( A1 => n27425, A2 => n26955, B1 => n26948, B2 => 
                           n22584, ZN => n6321);
   U23492 : OAI22_X1 port map( A1 => n27428, A2 => n26955, B1 => n26949, B2 => 
                           n22583, ZN => n6322);
   U23493 : OAI22_X1 port map( A1 => n27431, A2 => n26955, B1 => n26949, B2 => 
                           n22582, ZN => n6323);
   U23494 : OAI22_X1 port map( A1 => n27434, A2 => n26955, B1 => n26949, B2 => 
                           n22581, ZN => n6324);
   U23495 : OAI22_X1 port map( A1 => n27437, A2 => n26955, B1 => n26949, B2 => 
                           n22580, ZN => n6325);
   U23496 : OAI22_X1 port map( A1 => n27440, A2 => n26955, B1 => n26949, B2 => 
                           n22579, ZN => n6326);
   U23497 : OAI22_X1 port map( A1 => n27443, A2 => n26955, B1 => n26949, B2 => 
                           n22578, ZN => n6327);
   U23498 : OAI22_X1 port map( A1 => n27446, A2 => n26955, B1 => n26949, B2 => 
                           n22577, ZN => n6328);
   U23499 : OAI22_X1 port map( A1 => n27449, A2 => n26955, B1 => n26949, B2 => 
                           n22576, ZN => n6329);
   U23500 : OAI22_X1 port map( A1 => n27452, A2 => n26955, B1 => n26949, B2 => 
                           n22575, ZN => n6330);
   U23501 : OAI22_X1 port map( A1 => n27455, A2 => n26955, B1 => n26949, B2 => 
                           n22574, ZN => n6331);
   U23502 : OAI22_X1 port map( A1 => n27458, A2 => n26955, B1 => n26949, B2 => 
                           n22573, ZN => n6332);
   U23503 : OAI22_X1 port map( A1 => n27461, A2 => n26956, B1 => n26949, B2 => 
                           n22572, ZN => n6333);
   U23504 : OAI22_X1 port map( A1 => n27318, A2 => n27156, B1 => n27150, B2 => 
                           n22427, ZN => n7374);
   U23505 : OAI22_X1 port map( A1 => n27321, A2 => n27156, B1 => n27150, B2 => 
                           n22426, ZN => n7375);
   U23506 : OAI22_X1 port map( A1 => n27324, A2 => n27156, B1 => n27150, B2 => 
                           n22425, ZN => n7376);
   U23507 : OAI22_X1 port map( A1 => n27327, A2 => n27156, B1 => n27150, B2 => 
                           n22424, ZN => n7377);
   U23508 : OAI22_X1 port map( A1 => n27330, A2 => n27156, B1 => n27150, B2 => 
                           n22423, ZN => n7378);
   U23509 : OAI22_X1 port map( A1 => n27333, A2 => n27156, B1 => n27150, B2 => 
                           n22422, ZN => n7379);
   U23510 : OAI22_X1 port map( A1 => n27336, A2 => n27156, B1 => n27150, B2 => 
                           n22421, ZN => n7380);
   U23511 : OAI22_X1 port map( A1 => n27339, A2 => n27156, B1 => n27150, B2 => 
                           n22420, ZN => n7381);
   U23512 : OAI22_X1 port map( A1 => n27342, A2 => n27156, B1 => n27150, B2 => 
                           n22419, ZN => n7382);
   U23513 : OAI22_X1 port map( A1 => n27345, A2 => n27156, B1 => n27150, B2 => 
                           n22418, ZN => n7383);
   U23514 : OAI22_X1 port map( A1 => n27348, A2 => n27156, B1 => n27150, B2 => 
                           n22417, ZN => n7384);
   U23515 : OAI22_X1 port map( A1 => n27351, A2 => n27157, B1 => n27150, B2 => 
                           n22416, ZN => n7385);
   U23516 : OAI22_X1 port map( A1 => n27354, A2 => n27157, B1 => n27151, B2 => 
                           n22415, ZN => n7386);
   U23517 : OAI22_X1 port map( A1 => n27357, A2 => n27157, B1 => n27151, B2 => 
                           n22414, ZN => n7387);
   U23518 : OAI22_X1 port map( A1 => n27360, A2 => n27157, B1 => n27151, B2 => 
                           n22413, ZN => n7388);
   U23519 : OAI22_X1 port map( A1 => n27363, A2 => n27157, B1 => n27151, B2 => 
                           n22412, ZN => n7389);
   U23520 : OAI22_X1 port map( A1 => n27366, A2 => n27157, B1 => n27151, B2 => 
                           n22411, ZN => n7390);
   U23521 : OAI22_X1 port map( A1 => n27369, A2 => n27157, B1 => n27151, B2 => 
                           n22410, ZN => n7391);
   U23522 : OAI22_X1 port map( A1 => n27372, A2 => n27157, B1 => n27151, B2 => 
                           n22409, ZN => n7392);
   U23523 : OAI22_X1 port map( A1 => n27375, A2 => n27157, B1 => n27151, B2 => 
                           n22408, ZN => n7393);
   U23524 : OAI22_X1 port map( A1 => n27378, A2 => n27157, B1 => n27151, B2 => 
                           n22407, ZN => n7394);
   U23525 : OAI22_X1 port map( A1 => n27381, A2 => n27157, B1 => n27151, B2 => 
                           n22406, ZN => n7395);
   U23526 : OAI22_X1 port map( A1 => n27384, A2 => n27157, B1 => n27151, B2 => 
                           n22405, ZN => n7396);
   U23527 : OAI22_X1 port map( A1 => n27387, A2 => n27158, B1 => n27151, B2 => 
                           n22404, ZN => n7397);
   U23528 : OAI22_X1 port map( A1 => n27390, A2 => n27158, B1 => n27152, B2 => 
                           n22403, ZN => n7398);
   U23529 : OAI22_X1 port map( A1 => n27393, A2 => n27158, B1 => n27152, B2 => 
                           n22402, ZN => n7399);
   U23530 : OAI22_X1 port map( A1 => n27396, A2 => n27158, B1 => n27152, B2 => 
                           n22401, ZN => n7400);
   U23531 : OAI22_X1 port map( A1 => n27399, A2 => n27158, B1 => n27152, B2 => 
                           n22400, ZN => n7401);
   U23532 : OAI22_X1 port map( A1 => n27402, A2 => n27158, B1 => n27152, B2 => 
                           n22399, ZN => n7402);
   U23533 : OAI22_X1 port map( A1 => n27405, A2 => n27158, B1 => n27152, B2 => 
                           n22398, ZN => n7403);
   U23534 : OAI22_X1 port map( A1 => n27408, A2 => n27158, B1 => n27152, B2 => 
                           n22397, ZN => n7404);
   U23535 : OAI22_X1 port map( A1 => n27411, A2 => n27158, B1 => n27152, B2 => 
                           n22396, ZN => n7405);
   U23536 : OAI22_X1 port map( A1 => n27414, A2 => n27158, B1 => n27152, B2 => 
                           n22395, ZN => n7406);
   U23537 : OAI22_X1 port map( A1 => n27417, A2 => n27158, B1 => n27152, B2 => 
                           n22394, ZN => n7407);
   U23538 : OAI22_X1 port map( A1 => n27420, A2 => n27158, B1 => n27152, B2 => 
                           n22393, ZN => n7408);
   U23539 : OAI22_X1 port map( A1 => n27423, A2 => n27159, B1 => n27152, B2 => 
                           n22392, ZN => n7409);
   U23540 : OAI22_X1 port map( A1 => n27426, A2 => n27159, B1 => n27153, B2 => 
                           n22391, ZN => n7410);
   U23541 : OAI22_X1 port map( A1 => n27429, A2 => n27159, B1 => n27153, B2 => 
                           n22390, ZN => n7411);
   U23542 : OAI22_X1 port map( A1 => n27432, A2 => n27159, B1 => n27153, B2 => 
                           n22389, ZN => n7412);
   U23543 : OAI22_X1 port map( A1 => n27435, A2 => n27159, B1 => n27153, B2 => 
                           n22388, ZN => n7413);
   U23544 : OAI22_X1 port map( A1 => n27438, A2 => n27159, B1 => n27153, B2 => 
                           n22387, ZN => n7414);
   U23545 : OAI22_X1 port map( A1 => n27441, A2 => n27159, B1 => n27153, B2 => 
                           n22386, ZN => n7415);
   U23546 : OAI22_X1 port map( A1 => n27444, A2 => n27159, B1 => n27153, B2 => 
                           n22385, ZN => n7416);
   U23547 : OAI22_X1 port map( A1 => n27447, A2 => n27159, B1 => n27153, B2 => 
                           n22384, ZN => n7417);
   U23548 : OAI22_X1 port map( A1 => n27450, A2 => n27159, B1 => n27153, B2 => 
                           n22383, ZN => n7418);
   U23549 : OAI22_X1 port map( A1 => n27453, A2 => n27159, B1 => n27153, B2 => 
                           n22382, ZN => n7419);
   U23550 : OAI22_X1 port map( A1 => n27456, A2 => n27159, B1 => n27153, B2 => 
                           n22381, ZN => n7420);
   U23551 : OAI22_X1 port map( A1 => n27459, A2 => n27160, B1 => n27153, B2 => 
                           n22380, ZN => n7421);
   U23552 : OAI22_X1 port map( A1 => n27320, A2 => n26928, B1 => n26922, B2 => 
                           n22307, ZN => n6158);
   U23553 : OAI22_X1 port map( A1 => n27323, A2 => n26928, B1 => n26922, B2 => 
                           n22306, ZN => n6159);
   U23554 : OAI22_X1 port map( A1 => n27326, A2 => n26928, B1 => n26922, B2 => 
                           n22305, ZN => n6160);
   U23555 : OAI22_X1 port map( A1 => n27329, A2 => n26928, B1 => n26922, B2 => 
                           n22304, ZN => n6161);
   U23556 : OAI22_X1 port map( A1 => n27332, A2 => n26928, B1 => n26922, B2 => 
                           n22303, ZN => n6162);
   U23557 : OAI22_X1 port map( A1 => n27335, A2 => n26928, B1 => n26922, B2 => 
                           n22302, ZN => n6163);
   U23558 : OAI22_X1 port map( A1 => n27338, A2 => n26928, B1 => n26922, B2 => 
                           n22301, ZN => n6164);
   U23559 : OAI22_X1 port map( A1 => n27341, A2 => n26928, B1 => n26922, B2 => 
                           n22300, ZN => n6165);
   U23560 : OAI22_X1 port map( A1 => n27344, A2 => n26928, B1 => n26922, B2 => 
                           n22299, ZN => n6166);
   U23561 : OAI22_X1 port map( A1 => n27347, A2 => n26928, B1 => n26922, B2 => 
                           n22298, ZN => n6167);
   U23562 : OAI22_X1 port map( A1 => n27350, A2 => n26928, B1 => n26922, B2 => 
                           n22297, ZN => n6168);
   U23563 : OAI22_X1 port map( A1 => n27353, A2 => n26929, B1 => n26922, B2 => 
                           n22296, ZN => n6169);
   U23564 : OAI22_X1 port map( A1 => n27356, A2 => n26929, B1 => n26923, B2 => 
                           n22295, ZN => n6170);
   U23565 : OAI22_X1 port map( A1 => n27359, A2 => n26929, B1 => n26923, B2 => 
                           n22294, ZN => n6171);
   U23566 : OAI22_X1 port map( A1 => n27362, A2 => n26929, B1 => n26923, B2 => 
                           n22293, ZN => n6172);
   U23567 : OAI22_X1 port map( A1 => n27365, A2 => n26929, B1 => n26923, B2 => 
                           n22292, ZN => n6173);
   U23568 : OAI22_X1 port map( A1 => n27368, A2 => n26929, B1 => n26923, B2 => 
                           n22291, ZN => n6174);
   U23569 : OAI22_X1 port map( A1 => n27371, A2 => n26929, B1 => n26923, B2 => 
                           n22290, ZN => n6175);
   U23570 : OAI22_X1 port map( A1 => n27374, A2 => n26929, B1 => n26923, B2 => 
                           n22289, ZN => n6176);
   U23571 : OAI22_X1 port map( A1 => n27377, A2 => n26929, B1 => n26923, B2 => 
                           n22288, ZN => n6177);
   U23572 : OAI22_X1 port map( A1 => n27380, A2 => n26929, B1 => n26923, B2 => 
                           n22287, ZN => n6178);
   U23573 : OAI22_X1 port map( A1 => n27383, A2 => n26929, B1 => n26923, B2 => 
                           n22286, ZN => n6179);
   U23574 : OAI22_X1 port map( A1 => n27386, A2 => n26929, B1 => n26923, B2 => 
                           n22285, ZN => n6180);
   U23575 : OAI22_X1 port map( A1 => n27389, A2 => n26930, B1 => n26923, B2 => 
                           n22284, ZN => n6181);
   U23576 : OAI22_X1 port map( A1 => n27392, A2 => n26930, B1 => n26924, B2 => 
                           n22283, ZN => n6182);
   U23577 : OAI22_X1 port map( A1 => n27395, A2 => n26930, B1 => n26924, B2 => 
                           n22282, ZN => n6183);
   U23578 : OAI22_X1 port map( A1 => n27398, A2 => n26930, B1 => n26924, B2 => 
                           n22281, ZN => n6184);
   U23579 : OAI22_X1 port map( A1 => n27401, A2 => n26930, B1 => n26924, B2 => 
                           n22280, ZN => n6185);
   U23580 : OAI22_X1 port map( A1 => n27404, A2 => n26930, B1 => n26924, B2 => 
                           n22279, ZN => n6186);
   U23581 : OAI22_X1 port map( A1 => n27407, A2 => n26930, B1 => n26924, B2 => 
                           n22278, ZN => n6187);
   U23582 : OAI22_X1 port map( A1 => n27410, A2 => n26930, B1 => n26924, B2 => 
                           n22277, ZN => n6188);
   U23583 : OAI22_X1 port map( A1 => n27413, A2 => n26930, B1 => n26924, B2 => 
                           n22276, ZN => n6189);
   U23584 : OAI22_X1 port map( A1 => n27416, A2 => n26930, B1 => n26924, B2 => 
                           n22275, ZN => n6190);
   U23585 : OAI22_X1 port map( A1 => n27419, A2 => n26930, B1 => n26924, B2 => 
                           n22274, ZN => n6191);
   U23586 : OAI22_X1 port map( A1 => n27422, A2 => n26930, B1 => n26924, B2 => 
                           n22273, ZN => n6192);
   U23587 : OAI22_X1 port map( A1 => n27425, A2 => n26931, B1 => n26924, B2 => 
                           n22272, ZN => n6193);
   U23588 : OAI22_X1 port map( A1 => n27428, A2 => n26931, B1 => n26925, B2 => 
                           n22271, ZN => n6194);
   U23589 : OAI22_X1 port map( A1 => n27431, A2 => n26931, B1 => n26925, B2 => 
                           n22270, ZN => n6195);
   U23590 : OAI22_X1 port map( A1 => n27434, A2 => n26931, B1 => n26925, B2 => 
                           n22269, ZN => n6196);
   U23591 : OAI22_X1 port map( A1 => n27437, A2 => n26931, B1 => n26925, B2 => 
                           n22268, ZN => n6197);
   U23592 : OAI22_X1 port map( A1 => n27440, A2 => n26931, B1 => n26925, B2 => 
                           n22267, ZN => n6198);
   U23593 : OAI22_X1 port map( A1 => n27443, A2 => n26931, B1 => n26925, B2 => 
                           n22266, ZN => n6199);
   U23594 : OAI22_X1 port map( A1 => n27446, A2 => n26931, B1 => n26925, B2 => 
                           n22265, ZN => n6200);
   U23595 : OAI22_X1 port map( A1 => n27449, A2 => n26931, B1 => n26925, B2 => 
                           n22264, ZN => n6201);
   U23596 : OAI22_X1 port map( A1 => n27452, A2 => n26931, B1 => n26925, B2 => 
                           n22263, ZN => n6202);
   U23597 : OAI22_X1 port map( A1 => n27455, A2 => n26931, B1 => n26925, B2 => 
                           n22262, ZN => n6203);
   U23598 : OAI22_X1 port map( A1 => n27458, A2 => n26931, B1 => n26925, B2 => 
                           n22261, ZN => n6204);
   U23599 : OAI22_X1 port map( A1 => n27461, A2 => n26932, B1 => n26925, B2 => 
                           n22260, ZN => n6205);
   U23600 : OAI22_X1 port map( A1 => n27320, A2 => n26940, B1 => n26934, B2 => 
                           n22231, ZN => n6222);
   U23601 : OAI22_X1 port map( A1 => n27323, A2 => n26940, B1 => n26934, B2 => 
                           n22230, ZN => n6223);
   U23602 : OAI22_X1 port map( A1 => n27326, A2 => n26940, B1 => n26934, B2 => 
                           n22229, ZN => n6224);
   U23603 : OAI22_X1 port map( A1 => n27329, A2 => n26940, B1 => n26934, B2 => 
                           n22228, ZN => n6225);
   U23604 : OAI22_X1 port map( A1 => n27332, A2 => n26940, B1 => n26934, B2 => 
                           n22227, ZN => n6226);
   U23605 : OAI22_X1 port map( A1 => n27335, A2 => n26940, B1 => n26934, B2 => 
                           n22226, ZN => n6227);
   U23606 : OAI22_X1 port map( A1 => n27338, A2 => n26940, B1 => n26934, B2 => 
                           n22225, ZN => n6228);
   U23607 : OAI22_X1 port map( A1 => n27341, A2 => n26940, B1 => n26934, B2 => 
                           n22224, ZN => n6229);
   U23608 : OAI22_X1 port map( A1 => n27344, A2 => n26940, B1 => n26934, B2 => 
                           n22223, ZN => n6230);
   U23609 : OAI22_X1 port map( A1 => n27347, A2 => n26940, B1 => n26934, B2 => 
                           n22222, ZN => n6231);
   U23610 : OAI22_X1 port map( A1 => n27350, A2 => n26940, B1 => n26934, B2 => 
                           n22221, ZN => n6232);
   U23611 : OAI22_X1 port map( A1 => n27353, A2 => n26941, B1 => n26934, B2 => 
                           n22220, ZN => n6233);
   U23612 : OAI22_X1 port map( A1 => n27356, A2 => n26941, B1 => n26935, B2 => 
                           n22219, ZN => n6234);
   U23613 : OAI22_X1 port map( A1 => n27359, A2 => n26941, B1 => n26935, B2 => 
                           n22218, ZN => n6235);
   U23614 : OAI22_X1 port map( A1 => n27362, A2 => n26941, B1 => n26935, B2 => 
                           n22217, ZN => n6236);
   U23615 : OAI22_X1 port map( A1 => n27365, A2 => n26941, B1 => n26935, B2 => 
                           n22216, ZN => n6237);
   U23616 : OAI22_X1 port map( A1 => n27368, A2 => n26941, B1 => n26935, B2 => 
                           n22215, ZN => n6238);
   U23617 : OAI22_X1 port map( A1 => n27371, A2 => n26941, B1 => n26935, B2 => 
                           n22214, ZN => n6239);
   U23618 : OAI22_X1 port map( A1 => n27374, A2 => n26941, B1 => n26935, B2 => 
                           n22213, ZN => n6240);
   U23619 : OAI22_X1 port map( A1 => n27377, A2 => n26941, B1 => n26935, B2 => 
                           n22212, ZN => n6241);
   U23620 : OAI22_X1 port map( A1 => n27380, A2 => n26941, B1 => n26935, B2 => 
                           n22211, ZN => n6242);
   U23621 : OAI22_X1 port map( A1 => n27383, A2 => n26941, B1 => n26935, B2 => 
                           n22210, ZN => n6243);
   U23622 : OAI22_X1 port map( A1 => n27386, A2 => n26941, B1 => n26935, B2 => 
                           n22209, ZN => n6244);
   U23623 : OAI22_X1 port map( A1 => n27389, A2 => n26942, B1 => n26935, B2 => 
                           n22208, ZN => n6245);
   U23624 : OAI22_X1 port map( A1 => n27392, A2 => n26942, B1 => n26936, B2 => 
                           n22207, ZN => n6246);
   U23625 : OAI22_X1 port map( A1 => n27395, A2 => n26942, B1 => n26936, B2 => 
                           n22206, ZN => n6247);
   U23626 : OAI22_X1 port map( A1 => n27398, A2 => n26942, B1 => n26936, B2 => 
                           n22205, ZN => n6248);
   U23627 : OAI22_X1 port map( A1 => n27401, A2 => n26942, B1 => n26936, B2 => 
                           n22204, ZN => n6249);
   U23628 : OAI22_X1 port map( A1 => n27404, A2 => n26942, B1 => n26936, B2 => 
                           n22203, ZN => n6250);
   U23629 : OAI22_X1 port map( A1 => n27407, A2 => n26942, B1 => n26936, B2 => 
                           n22202, ZN => n6251);
   U23630 : OAI22_X1 port map( A1 => n27410, A2 => n26942, B1 => n26936, B2 => 
                           n22201, ZN => n6252);
   U23631 : OAI22_X1 port map( A1 => n27413, A2 => n26942, B1 => n26936, B2 => 
                           n22200, ZN => n6253);
   U23632 : OAI22_X1 port map( A1 => n27416, A2 => n26942, B1 => n26936, B2 => 
                           n22199, ZN => n6254);
   U23633 : OAI22_X1 port map( A1 => n27419, A2 => n26942, B1 => n26936, B2 => 
                           n22198, ZN => n6255);
   U23634 : OAI22_X1 port map( A1 => n27422, A2 => n26942, B1 => n26936, B2 => 
                           n22197, ZN => n6256);
   U23635 : OAI22_X1 port map( A1 => n27425, A2 => n26943, B1 => n26936, B2 => 
                           n22196, ZN => n6257);
   U23636 : OAI22_X1 port map( A1 => n27428, A2 => n26943, B1 => n26937, B2 => 
                           n22195, ZN => n6258);
   U23637 : OAI22_X1 port map( A1 => n27431, A2 => n26943, B1 => n26937, B2 => 
                           n22194, ZN => n6259);
   U23638 : OAI22_X1 port map( A1 => n27434, A2 => n26943, B1 => n26937, B2 => 
                           n22193, ZN => n6260);
   U23639 : OAI22_X1 port map( A1 => n27437, A2 => n26943, B1 => n26937, B2 => 
                           n22192, ZN => n6261);
   U23640 : OAI22_X1 port map( A1 => n27440, A2 => n26943, B1 => n26937, B2 => 
                           n22191, ZN => n6262);
   U23641 : OAI22_X1 port map( A1 => n27443, A2 => n26943, B1 => n26937, B2 => 
                           n22190, ZN => n6263);
   U23642 : OAI22_X1 port map( A1 => n27446, A2 => n26943, B1 => n26937, B2 => 
                           n22189, ZN => n6264);
   U23643 : OAI22_X1 port map( A1 => n27449, A2 => n26943, B1 => n26937, B2 => 
                           n22188, ZN => n6265);
   U23644 : OAI22_X1 port map( A1 => n27452, A2 => n26943, B1 => n26937, B2 => 
                           n22187, ZN => n6266);
   U23645 : OAI22_X1 port map( A1 => n27455, A2 => n26943, B1 => n26937, B2 => 
                           n22186, ZN => n6267);
   U23646 : OAI22_X1 port map( A1 => n27458, A2 => n26943, B1 => n26937, B2 => 
                           n22185, ZN => n6268);
   U23647 : OAI22_X1 port map( A1 => n27461, A2 => n26944, B1 => n26937, B2 => 
                           n22184, ZN => n6269);
   U23648 : OAI22_X1 port map( A1 => n27278, A2 => n27318, B1 => n27270, B2 => 
                           n22167, ZN => n8014);
   U23649 : OAI22_X1 port map( A1 => n27278, A2 => n27321, B1 => n27270, B2 => 
                           n22166, ZN => n8015);
   U23650 : OAI22_X1 port map( A1 => n27278, A2 => n27324, B1 => n27270, B2 => 
                           n22165, ZN => n8016);
   U23651 : OAI22_X1 port map( A1 => n27278, A2 => n27327, B1 => n27270, B2 => 
                           n22164, ZN => n8017);
   U23652 : OAI22_X1 port map( A1 => n27278, A2 => n27330, B1 => n27270, B2 => 
                           n22163, ZN => n8018);
   U23653 : OAI22_X1 port map( A1 => n27278, A2 => n27333, B1 => n27270, B2 => 
                           n22162, ZN => n8019);
   U23654 : OAI22_X1 port map( A1 => n27278, A2 => n27336, B1 => n27270, B2 => 
                           n22161, ZN => n8020);
   U23655 : OAI22_X1 port map( A1 => n27278, A2 => n27339, B1 => n27270, B2 => 
                           n22160, ZN => n8021);
   U23656 : OAI22_X1 port map( A1 => n27278, A2 => n27342, B1 => n27270, B2 => 
                           n22159, ZN => n8022);
   U23657 : OAI22_X1 port map( A1 => n27278, A2 => n27345, B1 => n27270, B2 => 
                           n22158, ZN => n8023);
   U23658 : OAI22_X1 port map( A1 => n27278, A2 => n27348, B1 => n27270, B2 => 
                           n22157, ZN => n8024);
   U23659 : OAI22_X1 port map( A1 => n27278, A2 => n27351, B1 => n27270, B2 => 
                           n22156, ZN => n8025);
   U23660 : OAI22_X1 port map( A1 => n27278, A2 => n27354, B1 => n27271, B2 => 
                           n22155, ZN => n8026);
   U23661 : OAI22_X1 port map( A1 => n27279, A2 => n27357, B1 => n27271, B2 => 
                           n22154, ZN => n8027);
   U23662 : OAI22_X1 port map( A1 => n27279, A2 => n27360, B1 => n27271, B2 => 
                           n22153, ZN => n8028);
   U23663 : OAI22_X1 port map( A1 => n27279, A2 => n27363, B1 => n27271, B2 => 
                           n22152, ZN => n8029);
   U23664 : OAI22_X1 port map( A1 => n27279, A2 => n27366, B1 => n27271, B2 => 
                           n22151, ZN => n8030);
   U23665 : OAI22_X1 port map( A1 => n27279, A2 => n27369, B1 => n27271, B2 => 
                           n22150, ZN => n8031);
   U23666 : OAI22_X1 port map( A1 => n27279, A2 => n27372, B1 => n27271, B2 => 
                           n22149, ZN => n8032);
   U23667 : OAI22_X1 port map( A1 => n27279, A2 => n27375, B1 => n27271, B2 => 
                           n22148, ZN => n8033);
   U23668 : OAI22_X1 port map( A1 => n27279, A2 => n27378, B1 => n27271, B2 => 
                           n22147, ZN => n8034);
   U23669 : OAI22_X1 port map( A1 => n27279, A2 => n27381, B1 => n27271, B2 => 
                           n22146, ZN => n8035);
   U23670 : OAI22_X1 port map( A1 => n27279, A2 => n27384, B1 => n27271, B2 => 
                           n22145, ZN => n8036);
   U23671 : OAI22_X1 port map( A1 => n27279, A2 => n27387, B1 => n27271, B2 => 
                           n22144, ZN => n8037);
   U23672 : OAI22_X1 port map( A1 => n27279, A2 => n27390, B1 => n27272, B2 => 
                           n22143, ZN => n8038);
   U23673 : OAI22_X1 port map( A1 => n27279, A2 => n27393, B1 => n27272, B2 => 
                           n22142, ZN => n8039);
   U23674 : OAI22_X1 port map( A1 => n27280, A2 => n27396, B1 => n27272, B2 => 
                           n22141, ZN => n8040);
   U23675 : OAI22_X1 port map( A1 => n27280, A2 => n27399, B1 => n27272, B2 => 
                           n22140, ZN => n8041);
   U23676 : OAI22_X1 port map( A1 => n27280, A2 => n27402, B1 => n27272, B2 => 
                           n22139, ZN => n8042);
   U23677 : OAI22_X1 port map( A1 => n27280, A2 => n27405, B1 => n27272, B2 => 
                           n22138, ZN => n8043);
   U23678 : OAI22_X1 port map( A1 => n27280, A2 => n27408, B1 => n27272, B2 => 
                           n22137, ZN => n8044);
   U23679 : OAI22_X1 port map( A1 => n27280, A2 => n27411, B1 => n27272, B2 => 
                           n22136, ZN => n8045);
   U23680 : OAI22_X1 port map( A1 => n27280, A2 => n27414, B1 => n27272, B2 => 
                           n22135, ZN => n8046);
   U23681 : OAI22_X1 port map( A1 => n27280, A2 => n27417, B1 => n27272, B2 => 
                           n22134, ZN => n8047);
   U23682 : OAI22_X1 port map( A1 => n27280, A2 => n27420, B1 => n27272, B2 => 
                           n22133, ZN => n8048);
   U23683 : OAI22_X1 port map( A1 => n27280, A2 => n27423, B1 => n27272, B2 => 
                           n22132, ZN => n8049);
   U23684 : OAI22_X1 port map( A1 => n27280, A2 => n27426, B1 => n27273, B2 => 
                           n22131, ZN => n8050);
   U23685 : OAI22_X1 port map( A1 => n27280, A2 => n27429, B1 => n27273, B2 => 
                           n22130, ZN => n8051);
   U23686 : OAI22_X1 port map( A1 => n27280, A2 => n27432, B1 => n27273, B2 => 
                           n22129, ZN => n8052);
   U23687 : OAI22_X1 port map( A1 => n27281, A2 => n27435, B1 => n27273, B2 => 
                           n22128, ZN => n8053);
   U23688 : OAI22_X1 port map( A1 => n27281, A2 => n27438, B1 => n27273, B2 => 
                           n22127, ZN => n8054);
   U23689 : OAI22_X1 port map( A1 => n27281, A2 => n27441, B1 => n27273, B2 => 
                           n22126, ZN => n8055);
   U23690 : OAI22_X1 port map( A1 => n27281, A2 => n27444, B1 => n27273, B2 => 
                           n22125, ZN => n8056);
   U23691 : OAI22_X1 port map( A1 => n27281, A2 => n27447, B1 => n27273, B2 => 
                           n22124, ZN => n8057);
   U23692 : OAI22_X1 port map( A1 => n27281, A2 => n27450, B1 => n27273, B2 => 
                           n22123, ZN => n8058);
   U23693 : OAI22_X1 port map( A1 => n27281, A2 => n27453, B1 => n27273, B2 => 
                           n22122, ZN => n8059);
   U23694 : OAI22_X1 port map( A1 => n27281, A2 => n27456, B1 => n27273, B2 => 
                           n22121, ZN => n8060);
   U23695 : OAI22_X1 port map( A1 => n27281, A2 => n27459, B1 => n27273, B2 => 
                           n22120, ZN => n8061);
   U23696 : OAI22_X1 port map( A1 => n27318, A2 => n27264, B1 => n27258, B2 => 
                           n22107, ZN => n7950);
   U23697 : OAI22_X1 port map( A1 => n27321, A2 => n27264, B1 => n27258, B2 => 
                           n22106, ZN => n7951);
   U23698 : OAI22_X1 port map( A1 => n27324, A2 => n27264, B1 => n27258, B2 => 
                           n22105, ZN => n7952);
   U23699 : OAI22_X1 port map( A1 => n27327, A2 => n27264, B1 => n27258, B2 => 
                           n22104, ZN => n7953);
   U23700 : OAI22_X1 port map( A1 => n27330, A2 => n27264, B1 => n27258, B2 => 
                           n22103, ZN => n7954);
   U23701 : OAI22_X1 port map( A1 => n27333, A2 => n27264, B1 => n27258, B2 => 
                           n22102, ZN => n7955);
   U23702 : OAI22_X1 port map( A1 => n27336, A2 => n27264, B1 => n27258, B2 => 
                           n22101, ZN => n7956);
   U23703 : OAI22_X1 port map( A1 => n27339, A2 => n27264, B1 => n27258, B2 => 
                           n22100, ZN => n7957);
   U23704 : OAI22_X1 port map( A1 => n27342, A2 => n27264, B1 => n27258, B2 => 
                           n22099, ZN => n7958);
   U23705 : OAI22_X1 port map( A1 => n27345, A2 => n27264, B1 => n27258, B2 => 
                           n22098, ZN => n7959);
   U23706 : OAI22_X1 port map( A1 => n27348, A2 => n27264, B1 => n27258, B2 => 
                           n22097, ZN => n7960);
   U23707 : OAI22_X1 port map( A1 => n27351, A2 => n27265, B1 => n27258, B2 => 
                           n22096, ZN => n7961);
   U23708 : OAI22_X1 port map( A1 => n27354, A2 => n27265, B1 => n27259, B2 => 
                           n22095, ZN => n7962);
   U23709 : OAI22_X1 port map( A1 => n27357, A2 => n27265, B1 => n27259, B2 => 
                           n22094, ZN => n7963);
   U23710 : OAI22_X1 port map( A1 => n27360, A2 => n27265, B1 => n27259, B2 => 
                           n22093, ZN => n7964);
   U23711 : OAI22_X1 port map( A1 => n27363, A2 => n27265, B1 => n27259, B2 => 
                           n22092, ZN => n7965);
   U23712 : OAI22_X1 port map( A1 => n27366, A2 => n27265, B1 => n27259, B2 => 
                           n22091, ZN => n7966);
   U23713 : OAI22_X1 port map( A1 => n27369, A2 => n27265, B1 => n27259, B2 => 
                           n22090, ZN => n7967);
   U23714 : OAI22_X1 port map( A1 => n27372, A2 => n27265, B1 => n27259, B2 => 
                           n22089, ZN => n7968);
   U23715 : OAI22_X1 port map( A1 => n27375, A2 => n27265, B1 => n27259, B2 => 
                           n22088, ZN => n7969);
   U23716 : OAI22_X1 port map( A1 => n27378, A2 => n27265, B1 => n27259, B2 => 
                           n22087, ZN => n7970);
   U23717 : OAI22_X1 port map( A1 => n27381, A2 => n27265, B1 => n27259, B2 => 
                           n22086, ZN => n7971);
   U23718 : OAI22_X1 port map( A1 => n27384, A2 => n27265, B1 => n27259, B2 => 
                           n22085, ZN => n7972);
   U23719 : OAI22_X1 port map( A1 => n27387, A2 => n27266, B1 => n27259, B2 => 
                           n22084, ZN => n7973);
   U23720 : OAI22_X1 port map( A1 => n27390, A2 => n27266, B1 => n27260, B2 => 
                           n22083, ZN => n7974);
   U23721 : OAI22_X1 port map( A1 => n27393, A2 => n27266, B1 => n27260, B2 => 
                           n22082, ZN => n7975);
   U23722 : OAI22_X1 port map( A1 => n27396, A2 => n27266, B1 => n27260, B2 => 
                           n22081, ZN => n7976);
   U23723 : OAI22_X1 port map( A1 => n27399, A2 => n27266, B1 => n27260, B2 => 
                           n22080, ZN => n7977);
   U23724 : OAI22_X1 port map( A1 => n27402, A2 => n27266, B1 => n27260, B2 => 
                           n22079, ZN => n7978);
   U23725 : OAI22_X1 port map( A1 => n27405, A2 => n27266, B1 => n27260, B2 => 
                           n22078, ZN => n7979);
   U23726 : OAI22_X1 port map( A1 => n27408, A2 => n27266, B1 => n27260, B2 => 
                           n22077, ZN => n7980);
   U23727 : OAI22_X1 port map( A1 => n27411, A2 => n27266, B1 => n27260, B2 => 
                           n22076, ZN => n7981);
   U23728 : OAI22_X1 port map( A1 => n27414, A2 => n27266, B1 => n27260, B2 => 
                           n22075, ZN => n7982);
   U23729 : OAI22_X1 port map( A1 => n27417, A2 => n27266, B1 => n27260, B2 => 
                           n22074, ZN => n7983);
   U23730 : OAI22_X1 port map( A1 => n27420, A2 => n27266, B1 => n27260, B2 => 
                           n22073, ZN => n7984);
   U23731 : OAI22_X1 port map( A1 => n27423, A2 => n27267, B1 => n27260, B2 => 
                           n22072, ZN => n7985);
   U23732 : OAI22_X1 port map( A1 => n27426, A2 => n27267, B1 => n27261, B2 => 
                           n22071, ZN => n7986);
   U23733 : OAI22_X1 port map( A1 => n27429, A2 => n27267, B1 => n27261, B2 => 
                           n22070, ZN => n7987);
   U23734 : OAI22_X1 port map( A1 => n27432, A2 => n27267, B1 => n27261, B2 => 
                           n22069, ZN => n7988);
   U23735 : OAI22_X1 port map( A1 => n27435, A2 => n27267, B1 => n27261, B2 => 
                           n22068, ZN => n7989);
   U23736 : OAI22_X1 port map( A1 => n27438, A2 => n27267, B1 => n27261, B2 => 
                           n22067, ZN => n7990);
   U23737 : OAI22_X1 port map( A1 => n27441, A2 => n27267, B1 => n27261, B2 => 
                           n22066, ZN => n7991);
   U23738 : OAI22_X1 port map( A1 => n27444, A2 => n27267, B1 => n27261, B2 => 
                           n22065, ZN => n7992);
   U23739 : OAI22_X1 port map( A1 => n27447, A2 => n27267, B1 => n27261, B2 => 
                           n22064, ZN => n7993);
   U23740 : OAI22_X1 port map( A1 => n27450, A2 => n27267, B1 => n27261, B2 => 
                           n22063, ZN => n7994);
   U23741 : OAI22_X1 port map( A1 => n27453, A2 => n27267, B1 => n27261, B2 => 
                           n22062, ZN => n7995);
   U23742 : OAI22_X1 port map( A1 => n27456, A2 => n27267, B1 => n27261, B2 => 
                           n22061, ZN => n7996);
   U23743 : OAI22_X1 port map( A1 => n27459, A2 => n27268, B1 => n27261, B2 => 
                           n22060, ZN => n7997);
   U23744 : OAI22_X1 port map( A1 => n27318, A2 => n27228, B1 => n27222, B2 => 
                           n21927, ZN => n7758);
   U23745 : OAI22_X1 port map( A1 => n27321, A2 => n27228, B1 => n27222, B2 => 
                           n21926, ZN => n7759);
   U23746 : OAI22_X1 port map( A1 => n27324, A2 => n27228, B1 => n27222, B2 => 
                           n21925, ZN => n7760);
   U23747 : OAI22_X1 port map( A1 => n27327, A2 => n27228, B1 => n27222, B2 => 
                           n21924, ZN => n7761);
   U23748 : OAI22_X1 port map( A1 => n27330, A2 => n27228, B1 => n27222, B2 => 
                           n21923, ZN => n7762);
   U23749 : OAI22_X1 port map( A1 => n27333, A2 => n27228, B1 => n27222, B2 => 
                           n21922, ZN => n7763);
   U23750 : OAI22_X1 port map( A1 => n27336, A2 => n27228, B1 => n27222, B2 => 
                           n21921, ZN => n7764);
   U23751 : OAI22_X1 port map( A1 => n27339, A2 => n27228, B1 => n27222, B2 => 
                           n21920, ZN => n7765);
   U23752 : OAI22_X1 port map( A1 => n27342, A2 => n27228, B1 => n27222, B2 => 
                           n21919, ZN => n7766);
   U23753 : OAI22_X1 port map( A1 => n27345, A2 => n27228, B1 => n27222, B2 => 
                           n21918, ZN => n7767);
   U23754 : OAI22_X1 port map( A1 => n27348, A2 => n27228, B1 => n27222, B2 => 
                           n21917, ZN => n7768);
   U23755 : OAI22_X1 port map( A1 => n27351, A2 => n27229, B1 => n27222, B2 => 
                           n21916, ZN => n7769);
   U23756 : OAI22_X1 port map( A1 => n27354, A2 => n27229, B1 => n27223, B2 => 
                           n21915, ZN => n7770);
   U23757 : OAI22_X1 port map( A1 => n27357, A2 => n27229, B1 => n27223, B2 => 
                           n21914, ZN => n7771);
   U23758 : OAI22_X1 port map( A1 => n27360, A2 => n27229, B1 => n27223, B2 => 
                           n21913, ZN => n7772);
   U23759 : OAI22_X1 port map( A1 => n27363, A2 => n27229, B1 => n27223, B2 => 
                           n21912, ZN => n7773);
   U23760 : OAI22_X1 port map( A1 => n27366, A2 => n27229, B1 => n27223, B2 => 
                           n21911, ZN => n7774);
   U23761 : OAI22_X1 port map( A1 => n27369, A2 => n27229, B1 => n27223, B2 => 
                           n21910, ZN => n7775);
   U23762 : OAI22_X1 port map( A1 => n27372, A2 => n27229, B1 => n27223, B2 => 
                           n21909, ZN => n7776);
   U23763 : OAI22_X1 port map( A1 => n27375, A2 => n27229, B1 => n27223, B2 => 
                           n21908, ZN => n7777);
   U23764 : OAI22_X1 port map( A1 => n27378, A2 => n27229, B1 => n27223, B2 => 
                           n21907, ZN => n7778);
   U23765 : OAI22_X1 port map( A1 => n27381, A2 => n27229, B1 => n27223, B2 => 
                           n21906, ZN => n7779);
   U23766 : OAI22_X1 port map( A1 => n27384, A2 => n27229, B1 => n27223, B2 => 
                           n21905, ZN => n7780);
   U23767 : OAI22_X1 port map( A1 => n27387, A2 => n27230, B1 => n27223, B2 => 
                           n21904, ZN => n7781);
   U23768 : OAI22_X1 port map( A1 => n27390, A2 => n27230, B1 => n27224, B2 => 
                           n21903, ZN => n7782);
   U23769 : OAI22_X1 port map( A1 => n27393, A2 => n27230, B1 => n27224, B2 => 
                           n21902, ZN => n7783);
   U23770 : OAI22_X1 port map( A1 => n27396, A2 => n27230, B1 => n27224, B2 => 
                           n21901, ZN => n7784);
   U23771 : OAI22_X1 port map( A1 => n27399, A2 => n27230, B1 => n27224, B2 => 
                           n21900, ZN => n7785);
   U23772 : OAI22_X1 port map( A1 => n27402, A2 => n27230, B1 => n27224, B2 => 
                           n21899, ZN => n7786);
   U23773 : OAI22_X1 port map( A1 => n27405, A2 => n27230, B1 => n27224, B2 => 
                           n21898, ZN => n7787);
   U23774 : OAI22_X1 port map( A1 => n27408, A2 => n27230, B1 => n27224, B2 => 
                           n21897, ZN => n7788);
   U23775 : OAI22_X1 port map( A1 => n27411, A2 => n27230, B1 => n27224, B2 => 
                           n21896, ZN => n7789);
   U23776 : OAI22_X1 port map( A1 => n27414, A2 => n27230, B1 => n27224, B2 => 
                           n21895, ZN => n7790);
   U23777 : OAI22_X1 port map( A1 => n27417, A2 => n27230, B1 => n27224, B2 => 
                           n21894, ZN => n7791);
   U23778 : OAI22_X1 port map( A1 => n27420, A2 => n27230, B1 => n27224, B2 => 
                           n21893, ZN => n7792);
   U23779 : OAI22_X1 port map( A1 => n27423, A2 => n27231, B1 => n27224, B2 => 
                           n21892, ZN => n7793);
   U23780 : OAI22_X1 port map( A1 => n27426, A2 => n27231, B1 => n27225, B2 => 
                           n21891, ZN => n7794);
   U23781 : OAI22_X1 port map( A1 => n27429, A2 => n27231, B1 => n27225, B2 => 
                           n21890, ZN => n7795);
   U23782 : OAI22_X1 port map( A1 => n27432, A2 => n27231, B1 => n27225, B2 => 
                           n21889, ZN => n7796);
   U23783 : OAI22_X1 port map( A1 => n27435, A2 => n27231, B1 => n27225, B2 => 
                           n21888, ZN => n7797);
   U23784 : OAI22_X1 port map( A1 => n27438, A2 => n27231, B1 => n27225, B2 => 
                           n21887, ZN => n7798);
   U23785 : OAI22_X1 port map( A1 => n27441, A2 => n27231, B1 => n27225, B2 => 
                           n21886, ZN => n7799);
   U23786 : OAI22_X1 port map( A1 => n27444, A2 => n27231, B1 => n27225, B2 => 
                           n21885, ZN => n7800);
   U23787 : OAI22_X1 port map( A1 => n27447, A2 => n27231, B1 => n27225, B2 => 
                           n21884, ZN => n7801);
   U23788 : OAI22_X1 port map( A1 => n27450, A2 => n27231, B1 => n27225, B2 => 
                           n21883, ZN => n7802);
   U23789 : OAI22_X1 port map( A1 => n27453, A2 => n27231, B1 => n27225, B2 => 
                           n21882, ZN => n7803);
   U23790 : OAI22_X1 port map( A1 => n27456, A2 => n27231, B1 => n27225, B2 => 
                           n21881, ZN => n7804);
   U23791 : OAI22_X1 port map( A1 => n27459, A2 => n27232, B1 => n27225, B2 => 
                           n21880, ZN => n7805);
   U23792 : OAI22_X1 port map( A1 => n27318, A2 => n27204, B1 => n27198, B2 => 
                           n21867, ZN => n7630);
   U23793 : OAI22_X1 port map( A1 => n27321, A2 => n27204, B1 => n27198, B2 => 
                           n21866, ZN => n7631);
   U23794 : OAI22_X1 port map( A1 => n27324, A2 => n27204, B1 => n27198, B2 => 
                           n21865, ZN => n7632);
   U23795 : OAI22_X1 port map( A1 => n27327, A2 => n27204, B1 => n27198, B2 => 
                           n21864, ZN => n7633);
   U23796 : OAI22_X1 port map( A1 => n27330, A2 => n27204, B1 => n27198, B2 => 
                           n21863, ZN => n7634);
   U23797 : OAI22_X1 port map( A1 => n27333, A2 => n27204, B1 => n27198, B2 => 
                           n21862, ZN => n7635);
   U23798 : OAI22_X1 port map( A1 => n27336, A2 => n27204, B1 => n27198, B2 => 
                           n21861, ZN => n7636);
   U23799 : OAI22_X1 port map( A1 => n27339, A2 => n27204, B1 => n27198, B2 => 
                           n21860, ZN => n7637);
   U23800 : OAI22_X1 port map( A1 => n27342, A2 => n27204, B1 => n27198, B2 => 
                           n21859, ZN => n7638);
   U23801 : OAI22_X1 port map( A1 => n27345, A2 => n27204, B1 => n27198, B2 => 
                           n21858, ZN => n7639);
   U23802 : OAI22_X1 port map( A1 => n27348, A2 => n27204, B1 => n27198, B2 => 
                           n21857, ZN => n7640);
   U23803 : OAI22_X1 port map( A1 => n27351, A2 => n27205, B1 => n27198, B2 => 
                           n21856, ZN => n7641);
   U23804 : OAI22_X1 port map( A1 => n27354, A2 => n27205, B1 => n27199, B2 => 
                           n21855, ZN => n7642);
   U23805 : OAI22_X1 port map( A1 => n27357, A2 => n27205, B1 => n27199, B2 => 
                           n21854, ZN => n7643);
   U23806 : OAI22_X1 port map( A1 => n27360, A2 => n27205, B1 => n27199, B2 => 
                           n21853, ZN => n7644);
   U23807 : OAI22_X1 port map( A1 => n27363, A2 => n27205, B1 => n27199, B2 => 
                           n21852, ZN => n7645);
   U23808 : OAI22_X1 port map( A1 => n27366, A2 => n27205, B1 => n27199, B2 => 
                           n21851, ZN => n7646);
   U23809 : OAI22_X1 port map( A1 => n27369, A2 => n27205, B1 => n27199, B2 => 
                           n21850, ZN => n7647);
   U23810 : OAI22_X1 port map( A1 => n27372, A2 => n27205, B1 => n27199, B2 => 
                           n21849, ZN => n7648);
   U23811 : OAI22_X1 port map( A1 => n27375, A2 => n27205, B1 => n27199, B2 => 
                           n21848, ZN => n7649);
   U23812 : OAI22_X1 port map( A1 => n27378, A2 => n27205, B1 => n27199, B2 => 
                           n21847, ZN => n7650);
   U23813 : OAI22_X1 port map( A1 => n27381, A2 => n27205, B1 => n27199, B2 => 
                           n21846, ZN => n7651);
   U23814 : OAI22_X1 port map( A1 => n27384, A2 => n27205, B1 => n27199, B2 => 
                           n21845, ZN => n7652);
   U23815 : OAI22_X1 port map( A1 => n27387, A2 => n27206, B1 => n27199, B2 => 
                           n21844, ZN => n7653);
   U23816 : OAI22_X1 port map( A1 => n27390, A2 => n27206, B1 => n27200, B2 => 
                           n21843, ZN => n7654);
   U23817 : OAI22_X1 port map( A1 => n27393, A2 => n27206, B1 => n27200, B2 => 
                           n21842, ZN => n7655);
   U23818 : OAI22_X1 port map( A1 => n27396, A2 => n27206, B1 => n27200, B2 => 
                           n21841, ZN => n7656);
   U23819 : OAI22_X1 port map( A1 => n27399, A2 => n27206, B1 => n27200, B2 => 
                           n21840, ZN => n7657);
   U23820 : OAI22_X1 port map( A1 => n27402, A2 => n27206, B1 => n27200, B2 => 
                           n21839, ZN => n7658);
   U23821 : OAI22_X1 port map( A1 => n27405, A2 => n27206, B1 => n27200, B2 => 
                           n21838, ZN => n7659);
   U23822 : OAI22_X1 port map( A1 => n27408, A2 => n27206, B1 => n27200, B2 => 
                           n21837, ZN => n7660);
   U23823 : OAI22_X1 port map( A1 => n27411, A2 => n27206, B1 => n27200, B2 => 
                           n21836, ZN => n7661);
   U23824 : OAI22_X1 port map( A1 => n27414, A2 => n27206, B1 => n27200, B2 => 
                           n21835, ZN => n7662);
   U23825 : OAI22_X1 port map( A1 => n27417, A2 => n27206, B1 => n27200, B2 => 
                           n21834, ZN => n7663);
   U23826 : OAI22_X1 port map( A1 => n27420, A2 => n27206, B1 => n27200, B2 => 
                           n21833, ZN => n7664);
   U23827 : OAI22_X1 port map( A1 => n27423, A2 => n27207, B1 => n27200, B2 => 
                           n21832, ZN => n7665);
   U23828 : OAI22_X1 port map( A1 => n27426, A2 => n27207, B1 => n27201, B2 => 
                           n21831, ZN => n7666);
   U23829 : OAI22_X1 port map( A1 => n27429, A2 => n27207, B1 => n27201, B2 => 
                           n21830, ZN => n7667);
   U23830 : OAI22_X1 port map( A1 => n27432, A2 => n27207, B1 => n27201, B2 => 
                           n21829, ZN => n7668);
   U23831 : OAI22_X1 port map( A1 => n27435, A2 => n27207, B1 => n27201, B2 => 
                           n21828, ZN => n7669);
   U23832 : OAI22_X1 port map( A1 => n27438, A2 => n27207, B1 => n27201, B2 => 
                           n21827, ZN => n7670);
   U23833 : OAI22_X1 port map( A1 => n27441, A2 => n27207, B1 => n27201, B2 => 
                           n21826, ZN => n7671);
   U23834 : OAI22_X1 port map( A1 => n27444, A2 => n27207, B1 => n27201, B2 => 
                           n21825, ZN => n7672);
   U23835 : OAI22_X1 port map( A1 => n27447, A2 => n27207, B1 => n27201, B2 => 
                           n21824, ZN => n7673);
   U23836 : OAI22_X1 port map( A1 => n27450, A2 => n27207, B1 => n27201, B2 => 
                           n21823, ZN => n7674);
   U23837 : OAI22_X1 port map( A1 => n27453, A2 => n27207, B1 => n27201, B2 => 
                           n21822, ZN => n7675);
   U23838 : OAI22_X1 port map( A1 => n27456, A2 => n27207, B1 => n27201, B2 => 
                           n21821, ZN => n7676);
   U23839 : OAI22_X1 port map( A1 => n27459, A2 => n27208, B1 => n27201, B2 => 
                           n21820, ZN => n7677);
   U23840 : OAI22_X1 port map( A1 => n27319, A2 => n27012, B1 => n27006, B2 => 
                           n21807, ZN => n6606);
   U23841 : OAI22_X1 port map( A1 => n27322, A2 => n27012, B1 => n27006, B2 => 
                           n21806, ZN => n6607);
   U23842 : OAI22_X1 port map( A1 => n27325, A2 => n27012, B1 => n27006, B2 => 
                           n21805, ZN => n6608);
   U23843 : OAI22_X1 port map( A1 => n27328, A2 => n27012, B1 => n27006, B2 => 
                           n21804, ZN => n6609);
   U23844 : OAI22_X1 port map( A1 => n27331, A2 => n27012, B1 => n27006, B2 => 
                           n21803, ZN => n6610);
   U23845 : OAI22_X1 port map( A1 => n27334, A2 => n27012, B1 => n27006, B2 => 
                           n21802, ZN => n6611);
   U23846 : OAI22_X1 port map( A1 => n27337, A2 => n27012, B1 => n27006, B2 => 
                           n21801, ZN => n6612);
   U23847 : OAI22_X1 port map( A1 => n27340, A2 => n27012, B1 => n27006, B2 => 
                           n21800, ZN => n6613);
   U23848 : OAI22_X1 port map( A1 => n27343, A2 => n27012, B1 => n27006, B2 => 
                           n21799, ZN => n6614);
   U23849 : OAI22_X1 port map( A1 => n27346, A2 => n27012, B1 => n27006, B2 => 
                           n21798, ZN => n6615);
   U23850 : OAI22_X1 port map( A1 => n27349, A2 => n27012, B1 => n27006, B2 => 
                           n21797, ZN => n6616);
   U23851 : OAI22_X1 port map( A1 => n27352, A2 => n27013, B1 => n27006, B2 => 
                           n21796, ZN => n6617);
   U23852 : OAI22_X1 port map( A1 => n27355, A2 => n27013, B1 => n27007, B2 => 
                           n21795, ZN => n6618);
   U23853 : OAI22_X1 port map( A1 => n27358, A2 => n27013, B1 => n27007, B2 => 
                           n21794, ZN => n6619);
   U23854 : OAI22_X1 port map( A1 => n27361, A2 => n27013, B1 => n27007, B2 => 
                           n21793, ZN => n6620);
   U23855 : OAI22_X1 port map( A1 => n27364, A2 => n27013, B1 => n27007, B2 => 
                           n21792, ZN => n6621);
   U23856 : OAI22_X1 port map( A1 => n27367, A2 => n27013, B1 => n27007, B2 => 
                           n21791, ZN => n6622);
   U23857 : OAI22_X1 port map( A1 => n27370, A2 => n27013, B1 => n27007, B2 => 
                           n21790, ZN => n6623);
   U23858 : OAI22_X1 port map( A1 => n27373, A2 => n27013, B1 => n27007, B2 => 
                           n21789, ZN => n6624);
   U23859 : OAI22_X1 port map( A1 => n27376, A2 => n27013, B1 => n27007, B2 => 
                           n21788, ZN => n6625);
   U23860 : OAI22_X1 port map( A1 => n27379, A2 => n27013, B1 => n27007, B2 => 
                           n21787, ZN => n6626);
   U23861 : OAI22_X1 port map( A1 => n27382, A2 => n27013, B1 => n27007, B2 => 
                           n21786, ZN => n6627);
   U23862 : OAI22_X1 port map( A1 => n27385, A2 => n27013, B1 => n27007, B2 => 
                           n21785, ZN => n6628);
   U23863 : OAI22_X1 port map( A1 => n27388, A2 => n27014, B1 => n27007, B2 => 
                           n21784, ZN => n6629);
   U23864 : OAI22_X1 port map( A1 => n27391, A2 => n27014, B1 => n27008, B2 => 
                           n21783, ZN => n6630);
   U23865 : OAI22_X1 port map( A1 => n27394, A2 => n27014, B1 => n27008, B2 => 
                           n21782, ZN => n6631);
   U23866 : OAI22_X1 port map( A1 => n27397, A2 => n27014, B1 => n27008, B2 => 
                           n21781, ZN => n6632);
   U23867 : OAI22_X1 port map( A1 => n27400, A2 => n27014, B1 => n27008, B2 => 
                           n21780, ZN => n6633);
   U23868 : OAI22_X1 port map( A1 => n27403, A2 => n27014, B1 => n27008, B2 => 
                           n21779, ZN => n6634);
   U23869 : OAI22_X1 port map( A1 => n27406, A2 => n27014, B1 => n27008, B2 => 
                           n21778, ZN => n6635);
   U23870 : OAI22_X1 port map( A1 => n27409, A2 => n27014, B1 => n27008, B2 => 
                           n21777, ZN => n6636);
   U23871 : OAI22_X1 port map( A1 => n27412, A2 => n27014, B1 => n27008, B2 => 
                           n21776, ZN => n6637);
   U23872 : OAI22_X1 port map( A1 => n27415, A2 => n27014, B1 => n27008, B2 => 
                           n21775, ZN => n6638);
   U23873 : OAI22_X1 port map( A1 => n27418, A2 => n27014, B1 => n27008, B2 => 
                           n21774, ZN => n6639);
   U23874 : OAI22_X1 port map( A1 => n27421, A2 => n27014, B1 => n27008, B2 => 
                           n21773, ZN => n6640);
   U23875 : OAI22_X1 port map( A1 => n27424, A2 => n27015, B1 => n27008, B2 => 
                           n21772, ZN => n6641);
   U23876 : OAI22_X1 port map( A1 => n27427, A2 => n27015, B1 => n27009, B2 => 
                           n21771, ZN => n6642);
   U23877 : OAI22_X1 port map( A1 => n27430, A2 => n27015, B1 => n27009, B2 => 
                           n21770, ZN => n6643);
   U23878 : OAI22_X1 port map( A1 => n27433, A2 => n27015, B1 => n27009, B2 => 
                           n21769, ZN => n6644);
   U23879 : OAI22_X1 port map( A1 => n27436, A2 => n27015, B1 => n27009, B2 => 
                           n21768, ZN => n6645);
   U23880 : OAI22_X1 port map( A1 => n27439, A2 => n27015, B1 => n27009, B2 => 
                           n21767, ZN => n6646);
   U23881 : OAI22_X1 port map( A1 => n27442, A2 => n27015, B1 => n27009, B2 => 
                           n21766, ZN => n6647);
   U23882 : OAI22_X1 port map( A1 => n27445, A2 => n27015, B1 => n27009, B2 => 
                           n21765, ZN => n6648);
   U23883 : OAI22_X1 port map( A1 => n27448, A2 => n27015, B1 => n27009, B2 => 
                           n21764, ZN => n6649);
   U23884 : OAI22_X1 port map( A1 => n27451, A2 => n27015, B1 => n27009, B2 => 
                           n21763, ZN => n6650);
   U23885 : OAI22_X1 port map( A1 => n27454, A2 => n27015, B1 => n27009, B2 => 
                           n21762, ZN => n6651);
   U23886 : OAI22_X1 port map( A1 => n27457, A2 => n27015, B1 => n27009, B2 => 
                           n21761, ZN => n6652);
   U23887 : OAI22_X1 port map( A1 => n27460, A2 => n27016, B1 => n27009, B2 => 
                           n21760, ZN => n6653);
   U23888 : OAI22_X1 port map( A1 => n27319, A2 => n27060, B1 => n27054, B2 => 
                           n21687, ZN => n6862);
   U23889 : OAI22_X1 port map( A1 => n27322, A2 => n27060, B1 => n27054, B2 => 
                           n21686, ZN => n6863);
   U23890 : OAI22_X1 port map( A1 => n27325, A2 => n27060, B1 => n27054, B2 => 
                           n21685, ZN => n6864);
   U23891 : OAI22_X1 port map( A1 => n27328, A2 => n27060, B1 => n27054, B2 => 
                           n21684, ZN => n6865);
   U23892 : OAI22_X1 port map( A1 => n27331, A2 => n27060, B1 => n27054, B2 => 
                           n21683, ZN => n6866);
   U23893 : OAI22_X1 port map( A1 => n27334, A2 => n27060, B1 => n27054, B2 => 
                           n21682, ZN => n6867);
   U23894 : OAI22_X1 port map( A1 => n27337, A2 => n27060, B1 => n27054, B2 => 
                           n21681, ZN => n6868);
   U23895 : OAI22_X1 port map( A1 => n27340, A2 => n27060, B1 => n27054, B2 => 
                           n21680, ZN => n6869);
   U23896 : OAI22_X1 port map( A1 => n27343, A2 => n27060, B1 => n27054, B2 => 
                           n21679, ZN => n6870);
   U23897 : OAI22_X1 port map( A1 => n27346, A2 => n27060, B1 => n27054, B2 => 
                           n21678, ZN => n6871);
   U23898 : OAI22_X1 port map( A1 => n27349, A2 => n27060, B1 => n27054, B2 => 
                           n21677, ZN => n6872);
   U23899 : OAI22_X1 port map( A1 => n27352, A2 => n27061, B1 => n27054, B2 => 
                           n21676, ZN => n6873);
   U23900 : OAI22_X1 port map( A1 => n27355, A2 => n27061, B1 => n27055, B2 => 
                           n21675, ZN => n6874);
   U23901 : OAI22_X1 port map( A1 => n27358, A2 => n27061, B1 => n27055, B2 => 
                           n21674, ZN => n6875);
   U23902 : OAI22_X1 port map( A1 => n27361, A2 => n27061, B1 => n27055, B2 => 
                           n21673, ZN => n6876);
   U23903 : OAI22_X1 port map( A1 => n27364, A2 => n27061, B1 => n27055, B2 => 
                           n21672, ZN => n6877);
   U23904 : OAI22_X1 port map( A1 => n27367, A2 => n27061, B1 => n27055, B2 => 
                           n21671, ZN => n6878);
   U23905 : OAI22_X1 port map( A1 => n27370, A2 => n27061, B1 => n27055, B2 => 
                           n21670, ZN => n6879);
   U23906 : OAI22_X1 port map( A1 => n27373, A2 => n27061, B1 => n27055, B2 => 
                           n21669, ZN => n6880);
   U23907 : OAI22_X1 port map( A1 => n27376, A2 => n27061, B1 => n27055, B2 => 
                           n21668, ZN => n6881);
   U23908 : OAI22_X1 port map( A1 => n27379, A2 => n27061, B1 => n27055, B2 => 
                           n21667, ZN => n6882);
   U23909 : OAI22_X1 port map( A1 => n27382, A2 => n27061, B1 => n27055, B2 => 
                           n21666, ZN => n6883);
   U23910 : OAI22_X1 port map( A1 => n27385, A2 => n27061, B1 => n27055, B2 => 
                           n21665, ZN => n6884);
   U23911 : OAI22_X1 port map( A1 => n27388, A2 => n27062, B1 => n27055, B2 => 
                           n21664, ZN => n6885);
   U23912 : OAI22_X1 port map( A1 => n27391, A2 => n27062, B1 => n27056, B2 => 
                           n21663, ZN => n6886);
   U23913 : OAI22_X1 port map( A1 => n27394, A2 => n27062, B1 => n27056, B2 => 
                           n21662, ZN => n6887);
   U23914 : OAI22_X1 port map( A1 => n27397, A2 => n27062, B1 => n27056, B2 => 
                           n21661, ZN => n6888);
   U23915 : OAI22_X1 port map( A1 => n27400, A2 => n27062, B1 => n27056, B2 => 
                           n21660, ZN => n6889);
   U23916 : OAI22_X1 port map( A1 => n27403, A2 => n27062, B1 => n27056, B2 => 
                           n21659, ZN => n6890);
   U23917 : OAI22_X1 port map( A1 => n27406, A2 => n27062, B1 => n27056, B2 => 
                           n21658, ZN => n6891);
   U23918 : OAI22_X1 port map( A1 => n27409, A2 => n27062, B1 => n27056, B2 => 
                           n21657, ZN => n6892);
   U23919 : OAI22_X1 port map( A1 => n27412, A2 => n27062, B1 => n27056, B2 => 
                           n21656, ZN => n6893);
   U23920 : OAI22_X1 port map( A1 => n27415, A2 => n27062, B1 => n27056, B2 => 
                           n21655, ZN => n6894);
   U23921 : OAI22_X1 port map( A1 => n27418, A2 => n27062, B1 => n27056, B2 => 
                           n21654, ZN => n6895);
   U23922 : OAI22_X1 port map( A1 => n27421, A2 => n27062, B1 => n27056, B2 => 
                           n21653, ZN => n6896);
   U23923 : OAI22_X1 port map( A1 => n27424, A2 => n27063, B1 => n27056, B2 => 
                           n21652, ZN => n6897);
   U23924 : OAI22_X1 port map( A1 => n27427, A2 => n27063, B1 => n27057, B2 => 
                           n21651, ZN => n6898);
   U23925 : OAI22_X1 port map( A1 => n27430, A2 => n27063, B1 => n27057, B2 => 
                           n21650, ZN => n6899);
   U23926 : OAI22_X1 port map( A1 => n27433, A2 => n27063, B1 => n27057, B2 => 
                           n21649, ZN => n6900);
   U23927 : OAI22_X1 port map( A1 => n27436, A2 => n27063, B1 => n27057, B2 => 
                           n21648, ZN => n6901);
   U23928 : OAI22_X1 port map( A1 => n27439, A2 => n27063, B1 => n27057, B2 => 
                           n21647, ZN => n6902);
   U23929 : OAI22_X1 port map( A1 => n27442, A2 => n27063, B1 => n27057, B2 => 
                           n21646, ZN => n6903);
   U23930 : OAI22_X1 port map( A1 => n27445, A2 => n27063, B1 => n27057, B2 => 
                           n21645, ZN => n6904);
   U23931 : OAI22_X1 port map( A1 => n27448, A2 => n27063, B1 => n27057, B2 => 
                           n21644, ZN => n6905);
   U23932 : OAI22_X1 port map( A1 => n27451, A2 => n27063, B1 => n27057, B2 => 
                           n21643, ZN => n6906);
   U23933 : OAI22_X1 port map( A1 => n27454, A2 => n27063, B1 => n27057, B2 => 
                           n21642, ZN => n6907);
   U23934 : OAI22_X1 port map( A1 => n27457, A2 => n27063, B1 => n27057, B2 => 
                           n21641, ZN => n6908);
   U23935 : OAI22_X1 port map( A1 => n27460, A2 => n27064, B1 => n27057, B2 => 
                           n21640, ZN => n6909);
   U23936 : OAI22_X1 port map( A1 => n27318, A2 => n27252, B1 => n27246, B2 => 
                           n21467, ZN => n7886);
   U23937 : OAI22_X1 port map( A1 => n27321, A2 => n27252, B1 => n27246, B2 => 
                           n21466, ZN => n7887);
   U23938 : OAI22_X1 port map( A1 => n27324, A2 => n27252, B1 => n27246, B2 => 
                           n21465, ZN => n7888);
   U23939 : OAI22_X1 port map( A1 => n27327, A2 => n27252, B1 => n27246, B2 => 
                           n21464, ZN => n7889);
   U23940 : OAI22_X1 port map( A1 => n27330, A2 => n27252, B1 => n27246, B2 => 
                           n21463, ZN => n7890);
   U23941 : OAI22_X1 port map( A1 => n27333, A2 => n27252, B1 => n27246, B2 => 
                           n21462, ZN => n7891);
   U23942 : OAI22_X1 port map( A1 => n27336, A2 => n27252, B1 => n27246, B2 => 
                           n21461, ZN => n7892);
   U23943 : OAI22_X1 port map( A1 => n27339, A2 => n27252, B1 => n27246, B2 => 
                           n21460, ZN => n7893);
   U23944 : OAI22_X1 port map( A1 => n27342, A2 => n27252, B1 => n27246, B2 => 
                           n21459, ZN => n7894);
   U23945 : OAI22_X1 port map( A1 => n27345, A2 => n27252, B1 => n27246, B2 => 
                           n21458, ZN => n7895);
   U23946 : OAI22_X1 port map( A1 => n27348, A2 => n27252, B1 => n27246, B2 => 
                           n21457, ZN => n7896);
   U23947 : OAI22_X1 port map( A1 => n27351, A2 => n27253, B1 => n27246, B2 => 
                           n21456, ZN => n7897);
   U23948 : OAI22_X1 port map( A1 => n27354, A2 => n27253, B1 => n27247, B2 => 
                           n21455, ZN => n7898);
   U23949 : OAI22_X1 port map( A1 => n27357, A2 => n27253, B1 => n27247, B2 => 
                           n21454, ZN => n7899);
   U23950 : OAI22_X1 port map( A1 => n27360, A2 => n27253, B1 => n27247, B2 => 
                           n21453, ZN => n7900);
   U23951 : OAI22_X1 port map( A1 => n27363, A2 => n27253, B1 => n27247, B2 => 
                           n21452, ZN => n7901);
   U23952 : OAI22_X1 port map( A1 => n27366, A2 => n27253, B1 => n27247, B2 => 
                           n21451, ZN => n7902);
   U23953 : OAI22_X1 port map( A1 => n27369, A2 => n27253, B1 => n27247, B2 => 
                           n21450, ZN => n7903);
   U23954 : OAI22_X1 port map( A1 => n27372, A2 => n27253, B1 => n27247, B2 => 
                           n21449, ZN => n7904);
   U23955 : OAI22_X1 port map( A1 => n27375, A2 => n27253, B1 => n27247, B2 => 
                           n21448, ZN => n7905);
   U23956 : OAI22_X1 port map( A1 => n27378, A2 => n27253, B1 => n27247, B2 => 
                           n21447, ZN => n7906);
   U23957 : OAI22_X1 port map( A1 => n27381, A2 => n27253, B1 => n27247, B2 => 
                           n21446, ZN => n7907);
   U23958 : OAI22_X1 port map( A1 => n27384, A2 => n27253, B1 => n27247, B2 => 
                           n21445, ZN => n7908);
   U23959 : OAI22_X1 port map( A1 => n27387, A2 => n27254, B1 => n27247, B2 => 
                           n21444, ZN => n7909);
   U23960 : OAI22_X1 port map( A1 => n27390, A2 => n27254, B1 => n27248, B2 => 
                           n21443, ZN => n7910);
   U23961 : OAI22_X1 port map( A1 => n27393, A2 => n27254, B1 => n27248, B2 => 
                           n21442, ZN => n7911);
   U23962 : OAI22_X1 port map( A1 => n27396, A2 => n27254, B1 => n27248, B2 => 
                           n21441, ZN => n7912);
   U23963 : OAI22_X1 port map( A1 => n27399, A2 => n27254, B1 => n27248, B2 => 
                           n21440, ZN => n7913);
   U23964 : OAI22_X1 port map( A1 => n27402, A2 => n27254, B1 => n27248, B2 => 
                           n21439, ZN => n7914);
   U23965 : OAI22_X1 port map( A1 => n27405, A2 => n27254, B1 => n27248, B2 => 
                           n21438, ZN => n7915);
   U23966 : OAI22_X1 port map( A1 => n27408, A2 => n27254, B1 => n27248, B2 => 
                           n21437, ZN => n7916);
   U23967 : OAI22_X1 port map( A1 => n27411, A2 => n27254, B1 => n27248, B2 => 
                           n21436, ZN => n7917);
   U23968 : OAI22_X1 port map( A1 => n27414, A2 => n27254, B1 => n27248, B2 => 
                           n21435, ZN => n7918);
   U23969 : OAI22_X1 port map( A1 => n27417, A2 => n27254, B1 => n27248, B2 => 
                           n21434, ZN => n7919);
   U23970 : OAI22_X1 port map( A1 => n27420, A2 => n27254, B1 => n27248, B2 => 
                           n21433, ZN => n7920);
   U23971 : OAI22_X1 port map( A1 => n27423, A2 => n27255, B1 => n27248, B2 => 
                           n21432, ZN => n7921);
   U23972 : OAI22_X1 port map( A1 => n27426, A2 => n27255, B1 => n27249, B2 => 
                           n21431, ZN => n7922);
   U23973 : OAI22_X1 port map( A1 => n27429, A2 => n27255, B1 => n27249, B2 => 
                           n21430, ZN => n7923);
   U23974 : OAI22_X1 port map( A1 => n27432, A2 => n27255, B1 => n27249, B2 => 
                           n21429, ZN => n7924);
   U23975 : OAI22_X1 port map( A1 => n27435, A2 => n27255, B1 => n27249, B2 => 
                           n21428, ZN => n7925);
   U23976 : OAI22_X1 port map( A1 => n27438, A2 => n27255, B1 => n27249, B2 => 
                           n21427, ZN => n7926);
   U23977 : OAI22_X1 port map( A1 => n27441, A2 => n27255, B1 => n27249, B2 => 
                           n21426, ZN => n7927);
   U23978 : OAI22_X1 port map( A1 => n27444, A2 => n27255, B1 => n27249, B2 => 
                           n21425, ZN => n7928);
   U23979 : OAI22_X1 port map( A1 => n27447, A2 => n27255, B1 => n27249, B2 => 
                           n21424, ZN => n7929);
   U23980 : OAI22_X1 port map( A1 => n27450, A2 => n27255, B1 => n27249, B2 => 
                           n21423, ZN => n7930);
   U23981 : OAI22_X1 port map( A1 => n27453, A2 => n27255, B1 => n27249, B2 => 
                           n21422, ZN => n7931);
   U23982 : OAI22_X1 port map( A1 => n27456, A2 => n27255, B1 => n27249, B2 => 
                           n21421, ZN => n7932);
   U23983 : OAI22_X1 port map( A1 => n27459, A2 => n27256, B1 => n27249, B2 => 
                           n21420, ZN => n7933);
   U23984 : OAI22_X1 port map( A1 => n27319, A2 => n27084, B1 => n27078, B2 => 
                           n21287, ZN => n6990);
   U23985 : OAI22_X1 port map( A1 => n27322, A2 => n27084, B1 => n27078, B2 => 
                           n21286, ZN => n6991);
   U23986 : OAI22_X1 port map( A1 => n27325, A2 => n27084, B1 => n27078, B2 => 
                           n21285, ZN => n6992);
   U23987 : OAI22_X1 port map( A1 => n27328, A2 => n27084, B1 => n27078, B2 => 
                           n21284, ZN => n6993);
   U23988 : OAI22_X1 port map( A1 => n27331, A2 => n27084, B1 => n27078, B2 => 
                           n21283, ZN => n6994);
   U23989 : OAI22_X1 port map( A1 => n27334, A2 => n27084, B1 => n27078, B2 => 
                           n21282, ZN => n6995);
   U23990 : OAI22_X1 port map( A1 => n27337, A2 => n27084, B1 => n27078, B2 => 
                           n21281, ZN => n6996);
   U23991 : OAI22_X1 port map( A1 => n27340, A2 => n27084, B1 => n27078, B2 => 
                           n21280, ZN => n6997);
   U23992 : OAI22_X1 port map( A1 => n27343, A2 => n27084, B1 => n27078, B2 => 
                           n21279, ZN => n6998);
   U23993 : OAI22_X1 port map( A1 => n27346, A2 => n27084, B1 => n27078, B2 => 
                           n21278, ZN => n6999);
   U23994 : OAI22_X1 port map( A1 => n27349, A2 => n27084, B1 => n27078, B2 => 
                           n21277, ZN => n7000);
   U23995 : OAI22_X1 port map( A1 => n27352, A2 => n27085, B1 => n27078, B2 => 
                           n21276, ZN => n7001);
   U23996 : OAI22_X1 port map( A1 => n27355, A2 => n27085, B1 => n27079, B2 => 
                           n21275, ZN => n7002);
   U23997 : OAI22_X1 port map( A1 => n27358, A2 => n27085, B1 => n27079, B2 => 
                           n21274, ZN => n7003);
   U23998 : OAI22_X1 port map( A1 => n27361, A2 => n27085, B1 => n27079, B2 => 
                           n21273, ZN => n7004);
   U23999 : OAI22_X1 port map( A1 => n27364, A2 => n27085, B1 => n27079, B2 => 
                           n21272, ZN => n7005);
   U24000 : OAI22_X1 port map( A1 => n27367, A2 => n27085, B1 => n27079, B2 => 
                           n21271, ZN => n7006);
   U24001 : OAI22_X1 port map( A1 => n27370, A2 => n27085, B1 => n27079, B2 => 
                           n21270, ZN => n7007);
   U24002 : OAI22_X1 port map( A1 => n27373, A2 => n27085, B1 => n27079, B2 => 
                           n21269, ZN => n7008);
   U24003 : OAI22_X1 port map( A1 => n27376, A2 => n27085, B1 => n27079, B2 => 
                           n21268, ZN => n7009);
   U24004 : OAI22_X1 port map( A1 => n27379, A2 => n27085, B1 => n27079, B2 => 
                           n21267, ZN => n7010);
   U24005 : OAI22_X1 port map( A1 => n27382, A2 => n27085, B1 => n27079, B2 => 
                           n21266, ZN => n7011);
   U24006 : OAI22_X1 port map( A1 => n27385, A2 => n27085, B1 => n27079, B2 => 
                           n21265, ZN => n7012);
   U24007 : OAI22_X1 port map( A1 => n27388, A2 => n27086, B1 => n27079, B2 => 
                           n21264, ZN => n7013);
   U24008 : OAI22_X1 port map( A1 => n27391, A2 => n27086, B1 => n27080, B2 => 
                           n21263, ZN => n7014);
   U24009 : OAI22_X1 port map( A1 => n27394, A2 => n27086, B1 => n27080, B2 => 
                           n21262, ZN => n7015);
   U24010 : OAI22_X1 port map( A1 => n27397, A2 => n27086, B1 => n27080, B2 => 
                           n21261, ZN => n7016);
   U24011 : OAI22_X1 port map( A1 => n27400, A2 => n27086, B1 => n27080, B2 => 
                           n21260, ZN => n7017);
   U24012 : OAI22_X1 port map( A1 => n27403, A2 => n27086, B1 => n27080, B2 => 
                           n21259, ZN => n7018);
   U24013 : OAI22_X1 port map( A1 => n27406, A2 => n27086, B1 => n27080, B2 => 
                           n21258, ZN => n7019);
   U24014 : OAI22_X1 port map( A1 => n27409, A2 => n27086, B1 => n27080, B2 => 
                           n21257, ZN => n7020);
   U24015 : OAI22_X1 port map( A1 => n27412, A2 => n27086, B1 => n27080, B2 => 
                           n21256, ZN => n7021);
   U24016 : OAI22_X1 port map( A1 => n27415, A2 => n27086, B1 => n27080, B2 => 
                           n21255, ZN => n7022);
   U24017 : OAI22_X1 port map( A1 => n27418, A2 => n27086, B1 => n27080, B2 => 
                           n21254, ZN => n7023);
   U24018 : OAI22_X1 port map( A1 => n27421, A2 => n27086, B1 => n27080, B2 => 
                           n21253, ZN => n7024);
   U24019 : OAI22_X1 port map( A1 => n27424, A2 => n27087, B1 => n27080, B2 => 
                           n21252, ZN => n7025);
   U24020 : OAI22_X1 port map( A1 => n27427, A2 => n27087, B1 => n27081, B2 => 
                           n21251, ZN => n7026);
   U24021 : OAI22_X1 port map( A1 => n27430, A2 => n27087, B1 => n27081, B2 => 
                           n21250, ZN => n7027);
   U24022 : OAI22_X1 port map( A1 => n27433, A2 => n27087, B1 => n27081, B2 => 
                           n21249, ZN => n7028);
   U24023 : OAI22_X1 port map( A1 => n27436, A2 => n27087, B1 => n27081, B2 => 
                           n21248, ZN => n7029);
   U24024 : OAI22_X1 port map( A1 => n27439, A2 => n27087, B1 => n27081, B2 => 
                           n21247, ZN => n7030);
   U24025 : OAI22_X1 port map( A1 => n27442, A2 => n27087, B1 => n27081, B2 => 
                           n21246, ZN => n7031);
   U24026 : OAI22_X1 port map( A1 => n27445, A2 => n27087, B1 => n27081, B2 => 
                           n21245, ZN => n7032);
   U24027 : OAI22_X1 port map( A1 => n27448, A2 => n27087, B1 => n27081, B2 => 
                           n21244, ZN => n7033);
   U24028 : OAI22_X1 port map( A1 => n27451, A2 => n27087, B1 => n27081, B2 => 
                           n21243, ZN => n7034);
   U24029 : OAI22_X1 port map( A1 => n27454, A2 => n27087, B1 => n27081, B2 => 
                           n21242, ZN => n7035);
   U24030 : OAI22_X1 port map( A1 => n27457, A2 => n27087, B1 => n27081, B2 => 
                           n21241, ZN => n7036);
   U24031 : OAI22_X1 port map( A1 => n27460, A2 => n27088, B1 => n27081, B2 => 
                           n21240, ZN => n7037);
   U24032 : OAI22_X1 port map( A1 => n27320, A2 => n26904, B1 => n26898, B2 => 
                           n20950, ZN => n6030);
   U24033 : OAI22_X1 port map( A1 => n27323, A2 => n26904, B1 => n26898, B2 => 
                           n20949, ZN => n6031);
   U24034 : OAI22_X1 port map( A1 => n27326, A2 => n26904, B1 => n26898, B2 => 
                           n20948, ZN => n6032);
   U24035 : OAI22_X1 port map( A1 => n27329, A2 => n26904, B1 => n26898, B2 => 
                           n20947, ZN => n6033);
   U24036 : OAI22_X1 port map( A1 => n27332, A2 => n26904, B1 => n26898, B2 => 
                           n20946, ZN => n6034);
   U24037 : OAI22_X1 port map( A1 => n27335, A2 => n26904, B1 => n26898, B2 => 
                           n20945, ZN => n6035);
   U24038 : OAI22_X1 port map( A1 => n27338, A2 => n26904, B1 => n26898, B2 => 
                           n20944, ZN => n6036);
   U24039 : OAI22_X1 port map( A1 => n27341, A2 => n26904, B1 => n26898, B2 => 
                           n20943, ZN => n6037);
   U24040 : OAI22_X1 port map( A1 => n27344, A2 => n26904, B1 => n26898, B2 => 
                           n20942, ZN => n6038);
   U24041 : OAI22_X1 port map( A1 => n27347, A2 => n26904, B1 => n26898, B2 => 
                           n20941, ZN => n6039);
   U24042 : OAI22_X1 port map( A1 => n27350, A2 => n26904, B1 => n26898, B2 => 
                           n20940, ZN => n6040);
   U24043 : OAI22_X1 port map( A1 => n27353, A2 => n26905, B1 => n26898, B2 => 
                           n20939, ZN => n6041);
   U24044 : OAI22_X1 port map( A1 => n27356, A2 => n26905, B1 => n26899, B2 => 
                           n20938, ZN => n6042);
   U24045 : OAI22_X1 port map( A1 => n27359, A2 => n26905, B1 => n26899, B2 => 
                           n20937, ZN => n6043);
   U24046 : OAI22_X1 port map( A1 => n27362, A2 => n26905, B1 => n26899, B2 => 
                           n20936, ZN => n6044);
   U24047 : OAI22_X1 port map( A1 => n27365, A2 => n26905, B1 => n26899, B2 => 
                           n20935, ZN => n6045);
   U24048 : OAI22_X1 port map( A1 => n27368, A2 => n26905, B1 => n26899, B2 => 
                           n20934, ZN => n6046);
   U24049 : OAI22_X1 port map( A1 => n27371, A2 => n26905, B1 => n26899, B2 => 
                           n20933, ZN => n6047);
   U24050 : OAI22_X1 port map( A1 => n27374, A2 => n26905, B1 => n26899, B2 => 
                           n20932, ZN => n6048);
   U24051 : OAI22_X1 port map( A1 => n27377, A2 => n26905, B1 => n26899, B2 => 
                           n20931, ZN => n6049);
   U24052 : OAI22_X1 port map( A1 => n27380, A2 => n26905, B1 => n26899, B2 => 
                           n20930, ZN => n6050);
   U24053 : OAI22_X1 port map( A1 => n27383, A2 => n26905, B1 => n26899, B2 => 
                           n20929, ZN => n6051);
   U24054 : OAI22_X1 port map( A1 => n27386, A2 => n26905, B1 => n26899, B2 => 
                           n20928, ZN => n6052);
   U24055 : OAI22_X1 port map( A1 => n27389, A2 => n26906, B1 => n26899, B2 => 
                           n20927, ZN => n6053);
   U24056 : OAI22_X1 port map( A1 => n27392, A2 => n26906, B1 => n26900, B2 => 
                           n20926, ZN => n6054);
   U24057 : OAI22_X1 port map( A1 => n27395, A2 => n26906, B1 => n26900, B2 => 
                           n20925, ZN => n6055);
   U24058 : OAI22_X1 port map( A1 => n27398, A2 => n26906, B1 => n26900, B2 => 
                           n20924, ZN => n6056);
   U24059 : OAI22_X1 port map( A1 => n27401, A2 => n26906, B1 => n26900, B2 => 
                           n20923, ZN => n6057);
   U24060 : OAI22_X1 port map( A1 => n27404, A2 => n26906, B1 => n26900, B2 => 
                           n20922, ZN => n6058);
   U24061 : OAI22_X1 port map( A1 => n27407, A2 => n26906, B1 => n26900, B2 => 
                           n20921, ZN => n6059);
   U24062 : OAI22_X1 port map( A1 => n27410, A2 => n26906, B1 => n26900, B2 => 
                           n20920, ZN => n6060);
   U24063 : OAI22_X1 port map( A1 => n27413, A2 => n26906, B1 => n26900, B2 => 
                           n20919, ZN => n6061);
   U24064 : OAI22_X1 port map( A1 => n27416, A2 => n26906, B1 => n26900, B2 => 
                           n20918, ZN => n6062);
   U24065 : OAI22_X1 port map( A1 => n27419, A2 => n26906, B1 => n26900, B2 => 
                           n20917, ZN => n6063);
   U24066 : OAI22_X1 port map( A1 => n27422, A2 => n26906, B1 => n26900, B2 => 
                           n20916, ZN => n6064);
   U24067 : OAI22_X1 port map( A1 => n27425, A2 => n26907, B1 => n26900, B2 => 
                           n20915, ZN => n6065);
   U24068 : OAI22_X1 port map( A1 => n27428, A2 => n26907, B1 => n26901, B2 => 
                           n20914, ZN => n6066);
   U24069 : OAI22_X1 port map( A1 => n27431, A2 => n26907, B1 => n26901, B2 => 
                           n20913, ZN => n6067);
   U24070 : OAI22_X1 port map( A1 => n27434, A2 => n26907, B1 => n26901, B2 => 
                           n20912, ZN => n6068);
   U24071 : OAI22_X1 port map( A1 => n27437, A2 => n26907, B1 => n26901, B2 => 
                           n20911, ZN => n6069);
   U24072 : OAI22_X1 port map( A1 => n27440, A2 => n26907, B1 => n26901, B2 => 
                           n20910, ZN => n6070);
   U24073 : OAI22_X1 port map( A1 => n27443, A2 => n26907, B1 => n26901, B2 => 
                           n20909, ZN => n6071);
   U24074 : OAI22_X1 port map( A1 => n27446, A2 => n26907, B1 => n26901, B2 => 
                           n20908, ZN => n6072);
   U24075 : OAI22_X1 port map( A1 => n27449, A2 => n26907, B1 => n26901, B2 => 
                           n20907, ZN => n6073);
   U24076 : OAI22_X1 port map( A1 => n27452, A2 => n26907, B1 => n26901, B2 => 
                           n20906, ZN => n6074);
   U24077 : OAI22_X1 port map( A1 => n27455, A2 => n26907, B1 => n26901, B2 => 
                           n20905, ZN => n6075);
   U24078 : OAI22_X1 port map( A1 => n27458, A2 => n26907, B1 => n26901, B2 => 
                           n20904, ZN => n6076);
   U24079 : OAI22_X1 port map( A1 => n27461, A2 => n26908, B1 => n26901, B2 => 
                           n20903, ZN => n6077);
   U24080 : OAI22_X1 port map( A1 => n27320, A2 => n26916, B1 => n26910, B2 => 
                           n20886, ZN => n6094);
   U24081 : OAI22_X1 port map( A1 => n27323, A2 => n26916, B1 => n26910, B2 => 
                           n20885, ZN => n6095);
   U24082 : OAI22_X1 port map( A1 => n27326, A2 => n26916, B1 => n26910, B2 => 
                           n20884, ZN => n6096);
   U24083 : OAI22_X1 port map( A1 => n27329, A2 => n26916, B1 => n26910, B2 => 
                           n20883, ZN => n6097);
   U24084 : OAI22_X1 port map( A1 => n27332, A2 => n26916, B1 => n26910, B2 => 
                           n20882, ZN => n6098);
   U24085 : OAI22_X1 port map( A1 => n27335, A2 => n26916, B1 => n26910, B2 => 
                           n20881, ZN => n6099);
   U24086 : OAI22_X1 port map( A1 => n27338, A2 => n26916, B1 => n26910, B2 => 
                           n20880, ZN => n6100);
   U24087 : OAI22_X1 port map( A1 => n27341, A2 => n26916, B1 => n26910, B2 => 
                           n20879, ZN => n6101);
   U24088 : OAI22_X1 port map( A1 => n27344, A2 => n26916, B1 => n26910, B2 => 
                           n20878, ZN => n6102);
   U24089 : OAI22_X1 port map( A1 => n27347, A2 => n26916, B1 => n26910, B2 => 
                           n20877, ZN => n6103);
   U24090 : OAI22_X1 port map( A1 => n27350, A2 => n26916, B1 => n26910, B2 => 
                           n20876, ZN => n6104);
   U24091 : OAI22_X1 port map( A1 => n27353, A2 => n26917, B1 => n26910, B2 => 
                           n20875, ZN => n6105);
   U24092 : OAI22_X1 port map( A1 => n27356, A2 => n26917, B1 => n26911, B2 => 
                           n20874, ZN => n6106);
   U24093 : OAI22_X1 port map( A1 => n27359, A2 => n26917, B1 => n26911, B2 => 
                           n20873, ZN => n6107);
   U24094 : OAI22_X1 port map( A1 => n27362, A2 => n26917, B1 => n26911, B2 => 
                           n20872, ZN => n6108);
   U24095 : OAI22_X1 port map( A1 => n27365, A2 => n26917, B1 => n26911, B2 => 
                           n20871, ZN => n6109);
   U24096 : OAI22_X1 port map( A1 => n27368, A2 => n26917, B1 => n26911, B2 => 
                           n20870, ZN => n6110);
   U24097 : OAI22_X1 port map( A1 => n27371, A2 => n26917, B1 => n26911, B2 => 
                           n20869, ZN => n6111);
   U24098 : OAI22_X1 port map( A1 => n27374, A2 => n26917, B1 => n26911, B2 => 
                           n20868, ZN => n6112);
   U24099 : OAI22_X1 port map( A1 => n27377, A2 => n26917, B1 => n26911, B2 => 
                           n20867, ZN => n6113);
   U24100 : OAI22_X1 port map( A1 => n27380, A2 => n26917, B1 => n26911, B2 => 
                           n20866, ZN => n6114);
   U24101 : OAI22_X1 port map( A1 => n27383, A2 => n26917, B1 => n26911, B2 => 
                           n20865, ZN => n6115);
   U24102 : OAI22_X1 port map( A1 => n27386, A2 => n26917, B1 => n26911, B2 => 
                           n20864, ZN => n6116);
   U24103 : OAI22_X1 port map( A1 => n27389, A2 => n26918, B1 => n26911, B2 => 
                           n20863, ZN => n6117);
   U24104 : OAI22_X1 port map( A1 => n27392, A2 => n26918, B1 => n26912, B2 => 
                           n20862, ZN => n6118);
   U24105 : OAI22_X1 port map( A1 => n27395, A2 => n26918, B1 => n26912, B2 => 
                           n20861, ZN => n6119);
   U24106 : OAI22_X1 port map( A1 => n27398, A2 => n26918, B1 => n26912, B2 => 
                           n20860, ZN => n6120);
   U24107 : OAI22_X1 port map( A1 => n27401, A2 => n26918, B1 => n26912, B2 => 
                           n20859, ZN => n6121);
   U24108 : OAI22_X1 port map( A1 => n27404, A2 => n26918, B1 => n26912, B2 => 
                           n20858, ZN => n6122);
   U24109 : OAI22_X1 port map( A1 => n27407, A2 => n26918, B1 => n26912, B2 => 
                           n20857, ZN => n6123);
   U24110 : OAI22_X1 port map( A1 => n27410, A2 => n26918, B1 => n26912, B2 => 
                           n20856, ZN => n6124);
   U24111 : OAI22_X1 port map( A1 => n27413, A2 => n26918, B1 => n26912, B2 => 
                           n20855, ZN => n6125);
   U24112 : OAI22_X1 port map( A1 => n27416, A2 => n26918, B1 => n26912, B2 => 
                           n20854, ZN => n6126);
   U24113 : OAI22_X1 port map( A1 => n27419, A2 => n26918, B1 => n26912, B2 => 
                           n20853, ZN => n6127);
   U24114 : OAI22_X1 port map( A1 => n27422, A2 => n26918, B1 => n26912, B2 => 
                           n20852, ZN => n6128);
   U24115 : OAI22_X1 port map( A1 => n27425, A2 => n26919, B1 => n26912, B2 => 
                           n20851, ZN => n6129);
   U24116 : OAI22_X1 port map( A1 => n27428, A2 => n26919, B1 => n26913, B2 => 
                           n20850, ZN => n6130);
   U24117 : OAI22_X1 port map( A1 => n27431, A2 => n26919, B1 => n26913, B2 => 
                           n20849, ZN => n6131);
   U24118 : OAI22_X1 port map( A1 => n27434, A2 => n26919, B1 => n26913, B2 => 
                           n20848, ZN => n6132);
   U24119 : OAI22_X1 port map( A1 => n27437, A2 => n26919, B1 => n26913, B2 => 
                           n20847, ZN => n6133);
   U24120 : OAI22_X1 port map( A1 => n27440, A2 => n26919, B1 => n26913, B2 => 
                           n20846, ZN => n6134);
   U24121 : OAI22_X1 port map( A1 => n27443, A2 => n26919, B1 => n26913, B2 => 
                           n20845, ZN => n6135);
   U24122 : OAI22_X1 port map( A1 => n27446, A2 => n26919, B1 => n26913, B2 => 
                           n20844, ZN => n6136);
   U24123 : OAI22_X1 port map( A1 => n27449, A2 => n26919, B1 => n26913, B2 => 
                           n20843, ZN => n6137);
   U24124 : OAI22_X1 port map( A1 => n27452, A2 => n26919, B1 => n26913, B2 => 
                           n20842, ZN => n6138);
   U24125 : OAI22_X1 port map( A1 => n27455, A2 => n26919, B1 => n26913, B2 => 
                           n20841, ZN => n6139);
   U24126 : OAI22_X1 port map( A1 => n27458, A2 => n26919, B1 => n26913, B2 => 
                           n20840, ZN => n6140);
   U24127 : OAI22_X1 port map( A1 => n27461, A2 => n26920, B1 => n26913, B2 => 
                           n20839, ZN => n6141);
   U24128 : OAI22_X1 port map( A1 => n27464, A2 => n26956, B1 => n26950, B2 => 
                           n22507, ZN => n6334);
   U24129 : OAI22_X1 port map( A1 => n27467, A2 => n26956, B1 => n26950, B2 => 
                           n22506, ZN => n6335);
   U24130 : OAI22_X1 port map( A1 => n27470, A2 => n26956, B1 => n26950, B2 => 
                           n22505, ZN => n6336);
   U24131 : OAI22_X1 port map( A1 => n27473, A2 => n26956, B1 => n26950, B2 => 
                           n22504, ZN => n6337);
   U24132 : OAI22_X1 port map( A1 => n27462, A2 => n27160, B1 => n27154, B2 => 
                           n22255, ZN => n7422);
   U24133 : OAI22_X1 port map( A1 => n27465, A2 => n27160, B1 => n27154, B2 => 
                           n22254, ZN => n7423);
   U24134 : OAI22_X1 port map( A1 => n27468, A2 => n27160, B1 => n27154, B2 => 
                           n22253, ZN => n7424);
   U24135 : OAI22_X1 port map( A1 => n27471, A2 => n27160, B1 => n27154, B2 => 
                           n22252, ZN => n7425);
   U24136 : OAI22_X1 port map( A1 => n27464, A2 => n26932, B1 => n26926, B2 => 
                           n22247, ZN => n6206);
   U24137 : OAI22_X1 port map( A1 => n27467, A2 => n26932, B1 => n26926, B2 => 
                           n22246, ZN => n6207);
   U24138 : OAI22_X1 port map( A1 => n27470, A2 => n26932, B1 => n26926, B2 => 
                           n22245, ZN => n6208);
   U24139 : OAI22_X1 port map( A1 => n27473, A2 => n26932, B1 => n26926, B2 => 
                           n22244, ZN => n6209);
   U24140 : OAI22_X1 port map( A1 => n27464, A2 => n26944, B1 => n26938, B2 => 
                           n22183, ZN => n6270);
   U24141 : OAI22_X1 port map( A1 => n27467, A2 => n26944, B1 => n26938, B2 => 
                           n22182, ZN => n6271);
   U24142 : OAI22_X1 port map( A1 => n27470, A2 => n26944, B1 => n26938, B2 => 
                           n22181, ZN => n6272);
   U24143 : OAI22_X1 port map( A1 => n27473, A2 => n26944, B1 => n26938, B2 => 
                           n22180, ZN => n6273);
   U24144 : OAI22_X1 port map( A1 => n27281, A2 => n27462, B1 => n27274, B2 => 
                           n21519, ZN => n8062);
   U24145 : OAI22_X1 port map( A1 => n27281, A2 => n27465, B1 => n27274, B2 => 
                           n21518, ZN => n8063);
   U24146 : OAI22_X1 port map( A1 => n27281, A2 => n27468, B1 => n27274, B2 => 
                           n21517, ZN => n8064);
   U24147 : OAI22_X1 port map( A1 => n27281, A2 => n27471, B1 => n27274, B2 => 
                           n21516, ZN => n8065);
   U24148 : OAI22_X1 port map( A1 => n27462, A2 => n27268, B1 => n27262, B2 => 
                           n21515, ZN => n7998);
   U24149 : OAI22_X1 port map( A1 => n27465, A2 => n27268, B1 => n27262, B2 => 
                           n21514, ZN => n7999);
   U24150 : OAI22_X1 port map( A1 => n27468, A2 => n27268, B1 => n27262, B2 => 
                           n21513, ZN => n8000);
   U24151 : OAI22_X1 port map( A1 => n27471, A2 => n27268, B1 => n27262, B2 => 
                           n21512, ZN => n8001);
   U24152 : OAI22_X1 port map( A1 => n27462, A2 => n27232, B1 => n27226, B2 => 
                           n21503, ZN => n7806);
   U24153 : OAI22_X1 port map( A1 => n27465, A2 => n27232, B1 => n27226, B2 => 
                           n21502, ZN => n7807);
   U24154 : OAI22_X1 port map( A1 => n27468, A2 => n27232, B1 => n27226, B2 => 
                           n21501, ZN => n7808);
   U24155 : OAI22_X1 port map( A1 => n27471, A2 => n27232, B1 => n27226, B2 => 
                           n21500, ZN => n7809);
   U24156 : OAI22_X1 port map( A1 => n27462, A2 => n27208, B1 => n27202, B2 => 
                           n21499, ZN => n7678);
   U24157 : OAI22_X1 port map( A1 => n27465, A2 => n27208, B1 => n27202, B2 => 
                           n21498, ZN => n7679);
   U24158 : OAI22_X1 port map( A1 => n27468, A2 => n27208, B1 => n27202, B2 => 
                           n21497, ZN => n7680);
   U24159 : OAI22_X1 port map( A1 => n27471, A2 => n27208, B1 => n27202, B2 => 
                           n21496, ZN => n7681);
   U24160 : OAI22_X1 port map( A1 => n27463, A2 => n27016, B1 => n27010, B2 => 
                           n21495, ZN => n6654);
   U24161 : OAI22_X1 port map( A1 => n27466, A2 => n27016, B1 => n27010, B2 => 
                           n21494, ZN => n6655);
   U24162 : OAI22_X1 port map( A1 => n27469, A2 => n27016, B1 => n27010, B2 => 
                           n21493, ZN => n6656);
   U24163 : OAI22_X1 port map( A1 => n27472, A2 => n27016, B1 => n27010, B2 => 
                           n21492, ZN => n6657);
   U24164 : OAI22_X1 port map( A1 => n27463, A2 => n27064, B1 => n27058, B2 => 
                           n21487, ZN => n6910);
   U24165 : OAI22_X1 port map( A1 => n27466, A2 => n27064, B1 => n27058, B2 => 
                           n21486, ZN => n6911);
   U24166 : OAI22_X1 port map( A1 => n27469, A2 => n27064, B1 => n27058, B2 => 
                           n21485, ZN => n6912);
   U24167 : OAI22_X1 port map( A1 => n27472, A2 => n27064, B1 => n27058, B2 => 
                           n21484, ZN => n6913);
   U24168 : OAI22_X1 port map( A1 => n27462, A2 => n27256, B1 => n27250, B2 => 
                           n21175, ZN => n7934);
   U24169 : OAI22_X1 port map( A1 => n27465, A2 => n27256, B1 => n27250, B2 => 
                           n21174, ZN => n7935);
   U24170 : OAI22_X1 port map( A1 => n27468, A2 => n27256, B1 => n27250, B2 => 
                           n21173, ZN => n7936);
   U24171 : OAI22_X1 port map( A1 => n27471, A2 => n27256, B1 => n27250, B2 => 
                           n21172, ZN => n7937);
   U24172 : OAI22_X1 port map( A1 => n27463, A2 => n27088, B1 => n27082, B2 => 
                           n21163, ZN => n7038);
   U24173 : OAI22_X1 port map( A1 => n27466, A2 => n27088, B1 => n27082, B2 => 
                           n21162, ZN => n7039);
   U24174 : OAI22_X1 port map( A1 => n27469, A2 => n27088, B1 => n27082, B2 => 
                           n21161, ZN => n7040);
   U24175 : OAI22_X1 port map( A1 => n27472, A2 => n27088, B1 => n27082, B2 => 
                           n21160, ZN => n7041);
   U24176 : OAI22_X1 port map( A1 => n27464, A2 => n26908, B1 => n26902, B2 => 
                           n20902, ZN => n6078);
   U24177 : OAI22_X1 port map( A1 => n27467, A2 => n26908, B1 => n26902, B2 => 
                           n20901, ZN => n6079);
   U24178 : OAI22_X1 port map( A1 => n27470, A2 => n26908, B1 => n26902, B2 => 
                           n20900, ZN => n6080);
   U24179 : OAI22_X1 port map( A1 => n27473, A2 => n26908, B1 => n26902, B2 => 
                           n20899, ZN => n6081);
   U24180 : OAI22_X1 port map( A1 => n27464, A2 => n26920, B1 => n26914, B2 => 
                           n20838, ZN => n6142);
   U24181 : OAI22_X1 port map( A1 => n27467, A2 => n26920, B1 => n26914, B2 => 
                           n20837, ZN => n6143);
   U24182 : OAI22_X1 port map( A1 => n27470, A2 => n26920, B1 => n26914, B2 => 
                           n20836, ZN => n6144);
   U24183 : OAI22_X1 port map( A1 => n27473, A2 => n26920, B1 => n26914, B2 => 
                           n20835, ZN => n6145);
   U24184 : OAI22_X1 port map( A1 => n27463, A2 => n27124, B1 => n9700, B2 => 
                           n27118, ZN => n7230);
   U24185 : OAI22_X1 port map( A1 => n27466, A2 => n27124, B1 => n9699, B2 => 
                           n27118, ZN => n7231);
   U24186 : OAI22_X1 port map( A1 => n27469, A2 => n27124, B1 => n9698, B2 => 
                           n27118, ZN => n7232);
   U24187 : OAI22_X1 port map( A1 => n27472, A2 => n27124, B1 => n9697, B2 => 
                           n27118, ZN => n7233);
   U24188 : OAI22_X1 port map( A1 => n27463, A2 => n27100, B1 => n9508, B2 => 
                           n27094, ZN => n7102);
   U24189 : OAI22_X1 port map( A1 => n27466, A2 => n27100, B1 => n9507, B2 => 
                           n27094, ZN => n7103);
   U24190 : OAI22_X1 port map( A1 => n27469, A2 => n27100, B1 => n9506, B2 => 
                           n27094, ZN => n7104);
   U24191 : OAI22_X1 port map( A1 => n27472, A2 => n27100, B1 => n9505, B2 => 
                           n27094, ZN => n7105);
   U24192 : OAI22_X1 port map( A1 => n27463, A2 => n27040, B1 => n9572, B2 => 
                           n27034, ZN => n6782);
   U24193 : OAI22_X1 port map( A1 => n27466, A2 => n27040, B1 => n9571, B2 => 
                           n27034, ZN => n6783);
   U24194 : OAI22_X1 port map( A1 => n27469, A2 => n27040, B1 => n9570, B2 => 
                           n27034, ZN => n6784);
   U24195 : OAI22_X1 port map( A1 => n27472, A2 => n27040, B1 => n9569, B2 => 
                           n27034, ZN => n6785);
   U24196 : OAI22_X1 port map( A1 => n27463, A2 => n27028, B1 => n9636, B2 => 
                           n27022, ZN => n6718);
   U24197 : OAI22_X1 port map( A1 => n27466, A2 => n27028, B1 => n9635, B2 => 
                           n27022, ZN => n6719);
   U24198 : OAI22_X1 port map( A1 => n27469, A2 => n27028, B1 => n9634, B2 => 
                           n27022, ZN => n6720);
   U24199 : OAI22_X1 port map( A1 => n27472, A2 => n27028, B1 => n9633, B2 => 
                           n27022, ZN => n6721);
   U24200 : AOI22_X1 port map( A1 => n26488, A2 => n25578, B1 => n26482, B2 => 
                           n25566, ZN => n24011);
   U24201 : AOI22_X1 port map( A1 => n26483, A2 => n25655, B1 => n26477, B2 => 
                           n25643, ZN => n25162);
   U24202 : AOI22_X1 port map( A1 => n26483, A2 => n25656, B1 => n26477, B2 => 
                           n25644, ZN => n25134);
   U24203 : AOI22_X1 port map( A1 => n26483, A2 => n25657, B1 => n26477, B2 => 
                           n25645, ZN => n25116);
   U24204 : AOI22_X1 port map( A1 => n26483, A2 => n25658, B1 => n26477, B2 => 
                           n25646, ZN => n25098);
   U24205 : AOI22_X1 port map( A1 => n26483, A2 => n25659, B1 => n26477, B2 => 
                           n25647, ZN => n25080);
   U24206 : AOI22_X1 port map( A1 => n26483, A2 => n25660, B1 => n26477, B2 => 
                           n25648, ZN => n25062);
   U24207 : AOI22_X1 port map( A1 => n26483, A2 => n25661, B1 => n26477, B2 => 
                           n25649, ZN => n25044);
   U24208 : AOI22_X1 port map( A1 => n26483, A2 => n25662, B1 => n26477, B2 => 
                           n25650, ZN => n25026);
   U24209 : AOI22_X1 port map( A1 => n26483, A2 => n25663, B1 => n26477, B2 => 
                           n25651, ZN => n25008);
   U24210 : AOI22_X1 port map( A1 => n26483, A2 => n25664, B1 => n26477, B2 => 
                           n25652, ZN => n24990);
   U24211 : AOI22_X1 port map( A1 => n26483, A2 => n25665, B1 => n26477, B2 => 
                           n25653, ZN => n24972);
   U24212 : AOI22_X1 port map( A1 => n26483, A2 => n25666, B1 => n26477, B2 => 
                           n25654, ZN => n24954);
   U24213 : AOI22_X1 port map( A1 => n26484, A2 => n25455, B1 => n26478, B2 => 
                           n25311, ZN => n24936);
   U24214 : AOI22_X1 port map( A1 => n26484, A2 => n25456, B1 => n26478, B2 => 
                           n25312, ZN => n24918);
   U24215 : AOI22_X1 port map( A1 => n26484, A2 => n25457, B1 => n26478, B2 => 
                           n25313, ZN => n24900);
   U24216 : AOI22_X1 port map( A1 => n26484, A2 => n25458, B1 => n26478, B2 => 
                           n25314, ZN => n24882);
   U24217 : AOI22_X1 port map( A1 => n26484, A2 => n25459, B1 => n26478, B2 => 
                           n25315, ZN => n24864);
   U24218 : AOI22_X1 port map( A1 => n26484, A2 => n25460, B1 => n26478, B2 => 
                           n25316, ZN => n24846);
   U24219 : AOI22_X1 port map( A1 => n26484, A2 => n25461, B1 => n26478, B2 => 
                           n25317, ZN => n24828);
   U24220 : AOI22_X1 port map( A1 => n26484, A2 => n25462, B1 => n26478, B2 => 
                           n25318, ZN => n24810);
   U24221 : AOI22_X1 port map( A1 => n26484, A2 => n25463, B1 => n26478, B2 => 
                           n25319, ZN => n24792);
   U24222 : AOI22_X1 port map( A1 => n26484, A2 => n25464, B1 => n26478, B2 => 
                           n25320, ZN => n24774);
   U24223 : AOI22_X1 port map( A1 => n26484, A2 => n25465, B1 => n26478, B2 => 
                           n25321, ZN => n24756);
   U24224 : AOI22_X1 port map( A1 => n26484, A2 => n25466, B1 => n26478, B2 => 
                           n25322, ZN => n24738);
   U24225 : AOI22_X1 port map( A1 => n26485, A2 => n25467, B1 => n26479, B2 => 
                           n25323, ZN => n24720);
   U24226 : AOI22_X1 port map( A1 => n26485, A2 => n25468, B1 => n26479, B2 => 
                           n25324, ZN => n24702);
   U24227 : AOI22_X1 port map( A1 => n26485, A2 => n25469, B1 => n26479, B2 => 
                           n25325, ZN => n24684);
   U24228 : AOI22_X1 port map( A1 => n26485, A2 => n25470, B1 => n26479, B2 => 
                           n25326, ZN => n24666);
   U24229 : AOI22_X1 port map( A1 => n26485, A2 => n25471, B1 => n26479, B2 => 
                           n25327, ZN => n24648);
   U24230 : AOI22_X1 port map( A1 => n26485, A2 => n25472, B1 => n26479, B2 => 
                           n25328, ZN => n24630);
   U24231 : AOI22_X1 port map( A1 => n26485, A2 => n25473, B1 => n26479, B2 => 
                           n25329, ZN => n24612);
   U24232 : AOI22_X1 port map( A1 => n26485, A2 => n25474, B1 => n26479, B2 => 
                           n25330, ZN => n24594);
   U24233 : AOI22_X1 port map( A1 => n26485, A2 => n25475, B1 => n26479, B2 => 
                           n25331, ZN => n24576);
   U24234 : AOI22_X1 port map( A1 => n26485, A2 => n25476, B1 => n26479, B2 => 
                           n25332, ZN => n24558);
   U24235 : AOI22_X1 port map( A1 => n26485, A2 => n25477, B1 => n26479, B2 => 
                           n25333, ZN => n24540);
   U24236 : AOI22_X1 port map( A1 => n26485, A2 => n25478, B1 => n26479, B2 => 
                           n25334, ZN => n24522);
   U24237 : AOI22_X1 port map( A1 => n26486, A2 => n25479, B1 => n26480, B2 => 
                           n25335, ZN => n24504);
   U24238 : AOI22_X1 port map( A1 => n26486, A2 => n25480, B1 => n26480, B2 => 
                           n25336, ZN => n24486);
   U24239 : AOI22_X1 port map( A1 => n26486, A2 => n25481, B1 => n26480, B2 => 
                           n25337, ZN => n24468);
   U24240 : AOI22_X1 port map( A1 => n26486, A2 => n25482, B1 => n26480, B2 => 
                           n25338, ZN => n24450);
   U24241 : AOI22_X1 port map( A1 => n26486, A2 => n25483, B1 => n26480, B2 => 
                           n25339, ZN => n24432);
   U24242 : AOI22_X1 port map( A1 => n26486, A2 => n25484, B1 => n26480, B2 => 
                           n25340, ZN => n24414);
   U24243 : AOI22_X1 port map( A1 => n26486, A2 => n25485, B1 => n26480, B2 => 
                           n25341, ZN => n24396);
   U24244 : AOI22_X1 port map( A1 => n26486, A2 => n25486, B1 => n26480, B2 => 
                           n25342, ZN => n24378);
   U24245 : AOI22_X1 port map( A1 => n26486, A2 => n25487, B1 => n26480, B2 => 
                           n25343, ZN => n24360);
   U24246 : AOI22_X1 port map( A1 => n26486, A2 => n25488, B1 => n26480, B2 => 
                           n25344, ZN => n24342);
   U24247 : AOI22_X1 port map( A1 => n26486, A2 => n25489, B1 => n26480, B2 => 
                           n25345, ZN => n24324);
   U24248 : AOI22_X1 port map( A1 => n26486, A2 => n25490, B1 => n26480, B2 => 
                           n25346, ZN => n24306);
   U24249 : AOI22_X1 port map( A1 => n26487, A2 => n25491, B1 => n26481, B2 => 
                           n25347, ZN => n24288);
   U24250 : AOI22_X1 port map( A1 => n26487, A2 => n25492, B1 => n26481, B2 => 
                           n25348, ZN => n24270);
   U24251 : AOI22_X1 port map( A1 => n26487, A2 => n25493, B1 => n26481, B2 => 
                           n25349, ZN => n24252);
   U24252 : AOI22_X1 port map( A1 => n26487, A2 => n25494, B1 => n26481, B2 => 
                           n25350, ZN => n24234);
   U24253 : AOI22_X1 port map( A1 => n26487, A2 => n25495, B1 => n26481, B2 => 
                           n25351, ZN => n24216);
   U24254 : AOI22_X1 port map( A1 => n26487, A2 => n25496, B1 => n26481, B2 => 
                           n25352, ZN => n24198);
   U24255 : AOI22_X1 port map( A1 => n26487, A2 => n25497, B1 => n26481, B2 => 
                           n25353, ZN => n24180);
   U24256 : AOI22_X1 port map( A1 => n26487, A2 => n25498, B1 => n26481, B2 => 
                           n25354, ZN => n24162);
   U24257 : AOI22_X1 port map( A1 => n26487, A2 => n25499, B1 => n26481, B2 => 
                           n25355, ZN => n24144);
   U24258 : AOI22_X1 port map( A1 => n26487, A2 => n25500, B1 => n26481, B2 => 
                           n25356, ZN => n24126);
   U24259 : AOI22_X1 port map( A1 => n26487, A2 => n25501, B1 => n26481, B2 => 
                           n25357, ZN => n24108);
   U24260 : AOI22_X1 port map( A1 => n26487, A2 => n25502, B1 => n26481, B2 => 
                           n25358, ZN => n24090);
   U24261 : AOI22_X1 port map( A1 => n26488, A2 => n25575, B1 => n26482, B2 => 
                           n25563, ZN => n24072);
   U24262 : AOI22_X1 port map( A1 => n26488, A2 => n25576, B1 => n26482, B2 => 
                           n25564, ZN => n24054);
   U24263 : AOI22_X1 port map( A1 => n26488, A2 => n25577, B1 => n26482, B2 => 
                           n25565, ZN => n24036);
   U24264 : AOI22_X1 port map( A1 => n26708, A2 => n25655, B1 => n26702, B2 => 
                           n25643, ZN => n23963);
   U24265 : AOI22_X1 port map( A1 => n26708, A2 => n25656, B1 => n26702, B2 => 
                           n25644, ZN => n23935);
   U24266 : AOI22_X1 port map( A1 => n26708, A2 => n25657, B1 => n26702, B2 => 
                           n25645, ZN => n23917);
   U24267 : AOI22_X1 port map( A1 => n26708, A2 => n25658, B1 => n26702, B2 => 
                           n25646, ZN => n23899);
   U24268 : AOI22_X1 port map( A1 => n26708, A2 => n25659, B1 => n26702, B2 => 
                           n25647, ZN => n23881);
   U24269 : AOI22_X1 port map( A1 => n26708, A2 => n25660, B1 => n26702, B2 => 
                           n25648, ZN => n23863);
   U24270 : AOI22_X1 port map( A1 => n26708, A2 => n25661, B1 => n26702, B2 => 
                           n25649, ZN => n23845);
   U24271 : AOI22_X1 port map( A1 => n26708, A2 => n25662, B1 => n26702, B2 => 
                           n25650, ZN => n23827);
   U24272 : AOI22_X1 port map( A1 => n26708, A2 => n25663, B1 => n26702, B2 => 
                           n25651, ZN => n23809);
   U24273 : AOI22_X1 port map( A1 => n26708, A2 => n25664, B1 => n26702, B2 => 
                           n25652, ZN => n23791);
   U24274 : AOI22_X1 port map( A1 => n26708, A2 => n25665, B1 => n26702, B2 => 
                           n25653, ZN => n23773);
   U24275 : AOI22_X1 port map( A1 => n26708, A2 => n25666, B1 => n26702, B2 => 
                           n25654, ZN => n23755);
   U24276 : AOI22_X1 port map( A1 => n26709, A2 => n25455, B1 => n26703, B2 => 
                           n25311, ZN => n23737);
   U24277 : AOI22_X1 port map( A1 => n26709, A2 => n25456, B1 => n26703, B2 => 
                           n25312, ZN => n23719);
   U24278 : AOI22_X1 port map( A1 => n26709, A2 => n25457, B1 => n26703, B2 => 
                           n25313, ZN => n23701);
   U24279 : AOI22_X1 port map( A1 => n26709, A2 => n25458, B1 => n26703, B2 => 
                           n25314, ZN => n23683);
   U24280 : AOI22_X1 port map( A1 => n26709, A2 => n25459, B1 => n26703, B2 => 
                           n25315, ZN => n23665);
   U24281 : AOI22_X1 port map( A1 => n26709, A2 => n25460, B1 => n26703, B2 => 
                           n25316, ZN => n23647);
   U24282 : AOI22_X1 port map( A1 => n26709, A2 => n25461, B1 => n26703, B2 => 
                           n25317, ZN => n23629);
   U24283 : AOI22_X1 port map( A1 => n26709, A2 => n25462, B1 => n26703, B2 => 
                           n25318, ZN => n23611);
   U24284 : AOI22_X1 port map( A1 => n26709, A2 => n25463, B1 => n26703, B2 => 
                           n25319, ZN => n23593);
   U24285 : AOI22_X1 port map( A1 => n26709, A2 => n25464, B1 => n26703, B2 => 
                           n25320, ZN => n23575);
   U24286 : AOI22_X1 port map( A1 => n26709, A2 => n25465, B1 => n26703, B2 => 
                           n25321, ZN => n23557);
   U24287 : AOI22_X1 port map( A1 => n26709, A2 => n25466, B1 => n26703, B2 => 
                           n25322, ZN => n23539);
   U24288 : AOI22_X1 port map( A1 => n26710, A2 => n25467, B1 => n26704, B2 => 
                           n25323, ZN => n23521);
   U24289 : AOI22_X1 port map( A1 => n26710, A2 => n25468, B1 => n26704, B2 => 
                           n25324, ZN => n23503);
   U24290 : AOI22_X1 port map( A1 => n26710, A2 => n25469, B1 => n26704, B2 => 
                           n25325, ZN => n23485);
   U24291 : AOI22_X1 port map( A1 => n26710, A2 => n25470, B1 => n26704, B2 => 
                           n25326, ZN => n23467);
   U24292 : AOI22_X1 port map( A1 => n26710, A2 => n25471, B1 => n26704, B2 => 
                           n25327, ZN => n23449);
   U24293 : AOI22_X1 port map( A1 => n26710, A2 => n25472, B1 => n26704, B2 => 
                           n25328, ZN => n23431);
   U24294 : AOI22_X1 port map( A1 => n26710, A2 => n25473, B1 => n26704, B2 => 
                           n25329, ZN => n23413);
   U24295 : AOI22_X1 port map( A1 => n26710, A2 => n25474, B1 => n26704, B2 => 
                           n25330, ZN => n23395);
   U24296 : AOI22_X1 port map( A1 => n26710, A2 => n25475, B1 => n26704, B2 => 
                           n25331, ZN => n23377);
   U24297 : AOI22_X1 port map( A1 => n26710, A2 => n25476, B1 => n26704, B2 => 
                           n25332, ZN => n23359);
   U24298 : AOI22_X1 port map( A1 => n26710, A2 => n25477, B1 => n26704, B2 => 
                           n25333, ZN => n23341);
   U24299 : AOI22_X1 port map( A1 => n26710, A2 => n25478, B1 => n26704, B2 => 
                           n25334, ZN => n23323);
   U24300 : AOI22_X1 port map( A1 => n26711, A2 => n25479, B1 => n26705, B2 => 
                           n25335, ZN => n23305);
   U24301 : AOI22_X1 port map( A1 => n26711, A2 => n25480, B1 => n26705, B2 => 
                           n25336, ZN => n23287);
   U24302 : AOI22_X1 port map( A1 => n26711, A2 => n25481, B1 => n26705, B2 => 
                           n25337, ZN => n23269);
   U24303 : AOI22_X1 port map( A1 => n26711, A2 => n25482, B1 => n26705, B2 => 
                           n25338, ZN => n23251);
   U24304 : AOI22_X1 port map( A1 => n26711, A2 => n25483, B1 => n26705, B2 => 
                           n25339, ZN => n23233);
   U24305 : AOI22_X1 port map( A1 => n26711, A2 => n25484, B1 => n26705, B2 => 
                           n25340, ZN => n23215);
   U24306 : AOI22_X1 port map( A1 => n26711, A2 => n25485, B1 => n26705, B2 => 
                           n25341, ZN => n23197);
   U24307 : AOI22_X1 port map( A1 => n26711, A2 => n25486, B1 => n26705, B2 => 
                           n25342, ZN => n23179);
   U24308 : AOI22_X1 port map( A1 => n26711, A2 => n25487, B1 => n26705, B2 => 
                           n25343, ZN => n23161);
   U24309 : AOI22_X1 port map( A1 => n26711, A2 => n25488, B1 => n26705, B2 => 
                           n25344, ZN => n23143);
   U24310 : AOI22_X1 port map( A1 => n26711, A2 => n25489, B1 => n26705, B2 => 
                           n25345, ZN => n23125);
   U24311 : AOI22_X1 port map( A1 => n26711, A2 => n25490, B1 => n26705, B2 => 
                           n25346, ZN => n23107);
   U24312 : AOI22_X1 port map( A1 => n26712, A2 => n25491, B1 => n26706, B2 => 
                           n25347, ZN => n23089);
   U24313 : AOI22_X1 port map( A1 => n26712, A2 => n25492, B1 => n26706, B2 => 
                           n25348, ZN => n23071);
   U24314 : AOI22_X1 port map( A1 => n26712, A2 => n25493, B1 => n26706, B2 => 
                           n25349, ZN => n23053);
   U24315 : AOI22_X1 port map( A1 => n26712, A2 => n25494, B1 => n26706, B2 => 
                           n25350, ZN => n23035);
   U24316 : AOI22_X1 port map( A1 => n26712, A2 => n25495, B1 => n26706, B2 => 
                           n25351, ZN => n23017);
   U24317 : AOI22_X1 port map( A1 => n26712, A2 => n25496, B1 => n26706, B2 => 
                           n25352, ZN => n22999);
   U24318 : AOI22_X1 port map( A1 => n26712, A2 => n25497, B1 => n26706, B2 => 
                           n25353, ZN => n22981);
   U24319 : AOI22_X1 port map( A1 => n26712, A2 => n25498, B1 => n26706, B2 => 
                           n25354, ZN => n22963);
   U24320 : AOI22_X1 port map( A1 => n26712, A2 => n25499, B1 => n26706, B2 => 
                           n25355, ZN => n22945);
   U24321 : AOI22_X1 port map( A1 => n26712, A2 => n25500, B1 => n26706, B2 => 
                           n25356, ZN => n22927);
   U24322 : AOI22_X1 port map( A1 => n26712, A2 => n25501, B1 => n26706, B2 => 
                           n25357, ZN => n22909);
   U24323 : AOI22_X1 port map( A1 => n26712, A2 => n25502, B1 => n26706, B2 => 
                           n25358, ZN => n22891);
   U24324 : AOI22_X1 port map( A1 => n26713, A2 => n25575, B1 => n26707, B2 => 
                           n25563, ZN => n22873);
   U24325 : AOI22_X1 port map( A1 => n26713, A2 => n25576, B1 => n26707, B2 => 
                           n25564, ZN => n22855);
   U24326 : AOI22_X1 port map( A1 => n26713, A2 => n25577, B1 => n26707, B2 => 
                           n25565, ZN => n22837);
   U24327 : AOI22_X1 port map( A1 => n26713, A2 => n25578, B1 => n26707, B2 => 
                           n25566, ZN => n22812);
   U24328 : OAI221_X1 port map( B1 => n9584, B2 => n26622, C1 => n20786, C2 => 
                           n26616, A => n24280, ZN => n24275);
   U24329 : AOI22_X1 port map( A1 => n26610, A2 => n25941, B1 => n26604, B2 => 
                           n20986, ZN => n24280);
   U24330 : OAI221_X1 port map( B1 => n9583, B2 => n26622, C1 => n20785, C2 => 
                           n26616, A => n24262, ZN => n24257);
   U24331 : AOI22_X1 port map( A1 => n26610, A2 => n25946, B1 => n26604, B2 => 
                           n20985, ZN => n24262);
   U24332 : OAI221_X1 port map( B1 => n9582, B2 => n26622, C1 => n20784, C2 => 
                           n26616, A => n24244, ZN => n24239);
   U24333 : AOI22_X1 port map( A1 => n26610, A2 => n25951, B1 => n26604, B2 => 
                           n20984, ZN => n24244);
   U24334 : OAI221_X1 port map( B1 => n9581, B2 => n26622, C1 => n20783, C2 => 
                           n26616, A => n24226, ZN => n24221);
   U24335 : AOI22_X1 port map( A1 => n26610, A2 => n25956, B1 => n26604, B2 => 
                           n20983, ZN => n24226);
   U24336 : OAI221_X1 port map( B1 => n9580, B2 => n26622, C1 => n20782, C2 => 
                           n26616, A => n24208, ZN => n24203);
   U24337 : AOI22_X1 port map( A1 => n26610, A2 => n25961, B1 => n26604, B2 => 
                           n20982, ZN => n24208);
   U24338 : OAI221_X1 port map( B1 => n9579, B2 => n26622, C1 => n20781, C2 => 
                           n26616, A => n24190, ZN => n24185);
   U24339 : AOI22_X1 port map( A1 => n26610, A2 => n25966, B1 => n26604, B2 => 
                           n20981, ZN => n24190);
   U24340 : OAI221_X1 port map( B1 => n9578, B2 => n26622, C1 => n20780, C2 => 
                           n26616, A => n24172, ZN => n24167);
   U24341 : AOI22_X1 port map( A1 => n26610, A2 => n25971, B1 => n26604, B2 => 
                           n20980, ZN => n24172);
   U24342 : OAI221_X1 port map( B1 => n9577, B2 => n26622, C1 => n20779, C2 => 
                           n26616, A => n24154, ZN => n24149);
   U24343 : AOI22_X1 port map( A1 => n26610, A2 => n25976, B1 => n26604, B2 => 
                           n20979, ZN => n24154);
   U24344 : OAI221_X1 port map( B1 => n9576, B2 => n26622, C1 => n20778, C2 => 
                           n26616, A => n24136, ZN => n24131);
   U24345 : AOI22_X1 port map( A1 => n26610, A2 => n25981, B1 => n26604, B2 => 
                           n20978, ZN => n24136);
   U24346 : OAI221_X1 port map( B1 => n9575, B2 => n26622, C1 => n20777, C2 => 
                           n26616, A => n24118, ZN => n24113);
   U24347 : AOI22_X1 port map( A1 => n26610, A2 => n25986, B1 => n26604, B2 => 
                           n20977, ZN => n24118);
   U24348 : OAI221_X1 port map( B1 => n9574, B2 => n26622, C1 => n20776, C2 => 
                           n26616, A => n24100, ZN => n24095);
   U24349 : AOI22_X1 port map( A1 => n26610, A2 => n25991, B1 => n26604, B2 => 
                           n20976, ZN => n24100);
   U24350 : OAI221_X1 port map( B1 => n9573, B2 => n26622, C1 => n20775, C2 => 
                           n26616, A => n24082, ZN => n24077);
   U24351 : AOI22_X1 port map( A1 => n26610, A2 => n25996, B1 => n26604, B2 => 
                           n20975, ZN => n24082);
   U24352 : OAI221_X1 port map( B1 => n9584, B2 => n26847, C1 => n20786, C2 => 
                           n26841, A => n23081, ZN => n23076);
   U24353 : AOI22_X1 port map( A1 => n26835, A2 => n25941, B1 => n26829, B2 => 
                           n20986, ZN => n23081);
   U24354 : OAI221_X1 port map( B1 => n9583, B2 => n26847, C1 => n20785, C2 => 
                           n26841, A => n23063, ZN => n23058);
   U24355 : AOI22_X1 port map( A1 => n26835, A2 => n25946, B1 => n26829, B2 => 
                           n20985, ZN => n23063);
   U24356 : OAI221_X1 port map( B1 => n9582, B2 => n26847, C1 => n20784, C2 => 
                           n26841, A => n23045, ZN => n23040);
   U24357 : AOI22_X1 port map( A1 => n26835, A2 => n25951, B1 => n26829, B2 => 
                           n20984, ZN => n23045);
   U24358 : OAI221_X1 port map( B1 => n9581, B2 => n26847, C1 => n20783, C2 => 
                           n26841, A => n23027, ZN => n23022);
   U24359 : AOI22_X1 port map( A1 => n26835, A2 => n25956, B1 => n26829, B2 => 
                           n20983, ZN => n23027);
   U24360 : OAI221_X1 port map( B1 => n9580, B2 => n26847, C1 => n20782, C2 => 
                           n26841, A => n23009, ZN => n23004);
   U24361 : AOI22_X1 port map( A1 => n26835, A2 => n25961, B1 => n26829, B2 => 
                           n20982, ZN => n23009);
   U24362 : OAI221_X1 port map( B1 => n9579, B2 => n26847, C1 => n20781, C2 => 
                           n26841, A => n22991, ZN => n22986);
   U24363 : AOI22_X1 port map( A1 => n26835, A2 => n25966, B1 => n26829, B2 => 
                           n20981, ZN => n22991);
   U24364 : OAI221_X1 port map( B1 => n9578, B2 => n26847, C1 => n20780, C2 => 
                           n26841, A => n22973, ZN => n22968);
   U24365 : AOI22_X1 port map( A1 => n26835, A2 => n25971, B1 => n26829, B2 => 
                           n20980, ZN => n22973);
   U24366 : OAI221_X1 port map( B1 => n9577, B2 => n26847, C1 => n20779, C2 => 
                           n26841, A => n22955, ZN => n22950);
   U24367 : AOI22_X1 port map( A1 => n26835, A2 => n25976, B1 => n26829, B2 => 
                           n20979, ZN => n22955);
   U24368 : OAI221_X1 port map( B1 => n9576, B2 => n26847, C1 => n20778, C2 => 
                           n26841, A => n22937, ZN => n22932);
   U24369 : AOI22_X1 port map( A1 => n26835, A2 => n25981, B1 => n26829, B2 => 
                           n20978, ZN => n22937);
   U24370 : OAI221_X1 port map( B1 => n9575, B2 => n26847, C1 => n20777, C2 => 
                           n26841, A => n22919, ZN => n22914);
   U24371 : AOI22_X1 port map( A1 => n26835, A2 => n25986, B1 => n26829, B2 => 
                           n20977, ZN => n22919);
   U24372 : OAI221_X1 port map( B1 => n9574, B2 => n26847, C1 => n20776, C2 => 
                           n26841, A => n22901, ZN => n22896);
   U24373 : AOI22_X1 port map( A1 => n26835, A2 => n25991, B1 => n26829, B2 => 
                           n20976, ZN => n22901);
   U24374 : OAI221_X1 port map( B1 => n9573, B2 => n26847, C1 => n20775, C2 => 
                           n26841, A => n22883, ZN => n22878);
   U24375 : AOI22_X1 port map( A1 => n26835, A2 => n25996, B1 => n26829, B2 => 
                           n20975, ZN => n22883);
   U24376 : OAI22_X1 port map( A1 => n27283, A2 => n27035, B1 => n9632, B2 => 
                           n27029, ZN => n6722);
   U24377 : OAI22_X1 port map( A1 => n27286, A2 => n27035, B1 => n9631, B2 => 
                           n27029, ZN => n6723);
   U24378 : OAI22_X1 port map( A1 => n27289, A2 => n27035, B1 => n9630, B2 => 
                           n27029, ZN => n6724);
   U24379 : OAI22_X1 port map( A1 => n27292, A2 => n27035, B1 => n9629, B2 => 
                           n27029, ZN => n6725);
   U24380 : OAI22_X1 port map( A1 => n27295, A2 => n27035, B1 => n9628, B2 => 
                           n27029, ZN => n6726);
   U24381 : OAI22_X1 port map( A1 => n27298, A2 => n27035, B1 => n9627, B2 => 
                           n27029, ZN => n6727);
   U24382 : OAI22_X1 port map( A1 => n27301, A2 => n27035, B1 => n9626, B2 => 
                           n27029, ZN => n6728);
   U24383 : OAI22_X1 port map( A1 => n27304, A2 => n27035, B1 => n9625, B2 => 
                           n27029, ZN => n6729);
   U24384 : OAI22_X1 port map( A1 => n27307, A2 => n27035, B1 => n9624, B2 => 
                           n27029, ZN => n6730);
   U24385 : OAI22_X1 port map( A1 => n27310, A2 => n27035, B1 => n9623, B2 => 
                           n27029, ZN => n6731);
   U24386 : OAI22_X1 port map( A1 => n27313, A2 => n27035, B1 => n9622, B2 => 
                           n27029, ZN => n6732);
   U24387 : OAI22_X1 port map( A1 => n27316, A2 => n27036, B1 => n9621, B2 => 
                           n27029, ZN => n6733);
   U24388 : OAI22_X1 port map( A1 => n27319, A2 => n27036, B1 => n9620, B2 => 
                           n27030, ZN => n6734);
   U24389 : OAI22_X1 port map( A1 => n27322, A2 => n27036, B1 => n9619, B2 => 
                           n27030, ZN => n6735);
   U24390 : OAI22_X1 port map( A1 => n27325, A2 => n27036, B1 => n9618, B2 => 
                           n27030, ZN => n6736);
   U24391 : OAI22_X1 port map( A1 => n27328, A2 => n27036, B1 => n9617, B2 => 
                           n27030, ZN => n6737);
   U24392 : OAI22_X1 port map( A1 => n27331, A2 => n27036, B1 => n9616, B2 => 
                           n27030, ZN => n6738);
   U24393 : OAI22_X1 port map( A1 => n27334, A2 => n27036, B1 => n9615, B2 => 
                           n27030, ZN => n6739);
   U24394 : OAI22_X1 port map( A1 => n27337, A2 => n27036, B1 => n9614, B2 => 
                           n27030, ZN => n6740);
   U24395 : OAI22_X1 port map( A1 => n27340, A2 => n27036, B1 => n9613, B2 => 
                           n27030, ZN => n6741);
   U24396 : OAI22_X1 port map( A1 => n27343, A2 => n27036, B1 => n9612, B2 => 
                           n27030, ZN => n6742);
   U24397 : OAI22_X1 port map( A1 => n27346, A2 => n27036, B1 => n9611, B2 => 
                           n27030, ZN => n6743);
   U24398 : OAI22_X1 port map( A1 => n27349, A2 => n27036, B1 => n9610, B2 => 
                           n27030, ZN => n6744);
   U24399 : OAI22_X1 port map( A1 => n27352, A2 => n27037, B1 => n9609, B2 => 
                           n27030, ZN => n6745);
   U24400 : OAI22_X1 port map( A1 => n27355, A2 => n27037, B1 => n9608, B2 => 
                           n27031, ZN => n6746);
   U24401 : OAI22_X1 port map( A1 => n27358, A2 => n27037, B1 => n9607, B2 => 
                           n27031, ZN => n6747);
   U24402 : OAI22_X1 port map( A1 => n27361, A2 => n27037, B1 => n9606, B2 => 
                           n27031, ZN => n6748);
   U24403 : OAI22_X1 port map( A1 => n27364, A2 => n27037, B1 => n9605, B2 => 
                           n27031, ZN => n6749);
   U24404 : OAI22_X1 port map( A1 => n27367, A2 => n27037, B1 => n9604, B2 => 
                           n27031, ZN => n6750);
   U24405 : OAI22_X1 port map( A1 => n27370, A2 => n27037, B1 => n9603, B2 => 
                           n27031, ZN => n6751);
   U24406 : OAI22_X1 port map( A1 => n27373, A2 => n27037, B1 => n9602, B2 => 
                           n27031, ZN => n6752);
   U24407 : OAI22_X1 port map( A1 => n27376, A2 => n27037, B1 => n9601, B2 => 
                           n27031, ZN => n6753);
   U24408 : OAI22_X1 port map( A1 => n27379, A2 => n27037, B1 => n9600, B2 => 
                           n27031, ZN => n6754);
   U24409 : OAI22_X1 port map( A1 => n27382, A2 => n27037, B1 => n9599, B2 => 
                           n27031, ZN => n6755);
   U24410 : OAI22_X1 port map( A1 => n27385, A2 => n27037, B1 => n9598, B2 => 
                           n27031, ZN => n6756);
   U24411 : OAI22_X1 port map( A1 => n27388, A2 => n27038, B1 => n9597, B2 => 
                           n27031, ZN => n6757);
   U24412 : OAI22_X1 port map( A1 => n27391, A2 => n27038, B1 => n9596, B2 => 
                           n27032, ZN => n6758);
   U24413 : OAI22_X1 port map( A1 => n27394, A2 => n27038, B1 => n9595, B2 => 
                           n27032, ZN => n6759);
   U24414 : OAI22_X1 port map( A1 => n27397, A2 => n27038, B1 => n9594, B2 => 
                           n27032, ZN => n6760);
   U24415 : OAI22_X1 port map( A1 => n27400, A2 => n27038, B1 => n9593, B2 => 
                           n27032, ZN => n6761);
   U24416 : OAI22_X1 port map( A1 => n27403, A2 => n27038, B1 => n9592, B2 => 
                           n27032, ZN => n6762);
   U24417 : OAI22_X1 port map( A1 => n27406, A2 => n27038, B1 => n9591, B2 => 
                           n27032, ZN => n6763);
   U24418 : OAI22_X1 port map( A1 => n27409, A2 => n27038, B1 => n9590, B2 => 
                           n27032, ZN => n6764);
   U24419 : OAI22_X1 port map( A1 => n27412, A2 => n27038, B1 => n9589, B2 => 
                           n27032, ZN => n6765);
   U24420 : OAI22_X1 port map( A1 => n27415, A2 => n27038, B1 => n9588, B2 => 
                           n27032, ZN => n6766);
   U24421 : OAI22_X1 port map( A1 => n27418, A2 => n27038, B1 => n9587, B2 => 
                           n27032, ZN => n6767);
   U24422 : OAI22_X1 port map( A1 => n27421, A2 => n27038, B1 => n9586, B2 => 
                           n27032, ZN => n6768);
   U24423 : OAI22_X1 port map( A1 => n27424, A2 => n27039, B1 => n9585, B2 => 
                           n27032, ZN => n6769);
   U24424 : OAI22_X1 port map( A1 => n27427, A2 => n27039, B1 => n9584, B2 => 
                           n27033, ZN => n6770);
   U24425 : OAI22_X1 port map( A1 => n27430, A2 => n27039, B1 => n9583, B2 => 
                           n27033, ZN => n6771);
   U24426 : OAI22_X1 port map( A1 => n27433, A2 => n27039, B1 => n9582, B2 => 
                           n27033, ZN => n6772);
   U24427 : OAI22_X1 port map( A1 => n27436, A2 => n27039, B1 => n9581, B2 => 
                           n27033, ZN => n6773);
   U24428 : OAI22_X1 port map( A1 => n27439, A2 => n27039, B1 => n9580, B2 => 
                           n27033, ZN => n6774);
   U24429 : OAI22_X1 port map( A1 => n27442, A2 => n27039, B1 => n9579, B2 => 
                           n27033, ZN => n6775);
   U24430 : OAI22_X1 port map( A1 => n27445, A2 => n27039, B1 => n9578, B2 => 
                           n27033, ZN => n6776);
   U24431 : OAI22_X1 port map( A1 => n27448, A2 => n27039, B1 => n9577, B2 => 
                           n27033, ZN => n6777);
   U24432 : OAI22_X1 port map( A1 => n27451, A2 => n27039, B1 => n9576, B2 => 
                           n27033, ZN => n6778);
   U24433 : OAI22_X1 port map( A1 => n27454, A2 => n27039, B1 => n9575, B2 => 
                           n27033, ZN => n6779);
   U24434 : OAI22_X1 port map( A1 => n27457, A2 => n27039, B1 => n9574, B2 => 
                           n27033, ZN => n6780);
   U24435 : OAI22_X1 port map( A1 => n27460, A2 => n27040, B1 => n9573, B2 => 
                           n27033, ZN => n6781);
   U24436 : OAI22_X1 port map( A1 => n27283, A2 => n27119, B1 => n9760, B2 => 
                           n27113, ZN => n7170);
   U24437 : OAI22_X1 port map( A1 => n27286, A2 => n27119, B1 => n9759, B2 => 
                           n27113, ZN => n7171);
   U24438 : OAI22_X1 port map( A1 => n27289, A2 => n27119, B1 => n9758, B2 => 
                           n27113, ZN => n7172);
   U24439 : OAI22_X1 port map( A1 => n27292, A2 => n27119, B1 => n9757, B2 => 
                           n27113, ZN => n7173);
   U24440 : OAI22_X1 port map( A1 => n27295, A2 => n27119, B1 => n9756, B2 => 
                           n27113, ZN => n7174);
   U24441 : OAI22_X1 port map( A1 => n27298, A2 => n27119, B1 => n9755, B2 => 
                           n27113, ZN => n7175);
   U24442 : OAI22_X1 port map( A1 => n27301, A2 => n27119, B1 => n9754, B2 => 
                           n27113, ZN => n7176);
   U24443 : OAI22_X1 port map( A1 => n27304, A2 => n27119, B1 => n9753, B2 => 
                           n27113, ZN => n7177);
   U24444 : OAI22_X1 port map( A1 => n27307, A2 => n27119, B1 => n9752, B2 => 
                           n27113, ZN => n7178);
   U24445 : OAI22_X1 port map( A1 => n27310, A2 => n27119, B1 => n9751, B2 => 
                           n27113, ZN => n7179);
   U24446 : OAI22_X1 port map( A1 => n27313, A2 => n27119, B1 => n9750, B2 => 
                           n27113, ZN => n7180);
   U24447 : OAI22_X1 port map( A1 => n27316, A2 => n27120, B1 => n9749, B2 => 
                           n27113, ZN => n7181);
   U24448 : OAI22_X1 port map( A1 => n27319, A2 => n27120, B1 => n9748, B2 => 
                           n27114, ZN => n7182);
   U24449 : OAI22_X1 port map( A1 => n27322, A2 => n27120, B1 => n9747, B2 => 
                           n27114, ZN => n7183);
   U24450 : OAI22_X1 port map( A1 => n27325, A2 => n27120, B1 => n9746, B2 => 
                           n27114, ZN => n7184);
   U24451 : OAI22_X1 port map( A1 => n27328, A2 => n27120, B1 => n9745, B2 => 
                           n27114, ZN => n7185);
   U24452 : OAI22_X1 port map( A1 => n27331, A2 => n27120, B1 => n9744, B2 => 
                           n27114, ZN => n7186);
   U24453 : OAI22_X1 port map( A1 => n27334, A2 => n27120, B1 => n9743, B2 => 
                           n27114, ZN => n7187);
   U24454 : OAI22_X1 port map( A1 => n27337, A2 => n27120, B1 => n9742, B2 => 
                           n27114, ZN => n7188);
   U24455 : OAI22_X1 port map( A1 => n27340, A2 => n27120, B1 => n9741, B2 => 
                           n27114, ZN => n7189);
   U24456 : OAI22_X1 port map( A1 => n27343, A2 => n27120, B1 => n9740, B2 => 
                           n27114, ZN => n7190);
   U24457 : OAI22_X1 port map( A1 => n27346, A2 => n27120, B1 => n9739, B2 => 
                           n27114, ZN => n7191);
   U24458 : OAI22_X1 port map( A1 => n27349, A2 => n27120, B1 => n9738, B2 => 
                           n27114, ZN => n7192);
   U24459 : OAI22_X1 port map( A1 => n27352, A2 => n27121, B1 => n9737, B2 => 
                           n27114, ZN => n7193);
   U24460 : OAI22_X1 port map( A1 => n27355, A2 => n27121, B1 => n9736, B2 => 
                           n27115, ZN => n7194);
   U24461 : OAI22_X1 port map( A1 => n27358, A2 => n27121, B1 => n9735, B2 => 
                           n27115, ZN => n7195);
   U24462 : OAI22_X1 port map( A1 => n27361, A2 => n27121, B1 => n9734, B2 => 
                           n27115, ZN => n7196);
   U24463 : OAI22_X1 port map( A1 => n27364, A2 => n27121, B1 => n9733, B2 => 
                           n27115, ZN => n7197);
   U24464 : OAI22_X1 port map( A1 => n27367, A2 => n27121, B1 => n9732, B2 => 
                           n27115, ZN => n7198);
   U24465 : OAI22_X1 port map( A1 => n27370, A2 => n27121, B1 => n9731, B2 => 
                           n27115, ZN => n7199);
   U24466 : OAI22_X1 port map( A1 => n27373, A2 => n27121, B1 => n9730, B2 => 
                           n27115, ZN => n7200);
   U24467 : OAI22_X1 port map( A1 => n27376, A2 => n27121, B1 => n9729, B2 => 
                           n27115, ZN => n7201);
   U24468 : OAI22_X1 port map( A1 => n27379, A2 => n27121, B1 => n9728, B2 => 
                           n27115, ZN => n7202);
   U24469 : OAI22_X1 port map( A1 => n27382, A2 => n27121, B1 => n9727, B2 => 
                           n27115, ZN => n7203);
   U24470 : OAI22_X1 port map( A1 => n27385, A2 => n27121, B1 => n9726, B2 => 
                           n27115, ZN => n7204);
   U24471 : OAI22_X1 port map( A1 => n27388, A2 => n27122, B1 => n9725, B2 => 
                           n27115, ZN => n7205);
   U24472 : OAI22_X1 port map( A1 => n27391, A2 => n27122, B1 => n9724, B2 => 
                           n27116, ZN => n7206);
   U24473 : OAI22_X1 port map( A1 => n27394, A2 => n27122, B1 => n9723, B2 => 
                           n27116, ZN => n7207);
   U24474 : OAI22_X1 port map( A1 => n27397, A2 => n27122, B1 => n9722, B2 => 
                           n27116, ZN => n7208);
   U24475 : OAI22_X1 port map( A1 => n27400, A2 => n27122, B1 => n9721, B2 => 
                           n27116, ZN => n7209);
   U24476 : OAI22_X1 port map( A1 => n27403, A2 => n27122, B1 => n9720, B2 => 
                           n27116, ZN => n7210);
   U24477 : OAI22_X1 port map( A1 => n27406, A2 => n27122, B1 => n9719, B2 => 
                           n27116, ZN => n7211);
   U24478 : OAI22_X1 port map( A1 => n27409, A2 => n27122, B1 => n9718, B2 => 
                           n27116, ZN => n7212);
   U24479 : OAI22_X1 port map( A1 => n27412, A2 => n27122, B1 => n9717, B2 => 
                           n27116, ZN => n7213);
   U24480 : OAI22_X1 port map( A1 => n27415, A2 => n27122, B1 => n9716, B2 => 
                           n27116, ZN => n7214);
   U24481 : OAI22_X1 port map( A1 => n27418, A2 => n27122, B1 => n9715, B2 => 
                           n27116, ZN => n7215);
   U24482 : OAI22_X1 port map( A1 => n27421, A2 => n27122, B1 => n9714, B2 => 
                           n27116, ZN => n7216);
   U24483 : OAI22_X1 port map( A1 => n27424, A2 => n27123, B1 => n9713, B2 => 
                           n27116, ZN => n7217);
   U24484 : OAI22_X1 port map( A1 => n27427, A2 => n27123, B1 => n9712, B2 => 
                           n27117, ZN => n7218);
   U24485 : OAI22_X1 port map( A1 => n27430, A2 => n27123, B1 => n9711, B2 => 
                           n27117, ZN => n7219);
   U24486 : OAI22_X1 port map( A1 => n27433, A2 => n27123, B1 => n9710, B2 => 
                           n27117, ZN => n7220);
   U24487 : OAI22_X1 port map( A1 => n27436, A2 => n27123, B1 => n9709, B2 => 
                           n27117, ZN => n7221);
   U24488 : OAI22_X1 port map( A1 => n27439, A2 => n27123, B1 => n9708, B2 => 
                           n27117, ZN => n7222);
   U24489 : OAI22_X1 port map( A1 => n27442, A2 => n27123, B1 => n9707, B2 => 
                           n27117, ZN => n7223);
   U24490 : OAI22_X1 port map( A1 => n27445, A2 => n27123, B1 => n9706, B2 => 
                           n27117, ZN => n7224);
   U24491 : OAI22_X1 port map( A1 => n27448, A2 => n27123, B1 => n9705, B2 => 
                           n27117, ZN => n7225);
   U24492 : OAI22_X1 port map( A1 => n27451, A2 => n27123, B1 => n9704, B2 => 
                           n27117, ZN => n7226);
   U24493 : OAI22_X1 port map( A1 => n27454, A2 => n27123, B1 => n9703, B2 => 
                           n27117, ZN => n7227);
   U24494 : OAI22_X1 port map( A1 => n27457, A2 => n27123, B1 => n9702, B2 => 
                           n27117, ZN => n7228);
   U24495 : OAI22_X1 port map( A1 => n27460, A2 => n27124, B1 => n9701, B2 => 
                           n27117, ZN => n7229);
   U24496 : OAI22_X1 port map( A1 => n27283, A2 => n27095, B1 => n9568, B2 => 
                           n27089, ZN => n7042);
   U24497 : OAI22_X1 port map( A1 => n27286, A2 => n27095, B1 => n9567, B2 => 
                           n27089, ZN => n7043);
   U24498 : OAI22_X1 port map( A1 => n27289, A2 => n27095, B1 => n9566, B2 => 
                           n27089, ZN => n7044);
   U24499 : OAI22_X1 port map( A1 => n27292, A2 => n27095, B1 => n9565, B2 => 
                           n27089, ZN => n7045);
   U24500 : OAI22_X1 port map( A1 => n27295, A2 => n27095, B1 => n9564, B2 => 
                           n27089, ZN => n7046);
   U24501 : OAI22_X1 port map( A1 => n27298, A2 => n27095, B1 => n9563, B2 => 
                           n27089, ZN => n7047);
   U24502 : OAI22_X1 port map( A1 => n27301, A2 => n27095, B1 => n9562, B2 => 
                           n27089, ZN => n7048);
   U24503 : OAI22_X1 port map( A1 => n27304, A2 => n27095, B1 => n9561, B2 => 
                           n27089, ZN => n7049);
   U24504 : OAI22_X1 port map( A1 => n27307, A2 => n27095, B1 => n9560, B2 => 
                           n27089, ZN => n7050);
   U24505 : OAI22_X1 port map( A1 => n27310, A2 => n27095, B1 => n9559, B2 => 
                           n27089, ZN => n7051);
   U24506 : OAI22_X1 port map( A1 => n27313, A2 => n27095, B1 => n9558, B2 => 
                           n27089, ZN => n7052);
   U24507 : OAI22_X1 port map( A1 => n27316, A2 => n27096, B1 => n9557, B2 => 
                           n27089, ZN => n7053);
   U24508 : OAI22_X1 port map( A1 => n27319, A2 => n27096, B1 => n9556, B2 => 
                           n27090, ZN => n7054);
   U24509 : OAI22_X1 port map( A1 => n27322, A2 => n27096, B1 => n9555, B2 => 
                           n27090, ZN => n7055);
   U24510 : OAI22_X1 port map( A1 => n27325, A2 => n27096, B1 => n9554, B2 => 
                           n27090, ZN => n7056);
   U24511 : OAI22_X1 port map( A1 => n27328, A2 => n27096, B1 => n9553, B2 => 
                           n27090, ZN => n7057);
   U24512 : OAI22_X1 port map( A1 => n27331, A2 => n27096, B1 => n9552, B2 => 
                           n27090, ZN => n7058);
   U24513 : OAI22_X1 port map( A1 => n27334, A2 => n27096, B1 => n9551, B2 => 
                           n27090, ZN => n7059);
   U24514 : OAI22_X1 port map( A1 => n27337, A2 => n27096, B1 => n9550, B2 => 
                           n27090, ZN => n7060);
   U24515 : OAI22_X1 port map( A1 => n27340, A2 => n27096, B1 => n9549, B2 => 
                           n27090, ZN => n7061);
   U24516 : OAI22_X1 port map( A1 => n27343, A2 => n27096, B1 => n9548, B2 => 
                           n27090, ZN => n7062);
   U24517 : OAI22_X1 port map( A1 => n27346, A2 => n27096, B1 => n9547, B2 => 
                           n27090, ZN => n7063);
   U24518 : OAI22_X1 port map( A1 => n27349, A2 => n27096, B1 => n9546, B2 => 
                           n27090, ZN => n7064);
   U24519 : OAI22_X1 port map( A1 => n27352, A2 => n27097, B1 => n9545, B2 => 
                           n27090, ZN => n7065);
   U24520 : OAI22_X1 port map( A1 => n27355, A2 => n27097, B1 => n9544, B2 => 
                           n27091, ZN => n7066);
   U24521 : OAI22_X1 port map( A1 => n27358, A2 => n27097, B1 => n9543, B2 => 
                           n27091, ZN => n7067);
   U24522 : OAI22_X1 port map( A1 => n27361, A2 => n27097, B1 => n9542, B2 => 
                           n27091, ZN => n7068);
   U24523 : OAI22_X1 port map( A1 => n27364, A2 => n27097, B1 => n9541, B2 => 
                           n27091, ZN => n7069);
   U24524 : OAI22_X1 port map( A1 => n27367, A2 => n27097, B1 => n9540, B2 => 
                           n27091, ZN => n7070);
   U24525 : OAI22_X1 port map( A1 => n27370, A2 => n27097, B1 => n9539, B2 => 
                           n27091, ZN => n7071);
   U24526 : OAI22_X1 port map( A1 => n27373, A2 => n27097, B1 => n9538, B2 => 
                           n27091, ZN => n7072);
   U24527 : OAI22_X1 port map( A1 => n27376, A2 => n27097, B1 => n9537, B2 => 
                           n27091, ZN => n7073);
   U24528 : OAI22_X1 port map( A1 => n27379, A2 => n27097, B1 => n9536, B2 => 
                           n27091, ZN => n7074);
   U24529 : OAI22_X1 port map( A1 => n27382, A2 => n27097, B1 => n9535, B2 => 
                           n27091, ZN => n7075);
   U24530 : OAI22_X1 port map( A1 => n27385, A2 => n27097, B1 => n9534, B2 => 
                           n27091, ZN => n7076);
   U24531 : OAI22_X1 port map( A1 => n27388, A2 => n27098, B1 => n9533, B2 => 
                           n27091, ZN => n7077);
   U24532 : OAI22_X1 port map( A1 => n27391, A2 => n27098, B1 => n9532, B2 => 
                           n27092, ZN => n7078);
   U24533 : OAI22_X1 port map( A1 => n27394, A2 => n27098, B1 => n9531, B2 => 
                           n27092, ZN => n7079);
   U24534 : OAI22_X1 port map( A1 => n27397, A2 => n27098, B1 => n9530, B2 => 
                           n27092, ZN => n7080);
   U24535 : OAI22_X1 port map( A1 => n27400, A2 => n27098, B1 => n9529, B2 => 
                           n27092, ZN => n7081);
   U24536 : OAI22_X1 port map( A1 => n27403, A2 => n27098, B1 => n9528, B2 => 
                           n27092, ZN => n7082);
   U24537 : OAI22_X1 port map( A1 => n27406, A2 => n27098, B1 => n9527, B2 => 
                           n27092, ZN => n7083);
   U24538 : OAI22_X1 port map( A1 => n27409, A2 => n27098, B1 => n9526, B2 => 
                           n27092, ZN => n7084);
   U24539 : OAI22_X1 port map( A1 => n27412, A2 => n27098, B1 => n9525, B2 => 
                           n27092, ZN => n7085);
   U24540 : OAI22_X1 port map( A1 => n27415, A2 => n27098, B1 => n9524, B2 => 
                           n27092, ZN => n7086);
   U24541 : OAI22_X1 port map( A1 => n27418, A2 => n27098, B1 => n9523, B2 => 
                           n27092, ZN => n7087);
   U24542 : OAI22_X1 port map( A1 => n27421, A2 => n27098, B1 => n9522, B2 => 
                           n27092, ZN => n7088);
   U24543 : OAI22_X1 port map( A1 => n27424, A2 => n27099, B1 => n9521, B2 => 
                           n27092, ZN => n7089);
   U24544 : OAI22_X1 port map( A1 => n27427, A2 => n27099, B1 => n9520, B2 => 
                           n27093, ZN => n7090);
   U24545 : OAI22_X1 port map( A1 => n27430, A2 => n27099, B1 => n9519, B2 => 
                           n27093, ZN => n7091);
   U24546 : OAI22_X1 port map( A1 => n27433, A2 => n27099, B1 => n9518, B2 => 
                           n27093, ZN => n7092);
   U24547 : OAI22_X1 port map( A1 => n27436, A2 => n27099, B1 => n9517, B2 => 
                           n27093, ZN => n7093);
   U24548 : OAI22_X1 port map( A1 => n27439, A2 => n27099, B1 => n9516, B2 => 
                           n27093, ZN => n7094);
   U24549 : OAI22_X1 port map( A1 => n27442, A2 => n27099, B1 => n9515, B2 => 
                           n27093, ZN => n7095);
   U24550 : OAI22_X1 port map( A1 => n27445, A2 => n27099, B1 => n9514, B2 => 
                           n27093, ZN => n7096);
   U24551 : OAI22_X1 port map( A1 => n27448, A2 => n27099, B1 => n9513, B2 => 
                           n27093, ZN => n7097);
   U24552 : OAI22_X1 port map( A1 => n27451, A2 => n27099, B1 => n9512, B2 => 
                           n27093, ZN => n7098);
   U24553 : OAI22_X1 port map( A1 => n27454, A2 => n27099, B1 => n9511, B2 => 
                           n27093, ZN => n7099);
   U24554 : OAI22_X1 port map( A1 => n27457, A2 => n27099, B1 => n9510, B2 => 
                           n27093, ZN => n7100);
   U24555 : OAI22_X1 port map( A1 => n27460, A2 => n27100, B1 => n9509, B2 => 
                           n27093, ZN => n7101);
   U24556 : OAI22_X1 port map( A1 => n27283, A2 => n27023, B1 => n9696, B2 => 
                           n27017, ZN => n6658);
   U24557 : OAI22_X1 port map( A1 => n27286, A2 => n27023, B1 => n9695, B2 => 
                           n27017, ZN => n6659);
   U24558 : OAI22_X1 port map( A1 => n27289, A2 => n27023, B1 => n9694, B2 => 
                           n27017, ZN => n6660);
   U24559 : OAI22_X1 port map( A1 => n27292, A2 => n27023, B1 => n9693, B2 => 
                           n27017, ZN => n6661);
   U24560 : OAI22_X1 port map( A1 => n27295, A2 => n27023, B1 => n9692, B2 => 
                           n27017, ZN => n6662);
   U24561 : OAI22_X1 port map( A1 => n27298, A2 => n27023, B1 => n9691, B2 => 
                           n27017, ZN => n6663);
   U24562 : OAI22_X1 port map( A1 => n27301, A2 => n27023, B1 => n9690, B2 => 
                           n27017, ZN => n6664);
   U24563 : OAI22_X1 port map( A1 => n27304, A2 => n27023, B1 => n9689, B2 => 
                           n27017, ZN => n6665);
   U24564 : OAI22_X1 port map( A1 => n27307, A2 => n27023, B1 => n9688, B2 => 
                           n27017, ZN => n6666);
   U24565 : OAI22_X1 port map( A1 => n27310, A2 => n27023, B1 => n9687, B2 => 
                           n27017, ZN => n6667);
   U24566 : OAI22_X1 port map( A1 => n27313, A2 => n27023, B1 => n9686, B2 => 
                           n27017, ZN => n6668);
   U24567 : OAI22_X1 port map( A1 => n27316, A2 => n27024, B1 => n9685, B2 => 
                           n27017, ZN => n6669);
   U24568 : OAI22_X1 port map( A1 => n27319, A2 => n27024, B1 => n9684, B2 => 
                           n27018, ZN => n6670);
   U24569 : OAI22_X1 port map( A1 => n27322, A2 => n27024, B1 => n9683, B2 => 
                           n27018, ZN => n6671);
   U24570 : OAI22_X1 port map( A1 => n27325, A2 => n27024, B1 => n9682, B2 => 
                           n27018, ZN => n6672);
   U24571 : OAI22_X1 port map( A1 => n27328, A2 => n27024, B1 => n9681, B2 => 
                           n27018, ZN => n6673);
   U24572 : OAI22_X1 port map( A1 => n27331, A2 => n27024, B1 => n9680, B2 => 
                           n27018, ZN => n6674);
   U24573 : OAI22_X1 port map( A1 => n27334, A2 => n27024, B1 => n9679, B2 => 
                           n27018, ZN => n6675);
   U24574 : OAI22_X1 port map( A1 => n27337, A2 => n27024, B1 => n9678, B2 => 
                           n27018, ZN => n6676);
   U24575 : OAI22_X1 port map( A1 => n27340, A2 => n27024, B1 => n9677, B2 => 
                           n27018, ZN => n6677);
   U24576 : OAI22_X1 port map( A1 => n27343, A2 => n27024, B1 => n9676, B2 => 
                           n27018, ZN => n6678);
   U24577 : OAI22_X1 port map( A1 => n27346, A2 => n27024, B1 => n9675, B2 => 
                           n27018, ZN => n6679);
   U24578 : OAI22_X1 port map( A1 => n27349, A2 => n27024, B1 => n9674, B2 => 
                           n27018, ZN => n6680);
   U24579 : OAI22_X1 port map( A1 => n27352, A2 => n27025, B1 => n9673, B2 => 
                           n27018, ZN => n6681);
   U24580 : OAI22_X1 port map( A1 => n27355, A2 => n27025, B1 => n9672, B2 => 
                           n27019, ZN => n6682);
   U24581 : OAI22_X1 port map( A1 => n27358, A2 => n27025, B1 => n9671, B2 => 
                           n27019, ZN => n6683);
   U24582 : OAI22_X1 port map( A1 => n27361, A2 => n27025, B1 => n9670, B2 => 
                           n27019, ZN => n6684);
   U24583 : OAI22_X1 port map( A1 => n27364, A2 => n27025, B1 => n9669, B2 => 
                           n27019, ZN => n6685);
   U24584 : OAI22_X1 port map( A1 => n27367, A2 => n27025, B1 => n9668, B2 => 
                           n27019, ZN => n6686);
   U24585 : OAI22_X1 port map( A1 => n27370, A2 => n27025, B1 => n9667, B2 => 
                           n27019, ZN => n6687);
   U24586 : OAI22_X1 port map( A1 => n27373, A2 => n27025, B1 => n9666, B2 => 
                           n27019, ZN => n6688);
   U24587 : OAI22_X1 port map( A1 => n27376, A2 => n27025, B1 => n9665, B2 => 
                           n27019, ZN => n6689);
   U24588 : OAI22_X1 port map( A1 => n27379, A2 => n27025, B1 => n9664, B2 => 
                           n27019, ZN => n6690);
   U24589 : OAI22_X1 port map( A1 => n27382, A2 => n27025, B1 => n9663, B2 => 
                           n27019, ZN => n6691);
   U24590 : OAI22_X1 port map( A1 => n27385, A2 => n27025, B1 => n9662, B2 => 
                           n27019, ZN => n6692);
   U24591 : OAI22_X1 port map( A1 => n27388, A2 => n27026, B1 => n9661, B2 => 
                           n27019, ZN => n6693);
   U24592 : OAI22_X1 port map( A1 => n27391, A2 => n27026, B1 => n9660, B2 => 
                           n27020, ZN => n6694);
   U24593 : OAI22_X1 port map( A1 => n27394, A2 => n27026, B1 => n9659, B2 => 
                           n27020, ZN => n6695);
   U24594 : OAI22_X1 port map( A1 => n27397, A2 => n27026, B1 => n9658, B2 => 
                           n27020, ZN => n6696);
   U24595 : OAI22_X1 port map( A1 => n27400, A2 => n27026, B1 => n9657, B2 => 
                           n27020, ZN => n6697);
   U24596 : OAI22_X1 port map( A1 => n27403, A2 => n27026, B1 => n9656, B2 => 
                           n27020, ZN => n6698);
   U24597 : OAI22_X1 port map( A1 => n27406, A2 => n27026, B1 => n9655, B2 => 
                           n27020, ZN => n6699);
   U24598 : OAI22_X1 port map( A1 => n27409, A2 => n27026, B1 => n9654, B2 => 
                           n27020, ZN => n6700);
   U24599 : OAI22_X1 port map( A1 => n27412, A2 => n27026, B1 => n9653, B2 => 
                           n27020, ZN => n6701);
   U24600 : OAI22_X1 port map( A1 => n27415, A2 => n27026, B1 => n9652, B2 => 
                           n27020, ZN => n6702);
   U24601 : OAI22_X1 port map( A1 => n27418, A2 => n27026, B1 => n9651, B2 => 
                           n27020, ZN => n6703);
   U24602 : OAI22_X1 port map( A1 => n27421, A2 => n27026, B1 => n9650, B2 => 
                           n27020, ZN => n6704);
   U24603 : OAI22_X1 port map( A1 => n27424, A2 => n27027, B1 => n9649, B2 => 
                           n27020, ZN => n6705);
   U24604 : OAI22_X1 port map( A1 => n27427, A2 => n27027, B1 => n9648, B2 => 
                           n27021, ZN => n6706);
   U24605 : OAI22_X1 port map( A1 => n27430, A2 => n27027, B1 => n9647, B2 => 
                           n27021, ZN => n6707);
   U24606 : OAI22_X1 port map( A1 => n27433, A2 => n27027, B1 => n9646, B2 => 
                           n27021, ZN => n6708);
   U24607 : OAI22_X1 port map( A1 => n27436, A2 => n27027, B1 => n9645, B2 => 
                           n27021, ZN => n6709);
   U24608 : OAI22_X1 port map( A1 => n27439, A2 => n27027, B1 => n9644, B2 => 
                           n27021, ZN => n6710);
   U24609 : OAI22_X1 port map( A1 => n27442, A2 => n27027, B1 => n9643, B2 => 
                           n27021, ZN => n6711);
   U24610 : OAI22_X1 port map( A1 => n27445, A2 => n27027, B1 => n9642, B2 => 
                           n27021, ZN => n6712);
   U24611 : OAI22_X1 port map( A1 => n27448, A2 => n27027, B1 => n9641, B2 => 
                           n27021, ZN => n6713);
   U24612 : OAI22_X1 port map( A1 => n27451, A2 => n27027, B1 => n9640, B2 => 
                           n27021, ZN => n6714);
   U24613 : OAI22_X1 port map( A1 => n27454, A2 => n27027, B1 => n9639, B2 => 
                           n27021, ZN => n6715);
   U24614 : OAI22_X1 port map( A1 => n27457, A2 => n27027, B1 => n9638, B2 => 
                           n27021, ZN => n6716);
   U24615 : OAI22_X1 port map( A1 => n27460, A2 => n27028, B1 => n9637, B2 => 
                           n27021, ZN => n6717);
   U24616 : OAI22_X1 port map( A1 => n27284, A2 => n26951, B1 => n26945, B2 => 
                           n22631, ZN => n6274);
   U24617 : OAI22_X1 port map( A1 => n27287, A2 => n26951, B1 => n26945, B2 => 
                           n22630, ZN => n6275);
   U24618 : OAI22_X1 port map( A1 => n27290, A2 => n26951, B1 => n26945, B2 => 
                           n22629, ZN => n6276);
   U24619 : OAI22_X1 port map( A1 => n27293, A2 => n26951, B1 => n26945, B2 => 
                           n22628, ZN => n6277);
   U24620 : OAI22_X1 port map( A1 => n27296, A2 => n26951, B1 => n26945, B2 => 
                           n22627, ZN => n6278);
   U24621 : OAI22_X1 port map( A1 => n27299, A2 => n26951, B1 => n26945, B2 => 
                           n22626, ZN => n6279);
   U24622 : OAI22_X1 port map( A1 => n27302, A2 => n26951, B1 => n26945, B2 => 
                           n22625, ZN => n6280);
   U24623 : OAI22_X1 port map( A1 => n27305, A2 => n26951, B1 => n26945, B2 => 
                           n22624, ZN => n6281);
   U24624 : OAI22_X1 port map( A1 => n27308, A2 => n26951, B1 => n26945, B2 => 
                           n22623, ZN => n6282);
   U24625 : OAI22_X1 port map( A1 => n27311, A2 => n26951, B1 => n26945, B2 => 
                           n22622, ZN => n6283);
   U24626 : OAI22_X1 port map( A1 => n27314, A2 => n26951, B1 => n26945, B2 => 
                           n22621, ZN => n6284);
   U24627 : OAI22_X1 port map( A1 => n27317, A2 => n26952, B1 => n26945, B2 => 
                           n22620, ZN => n6285);
   U24628 : OAI22_X1 port map( A1 => n27282, A2 => n27155, B1 => n27149, B2 => 
                           n22439, ZN => n7362);
   U24629 : OAI22_X1 port map( A1 => n27285, A2 => n27155, B1 => n27149, B2 => 
                           n22438, ZN => n7363);
   U24630 : OAI22_X1 port map( A1 => n27288, A2 => n27155, B1 => n27149, B2 => 
                           n22437, ZN => n7364);
   U24631 : OAI22_X1 port map( A1 => n27291, A2 => n27155, B1 => n27149, B2 => 
                           n22436, ZN => n7365);
   U24632 : OAI22_X1 port map( A1 => n27294, A2 => n27155, B1 => n27149, B2 => 
                           n22435, ZN => n7366);
   U24633 : OAI22_X1 port map( A1 => n27297, A2 => n27155, B1 => n27149, B2 => 
                           n22434, ZN => n7367);
   U24634 : OAI22_X1 port map( A1 => n27300, A2 => n27155, B1 => n27149, B2 => 
                           n22433, ZN => n7368);
   U24635 : OAI22_X1 port map( A1 => n27303, A2 => n27155, B1 => n27149, B2 => 
                           n22432, ZN => n7369);
   U24636 : OAI22_X1 port map( A1 => n27306, A2 => n27155, B1 => n27149, B2 => 
                           n22431, ZN => n7370);
   U24637 : OAI22_X1 port map( A1 => n27309, A2 => n27155, B1 => n27149, B2 => 
                           n22430, ZN => n7371);
   U24638 : OAI22_X1 port map( A1 => n27312, A2 => n27155, B1 => n27149, B2 => 
                           n22429, ZN => n7372);
   U24639 : OAI22_X1 port map( A1 => n27315, A2 => n27156, B1 => n27149, B2 => 
                           n22428, ZN => n7373);
   U24640 : OAI22_X1 port map( A1 => n27284, A2 => n26927, B1 => n26921, B2 => 
                           n22319, ZN => n6146);
   U24641 : OAI22_X1 port map( A1 => n27287, A2 => n26927, B1 => n26921, B2 => 
                           n22318, ZN => n6147);
   U24642 : OAI22_X1 port map( A1 => n27290, A2 => n26927, B1 => n26921, B2 => 
                           n22317, ZN => n6148);
   U24643 : OAI22_X1 port map( A1 => n27293, A2 => n26927, B1 => n26921, B2 => 
                           n22316, ZN => n6149);
   U24644 : OAI22_X1 port map( A1 => n27296, A2 => n26927, B1 => n26921, B2 => 
                           n22315, ZN => n6150);
   U24645 : OAI22_X1 port map( A1 => n27299, A2 => n26927, B1 => n26921, B2 => 
                           n22314, ZN => n6151);
   U24646 : OAI22_X1 port map( A1 => n27302, A2 => n26927, B1 => n26921, B2 => 
                           n22313, ZN => n6152);
   U24647 : OAI22_X1 port map( A1 => n27305, A2 => n26927, B1 => n26921, B2 => 
                           n22312, ZN => n6153);
   U24648 : OAI22_X1 port map( A1 => n27308, A2 => n26927, B1 => n26921, B2 => 
                           n22311, ZN => n6154);
   U24649 : OAI22_X1 port map( A1 => n27311, A2 => n26927, B1 => n26921, B2 => 
                           n22310, ZN => n6155);
   U24650 : OAI22_X1 port map( A1 => n27314, A2 => n26927, B1 => n26921, B2 => 
                           n22309, ZN => n6156);
   U24651 : OAI22_X1 port map( A1 => n27317, A2 => n26928, B1 => n26921, B2 => 
                           n22308, ZN => n6157);
   U24652 : OAI22_X1 port map( A1 => n27284, A2 => n26939, B1 => n26933, B2 => 
                           n22243, ZN => n6210);
   U24653 : OAI22_X1 port map( A1 => n27287, A2 => n26939, B1 => n26933, B2 => 
                           n22242, ZN => n6211);
   U24654 : OAI22_X1 port map( A1 => n27290, A2 => n26939, B1 => n26933, B2 => 
                           n22241, ZN => n6212);
   U24655 : OAI22_X1 port map( A1 => n27293, A2 => n26939, B1 => n26933, B2 => 
                           n22240, ZN => n6213);
   U24656 : OAI22_X1 port map( A1 => n27296, A2 => n26939, B1 => n26933, B2 => 
                           n22239, ZN => n6214);
   U24657 : OAI22_X1 port map( A1 => n27299, A2 => n26939, B1 => n26933, B2 => 
                           n22238, ZN => n6215);
   U24658 : OAI22_X1 port map( A1 => n27302, A2 => n26939, B1 => n26933, B2 => 
                           n22237, ZN => n6216);
   U24659 : OAI22_X1 port map( A1 => n27305, A2 => n26939, B1 => n26933, B2 => 
                           n22236, ZN => n6217);
   U24660 : OAI22_X1 port map( A1 => n27308, A2 => n26939, B1 => n26933, B2 => 
                           n22235, ZN => n6218);
   U24661 : OAI22_X1 port map( A1 => n27311, A2 => n26939, B1 => n26933, B2 => 
                           n22234, ZN => n6219);
   U24662 : OAI22_X1 port map( A1 => n27314, A2 => n26939, B1 => n26933, B2 => 
                           n22233, ZN => n6220);
   U24663 : OAI22_X1 port map( A1 => n27317, A2 => n26940, B1 => n26933, B2 => 
                           n22232, ZN => n6221);
   U24664 : OAI22_X1 port map( A1 => n27277, A2 => n27282, B1 => n27269, B2 => 
                           n22179, ZN => n8002);
   U24665 : OAI22_X1 port map( A1 => n27277, A2 => n27285, B1 => n27269, B2 => 
                           n22178, ZN => n8003);
   U24666 : OAI22_X1 port map( A1 => n27277, A2 => n27288, B1 => n27269, B2 => 
                           n22177, ZN => n8004);
   U24667 : OAI22_X1 port map( A1 => n27277, A2 => n27291, B1 => n27269, B2 => 
                           n22176, ZN => n8005);
   U24668 : OAI22_X1 port map( A1 => n27277, A2 => n27294, B1 => n27269, B2 => 
                           n22175, ZN => n8006);
   U24669 : OAI22_X1 port map( A1 => n27277, A2 => n27297, B1 => n27269, B2 => 
                           n22174, ZN => n8007);
   U24670 : OAI22_X1 port map( A1 => n27277, A2 => n27300, B1 => n27269, B2 => 
                           n22173, ZN => n8008);
   U24671 : OAI22_X1 port map( A1 => n27277, A2 => n27303, B1 => n27269, B2 => 
                           n22172, ZN => n8009);
   U24672 : OAI22_X1 port map( A1 => n27277, A2 => n27306, B1 => n27269, B2 => 
                           n22171, ZN => n8010);
   U24673 : OAI22_X1 port map( A1 => n27277, A2 => n27309, B1 => n27269, B2 => 
                           n22170, ZN => n8011);
   U24674 : OAI22_X1 port map( A1 => n27277, A2 => n27312, B1 => n27269, B2 => 
                           n22169, ZN => n8012);
   U24675 : OAI22_X1 port map( A1 => n27277, A2 => n27315, B1 => n27269, B2 => 
                           n22168, ZN => n8013);
   U24676 : OAI22_X1 port map( A1 => n27282, A2 => n27263, B1 => n27257, B2 => 
                           n22119, ZN => n7938);
   U24677 : OAI22_X1 port map( A1 => n27285, A2 => n27263, B1 => n27257, B2 => 
                           n22118, ZN => n7939);
   U24678 : OAI22_X1 port map( A1 => n27288, A2 => n27263, B1 => n27257, B2 => 
                           n22117, ZN => n7940);
   U24679 : OAI22_X1 port map( A1 => n27291, A2 => n27263, B1 => n27257, B2 => 
                           n22116, ZN => n7941);
   U24680 : OAI22_X1 port map( A1 => n27294, A2 => n27263, B1 => n27257, B2 => 
                           n22115, ZN => n7942);
   U24681 : OAI22_X1 port map( A1 => n27297, A2 => n27263, B1 => n27257, B2 => 
                           n22114, ZN => n7943);
   U24682 : OAI22_X1 port map( A1 => n27300, A2 => n27263, B1 => n27257, B2 => 
                           n22113, ZN => n7944);
   U24683 : OAI22_X1 port map( A1 => n27303, A2 => n27263, B1 => n27257, B2 => 
                           n22112, ZN => n7945);
   U24684 : OAI22_X1 port map( A1 => n27306, A2 => n27263, B1 => n27257, B2 => 
                           n22111, ZN => n7946);
   U24685 : OAI22_X1 port map( A1 => n27309, A2 => n27263, B1 => n27257, B2 => 
                           n22110, ZN => n7947);
   U24686 : OAI22_X1 port map( A1 => n27312, A2 => n27263, B1 => n27257, B2 => 
                           n22109, ZN => n7948);
   U24687 : OAI22_X1 port map( A1 => n27315, A2 => n27264, B1 => n27257, B2 => 
                           n22108, ZN => n7949);
   U24688 : OAI22_X1 port map( A1 => n27282, A2 => n27227, B1 => n27221, B2 => 
                           n21939, ZN => n7746);
   U24689 : OAI22_X1 port map( A1 => n27285, A2 => n27227, B1 => n27221, B2 => 
                           n21938, ZN => n7747);
   U24690 : OAI22_X1 port map( A1 => n27288, A2 => n27227, B1 => n27221, B2 => 
                           n21937, ZN => n7748);
   U24691 : OAI22_X1 port map( A1 => n27291, A2 => n27227, B1 => n27221, B2 => 
                           n21936, ZN => n7749);
   U24692 : OAI22_X1 port map( A1 => n27294, A2 => n27227, B1 => n27221, B2 => 
                           n21935, ZN => n7750);
   U24693 : OAI22_X1 port map( A1 => n27297, A2 => n27227, B1 => n27221, B2 => 
                           n21934, ZN => n7751);
   U24694 : OAI22_X1 port map( A1 => n27300, A2 => n27227, B1 => n27221, B2 => 
                           n21933, ZN => n7752);
   U24695 : OAI22_X1 port map( A1 => n27303, A2 => n27227, B1 => n27221, B2 => 
                           n21932, ZN => n7753);
   U24696 : OAI22_X1 port map( A1 => n27306, A2 => n27227, B1 => n27221, B2 => 
                           n21931, ZN => n7754);
   U24697 : OAI22_X1 port map( A1 => n27309, A2 => n27227, B1 => n27221, B2 => 
                           n21930, ZN => n7755);
   U24698 : OAI22_X1 port map( A1 => n27312, A2 => n27227, B1 => n27221, B2 => 
                           n21929, ZN => n7756);
   U24699 : OAI22_X1 port map( A1 => n27315, A2 => n27228, B1 => n27221, B2 => 
                           n21928, ZN => n7757);
   U24700 : OAI22_X1 port map( A1 => n27282, A2 => n27203, B1 => n27197, B2 => 
                           n21879, ZN => n7618);
   U24701 : OAI22_X1 port map( A1 => n27285, A2 => n27203, B1 => n27197, B2 => 
                           n21878, ZN => n7619);
   U24702 : OAI22_X1 port map( A1 => n27288, A2 => n27203, B1 => n27197, B2 => 
                           n21877, ZN => n7620);
   U24703 : OAI22_X1 port map( A1 => n27291, A2 => n27203, B1 => n27197, B2 => 
                           n21876, ZN => n7621);
   U24704 : OAI22_X1 port map( A1 => n27294, A2 => n27203, B1 => n27197, B2 => 
                           n21875, ZN => n7622);
   U24705 : OAI22_X1 port map( A1 => n27297, A2 => n27203, B1 => n27197, B2 => 
                           n21874, ZN => n7623);
   U24706 : OAI22_X1 port map( A1 => n27300, A2 => n27203, B1 => n27197, B2 => 
                           n21873, ZN => n7624);
   U24707 : OAI22_X1 port map( A1 => n27303, A2 => n27203, B1 => n27197, B2 => 
                           n21872, ZN => n7625);
   U24708 : OAI22_X1 port map( A1 => n27306, A2 => n27203, B1 => n27197, B2 => 
                           n21871, ZN => n7626);
   U24709 : OAI22_X1 port map( A1 => n27309, A2 => n27203, B1 => n27197, B2 => 
                           n21870, ZN => n7627);
   U24710 : OAI22_X1 port map( A1 => n27312, A2 => n27203, B1 => n27197, B2 => 
                           n21869, ZN => n7628);
   U24711 : OAI22_X1 port map( A1 => n27315, A2 => n27204, B1 => n27197, B2 => 
                           n21868, ZN => n7629);
   U24712 : OAI22_X1 port map( A1 => n27283, A2 => n27011, B1 => n27005, B2 => 
                           n21819, ZN => n6594);
   U24713 : OAI22_X1 port map( A1 => n27286, A2 => n27011, B1 => n27005, B2 => 
                           n21818, ZN => n6595);
   U24714 : OAI22_X1 port map( A1 => n27289, A2 => n27011, B1 => n27005, B2 => 
                           n21817, ZN => n6596);
   U24715 : OAI22_X1 port map( A1 => n27292, A2 => n27011, B1 => n27005, B2 => 
                           n21816, ZN => n6597);
   U24716 : OAI22_X1 port map( A1 => n27295, A2 => n27011, B1 => n27005, B2 => 
                           n21815, ZN => n6598);
   U24717 : OAI22_X1 port map( A1 => n27298, A2 => n27011, B1 => n27005, B2 => 
                           n21814, ZN => n6599);
   U24718 : OAI22_X1 port map( A1 => n27301, A2 => n27011, B1 => n27005, B2 => 
                           n21813, ZN => n6600);
   U24719 : OAI22_X1 port map( A1 => n27304, A2 => n27011, B1 => n27005, B2 => 
                           n21812, ZN => n6601);
   U24720 : OAI22_X1 port map( A1 => n27307, A2 => n27011, B1 => n27005, B2 => 
                           n21811, ZN => n6602);
   U24721 : OAI22_X1 port map( A1 => n27310, A2 => n27011, B1 => n27005, B2 => 
                           n21810, ZN => n6603);
   U24722 : OAI22_X1 port map( A1 => n27313, A2 => n27011, B1 => n27005, B2 => 
                           n21809, ZN => n6604);
   U24723 : OAI22_X1 port map( A1 => n27316, A2 => n27012, B1 => n27005, B2 => 
                           n21808, ZN => n6605);
   U24724 : OAI22_X1 port map( A1 => n27283, A2 => n27059, B1 => n27053, B2 => 
                           n21699, ZN => n6850);
   U24725 : OAI22_X1 port map( A1 => n27286, A2 => n27059, B1 => n27053, B2 => 
                           n21698, ZN => n6851);
   U24726 : OAI22_X1 port map( A1 => n27289, A2 => n27059, B1 => n27053, B2 => 
                           n21697, ZN => n6852);
   U24727 : OAI22_X1 port map( A1 => n27292, A2 => n27059, B1 => n27053, B2 => 
                           n21696, ZN => n6853);
   U24728 : OAI22_X1 port map( A1 => n27295, A2 => n27059, B1 => n27053, B2 => 
                           n21695, ZN => n6854);
   U24729 : OAI22_X1 port map( A1 => n27298, A2 => n27059, B1 => n27053, B2 => 
                           n21694, ZN => n6855);
   U24730 : OAI22_X1 port map( A1 => n27301, A2 => n27059, B1 => n27053, B2 => 
                           n21693, ZN => n6856);
   U24731 : OAI22_X1 port map( A1 => n27304, A2 => n27059, B1 => n27053, B2 => 
                           n21692, ZN => n6857);
   U24732 : OAI22_X1 port map( A1 => n27307, A2 => n27059, B1 => n27053, B2 => 
                           n21691, ZN => n6858);
   U24733 : OAI22_X1 port map( A1 => n27310, A2 => n27059, B1 => n27053, B2 => 
                           n21690, ZN => n6859);
   U24734 : OAI22_X1 port map( A1 => n27313, A2 => n27059, B1 => n27053, B2 => 
                           n21689, ZN => n6860);
   U24735 : OAI22_X1 port map( A1 => n27316, A2 => n27060, B1 => n27053, B2 => 
                           n21688, ZN => n6861);
   U24736 : OAI22_X1 port map( A1 => n27282, A2 => n27251, B1 => n27245, B2 => 
                           n21479, ZN => n7874);
   U24737 : OAI22_X1 port map( A1 => n27285, A2 => n27251, B1 => n27245, B2 => 
                           n21478, ZN => n7875);
   U24738 : OAI22_X1 port map( A1 => n27288, A2 => n27251, B1 => n27245, B2 => 
                           n21477, ZN => n7876);
   U24739 : OAI22_X1 port map( A1 => n27291, A2 => n27251, B1 => n27245, B2 => 
                           n21476, ZN => n7877);
   U24740 : OAI22_X1 port map( A1 => n27294, A2 => n27251, B1 => n27245, B2 => 
                           n21475, ZN => n7878);
   U24741 : OAI22_X1 port map( A1 => n27297, A2 => n27251, B1 => n27245, B2 => 
                           n21474, ZN => n7879);
   U24742 : OAI22_X1 port map( A1 => n27300, A2 => n27251, B1 => n27245, B2 => 
                           n21473, ZN => n7880);
   U24743 : OAI22_X1 port map( A1 => n27303, A2 => n27251, B1 => n27245, B2 => 
                           n21472, ZN => n7881);
   U24744 : OAI22_X1 port map( A1 => n27306, A2 => n27251, B1 => n27245, B2 => 
                           n21471, ZN => n7882);
   U24745 : OAI22_X1 port map( A1 => n27309, A2 => n27251, B1 => n27245, B2 => 
                           n21470, ZN => n7883);
   U24746 : OAI22_X1 port map( A1 => n27312, A2 => n27251, B1 => n27245, B2 => 
                           n21469, ZN => n7884);
   U24747 : OAI22_X1 port map( A1 => n27315, A2 => n27252, B1 => n27245, B2 => 
                           n21468, ZN => n7885);
   U24748 : OAI22_X1 port map( A1 => n27283, A2 => n27083, B1 => n27077, B2 => 
                           n21299, ZN => n6978);
   U24749 : OAI22_X1 port map( A1 => n27286, A2 => n27083, B1 => n27077, B2 => 
                           n21298, ZN => n6979);
   U24750 : OAI22_X1 port map( A1 => n27289, A2 => n27083, B1 => n27077, B2 => 
                           n21297, ZN => n6980);
   U24751 : OAI22_X1 port map( A1 => n27292, A2 => n27083, B1 => n27077, B2 => 
                           n21296, ZN => n6981);
   U24752 : OAI22_X1 port map( A1 => n27295, A2 => n27083, B1 => n27077, B2 => 
                           n21295, ZN => n6982);
   U24753 : OAI22_X1 port map( A1 => n27298, A2 => n27083, B1 => n27077, B2 => 
                           n21294, ZN => n6983);
   U24754 : OAI22_X1 port map( A1 => n27301, A2 => n27083, B1 => n27077, B2 => 
                           n21293, ZN => n6984);
   U24755 : OAI22_X1 port map( A1 => n27304, A2 => n27083, B1 => n27077, B2 => 
                           n21292, ZN => n6985);
   U24756 : OAI22_X1 port map( A1 => n27307, A2 => n27083, B1 => n27077, B2 => 
                           n21291, ZN => n6986);
   U24757 : OAI22_X1 port map( A1 => n27310, A2 => n27083, B1 => n27077, B2 => 
                           n21290, ZN => n6987);
   U24758 : OAI22_X1 port map( A1 => n27313, A2 => n27083, B1 => n27077, B2 => 
                           n21289, ZN => n6988);
   U24759 : OAI22_X1 port map( A1 => n27316, A2 => n27084, B1 => n27077, B2 => 
                           n21288, ZN => n6989);
   U24760 : OAI22_X1 port map( A1 => n27284, A2 => n26903, B1 => n26897, B2 => 
                           n20962, ZN => n6018);
   U24761 : OAI22_X1 port map( A1 => n27287, A2 => n26903, B1 => n26897, B2 => 
                           n20961, ZN => n6019);
   U24762 : OAI22_X1 port map( A1 => n27290, A2 => n26903, B1 => n26897, B2 => 
                           n20960, ZN => n6020);
   U24763 : OAI22_X1 port map( A1 => n27293, A2 => n26903, B1 => n26897, B2 => 
                           n20959, ZN => n6021);
   U24764 : OAI22_X1 port map( A1 => n27296, A2 => n26903, B1 => n26897, B2 => 
                           n20958, ZN => n6022);
   U24765 : OAI22_X1 port map( A1 => n27299, A2 => n26903, B1 => n26897, B2 => 
                           n20957, ZN => n6023);
   U24766 : OAI22_X1 port map( A1 => n27302, A2 => n26903, B1 => n26897, B2 => 
                           n20956, ZN => n6024);
   U24767 : OAI22_X1 port map( A1 => n27305, A2 => n26903, B1 => n26897, B2 => 
                           n20955, ZN => n6025);
   U24768 : OAI22_X1 port map( A1 => n27308, A2 => n26903, B1 => n26897, B2 => 
                           n20954, ZN => n6026);
   U24769 : OAI22_X1 port map( A1 => n27311, A2 => n26903, B1 => n26897, B2 => 
                           n20953, ZN => n6027);
   U24770 : OAI22_X1 port map( A1 => n27314, A2 => n26903, B1 => n26897, B2 => 
                           n20952, ZN => n6028);
   U24771 : OAI22_X1 port map( A1 => n27317, A2 => n26904, B1 => n26897, B2 => 
                           n20951, ZN => n6029);
   U24772 : OAI22_X1 port map( A1 => n27284, A2 => n26915, B1 => n26909, B2 => 
                           n20898, ZN => n6082);
   U24773 : OAI22_X1 port map( A1 => n27287, A2 => n26915, B1 => n26909, B2 => 
                           n20897, ZN => n6083);
   U24774 : OAI22_X1 port map( A1 => n27290, A2 => n26915, B1 => n26909, B2 => 
                           n20896, ZN => n6084);
   U24775 : OAI22_X1 port map( A1 => n27293, A2 => n26915, B1 => n26909, B2 => 
                           n20895, ZN => n6085);
   U24776 : OAI22_X1 port map( A1 => n27296, A2 => n26915, B1 => n26909, B2 => 
                           n20894, ZN => n6086);
   U24777 : OAI22_X1 port map( A1 => n27299, A2 => n26915, B1 => n26909, B2 => 
                           n20893, ZN => n6087);
   U24778 : OAI22_X1 port map( A1 => n27302, A2 => n26915, B1 => n26909, B2 => 
                           n20892, ZN => n6088);
   U24779 : OAI22_X1 port map( A1 => n27305, A2 => n26915, B1 => n26909, B2 => 
                           n20891, ZN => n6089);
   U24780 : OAI22_X1 port map( A1 => n27308, A2 => n26915, B1 => n26909, B2 => 
                           n20890, ZN => n6090);
   U24781 : OAI22_X1 port map( A1 => n27311, A2 => n26915, B1 => n26909, B2 => 
                           n20889, ZN => n6091);
   U24782 : OAI22_X1 port map( A1 => n27314, A2 => n26915, B1 => n26909, B2 => 
                           n20888, ZN => n6092);
   U24783 : OAI22_X1 port map( A1 => n27317, A2 => n26916, B1 => n26909, B2 => 
                           n20887, ZN => n6093);
   U24784 : OAI21_X1 port map( B1 => n26533, B2 => n19454, A => ENABLE, ZN => 
                           n19580);
   U24785 : OAI21_X1 port map( B1 => n26533, B2 => n18553, A => n27481, ZN => 
                           n19507);
   U24786 : OAI21_X1 port map( B1 => n26533, B2 => n18536, A => n27481, ZN => 
                           n19508);
   U24787 : OAI21_X1 port map( B1 => n26533, B2 => n18519, A => n27481, ZN => 
                           n19509);
   U24788 : OAI21_X1 port map( B1 => n26533, B2 => n18502, A => n27481, ZN => 
                           n19510);
   U24789 : OAI21_X1 port map( B1 => n26533, B2 => n18485, A => n27481, ZN => 
                           n19511);
   U24790 : OAI21_X1 port map( B1 => n26533, B2 => n18468, A => n27481, ZN => 
                           n19512);
   U24791 : OAI21_X1 port map( B1 => n26533, B2 => n18451, A => n27481, ZN => 
                           n19513);
   U24792 : OAI21_X1 port map( B1 => n26533, B2 => n18434, A => n27481, ZN => 
                           n19514);
   U24793 : OAI21_X1 port map( B1 => n26533, B2 => n18417, A => n27482, ZN => 
                           n19515);
   U24794 : OAI21_X1 port map( B1 => n26533, B2 => n18400, A => n27482, ZN => 
                           n19516);
   U24795 : OAI21_X1 port map( B1 => n26533, B2 => n18383, A => n27482, ZN => 
                           n19517);
   U24796 : OAI21_X1 port map( B1 => n26758, B2 => n18315, A => n27486, ZN => 
                           n19571);
   U24797 : OAI21_X1 port map( B1 => n26758, B2 => n18314, A => n27486, ZN => 
                           n19570);
   U24798 : OAI21_X1 port map( B1 => n26758, B2 => n18313, A => n27486, ZN => 
                           n19573);
   U24799 : OAI21_X1 port map( B1 => n26758, B2 => n18312, A => n27486, ZN => 
                           n19572);
   U24800 : OAI21_X1 port map( B1 => n26758, B2 => n18311, A => ENABLE, ZN => 
                           n19575);
   U24801 : OAI21_X1 port map( B1 => n26758, B2 => n18310, A => n27486, ZN => 
                           n19574);
   U24802 : OAI21_X1 port map( B1 => n26758, B2 => n18309, A => ENABLE, ZN => 
                           n19577);
   U24803 : OAI21_X1 port map( B1 => n26758, B2 => n18307, A => ENABLE, ZN => 
                           n19579);
   U24804 : OAI21_X1 port map( B1 => n26758, B2 => n18306, A => ENABLE, ZN => 
                           n19576);
   U24805 : OAI21_X1 port map( B1 => n26758, B2 => n18305, A => ENABLE, ZN => 
                           n19581);
   U24806 : OAI21_X1 port map( B1 => n26758, B2 => n18304, A => ENABLE, ZN => 
                           n19578);
   U24807 : OAI21_X1 port map( B1 => n26758, B2 => n18303, A => ENABLE, ZN => 
                           n19582);
   U24808 : OAI21_X1 port map( B1 => n26535, B2 => n19437, A => n27477, ZN => 
                           n19455);
   U24809 : OAI21_X1 port map( B1 => n26535, B2 => n19420, A => n27477, ZN => 
                           n19456);
   U24810 : OAI21_X1 port map( B1 => n26535, B2 => n19403, A => n27477, ZN => 
                           n19457);
   U24811 : OAI21_X1 port map( B1 => n26535, B2 => n19386, A => n27477, ZN => 
                           n19458);
   U24812 : OAI21_X1 port map( B1 => n26535, B2 => n19369, A => n27477, ZN => 
                           n19459);
   U24813 : OAI21_X1 port map( B1 => n26535, B2 => n19352, A => n27477, ZN => 
                           n19460);
   U24814 : OAI21_X1 port map( B1 => n26535, B2 => n19335, A => n27477, ZN => 
                           n19461);
   U24815 : OAI21_X1 port map( B1 => n26535, B2 => n19318, A => n27477, ZN => 
                           n19462);
   U24816 : OAI21_X1 port map( B1 => n26535, B2 => n19301, A => n27477, ZN => 
                           n19463);
   U24817 : OAI21_X1 port map( B1 => n26535, B2 => n19284, A => n27477, ZN => 
                           n19464);
   U24818 : OAI21_X1 port map( B1 => n26535, B2 => n19267, A => n27477, ZN => 
                           n19465);
   U24819 : OAI21_X1 port map( B1 => n26535, B2 => n19250, A => n27477, ZN => 
                           n19466);
   U24820 : OAI21_X1 port map( B1 => n26535, B2 => n19233, A => n27478, ZN => 
                           n19467);
   U24821 : OAI21_X1 port map( B1 => n26534, B2 => n19216, A => n27478, ZN => 
                           n19468);
   U24822 : OAI21_X1 port map( B1 => n26534, B2 => n19199, A => n27478, ZN => 
                           n19469);
   U24823 : OAI21_X1 port map( B1 => n26534, B2 => n19182, A => n27478, ZN => 
                           n19470);
   U24824 : OAI21_X1 port map( B1 => n26534, B2 => n19165, A => n27478, ZN => 
                           n19471);
   U24825 : OAI21_X1 port map( B1 => n26534, B2 => n19148, A => n27478, ZN => 
                           n19472);
   U24826 : OAI21_X1 port map( B1 => n26534, B2 => n19131, A => n27478, ZN => 
                           n19473);
   U24827 : OAI21_X1 port map( B1 => n26534, B2 => n19114, A => n27478, ZN => 
                           n19474);
   U24828 : OAI21_X1 port map( B1 => n26534, B2 => n19097, A => n27478, ZN => 
                           n19475);
   U24829 : OAI21_X1 port map( B1 => n26534, B2 => n19080, A => n27478, ZN => 
                           n19476);
   U24830 : OAI21_X1 port map( B1 => n26534, B2 => n19063, A => n27478, ZN => 
                           n19477);
   U24831 : OAI21_X1 port map( B1 => n26534, B2 => n19046, A => n27478, ZN => 
                           n19478);
   U24832 : OAI21_X1 port map( B1 => n26534, B2 => n19029, A => n27479, ZN => 
                           n19479);
   U24833 : OAI21_X1 port map( B1 => n26534, B2 => n19012, A => n27479, ZN => 
                           n19480);
   U24834 : OAI21_X1 port map( B1 => n26534, B2 => n18995, A => n27479, ZN => 
                           n19481);
   U24835 : OAI21_X1 port map( B1 => n26533, B2 => n18978, A => n27479, ZN => 
                           n19482);
   U24836 : OAI21_X1 port map( B1 => n26535, B2 => n18961, A => n27479, ZN => 
                           n19483);
   U24837 : OAI21_X1 port map( B1 => n26534, B2 => n18944, A => n27479, ZN => 
                           n19484);
   U24838 : OAI21_X1 port map( B1 => n26533, B2 => n18927, A => n27479, ZN => 
                           n19485);
   U24839 : OAI21_X1 port map( B1 => n26535, B2 => n18910, A => n27479, ZN => 
                           n19486);
   U24840 : OAI21_X1 port map( B1 => n26534, B2 => n18893, A => n27479, ZN => 
                           n19487);
   U24841 : OAI21_X1 port map( B1 => n26533, B2 => n18876, A => n27479, ZN => 
                           n19488);
   U24842 : OAI21_X1 port map( B1 => n26535, B2 => n18859, A => n27479, ZN => 
                           n19489);
   U24843 : OAI21_X1 port map( B1 => n26534, B2 => n18842, A => n27479, ZN => 
                           n19490);
   U24844 : OAI21_X1 port map( B1 => n26533, B2 => n18825, A => n27480, ZN => 
                           n19491);
   U24845 : OAI21_X1 port map( B1 => n26535, B2 => n18808, A => n27480, ZN => 
                           n19492);
   U24846 : OAI21_X1 port map( B1 => n26534, B2 => n18791, A => n27480, ZN => 
                           n19493);
   U24847 : OAI21_X1 port map( B1 => n26535, B2 => n18774, A => n27480, ZN => 
                           n19494);
   U24848 : OAI21_X1 port map( B1 => n26534, B2 => n18757, A => n27480, ZN => 
                           n19495);
   U24849 : OAI21_X1 port map( B1 => n26534, B2 => n18740, A => n27480, ZN => 
                           n19496);
   U24850 : OAI21_X1 port map( B1 => n26533, B2 => n18723, A => n27480, ZN => 
                           n19497);
   U24851 : OAI21_X1 port map( B1 => n26535, B2 => n18706, A => n27480, ZN => 
                           n19498);
   U24852 : OAI21_X1 port map( B1 => n26534, B2 => n18689, A => n27480, ZN => 
                           n19499);
   U24853 : OAI21_X1 port map( B1 => n26533, B2 => n18672, A => n27480, ZN => 
                           n19500);
   U24854 : OAI21_X1 port map( B1 => n26533, B2 => n18655, A => n27480, ZN => 
                           n19501);
   U24855 : OAI21_X1 port map( B1 => n26535, B2 => n18638, A => n27480, ZN => 
                           n19502);
   U24856 : OAI21_X1 port map( B1 => n26534, B2 => n18621, A => n27481, ZN => 
                           n19503);
   U24857 : OAI21_X1 port map( B1 => n26535, B2 => n18604, A => n27481, ZN => 
                           n19504);
   U24858 : OAI21_X1 port map( B1 => n26533, B2 => n18587, A => n27481, ZN => 
                           n19505);
   U24859 : OAI21_X1 port map( B1 => n26535, B2 => n18570, A => n27481, ZN => 
                           n19506);
   U24860 : OAI21_X1 port map( B1 => n26760, B2 => n18366, A => n27482, ZN => 
                           n19518);
   U24861 : OAI21_X1 port map( B1 => n26758, B2 => n18365, A => n27482, ZN => 
                           n19521);
   U24862 : OAI21_X1 port map( B1 => n26759, B2 => n18364, A => n27482, ZN => 
                           n19522);
   U24863 : OAI21_X1 port map( B1 => n26760, B2 => n18363, A => n27482, ZN => 
                           n19523);
   U24864 : OAI21_X1 port map( B1 => n26758, B2 => n18362, A => n27482, ZN => 
                           n19524);
   U24865 : OAI21_X1 port map( B1 => n26759, B2 => n18361, A => n27482, ZN => 
                           n19525);
   U24866 : OAI21_X1 port map( B1 => n26760, B2 => n18360, A => n27482, ZN => 
                           n19526);
   U24867 : OAI21_X1 port map( B1 => n26758, B2 => n18359, A => n27483, ZN => 
                           n19527);
   U24868 : OAI21_X1 port map( B1 => n26759, B2 => n18358, A => n27483, ZN => 
                           n19528);
   U24869 : OAI21_X1 port map( B1 => n26760, B2 => n18357, A => n27483, ZN => 
                           n19529);
   U24870 : OAI21_X1 port map( B1 => n26758, B2 => n18356, A => n27483, ZN => 
                           n19530);
   U24871 : OAI21_X1 port map( B1 => n26760, B2 => n18355, A => n27483, ZN => 
                           n19531);
   U24872 : OAI21_X1 port map( B1 => n26760, B2 => n18354, A => n27483, ZN => 
                           n19532);
   U24873 : OAI21_X1 port map( B1 => n26760, B2 => n18353, A => n27483, ZN => 
                           n19533);
   U24874 : OAI21_X1 port map( B1 => n26760, B2 => n18352, A => n27483, ZN => 
                           n19534);
   U24875 : OAI21_X1 port map( B1 => n26760, B2 => n18351, A => n27483, ZN => 
                           n19535);
   U24876 : OAI21_X1 port map( B1 => n26760, B2 => n18350, A => n27483, ZN => 
                           n19536);
   U24877 : OAI21_X1 port map( B1 => n26760, B2 => n18349, A => n27483, ZN => 
                           n19537);
   U24878 : OAI21_X1 port map( B1 => n26760, B2 => n18348, A => n27483, ZN => 
                           n19538);
   U24879 : OAI21_X1 port map( B1 => n26760, B2 => n18347, A => n27484, ZN => 
                           n19539);
   U24880 : OAI21_X1 port map( B1 => n26760, B2 => n18346, A => n27484, ZN => 
                           n19540);
   U24881 : OAI21_X1 port map( B1 => n26760, B2 => n18345, A => n27484, ZN => 
                           n19541);
   U24882 : OAI21_X1 port map( B1 => n26760, B2 => n18344, A => n27484, ZN => 
                           n19542);
   U24883 : OAI21_X1 port map( B1 => n26760, B2 => n18343, A => n27484, ZN => 
                           n19543);
   U24884 : OAI21_X1 port map( B1 => n26759, B2 => n18342, A => n27484, ZN => 
                           n19544);
   U24885 : OAI21_X1 port map( B1 => n26760, B2 => n18341, A => n27484, ZN => 
                           n19545);
   U24886 : OAI21_X1 port map( B1 => n26760, B2 => n18340, A => n27484, ZN => 
                           n19546);
   U24887 : OAI21_X1 port map( B1 => n26758, B2 => n18339, A => n27484, ZN => 
                           n19547);
   U24888 : OAI21_X1 port map( B1 => n26759, B2 => n18338, A => n27484, ZN => 
                           n19548);
   U24889 : OAI21_X1 port map( B1 => n26759, B2 => n18337, A => n27482, ZN => 
                           n19520);
   U24890 : OAI21_X1 port map( B1 => n26758, B2 => n18336, A => n27484, ZN => 
                           n19550);
   U24891 : OAI21_X1 port map( B1 => n26760, B2 => n18335, A => n27485, ZN => 
                           n19551);
   U24892 : OAI21_X1 port map( B1 => n26760, B2 => n18334, A => n27482, ZN => 
                           n19519);
   U24893 : OAI21_X1 port map( B1 => n26758, B2 => n18333, A => n27485, ZN => 
                           n19553);
   U24894 : OAI21_X1 port map( B1 => n26759, B2 => n18332, A => n27485, ZN => 
                           n19552);
   U24895 : OAI21_X1 port map( B1 => n26759, B2 => n18331, A => n27485, ZN => 
                           n19555);
   U24896 : OAI21_X1 port map( B1 => n26760, B2 => n18330, A => n27485, ZN => 
                           n19554);
   U24897 : OAI21_X1 port map( B1 => n26759, B2 => n18329, A => n27485, ZN => 
                           n19557);
   U24898 : OAI21_X1 port map( B1 => n26758, B2 => n18328, A => n27485, ZN => 
                           n19556);
   U24899 : OAI21_X1 port map( B1 => n26759, B2 => n18327, A => n27485, ZN => 
                           n19559);
   U24900 : OAI21_X1 port map( B1 => n26759, B2 => n18326, A => n27485, ZN => 
                           n19558);
   U24901 : OAI21_X1 port map( B1 => n26759, B2 => n18325, A => n27485, ZN => 
                           n19561);
   U24902 : OAI21_X1 port map( B1 => n26759, B2 => n18324, A => n27485, ZN => 
                           n19560);
   U24903 : OAI21_X1 port map( B1 => n26759, B2 => n18323, A => n27486, ZN => 
                           n19563);
   U24904 : OAI21_X1 port map( B1 => n26759, B2 => n18322, A => n27485, ZN => 
                           n19562);
   U24905 : OAI21_X1 port map( B1 => n26759, B2 => n18321, A => n27486, ZN => 
                           n19565);
   U24906 : OAI21_X1 port map( B1 => n26759, B2 => n18320, A => n27486, ZN => 
                           n19564);
   U24907 : OAI21_X1 port map( B1 => n26759, B2 => n18319, A => n27486, ZN => 
                           n19567);
   U24908 : OAI21_X1 port map( B1 => n26759, B2 => n18318, A => n27486, ZN => 
                           n19566);
   U24909 : OAI21_X1 port map( B1 => n26759, B2 => n18317, A => n27486, ZN => 
                           n19569);
   U24910 : OAI21_X1 port map( B1 => n26759, B2 => n18316, A => n27486, ZN => 
                           n19568);
   U24911 : OAI21_X1 port map( B1 => n26759, B2 => n18308, A => n27484, ZN => 
                           n19549);
   U24912 : NOR3_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(2), A3 => ADD_WR(0)
                           , ZN => n22694);
   U24913 : NOR3_X1 port map( A1 => n20633, A2 => ADD_WR(2), A3 => n20632, ZN 
                           => n22704);
   U24914 : NOR3_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(2), A3 => n20632, 
                           ZN => n22701);
   U24915 : NOR3_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(2), A3 => n20633, 
                           ZN => n22698);
   U24916 : NOR3_X1 port map( A1 => n20643, A2 => ADD_RD2(3), A3 => n20639, ZN 
                           => n25147);
   U24917 : NOR3_X1 port map( A1 => n20638, A2 => ADD_RD1(3), A3 => n20634, ZN 
                           => n23948);
   U24918 : NOR3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(4), A3 => n20640,
                           ZN => n25153);
   U24919 : NOR3_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(4), A3 => n20635,
                           ZN => n23954);
   U24920 : NOR3_X1 port map( A1 => n20643, A2 => ADD_RD2(4), A3 => n20640, ZN 
                           => n25155);
   U24921 : NOR3_X1 port map( A1 => n20638, A2 => ADD_RD1(4), A3 => n20635, ZN 
                           => n23956);
   U24922 : NOR3_X1 port map( A1 => n20640, A2 => ADD_RD2(0), A3 => n20639, ZN 
                           => n25146);
   U24923 : NOR3_X1 port map( A1 => n20635, A2 => ADD_RD1(0), A3 => n20634, ZN 
                           => n23947);
   U24924 : NOR3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(3), A3 => n20639,
                           ZN => n25150);
   U24925 : NOR3_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(3), A3 => n20634,
                           ZN => n23951);
   U24926 : NOR3_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), A3 => 
                           ADD_RD2(0), ZN => n25163);
   U24927 : NOR3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), A3 => 
                           ADD_RD1(0), ZN => n23964);
   U24928 : AND3_X1 port map( A1 => n22717, A2 => n20631, A3 => ADD_WR(4), ZN 
                           => n22737);
   U24929 : AND3_X1 port map( A1 => ADD_WR(3), A2 => n22717, A3 => ADD_WR(4), 
                           ZN => n22754);
   U24930 : AND3_X1 port map( A1 => n22717, A2 => n20630, A3 => ADD_WR(3), ZN 
                           => n22720);
   U24931 : NOR2_X1 port map( A1 => n26536, A2 => WR, ZN => n25164);
   U24932 : NOR2_X1 port map( A1 => n26761, A2 => WR, ZN => n23965);
   U24933 : NAND2_X1 port map( A1 => WR, A2 => n26533, ZN => n24015);
   U24934 : NAND2_X1 port map( A1 => WR, A2 => n26758, ZN => n22816);
   U24935 : AND3_X1 port map( A1 => n25164, A2 => n20641, A3 => ADD_RD2(1), ZN 
                           => n25144);
   U24936 : AND3_X1 port map( A1 => n23965, A2 => n20636, A3 => ADD_RD1(1), ZN 
                           => n23945);
   U24937 : AND3_X1 port map( A1 => ADD_RD2(1), A2 => n25164, A3 => ADD_RD2(2),
                           ZN => n25148);
   U24938 : AND3_X1 port map( A1 => ADD_RD1(1), A2 => n23965, A3 => ADD_RD1(2),
                           ZN => n23949);
   U24939 : AND3_X1 port map( A1 => n25164, A2 => n20642, A3 => ADD_RD2(2), ZN 
                           => n25145);
   U24940 : AND3_X1 port map( A1 => n23965, A2 => n20637, A3 => ADD_RD1(2), ZN 
                           => n23946);
   U24941 : INV_X1 port map( A => ADD_RD2(4), ZN => n20639);
   U24942 : INV_X1 port map( A => ADD_RD1(4), ZN => n20634);
   U24943 : INV_X1 port map( A => ADD_RD2(3), ZN => n20640);
   U24944 : INV_X1 port map( A => ADD_RD1(3), ZN => n20635);
   U24945 : AND3_X1 port map( A1 => n20633, A2 => n20632, A3 => ADD_WR(2), ZN 
                           => n22707);
   U24946 : AND3_X1 port map( A1 => ADD_WR(0), A2 => n20632, A3 => ADD_WR(2), 
                           ZN => n22710);
   U24947 : AND3_X1 port map( A1 => ADD_WR(1), A2 => n20633, A3 => ADD_WR(2), 
                           ZN => n22713);
   U24948 : AND3_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(0), A3 => ADD_WR(2)
                           , ZN => n22716);
   U24949 : INV_X1 port map( A => ADD_WR(1), ZN => n20632);
   U24950 : INV_X1 port map( A => ADD_WR(0), ZN => n20633);
   U24951 : NOR2_X1 port map( A1 => RD2, A2 => n27487, ZN => n24003);
   U24952 : NOR2_X1 port map( A1 => RD1, A2 => n27487, ZN => n22804);
   U24953 : INV_X1 port map( A => ADD_RD2(0), ZN => n20643);
   U24954 : INV_X1 port map( A => ADD_RD1(0), ZN => n20638);
   U24955 : AND2_X1 port map( A1 => WR, A2 => ENABLE, ZN => n22717);
   U24956 : INV_X1 port map( A => RESET, ZN => n20626);
   U24957 : INV_X1 port map( A => DATAIN(0), ZN => n20707);
   U24958 : INV_X1 port map( A => DATAIN(1), ZN => n20706);
   U24959 : INV_X1 port map( A => DATAIN(2), ZN => n20705);
   U24960 : INV_X1 port map( A => DATAIN(3), ZN => n20704);
   U24961 : INV_X1 port map( A => DATAIN(4), ZN => n20703);
   U24962 : INV_X1 port map( A => DATAIN(5), ZN => n20702);
   U24963 : INV_X1 port map( A => DATAIN(6), ZN => n20701);
   U24964 : INV_X1 port map( A => DATAIN(7), ZN => n20700);
   U24965 : INV_X1 port map( A => DATAIN(8), ZN => n20699);
   U24966 : INV_X1 port map( A => DATAIN(9), ZN => n20698);
   U24967 : INV_X1 port map( A => DATAIN(10), ZN => n20697);
   U24968 : INV_X1 port map( A => DATAIN(11), ZN => n20696);
   U24969 : INV_X1 port map( A => DATAIN(12), ZN => n20695);
   U24970 : INV_X1 port map( A => DATAIN(13), ZN => n20694);
   U24971 : INV_X1 port map( A => DATAIN(14), ZN => n20693);
   U24972 : INV_X1 port map( A => DATAIN(15), ZN => n20692);
   U24973 : INV_X1 port map( A => DATAIN(16), ZN => n20691);
   U24974 : INV_X1 port map( A => DATAIN(17), ZN => n20690);
   U24975 : INV_X1 port map( A => DATAIN(18), ZN => n20689);
   U24976 : INV_X1 port map( A => DATAIN(19), ZN => n20688);
   U24977 : INV_X1 port map( A => DATAIN(20), ZN => n20687);
   U24978 : INV_X1 port map( A => DATAIN(21), ZN => n20686);
   U24979 : INV_X1 port map( A => DATAIN(22), ZN => n20685);
   U24980 : INV_X1 port map( A => DATAIN(23), ZN => n20684);
   U24981 : INV_X1 port map( A => DATAIN(24), ZN => n20683);
   U24982 : INV_X1 port map( A => DATAIN(25), ZN => n20682);
   U24983 : INV_X1 port map( A => DATAIN(26), ZN => n20681);
   U24984 : INV_X1 port map( A => DATAIN(27), ZN => n20680);
   U24985 : INV_X1 port map( A => DATAIN(28), ZN => n20679);
   U24986 : INV_X1 port map( A => DATAIN(29), ZN => n20678);
   U24987 : INV_X1 port map( A => DATAIN(30), ZN => n20677);
   U24988 : INV_X1 port map( A => DATAIN(31), ZN => n20676);
   U24989 : INV_X1 port map( A => DATAIN(32), ZN => n20675);
   U24990 : INV_X1 port map( A => DATAIN(33), ZN => n20674);
   U24991 : INV_X1 port map( A => DATAIN(34), ZN => n20673);
   U24992 : INV_X1 port map( A => DATAIN(35), ZN => n20672);
   U24993 : INV_X1 port map( A => DATAIN(36), ZN => n20671);
   U24994 : INV_X1 port map( A => DATAIN(37), ZN => n20670);
   U24995 : INV_X1 port map( A => DATAIN(38), ZN => n20669);
   U24996 : INV_X1 port map( A => DATAIN(39), ZN => n20668);
   U24997 : INV_X1 port map( A => DATAIN(40), ZN => n20667);
   U24998 : INV_X1 port map( A => DATAIN(41), ZN => n20666);
   U24999 : INV_X1 port map( A => DATAIN(42), ZN => n20665);
   U25000 : INV_X1 port map( A => DATAIN(43), ZN => n20664);
   U25001 : INV_X1 port map( A => DATAIN(44), ZN => n20663);
   U25002 : INV_X1 port map( A => DATAIN(45), ZN => n20662);
   U25003 : INV_X1 port map( A => DATAIN(46), ZN => n20661);
   U25004 : INV_X1 port map( A => DATAIN(47), ZN => n20660);
   U25005 : INV_X1 port map( A => DATAIN(48), ZN => n20659);
   U25006 : INV_X1 port map( A => DATAIN(49), ZN => n20658);
   U25007 : INV_X1 port map( A => DATAIN(50), ZN => n20657);
   U25008 : INV_X1 port map( A => DATAIN(51), ZN => n20656);
   U25009 : INV_X1 port map( A => DATAIN(52), ZN => n20655);
   U25010 : INV_X1 port map( A => DATAIN(53), ZN => n20654);
   U25011 : INV_X1 port map( A => DATAIN(54), ZN => n20653);
   U25012 : INV_X1 port map( A => DATAIN(55), ZN => n20652);
   U25013 : INV_X1 port map( A => DATAIN(56), ZN => n20651);
   U25014 : INV_X1 port map( A => DATAIN(57), ZN => n20650);
   U25015 : INV_X1 port map( A => DATAIN(58), ZN => n20649);
   U25016 : INV_X1 port map( A => DATAIN(59), ZN => n20648);
   U25017 : INV_X1 port map( A => DATAIN(60), ZN => n20647);
   U25018 : INV_X1 port map( A => DATAIN(61), ZN => n20646);
   U25019 : INV_X1 port map( A => DATAIN(62), ZN => n20645);
   U25020 : INV_X1 port map( A => DATAIN(63), ZN => n20644);
   U25021 : AND4_X1 port map( A1 => n25164, A2 => ADD_RD2(0), A3 => n20640, A4 
                           => n20639, ZN => n25165);
   U25022 : AND4_X1 port map( A1 => n23965, A2 => ADD_RD1(0), A3 => n20635, A4 
                           => n20634, ZN => n23966);
   U25023 : INV_X1 port map( A => ADD_RD2(2), ZN => n20641);
   U25024 : INV_X1 port map( A => ADD_RD1(2), ZN => n20636);
   U25025 : INV_X1 port map( A => ADD_RD2(1), ZN => n20642);
   U25026 : INV_X1 port map( A => ADD_RD1(1), ZN => n20637);
   U25027 : INV_X1 port map( A => ADD_WR(4), ZN => n20630);
   U25028 : INV_X1 port map( A => ADD_WR(3), ZN => n20631);
   U25029 : CLKBUF_X1 port map( A => n24019, Z => n26452);
   U25030 : CLKBUF_X1 port map( A => n24018, Z => n26458);
   U25031 : CLKBUF_X1 port map( A => n24017, Z => n26464);
   U25032 : CLKBUF_X1 port map( A => n24015, Z => n26470);
   U25033 : CLKBUF_X1 port map( A => n24014, Z => n26476);
   U25034 : CLKBUF_X1 port map( A => n24013, Z => n26482);
   U25035 : CLKBUF_X1 port map( A => n24012, Z => n26488);
   U25036 : CLKBUF_X1 port map( A => n24010, Z => n26494);
   U25037 : CLKBUF_X1 port map( A => n24009, Z => n26500);
   U25038 : CLKBUF_X1 port map( A => n24008, Z => n26506);
   U25039 : CLKBUF_X1 port map( A => n24007, Z => n26512);
   U25040 : CLKBUF_X1 port map( A => n24005, Z => n26518);
   U25041 : CLKBUF_X1 port map( A => n24004, Z => n26524);
   U25042 : CLKBUF_X1 port map( A => n24002, Z => n26557);
   U25043 : CLKBUF_X1 port map( A => n24000, Z => n26563);
   U25044 : CLKBUF_X1 port map( A => n23999, Z => n26569);
   U25045 : CLKBUF_X1 port map( A => n23994, Z => n26575);
   U25046 : CLKBUF_X1 port map( A => n23993, Z => n26581);
   U25047 : CLKBUF_X1 port map( A => n23992, Z => n26587);
   U25048 : CLKBUF_X1 port map( A => n23990, Z => n26593);
   U25049 : CLKBUF_X1 port map( A => n23989, Z => n26599);
   U25050 : CLKBUF_X1 port map( A => n23988, Z => n26605);
   U25051 : CLKBUF_X1 port map( A => n23987, Z => n26611);
   U25052 : CLKBUF_X1 port map( A => n23985, Z => n26617);
   U25053 : CLKBUF_X1 port map( A => n23984, Z => n26623);
   U25054 : CLKBUF_X1 port map( A => n23983, Z => n26629);
   U25055 : CLKBUF_X1 port map( A => n23982, Z => n26635);
   U25056 : CLKBUF_X1 port map( A => n23980, Z => n26641);
   U25057 : CLKBUF_X1 port map( A => n23979, Z => n26647);
   U25058 : CLKBUF_X1 port map( A => n23978, Z => n26653);
   U25059 : CLKBUF_X1 port map( A => n23977, Z => n26659);
   U25060 : CLKBUF_X1 port map( A => n23975, Z => n26665);
   U25061 : CLKBUF_X1 port map( A => n23974, Z => n26671);
   U25062 : CLKBUF_X1 port map( A => n22820, Z => n26677);
   U25063 : CLKBUF_X1 port map( A => n22819, Z => n26683);
   U25064 : CLKBUF_X1 port map( A => n22818, Z => n26689);
   U25065 : CLKBUF_X1 port map( A => n22816, Z => n26695);
   U25066 : CLKBUF_X1 port map( A => n22815, Z => n26701);
   U25067 : CLKBUF_X1 port map( A => n22814, Z => n26707);
   U25068 : CLKBUF_X1 port map( A => n22813, Z => n26713);
   U25069 : CLKBUF_X1 port map( A => n22811, Z => n26719);
   U25070 : CLKBUF_X1 port map( A => n22810, Z => n26725);
   U25071 : CLKBUF_X1 port map( A => n22809, Z => n26731);
   U25072 : CLKBUF_X1 port map( A => n22808, Z => n26737);
   U25073 : CLKBUF_X1 port map( A => n22806, Z => n26743);
   U25074 : CLKBUF_X1 port map( A => n22805, Z => n26749);
   U25075 : CLKBUF_X1 port map( A => n22803, Z => n26782);
   U25076 : CLKBUF_X1 port map( A => n22801, Z => n26788);
   U25077 : CLKBUF_X1 port map( A => n22800, Z => n26794);
   U25078 : CLKBUF_X1 port map( A => n22795, Z => n26800);
   U25079 : CLKBUF_X1 port map( A => n22794, Z => n26806);
   U25080 : CLKBUF_X1 port map( A => n22793, Z => n26812);
   U25081 : CLKBUF_X1 port map( A => n22791, Z => n26818);
   U25082 : CLKBUF_X1 port map( A => n22790, Z => n26824);
   U25083 : CLKBUF_X1 port map( A => n22789, Z => n26830);
   U25084 : CLKBUF_X1 port map( A => n22788, Z => n26836);
   U25085 : CLKBUF_X1 port map( A => n22786, Z => n26842);
   U25086 : CLKBUF_X1 port map( A => n22785, Z => n26848);
   U25087 : CLKBUF_X1 port map( A => n22784, Z => n26854);
   U25088 : CLKBUF_X1 port map( A => n22783, Z => n26860);
   U25089 : CLKBUF_X1 port map( A => n22781, Z => n26866);
   U25090 : CLKBUF_X1 port map( A => n22780, Z => n26872);
   U25091 : CLKBUF_X1 port map( A => n22779, Z => n26878);
   U25092 : CLKBUF_X1 port map( A => n22778, Z => n26884);
   U25093 : CLKBUF_X1 port map( A => n22776, Z => n26890);
   U25094 : CLKBUF_X1 port map( A => n22775, Z => n26896);
   U25095 : CLKBUF_X1 port map( A => n22768, Z => n26902);
   U25096 : CLKBUF_X1 port map( A => n22767, Z => n26908);
   U25097 : CLKBUF_X1 port map( A => n22766, Z => n26914);
   U25098 : CLKBUF_X1 port map( A => n22765, Z => n26920);
   U25099 : CLKBUF_X1 port map( A => n22764, Z => n26926);
   U25100 : CLKBUF_X1 port map( A => n22763, Z => n26932);
   U25101 : CLKBUF_X1 port map( A => n22762, Z => n26938);
   U25102 : CLKBUF_X1 port map( A => n22761, Z => n26944);
   U25103 : CLKBUF_X1 port map( A => n22760, Z => n26950);
   U25104 : CLKBUF_X1 port map( A => n22759, Z => n26956);
   U25105 : CLKBUF_X1 port map( A => n22758, Z => n26962);
   U25106 : CLKBUF_X1 port map( A => n22757, Z => n26968);
   U25107 : CLKBUF_X1 port map( A => n22756, Z => n26974);
   U25108 : CLKBUF_X1 port map( A => n22755, Z => n26980);
   U25109 : CLKBUF_X1 port map( A => n22753, Z => n26986);
   U25110 : CLKBUF_X1 port map( A => n22752, Z => n26992);
   U25111 : CLKBUF_X1 port map( A => n22751, Z => n26998);
   U25112 : CLKBUF_X1 port map( A => n22750, Z => n27004);
   U25113 : CLKBUF_X1 port map( A => n22749, Z => n27010);
   U25114 : CLKBUF_X1 port map( A => n22748, Z => n27016);
   U25115 : CLKBUF_X1 port map( A => n22747, Z => n27022);
   U25116 : CLKBUF_X1 port map( A => n22746, Z => n27028);
   U25117 : CLKBUF_X1 port map( A => n22745, Z => n27034);
   U25118 : CLKBUF_X1 port map( A => n22744, Z => n27040);
   U25119 : CLKBUF_X1 port map( A => n22743, Z => n27046);
   U25120 : CLKBUF_X1 port map( A => n22742, Z => n27052);
   U25121 : CLKBUF_X1 port map( A => n22741, Z => n27058);
   U25122 : CLKBUF_X1 port map( A => n22740, Z => n27064);
   U25123 : CLKBUF_X1 port map( A => n22739, Z => n27070);
   U25124 : CLKBUF_X1 port map( A => n22738, Z => n27076);
   U25125 : CLKBUF_X1 port map( A => n22736, Z => n27082);
   U25126 : CLKBUF_X1 port map( A => n22735, Z => n27088);
   U25127 : CLKBUF_X1 port map( A => n22734, Z => n27094);
   U25128 : CLKBUF_X1 port map( A => n22733, Z => n27100);
   U25129 : CLKBUF_X1 port map( A => n22732, Z => n27106);
   U25130 : CLKBUF_X1 port map( A => n22731, Z => n27112);
   U25131 : CLKBUF_X1 port map( A => n22730, Z => n27118);
   U25132 : CLKBUF_X1 port map( A => n22729, Z => n27124);
   U25133 : CLKBUF_X1 port map( A => n22728, Z => n27130);
   U25134 : CLKBUF_X1 port map( A => n22727, Z => n27136);
   U25135 : CLKBUF_X1 port map( A => n22726, Z => n27142);
   U25136 : CLKBUF_X1 port map( A => n22725, Z => n27148);
   U25137 : CLKBUF_X1 port map( A => n22724, Z => n27154);
   U25138 : CLKBUF_X1 port map( A => n22723, Z => n27160);
   U25139 : CLKBUF_X1 port map( A => n22722, Z => n27166);
   U25140 : CLKBUF_X1 port map( A => n22721, Z => n27172);
   U25141 : CLKBUF_X1 port map( A => n22719, Z => n27178);
   U25142 : CLKBUF_X1 port map( A => n22718, Z => n27184);
   U25143 : CLKBUF_X1 port map( A => n22715, Z => n27190);
   U25144 : CLKBUF_X1 port map( A => n22714, Z => n27196);
   U25145 : CLKBUF_X1 port map( A => n22712, Z => n27202);
   U25146 : CLKBUF_X1 port map( A => n22711, Z => n27208);
   U25147 : CLKBUF_X1 port map( A => n22709, Z => n27214);
   U25148 : CLKBUF_X1 port map( A => n22708, Z => n27220);
   U25149 : CLKBUF_X1 port map( A => n22706, Z => n27226);
   U25150 : CLKBUF_X1 port map( A => n22705, Z => n27232);
   U25151 : CLKBUF_X1 port map( A => n22703, Z => n27238);
   U25152 : CLKBUF_X1 port map( A => n22702, Z => n27244);
   U25153 : CLKBUF_X1 port map( A => n22700, Z => n27250);
   U25154 : CLKBUF_X1 port map( A => n22699, Z => n27256);
   U25155 : CLKBUF_X1 port map( A => n22697, Z => n27262);
   U25156 : CLKBUF_X1 port map( A => n22696, Z => n27268);
   U25157 : CLKBUF_X1 port map( A => n22693, Z => n27274);
   U25158 : INV_X1 port map( A => ENABLE, ZN => n27487);

end SYN_beh;
