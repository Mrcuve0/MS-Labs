
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_Booth is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_Booth;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_959 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_959;

architecture SYN_BEHAVIORAL of FA_959 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net90527, n2, n4, n5 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => Ci, B2 => n4, A => n5, ZN => n2);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : OR2_X1 port map( A1 => B, A2 => A, ZN => n4);
   U5 : XNOR2_X1 port map( A => Ci, B => net90527, ZN => S);
   U6 : XNOR2_X1 port map( A => B, B => A, ZN => net90527);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_958 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_958;

architecture SYN_BEHAVIORAL of FA_958 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net121879, net121878, n4 : std_logic;

begin
   
   U1 : NOR2_X1 port map( A1 => A, A2 => B, ZN => net121878);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U4 : AOI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => net121879);
   U5 : NOR2_X1 port map( A1 => net121879, A2 => net121878, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_957 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_957;

architecture SYN_BEHAVIORAL of FA_957 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U5 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_956 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_956;

architecture SYN_BEHAVIORAL of FA_956 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_955 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_955;

architecture SYN_BEHAVIORAL of FA_955 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_954 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_954;

architecture SYN_BEHAVIORAL of FA_954 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_953 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_953;

architecture SYN_BEHAVIORAL of FA_953 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_952 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_952;

architecture SYN_BEHAVIORAL of FA_952 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_951 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_951;

architecture SYN_BEHAVIORAL of FA_951 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_950 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_950;

architecture SYN_BEHAVIORAL of FA_950 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_949 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_949;

architecture SYN_BEHAVIORAL of FA_949 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_948 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_948;

architecture SYN_BEHAVIORAL of FA_948 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_947 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_947;

architecture SYN_BEHAVIORAL of FA_947 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_946 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_946;

architecture SYN_BEHAVIORAL of FA_946 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_945 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_945;

architecture SYN_BEHAVIORAL of FA_945 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U2 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U4 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_944 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_944;

architecture SYN_BEHAVIORAL of FA_944 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_943 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_943;

architecture SYN_BEHAVIORAL of FA_943 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_942 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_942;

architecture SYN_BEHAVIORAL of FA_942 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_941 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_941;

architecture SYN_BEHAVIORAL of FA_941 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_940 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_940;

architecture SYN_BEHAVIORAL of FA_940 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_939 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_939;

architecture SYN_BEHAVIORAL of FA_939 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_938 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_938;

architecture SYN_BEHAVIORAL of FA_938 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_937 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_937;

architecture SYN_BEHAVIORAL of FA_937 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_936 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_936;

architecture SYN_BEHAVIORAL of FA_936 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_935 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_935;

architecture SYN_BEHAVIORAL of FA_935 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_934 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_934;

architecture SYN_BEHAVIORAL of FA_934 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_933 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_933;

architecture SYN_BEHAVIORAL of FA_933 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_932 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_932;

architecture SYN_BEHAVIORAL of FA_932 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_931 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_931;

architecture SYN_BEHAVIORAL of FA_931 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_930 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_930;

architecture SYN_BEHAVIORAL of FA_930 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U2 : INV_X1 port map( A => n6, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_929 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_929;

architecture SYN_BEHAVIORAL of FA_929 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_928 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_928;

architecture SYN_BEHAVIORAL of FA_928 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_927 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_927;

architecture SYN_BEHAVIORAL of FA_927 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_926 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_926;

architecture SYN_BEHAVIORAL of FA_926 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_925 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_925;

architecture SYN_BEHAVIORAL of FA_925 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U2 : INV_X1 port map( A => n6, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_924 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_924;

architecture SYN_BEHAVIORAL of FA_924 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_923 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_923;

architecture SYN_BEHAVIORAL of FA_923 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_922 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_922;

architecture SYN_BEHAVIORAL of FA_922 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_921 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_921;

architecture SYN_BEHAVIORAL of FA_921 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_920 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_920;

architecture SYN_BEHAVIORAL of FA_920 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_919 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_919;

architecture SYN_BEHAVIORAL of FA_919 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_918 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_918;

architecture SYN_BEHAVIORAL of FA_918 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_917 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_917;

architecture SYN_BEHAVIORAL of FA_917 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_916 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_916;

architecture SYN_BEHAVIORAL of FA_916 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_915 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_915;

architecture SYN_BEHAVIORAL of FA_915 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_914 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_914;

architecture SYN_BEHAVIORAL of FA_914 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_913 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_913;

architecture SYN_BEHAVIORAL of FA_913 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_912 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_912;

architecture SYN_BEHAVIORAL of FA_912 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_911 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_911;

architecture SYN_BEHAVIORAL of FA_911 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_910 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_910;

architecture SYN_BEHAVIORAL of FA_910 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_909 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_909;

architecture SYN_BEHAVIORAL of FA_909 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_908 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_908;

architecture SYN_BEHAVIORAL of FA_908 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : INV_X1 port map( A => n6, ZN => n4);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_907 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_907;

architecture SYN_BEHAVIORAL of FA_907 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_906 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_906;

architecture SYN_BEHAVIORAL of FA_906 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_905 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_905;

architecture SYN_BEHAVIORAL of FA_905 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_904 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_904;

architecture SYN_BEHAVIORAL of FA_904 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_903 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_903;

architecture SYN_BEHAVIORAL of FA_903 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_902 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_902;

architecture SYN_BEHAVIORAL of FA_902 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_901 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_901;

architecture SYN_BEHAVIORAL of FA_901 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_900 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_900;

architecture SYN_BEHAVIORAL of FA_900 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_899 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_899;

architecture SYN_BEHAVIORAL of FA_899 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_898 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_898;

architecture SYN_BEHAVIORAL of FA_898 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_897 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_897;

architecture SYN_BEHAVIORAL of FA_897 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_896 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_896;

architecture SYN_BEHAVIORAL of FA_896 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, net90553, n4 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => Ci, ZN => net90553);
   U2 : XNOR2_X1 port map( A => net90553, B => n4, ZN => S);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n2);
   U5 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_895 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_895;

architecture SYN_BEHAVIORAL of FA_895 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : AOI21_X1 port map( B1 => A, B2 => n7, A => Ci, ZN => n5);
   U4 : NOR2_X1 port map( A1 => A, A2 => n7, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : NOR2_X1 port map( A1 => n5, A2 => n4, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_894 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_894;

architecture SYN_BEHAVIORAL of FA_894 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U3 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n5, B2 => Ci, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_893 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_893;

architecture SYN_BEHAVIORAL of FA_893 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U2 : XNOR2_X1 port map( A => n5, B => Ci, ZN => S);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n5);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n4, B2 => Ci, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_892 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_892;

architecture SYN_BEHAVIORAL of FA_892 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_891 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_891;

architecture SYN_BEHAVIORAL of FA_891 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_890 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_890;

architecture SYN_BEHAVIORAL of FA_890 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_889 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_889;

architecture SYN_BEHAVIORAL of FA_889 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_888 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_888;

architecture SYN_BEHAVIORAL of FA_888 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => A, A2 => B, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_887 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_887;

architecture SYN_BEHAVIORAL of FA_887 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_886 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_886;

architecture SYN_BEHAVIORAL of FA_886 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_885 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_885;

architecture SYN_BEHAVIORAL of FA_885 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_884 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_884;

architecture SYN_BEHAVIORAL of FA_884 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_883 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_883;

architecture SYN_BEHAVIORAL of FA_883 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_882 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_882;

architecture SYN_BEHAVIORAL of FA_882 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_881 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_881;

architecture SYN_BEHAVIORAL of FA_881 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_880 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_880;

architecture SYN_BEHAVIORAL of FA_880 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_879 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_879;

architecture SYN_BEHAVIORAL of FA_879 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_878 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_878;

architecture SYN_BEHAVIORAL of FA_878 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_877 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_877;

architecture SYN_BEHAVIORAL of FA_877 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n8);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n9, ZN => Co);
   U7 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_876 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_876;

architecture SYN_BEHAVIORAL of FA_876 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_875 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_875;

architecture SYN_BEHAVIORAL of FA_875 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_874 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_874;

architecture SYN_BEHAVIORAL of FA_874 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_873 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_873;

architecture SYN_BEHAVIORAL of FA_873 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_872 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_872;

architecture SYN_BEHAVIORAL of FA_872 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_871 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_871;

architecture SYN_BEHAVIORAL of FA_871 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_870 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_870;

architecture SYN_BEHAVIORAL of FA_870 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_869 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_869;

architecture SYN_BEHAVIORAL of FA_869 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_868 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_868;

architecture SYN_BEHAVIORAL of FA_868 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_867 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_867;

architecture SYN_BEHAVIORAL of FA_867 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_866 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_866;

architecture SYN_BEHAVIORAL of FA_866 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_865 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_865;

architecture SYN_BEHAVIORAL of FA_865 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_864 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_864;

architecture SYN_BEHAVIORAL of FA_864 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_863 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_863;

architecture SYN_BEHAVIORAL of FA_863 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_862 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_862;

architecture SYN_BEHAVIORAL of FA_862 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_861 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_861;

architecture SYN_BEHAVIORAL of FA_861 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_860 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_860;

architecture SYN_BEHAVIORAL of FA_860 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_859 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_859;

architecture SYN_BEHAVIORAL of FA_859 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_858 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_858;

architecture SYN_BEHAVIORAL of FA_858 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_857 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_857;

architecture SYN_BEHAVIORAL of FA_857 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_856 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_856;

architecture SYN_BEHAVIORAL of FA_856 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_855 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_855;

architecture SYN_BEHAVIORAL of FA_855 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_854 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_854;

architecture SYN_BEHAVIORAL of FA_854 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_853 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_853;

architecture SYN_BEHAVIORAL of FA_853 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_852 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_852;

architecture SYN_BEHAVIORAL of FA_852 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_851 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_851;

architecture SYN_BEHAVIORAL of FA_851 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_850 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_850;

architecture SYN_BEHAVIORAL of FA_850 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_849 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_849;

architecture SYN_BEHAVIORAL of FA_849 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_848 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_848;

architecture SYN_BEHAVIORAL of FA_848 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_847 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_847;

architecture SYN_BEHAVIORAL of FA_847 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_846 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_846;

architecture SYN_BEHAVIORAL of FA_846 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_845 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_845;

architecture SYN_BEHAVIORAL of FA_845 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_844 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_844;

architecture SYN_BEHAVIORAL of FA_844 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_843 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_843;

architecture SYN_BEHAVIORAL of FA_843 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_842 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_842;

architecture SYN_BEHAVIORAL of FA_842 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_841 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_841;

architecture SYN_BEHAVIORAL of FA_841 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_840 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_840;

architecture SYN_BEHAVIORAL of FA_840 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_839 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_839;

architecture SYN_BEHAVIORAL of FA_839 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_838 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_838;

architecture SYN_BEHAVIORAL of FA_838 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_837 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_837;

architecture SYN_BEHAVIORAL of FA_837 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_836 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_836;

architecture SYN_BEHAVIORAL of FA_836 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_835 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_835;

architecture SYN_BEHAVIORAL of FA_835 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_834 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_834;

architecture SYN_BEHAVIORAL of FA_834 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_833 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_833;

architecture SYN_BEHAVIORAL of FA_833 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U4 : XNOR2_X1 port map( A => n5, B => B, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => n4, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_832 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_832;

architecture SYN_BEHAVIORAL of FA_832 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, net90513, n4 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : INV_X1 port map( A => Ci, ZN => net90513);
   U2 : XNOR2_X1 port map( A => net90513, B => n4, ZN => S);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n2);
   U5 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_831 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_831;

architecture SYN_BEHAVIORAL of FA_831 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n6, B2 => Ci, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_830 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_830;

architecture SYN_BEHAVIORAL of FA_830 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n4, B2 => Ci, ZN => n2);
   U2 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_829 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_829;

architecture SYN_BEHAVIORAL of FA_829 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n4, B2 => Ci, ZN => n2);
   U2 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_828 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_828;

architecture SYN_BEHAVIORAL of FA_828 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_827 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_827;

architecture SYN_BEHAVIORAL of FA_827 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_826 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_826;

architecture SYN_BEHAVIORAL of FA_826 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_825 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_825;

architecture SYN_BEHAVIORAL of FA_825 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_824 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_824;

architecture SYN_BEHAVIORAL of FA_824 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_823 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_823;

architecture SYN_BEHAVIORAL of FA_823 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_822 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_822;

architecture SYN_BEHAVIORAL of FA_822 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : AOI22_X1 port map( A1 => A, A2 => n4, B1 => Ci, B2 => n6, ZN => n5);
   U5 : INV_X1 port map( A => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_821 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_821;

architecture SYN_BEHAVIORAL of FA_821 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U3 : CLKBUF_X1 port map( A => B, Z => n5);
   U4 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_820 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_820;

architecture SYN_BEHAVIORAL of FA_820 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_819 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_819;

architecture SYN_BEHAVIORAL of FA_819 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n7);
   U4 : AOI22_X1 port map( A1 => A, A2 => n4, B1 => Ci, B2 => n6, ZN => n5);
   U5 : INV_X1 port map( A => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_818 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_818;

architecture SYN_BEHAVIORAL of FA_818 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_817 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_817;

architecture SYN_BEHAVIORAL of FA_817 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_816 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_816;

architecture SYN_BEHAVIORAL of FA_816 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_815 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_815;

architecture SYN_BEHAVIORAL of FA_815 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_814 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_814;

architecture SYN_BEHAVIORAL of FA_814 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_813 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_813;

architecture SYN_BEHAVIORAL of FA_813 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U3 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n6, B2 => Ci, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_812 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_812;

architecture SYN_BEHAVIORAL of FA_812 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_811 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_811;

architecture SYN_BEHAVIORAL of FA_811 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_810 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_810;

architecture SYN_BEHAVIORAL of FA_810 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_809 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_809;

architecture SYN_BEHAVIORAL of FA_809 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_808 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_808;

architecture SYN_BEHAVIORAL of FA_808 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n6, B2 => Ci, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_807 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_807;

architecture SYN_BEHAVIORAL of FA_807 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_806 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_806;

architecture SYN_BEHAVIORAL of FA_806 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_805 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_805;

architecture SYN_BEHAVIORAL of FA_805 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_804 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_804;

architecture SYN_BEHAVIORAL of FA_804 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_803 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_803;

architecture SYN_BEHAVIORAL of FA_803 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_802 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_802;

architecture SYN_BEHAVIORAL of FA_802 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_801 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_801;

architecture SYN_BEHAVIORAL of FA_801 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : AOI22_X1 port map( A1 => A, A2 => B, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_800 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_800;

architecture SYN_BEHAVIORAL of FA_800 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_799 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_799;

architecture SYN_BEHAVIORAL of FA_799 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_798 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_798;

architecture SYN_BEHAVIORAL of FA_798 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_797 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_797;

architecture SYN_BEHAVIORAL of FA_797 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_796 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_796;

architecture SYN_BEHAVIORAL of FA_796 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n8 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U3 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);
   U4 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_795 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_795;

architecture SYN_BEHAVIORAL of FA_795 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_794 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_794;

architecture SYN_BEHAVIORAL of FA_794 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_793 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_793;

architecture SYN_BEHAVIORAL of FA_793 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_792 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_792;

architecture SYN_BEHAVIORAL of FA_792 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_791 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_791;

architecture SYN_BEHAVIORAL of FA_791 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_790 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_790;

architecture SYN_BEHAVIORAL of FA_790 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_789 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_789;

architecture SYN_BEHAVIORAL of FA_789 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_788 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_788;

architecture SYN_BEHAVIORAL of FA_788 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_787 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_787;

architecture SYN_BEHAVIORAL of FA_787 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_786 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_786;

architecture SYN_BEHAVIORAL of FA_786 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_785 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_785;

architecture SYN_BEHAVIORAL of FA_785 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_784 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_784;

architecture SYN_BEHAVIORAL of FA_784 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n6, B2 => Ci, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_783 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_783;

architecture SYN_BEHAVIORAL of FA_783 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_782 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_782;

architecture SYN_BEHAVIORAL of FA_782 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_781 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_781;

architecture SYN_BEHAVIORAL of FA_781 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => A, A2 => B, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_780 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_780;

architecture SYN_BEHAVIORAL of FA_780 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_779 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_779;

architecture SYN_BEHAVIORAL of FA_779 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_778 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_778;

architecture SYN_BEHAVIORAL of FA_778 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n6, B2 => Ci, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_777 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_777;

architecture SYN_BEHAVIORAL of FA_777 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_776 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_776;

architecture SYN_BEHAVIORAL of FA_776 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_775 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_775;

architecture SYN_BEHAVIORAL of FA_775 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_774 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_774;

architecture SYN_BEHAVIORAL of FA_774 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_773 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_773;

architecture SYN_BEHAVIORAL of FA_773 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_772 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_772;

architecture SYN_BEHAVIORAL of FA_772 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_771 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_771;

architecture SYN_BEHAVIORAL of FA_771 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_770 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_770;

architecture SYN_BEHAVIORAL of FA_770 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n6, B2 => Ci, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_769 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_769;

architecture SYN_BEHAVIORAL of FA_769 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : CLKBUF_X1 port map( A => n7, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U4 : XNOR2_X1 port map( A => n5, B => B, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_768 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_768;

architecture SYN_BEHAVIORAL of FA_768 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => Ci, ZN => n5);
   U2 : INV_X1 port map( A => A, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : XNOR2_X1 port map( A => n7, B => n5, ZN => S);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_767 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_767;

architecture SYN_BEHAVIORAL of FA_767 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_766 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_766;

architecture SYN_BEHAVIORAL of FA_766 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n4, B2 => Ci, ZN => n2);
   U4 : INV_X1 port map( A => A, ZN => n5);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_765 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_765;

architecture SYN_BEHAVIORAL of FA_765 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n4, B2 => Ci, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_764 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_764;

architecture SYN_BEHAVIORAL of FA_764 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_763 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_763;

architecture SYN_BEHAVIORAL of FA_763 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_762 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_762;

architecture SYN_BEHAVIORAL of FA_762 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_761 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_761;

architecture SYN_BEHAVIORAL of FA_761 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_760 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_760;

architecture SYN_BEHAVIORAL of FA_760 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => A, A2 => n4, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_759 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_759;

architecture SYN_BEHAVIORAL of FA_759 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_758 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_758;

architecture SYN_BEHAVIORAL of FA_758 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => A, A2 => n4, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_757 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_757;

architecture SYN_BEHAVIORAL of FA_757 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_756 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_756;

architecture SYN_BEHAVIORAL of FA_756 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => A, A2 => n4, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_755 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_755;

architecture SYN_BEHAVIORAL of FA_755 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_754 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_754;

architecture SYN_BEHAVIORAL of FA_754 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_753 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_753;

architecture SYN_BEHAVIORAL of FA_753 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_752 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_752;

architecture SYN_BEHAVIORAL of FA_752 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => A, A2 => n4, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_751 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_751;

architecture SYN_BEHAVIORAL of FA_751 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_750 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_750;

architecture SYN_BEHAVIORAL of FA_750 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_749 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_749;

architecture SYN_BEHAVIORAL of FA_749 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_748 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_748;

architecture SYN_BEHAVIORAL of FA_748 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_747 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_747;

architecture SYN_BEHAVIORAL of FA_747 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_746 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_746;

architecture SYN_BEHAVIORAL of FA_746 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_745 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_745;

architecture SYN_BEHAVIORAL of FA_745 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_744 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_744;

architecture SYN_BEHAVIORAL of FA_744 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_743 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_743;

architecture SYN_BEHAVIORAL of FA_743 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_742 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_742;

architecture SYN_BEHAVIORAL of FA_742 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_741 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_741;

architecture SYN_BEHAVIORAL of FA_741 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => A, A2 => n4, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_740 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_740;

architecture SYN_BEHAVIORAL of FA_740 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_739 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_739;

architecture SYN_BEHAVIORAL of FA_739 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_738 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_738;

architecture SYN_BEHAVIORAL of FA_738 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_737 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_737;

architecture SYN_BEHAVIORAL of FA_737 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_736 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_736;

architecture SYN_BEHAVIORAL of FA_736 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_735 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_735;

architecture SYN_BEHAVIORAL of FA_735 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_734 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_734;

architecture SYN_BEHAVIORAL of FA_734 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_733 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_733;

architecture SYN_BEHAVIORAL of FA_733 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_732 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_732;

architecture SYN_BEHAVIORAL of FA_732 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_731 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_731;

architecture SYN_BEHAVIORAL of FA_731 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_730 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_730;

architecture SYN_BEHAVIORAL of FA_730 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => A, A2 => n4, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_729 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_729;

architecture SYN_BEHAVIORAL of FA_729 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => A, A2 => n4, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_728 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_728;

architecture SYN_BEHAVIORAL of FA_728 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_727 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_727;

architecture SYN_BEHAVIORAL of FA_727 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_726 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_726;

architecture SYN_BEHAVIORAL of FA_726 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_725 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_725;

architecture SYN_BEHAVIORAL of FA_725 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => A, A2 => n4, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_724 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_724;

architecture SYN_BEHAVIORAL of FA_724 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => A, A2 => n4, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_723 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_723;

architecture SYN_BEHAVIORAL of FA_723 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_722 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_722;

architecture SYN_BEHAVIORAL of FA_722 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n8, n9 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : XOR2_X1 port map( A => n5, B => B, Z => n4);
   U3 : INV_X1 port map( A => A, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n8);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n9, ZN => Co);
   U7 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n8, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_721 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_721;

architecture SYN_BEHAVIORAL of FA_721 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_720 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_720;

architecture SYN_BEHAVIORAL of FA_720 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_719 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_719;

architecture SYN_BEHAVIORAL of FA_719 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n10 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => n4);
   U2 : INV_X1 port map( A => A, ZN => n7);
   U3 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : XNOR2_X1 port map( A => Ci, B => n5, ZN => S);
   U5 : XNOR2_X1 port map( A => n7, B => B, ZN => n6);
   U6 : CLKBUF_X1 port map( A => B, Z => n8);
   U7 : INV_X1 port map( A => n10, ZN => Co);
   U8 : AOI22_X1 port map( A1 => n8, A2 => A, B1 => n6, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_718 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_718;

architecture SYN_BEHAVIORAL of FA_718 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_717 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_717;

architecture SYN_BEHAVIORAL of FA_717 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_716 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_716;

architecture SYN_BEHAVIORAL of FA_716 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_715 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_715;

architecture SYN_BEHAVIORAL of FA_715 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_714 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_714;

architecture SYN_BEHAVIORAL of FA_714 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_713 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_713;

architecture SYN_BEHAVIORAL of FA_713 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_712 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_712;

architecture SYN_BEHAVIORAL of FA_712 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_711 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_711;

architecture SYN_BEHAVIORAL of FA_711 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_710 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_710;

architecture SYN_BEHAVIORAL of FA_710 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => A, A2 => n4, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_709 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_709;

architecture SYN_BEHAVIORAL of FA_709 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_708 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_708;

architecture SYN_BEHAVIORAL of FA_708 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_707 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_707;

architecture SYN_BEHAVIORAL of FA_707 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_706 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_706;

architecture SYN_BEHAVIORAL of FA_706 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_705 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_705;

architecture SYN_BEHAVIORAL of FA_705 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n8, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n8);
   U4 : CLKBUF_X1 port map( A => n8, Z => n5);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n9, ZN => Co);
   U7 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n5, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_704 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_704;

architecture SYN_BEHAVIORAL of FA_704 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : INV_X1 port map( A => Ci, ZN => n4);
   U3 : XNOR2_X1 port map( A => n4, B => n7, ZN => S);
   U4 : XNOR2_X1 port map( A => n5, B => B, ZN => n7);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_703 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_703;

architecture SYN_BEHAVIORAL of FA_703 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : XNOR2_X1 port map( A => B, B => n6, ZN => n4);
   U4 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n4, B2 => Ci, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_702 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_702;

architecture SYN_BEHAVIORAL of FA_702 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n4, B2 => Ci, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_701 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_701;

architecture SYN_BEHAVIORAL of FA_701 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n4, B2 => Ci, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_700 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_700;

architecture SYN_BEHAVIORAL of FA_700 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n4, B2 => Ci, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_699 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_699;

architecture SYN_BEHAVIORAL of FA_699 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_698 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_698;

architecture SYN_BEHAVIORAL of FA_698 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_697 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_697;

architecture SYN_BEHAVIORAL of FA_697 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_696 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_696;

architecture SYN_BEHAVIORAL of FA_696 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_695 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_695;

architecture SYN_BEHAVIORAL of FA_695 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_694 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_694;

architecture SYN_BEHAVIORAL of FA_694 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_693 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_693;

architecture SYN_BEHAVIORAL of FA_693 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_692 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_692;

architecture SYN_BEHAVIORAL of FA_692 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_691 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_691;

architecture SYN_BEHAVIORAL of FA_691 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_690 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_690;

architecture SYN_BEHAVIORAL of FA_690 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_689 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_689;

architecture SYN_BEHAVIORAL of FA_689 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U3 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_688 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_688;

architecture SYN_BEHAVIORAL of FA_688 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_687 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_687;

architecture SYN_BEHAVIORAL of FA_687 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_686 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_686;

architecture SYN_BEHAVIORAL of FA_686 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_685 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_685;

architecture SYN_BEHAVIORAL of FA_685 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => A, A2 => n4, B1 => n7, B2 => Ci, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_684 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_684;

architecture SYN_BEHAVIORAL of FA_684 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_683 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_683;

architecture SYN_BEHAVIORAL of FA_683 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => A, A2 => n4, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_682 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_682;

architecture SYN_BEHAVIORAL of FA_682 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_681 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_681;

architecture SYN_BEHAVIORAL of FA_681 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_680 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_680;

architecture SYN_BEHAVIORAL of FA_680 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => A, A2 => n4, B1 => n7, B2 => Ci, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_679 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_679;

architecture SYN_BEHAVIORAL of FA_679 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_678 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_678;

architecture SYN_BEHAVIORAL of FA_678 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_677 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_677;

architecture SYN_BEHAVIORAL of FA_677 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_676 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_676;

architecture SYN_BEHAVIORAL of FA_676 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_675 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_675;

architecture SYN_BEHAVIORAL of FA_675 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_674 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_674;

architecture SYN_BEHAVIORAL of FA_674 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_673 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_673;

architecture SYN_BEHAVIORAL of FA_673 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_672 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_672;

architecture SYN_BEHAVIORAL of FA_672 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_671 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_671;

architecture SYN_BEHAVIORAL of FA_671 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_670 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_670;

architecture SYN_BEHAVIORAL of FA_670 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_669 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_669;

architecture SYN_BEHAVIORAL of FA_669 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_668 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_668;

architecture SYN_BEHAVIORAL of FA_668 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_667 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_667;

architecture SYN_BEHAVIORAL of FA_667 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_666 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_666;

architecture SYN_BEHAVIORAL of FA_666 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => A, A2 => n4, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_665 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_665;

architecture SYN_BEHAVIORAL of FA_665 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n9, n10 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : INV_X1 port map( A => n7, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n9);
   U7 : INV_X1 port map( A => n10, ZN => Co);
   U8 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n9, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_664 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_664;

architecture SYN_BEHAVIORAL of FA_664 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n9, n10 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => n4);
   U2 : INV_X1 port map( A => A, ZN => n7);
   U3 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n9);
   U7 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n9, ZN => n10);
   U8 : INV_X1 port map( A => n10, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_663 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_663;

architecture SYN_BEHAVIORAL of FA_663 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_662 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_662;

architecture SYN_BEHAVIORAL of FA_662 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_661 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_661;

architecture SYN_BEHAVIORAL of FA_661 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_660 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_660;

architecture SYN_BEHAVIORAL of FA_660 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => A, A2 => n4, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_659 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_659;

architecture SYN_BEHAVIORAL of FA_659 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_658 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_658;

architecture SYN_BEHAVIORAL of FA_658 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_657 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_657;

architecture SYN_BEHAVIORAL of FA_657 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_656 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_656;

architecture SYN_BEHAVIORAL of FA_656 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_655 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_655;

architecture SYN_BEHAVIORAL of FA_655 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_654 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_654;

architecture SYN_BEHAVIORAL of FA_654 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_653 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_653;

architecture SYN_BEHAVIORAL of FA_653 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_652 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_652;

architecture SYN_BEHAVIORAL of FA_652 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_651 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_651;

architecture SYN_BEHAVIORAL of FA_651 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_650 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_650;

architecture SYN_BEHAVIORAL of FA_650 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_649 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_649;

architecture SYN_BEHAVIORAL of FA_649 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_648 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_648;

architecture SYN_BEHAVIORAL of FA_648 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => A, A2 => n4, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_647 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_647;

architecture SYN_BEHAVIORAL of FA_647 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_646 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_646;

architecture SYN_BEHAVIORAL of FA_646 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_645 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_645;

architecture SYN_BEHAVIORAL of FA_645 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_644 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_644;

architecture SYN_BEHAVIORAL of FA_644 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_643 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_643;

architecture SYN_BEHAVIORAL of FA_643 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_642 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_642;

architecture SYN_BEHAVIORAL of FA_642 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_641 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_641;

architecture SYN_BEHAVIORAL of FA_641 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : CLKBUF_X1 port map( A => n7, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_640 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_640;

architecture SYN_BEHAVIORAL of FA_640 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => Ci, ZN => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U3 : XNOR2_X1 port map( A => n4, B => n7, ZN => S);
   U4 : XNOR2_X1 port map( A => n5, B => B, ZN => n7);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_639 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_639;

architecture SYN_BEHAVIORAL of FA_639 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_638 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_638;

architecture SYN_BEHAVIORAL of FA_638 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n4, B2 => Ci, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_637 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_637;

architecture SYN_BEHAVIORAL of FA_637 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n4, B2 => Ci, ZN => n2);
   U4 : INV_X1 port map( A => n2, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_636 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_636;

architecture SYN_BEHAVIORAL of FA_636 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n4, B2 => Ci, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_635 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_635;

architecture SYN_BEHAVIORAL of FA_635 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_634 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_634;

architecture SYN_BEHAVIORAL of FA_634 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_633 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_633;

architecture SYN_BEHAVIORAL of FA_633 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_632 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_632;

architecture SYN_BEHAVIORAL of FA_632 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_631 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_631;

architecture SYN_BEHAVIORAL of FA_631 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_630 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_630;

architecture SYN_BEHAVIORAL of FA_630 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_629 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_629;

architecture SYN_BEHAVIORAL of FA_629 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_628 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_628;

architecture SYN_BEHAVIORAL of FA_628 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_627 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_627;

architecture SYN_BEHAVIORAL of FA_627 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_626 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_626;

architecture SYN_BEHAVIORAL of FA_626 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_625 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_625;

architecture SYN_BEHAVIORAL of FA_625 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_624 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_624;

architecture SYN_BEHAVIORAL of FA_624 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_623 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_623;

architecture SYN_BEHAVIORAL of FA_623 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_622 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_622;

architecture SYN_BEHAVIORAL of FA_622 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_621 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_621;

architecture SYN_BEHAVIORAL of FA_621 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_620 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_620;

architecture SYN_BEHAVIORAL of FA_620 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_619 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_619;

architecture SYN_BEHAVIORAL of FA_619 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_618 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_618;

architecture SYN_BEHAVIORAL of FA_618 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : INV_X1 port map( A => n2, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_617 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_617;

architecture SYN_BEHAVIORAL of FA_617 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : INV_X1 port map( A => n2, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_616 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_616;

architecture SYN_BEHAVIORAL of FA_616 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_615 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_615;

architecture SYN_BEHAVIORAL of FA_615 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_614 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_614;

architecture SYN_BEHAVIORAL of FA_614 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_613 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_613;

architecture SYN_BEHAVIORAL of FA_613 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_612 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_612;

architecture SYN_BEHAVIORAL of FA_612 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => A, A2 => n7, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_611 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_611;

architecture SYN_BEHAVIORAL of FA_611 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_610 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_610;

architecture SYN_BEHAVIORAL of FA_610 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_609 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_609;

architecture SYN_BEHAVIORAL of FA_609 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => A, A2 => n7, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_608 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_608;

architecture SYN_BEHAVIORAL of FA_608 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_607 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_607;

architecture SYN_BEHAVIORAL of FA_607 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_606 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_606;

architecture SYN_BEHAVIORAL of FA_606 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => A, A2 => n7, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_605 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_605;

architecture SYN_BEHAVIORAL of FA_605 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_604 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_604;

architecture SYN_BEHAVIORAL of FA_604 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_603 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_603;

architecture SYN_BEHAVIORAL of FA_603 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_602 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_602;

architecture SYN_BEHAVIORAL of FA_602 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => A, A2 => n7, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_601 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_601;

architecture SYN_BEHAVIORAL of FA_601 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_600 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_600;

architecture SYN_BEHAVIORAL of FA_600 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_599 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_599;

architecture SYN_BEHAVIORAL of FA_599 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_598 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_598;

architecture SYN_BEHAVIORAL of FA_598 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_597 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_597;

architecture SYN_BEHAVIORAL of FA_597 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_596 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_596;

architecture SYN_BEHAVIORAL of FA_596 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_595 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_595;

architecture SYN_BEHAVIORAL of FA_595 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_594 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_594;

architecture SYN_BEHAVIORAL of FA_594 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_593 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_593;

architecture SYN_BEHAVIORAL of FA_593 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_592 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_592;

architecture SYN_BEHAVIORAL of FA_592 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_591 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_591;

architecture SYN_BEHAVIORAL of FA_591 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_590 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_590;

architecture SYN_BEHAVIORAL of FA_590 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_589 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_589;

architecture SYN_BEHAVIORAL of FA_589 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_588 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_588;

architecture SYN_BEHAVIORAL of FA_588 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_587 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_587;

architecture SYN_BEHAVIORAL of FA_587 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => A, A2 => n7, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_586 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_586;

architecture SYN_BEHAVIORAL of FA_586 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => A, A2 => n6, B1 => n5, B2 => Ci, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_585 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_585;

architecture SYN_BEHAVIORAL of FA_585 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_584 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_584;

architecture SYN_BEHAVIORAL of FA_584 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_583 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_583;

architecture SYN_BEHAVIORAL of FA_583 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_582 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_582;

architecture SYN_BEHAVIORAL of FA_582 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_581 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_581;

architecture SYN_BEHAVIORAL of FA_581 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => A, A2 => n6, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_580 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_580;

architecture SYN_BEHAVIORAL of FA_580 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_579 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_579;

architecture SYN_BEHAVIORAL of FA_579 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_578 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_578;

architecture SYN_BEHAVIORAL of FA_578 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_577 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_577;

architecture SYN_BEHAVIORAL of FA_577 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n8, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : CLKBUF_X1 port map( A => n8, Z => n5);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n8);
   U6 : INV_X1 port map( A => n9, ZN => Co);
   U7 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n5, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_576 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_576;

architecture SYN_BEHAVIORAL of FA_576 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => Ci, ZN => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U3 : XNOR2_X1 port map( A => n4, B => n7, ZN => S);
   U4 : XNOR2_X1 port map( A => n5, B => B, ZN => n7);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_575 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_575;

architecture SYN_BEHAVIORAL of FA_575 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_574 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_574;

architecture SYN_BEHAVIORAL of FA_574 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n4, B2 => Ci, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_573 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_573;

architecture SYN_BEHAVIORAL of FA_573 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : INV_X1 port map( A => n8, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_572 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_572;

architecture SYN_BEHAVIORAL of FA_572 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n4, B2 => Ci, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_571 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_571;

architecture SYN_BEHAVIORAL of FA_571 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_570 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_570;

architecture SYN_BEHAVIORAL of FA_570 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_569 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_569;

architecture SYN_BEHAVIORAL of FA_569 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_568 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_568;

architecture SYN_BEHAVIORAL of FA_568 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => A, A2 => n7, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_567 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_567;

architecture SYN_BEHAVIORAL of FA_567 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_566 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_566;

architecture SYN_BEHAVIORAL of FA_566 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_565 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_565;

architecture SYN_BEHAVIORAL of FA_565 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => A, A2 => n7, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_564 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_564;

architecture SYN_BEHAVIORAL of FA_564 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U3 : INV_X1 port map( A => n4, ZN => Co);
   U4 : CLKBUF_X1 port map( A => B, Z => n7);
   U5 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_563 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_563;

architecture SYN_BEHAVIORAL of FA_563 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_562 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_562;

architecture SYN_BEHAVIORAL of FA_562 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_561 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_561;

architecture SYN_BEHAVIORAL of FA_561 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => A, A2 => n7, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_560 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_560;

architecture SYN_BEHAVIORAL of FA_560 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => A, A2 => n7, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_559 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_559;

architecture SYN_BEHAVIORAL of FA_559 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_558 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_558;

architecture SYN_BEHAVIORAL of FA_558 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_557 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_557;

architecture SYN_BEHAVIORAL of FA_557 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => A, A2 => n7, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_556 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_556;

architecture SYN_BEHAVIORAL of FA_556 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_555 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_555;

architecture SYN_BEHAVIORAL of FA_555 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => A, A2 => n7, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_554 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_554;

architecture SYN_BEHAVIORAL of FA_554 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => A, A2 => n6, B1 => Ci, B2 => n4, ZN => n2);
   U4 : INV_X1 port map( A => n2, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_553 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_553;

architecture SYN_BEHAVIORAL of FA_553 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_552 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_552;

architecture SYN_BEHAVIORAL of FA_552 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_551 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_551;

architecture SYN_BEHAVIORAL of FA_551 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_550 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_550;

architecture SYN_BEHAVIORAL of FA_550 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_549 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_549;

architecture SYN_BEHAVIORAL of FA_549 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_548 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_548;

architecture SYN_BEHAVIORAL of FA_548 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_547 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_547;

architecture SYN_BEHAVIORAL of FA_547 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_546 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_546;

architecture SYN_BEHAVIORAL of FA_546 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => A, A2 => n4, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_545 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_545;

architecture SYN_BEHAVIORAL of FA_545 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_544 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_544;

architecture SYN_BEHAVIORAL of FA_544 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_543 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_543;

architecture SYN_BEHAVIORAL of FA_543 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_542 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_542;

architecture SYN_BEHAVIORAL of FA_542 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => A, A2 => n4, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_541 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_541;

architecture SYN_BEHAVIORAL of FA_541 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_540 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_540;

architecture SYN_BEHAVIORAL of FA_540 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_539 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_539;

architecture SYN_BEHAVIORAL of FA_539 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_538 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_538;

architecture SYN_BEHAVIORAL of FA_538 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_537 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_537;

architecture SYN_BEHAVIORAL of FA_537 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_536 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_536;

architecture SYN_BEHAVIORAL of FA_536 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_535 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_535;

architecture SYN_BEHAVIORAL of FA_535 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => A, A2 => n4, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_534 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_534;

architecture SYN_BEHAVIORAL of FA_534 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_533 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_533;

architecture SYN_BEHAVIORAL of FA_533 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_532 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_532;

architecture SYN_BEHAVIORAL of FA_532 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_531 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_531;

architecture SYN_BEHAVIORAL of FA_531 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_530 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_530;

architecture SYN_BEHAVIORAL of FA_530 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_529 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_529;

architecture SYN_BEHAVIORAL of FA_529 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U3 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_528 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_528;

architecture SYN_BEHAVIORAL of FA_528 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_527 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_527;

architecture SYN_BEHAVIORAL of FA_527 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_526 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_526;

architecture SYN_BEHAVIORAL of FA_526 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n9, n10 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : INV_X1 port map( A => n7, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : XNOR2_X1 port map( A => Ci, B => n5, ZN => S);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n9);
   U7 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n9, ZN => n10);
   U8 : INV_X1 port map( A => n10, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_525 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_525;

architecture SYN_BEHAVIORAL of FA_525 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_524 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_524;

architecture SYN_BEHAVIORAL of FA_524 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_523 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_523;

architecture SYN_BEHAVIORAL of FA_523 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_522 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_522;

architecture SYN_BEHAVIORAL of FA_522 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_521 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_521;

architecture SYN_BEHAVIORAL of FA_521 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_520 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_520;

architecture SYN_BEHAVIORAL of FA_520 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_519 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_519;

architecture SYN_BEHAVIORAL of FA_519 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_518 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_518;

architecture SYN_BEHAVIORAL of FA_518 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_517 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_517;

architecture SYN_BEHAVIORAL of FA_517 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_516 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_516;

architecture SYN_BEHAVIORAL of FA_516 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => A, A2 => n4, B1 => n7, B2 => Ci, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_515 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_515;

architecture SYN_BEHAVIORAL of FA_515 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : INV_X1 port map( A => n2, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_514 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_514;

architecture SYN_BEHAVIORAL of FA_514 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_513 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_513;

architecture SYN_BEHAVIORAL of FA_513 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n8, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U4 : CLKBUF_X1 port map( A => n8, Z => n5);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n8);
   U6 : INV_X1 port map( A => n9, ZN => Co);
   U7 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => n4, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_512 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_512;

architecture SYN_BEHAVIORAL of FA_512 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n6, B2 => Ci, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_511 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_511;

architecture SYN_BEHAVIORAL of FA_511 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_510 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_510;

architecture SYN_BEHAVIORAL of FA_510 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n4, B2 => Ci, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_509 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_509;

architecture SYN_BEHAVIORAL of FA_509 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n4, B2 => Ci, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_508 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_508;

architecture SYN_BEHAVIORAL of FA_508 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_507 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_507;

architecture SYN_BEHAVIORAL of FA_507 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_506 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_506;

architecture SYN_BEHAVIORAL of FA_506 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_505 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_505;

architecture SYN_BEHAVIORAL of FA_505 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_504 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_504;

architecture SYN_BEHAVIORAL of FA_504 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_503 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_503;

architecture SYN_BEHAVIORAL of FA_503 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_502 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_502;

architecture SYN_BEHAVIORAL of FA_502 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_501 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_501;

architecture SYN_BEHAVIORAL of FA_501 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_500 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_500;

architecture SYN_BEHAVIORAL of FA_500 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_499 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_499;

architecture SYN_BEHAVIORAL of FA_499 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_498 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_498;

architecture SYN_BEHAVIORAL of FA_498 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_497 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_497;

architecture SYN_BEHAVIORAL of FA_497 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U2 : AOI21_X1 port map( B1 => n7, B2 => A, A => Ci, ZN => n5);
   U3 : NOR2_X1 port map( A1 => n7, A2 => A, ZN => n4);
   U4 : NOR2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_496 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_496;

architecture SYN_BEHAVIORAL of FA_496 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_495 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_495;

architecture SYN_BEHAVIORAL of FA_495 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_494 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_494;

architecture SYN_BEHAVIORAL of FA_494 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => A, A2 => n7, B1 => n5, B2 => Ci, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_493 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_493;

architecture SYN_BEHAVIORAL of FA_493 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_492 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_492;

architecture SYN_BEHAVIORAL of FA_492 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_491 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_491;

architecture SYN_BEHAVIORAL of FA_491 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_490 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_490;

architecture SYN_BEHAVIORAL of FA_490 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_489 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_489;

architecture SYN_BEHAVIORAL of FA_489 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net92921, net92920, net93797, net92919, n2, n4, n5, n6 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n4, B2 => Ci, ZN => n2);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : CLKBUF_X1 port map( A => B, Z => n6);
   U4 : INV_X1 port map( A => A, ZN => n5);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => net93797, ZN => net92921);
   U6 : INV_X1 port map( A => Ci, ZN => net92919);
   U7 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U8 : NAND2_X1 port map( A1 => n4, A2 => net92919, ZN => net92920);
   U9 : XOR2_X1 port map( A => B, B => n5, Z => net93797);
   U10 : NAND2_X1 port map( A1 => net92920, A2 => net92921, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_488 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_488;

architecture SYN_BEHAVIORAL of FA_488 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n5);
   U5 : INV_X1 port map( A => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_487 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_487;

architecture SYN_BEHAVIORAL of FA_487 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : AOI22_X1 port map( A1 => A, A2 => n4, B1 => Ci, B2 => n6, ZN => n5);
   U5 : INV_X1 port map( A => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_486 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_486;

architecture SYN_BEHAVIORAL of FA_486 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_485 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_485;

architecture SYN_BEHAVIORAL of FA_485 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => A, A2 => n7, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_484 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_484;

architecture SYN_BEHAVIORAL of FA_484 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n6, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_483 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_483;

architecture SYN_BEHAVIORAL of FA_483 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_482 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_482;

architecture SYN_BEHAVIORAL of FA_482 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_481 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_481;

architecture SYN_BEHAVIORAL of FA_481 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_480 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_480;

architecture SYN_BEHAVIORAL of FA_480 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_479 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_479;

architecture SYN_BEHAVIORAL of FA_479 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_478 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_478;

architecture SYN_BEHAVIORAL of FA_478 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_477 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_477;

architecture SYN_BEHAVIORAL of FA_477 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_476 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_476;

architecture SYN_BEHAVIORAL of FA_476 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_475 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_475;

architecture SYN_BEHAVIORAL of FA_475 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_474 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_474;

architecture SYN_BEHAVIORAL of FA_474 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_473 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_473;

architecture SYN_BEHAVIORAL of FA_473 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_472 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_472;

architecture SYN_BEHAVIORAL of FA_472 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_471 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_471;

architecture SYN_BEHAVIORAL of FA_471 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : AOI22_X1 port map( A1 => A, A2 => B, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_470 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_470;

architecture SYN_BEHAVIORAL of FA_470 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_469 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_469;

architecture SYN_BEHAVIORAL of FA_469 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_468 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_468;

architecture SYN_BEHAVIORAL of FA_468 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_467 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_467;

architecture SYN_BEHAVIORAL of FA_467 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_466 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_466;

architecture SYN_BEHAVIORAL of FA_466 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : AOI22_X1 port map( A1 => A, A2 => B, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_465 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_465;

architecture SYN_BEHAVIORAL of FA_465 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_464 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_464;

architecture SYN_BEHAVIORAL of FA_464 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_463 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_463;

architecture SYN_BEHAVIORAL of FA_463 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_462 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_462;

architecture SYN_BEHAVIORAL of FA_462 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_461 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_461;

architecture SYN_BEHAVIORAL of FA_461 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_460 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_460;

architecture SYN_BEHAVIORAL of FA_460 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_459 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_459;

architecture SYN_BEHAVIORAL of FA_459 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_458 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_458;

architecture SYN_BEHAVIORAL of FA_458 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => n5, B => B, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_457 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_457;

architecture SYN_BEHAVIORAL of FA_457 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_456 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_456;

architecture SYN_BEHAVIORAL of FA_456 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_455 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_455;

architecture SYN_BEHAVIORAL of FA_455 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_454 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_454;

architecture SYN_BEHAVIORAL of FA_454 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_453 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_453;

architecture SYN_BEHAVIORAL of FA_453 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_452 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_452;

architecture SYN_BEHAVIORAL of FA_452 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_451 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_451;

architecture SYN_BEHAVIORAL of FA_451 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_450 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_450;

architecture SYN_BEHAVIORAL of FA_450 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n4, B2 => Ci, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_449 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_449;

architecture SYN_BEHAVIORAL of FA_449 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n9, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U4 : CLKBUF_X1 port map( A => n9, Z => n5);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n9);
   U6 : CLKBUF_X1 port map( A => B, Z => n7);
   U7 : INV_X1 port map( A => n10, ZN => Co);
   U8 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => n5, B2 => n4, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_448 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_448;

architecture SYN_BEHAVIORAL of FA_448 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => Ci, ZN => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U3 : XNOR2_X1 port map( A => n4, B => n7, ZN => S);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_447 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_447;

architecture SYN_BEHAVIORAL of FA_447 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_446 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_446;

architecture SYN_BEHAVIORAL of FA_446 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n4, B2 => Ci, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_445 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_445;

architecture SYN_BEHAVIORAL of FA_445 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_444 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_444;

architecture SYN_BEHAVIORAL of FA_444 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n6, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_443 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_443;

architecture SYN_BEHAVIORAL of FA_443 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_442 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_442;

architecture SYN_BEHAVIORAL of FA_442 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_441 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_441;

architecture SYN_BEHAVIORAL of FA_441 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_440 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_440;

architecture SYN_BEHAVIORAL of FA_440 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_439 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_439;

architecture SYN_BEHAVIORAL of FA_439 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_438 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_438;

architecture SYN_BEHAVIORAL of FA_438 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_437 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_437;

architecture SYN_BEHAVIORAL of FA_437 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_436 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_436;

architecture SYN_BEHAVIORAL of FA_436 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_435 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_435;

architecture SYN_BEHAVIORAL of FA_435 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_434 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_434;

architecture SYN_BEHAVIORAL of FA_434 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_433 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_433;

architecture SYN_BEHAVIORAL of FA_433 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_432 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_432;

architecture SYN_BEHAVIORAL of FA_432 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_431 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_431;

architecture SYN_BEHAVIORAL of FA_431 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_430 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_430;

architecture SYN_BEHAVIORAL of FA_430 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_429 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_429;

architecture SYN_BEHAVIORAL of FA_429 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_428 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_428;

architecture SYN_BEHAVIORAL of FA_428 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_427 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_427;

architecture SYN_BEHAVIORAL of FA_427 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_426 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_426;

architecture SYN_BEHAVIORAL of FA_426 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_425 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_425;

architecture SYN_BEHAVIORAL of FA_425 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : AOI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n5);
   U3 : NOR2_X1 port map( A1 => B, A2 => A, ZN => n4);
   U4 : NOR2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U5 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_424 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_424;

architecture SYN_BEHAVIORAL of FA_424 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => A, A2 => n7, B1 => n5, B2 => Ci, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_423 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_423;

architecture SYN_BEHAVIORAL of FA_423 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_422 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_422;

architecture SYN_BEHAVIORAL of FA_422 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_421 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_421;

architecture SYN_BEHAVIORAL of FA_421 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => A, A2 => n7, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_420 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_420;

architecture SYN_BEHAVIORAL of FA_420 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n6, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_419 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_419;

architecture SYN_BEHAVIORAL of FA_419 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_418 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_418;

architecture SYN_BEHAVIORAL of FA_418 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_417 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_417;

architecture SYN_BEHAVIORAL of FA_417 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_416 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_416;

architecture SYN_BEHAVIORAL of FA_416 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_415 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_415;

architecture SYN_BEHAVIORAL of FA_415 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_414 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_414;

architecture SYN_BEHAVIORAL of FA_414 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_413 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_413;

architecture SYN_BEHAVIORAL of FA_413 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_412 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_412;

architecture SYN_BEHAVIORAL of FA_412 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_411 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_411;

architecture SYN_BEHAVIORAL of FA_411 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n9, n10 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : XNOR2_X1 port map( A => Ci, B => n5, ZN => S);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n9);
   U6 : CLKBUF_X1 port map( A => B, Z => n7);
   U7 : INV_X1 port map( A => n10, ZN => Co);
   U8 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n9, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_410 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_410;

architecture SYN_BEHAVIORAL of FA_410 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => A, A2 => n4, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_409 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_409;

architecture SYN_BEHAVIORAL of FA_409 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_408 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_408;

architecture SYN_BEHAVIORAL of FA_408 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_407 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_407;

architecture SYN_BEHAVIORAL of FA_407 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_406 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_406;

architecture SYN_BEHAVIORAL of FA_406 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_405 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_405;

architecture SYN_BEHAVIORAL of FA_405 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_404 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_404;

architecture SYN_BEHAVIORAL of FA_404 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => A, A2 => n4, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_403 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_403;

architecture SYN_BEHAVIORAL of FA_403 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_402 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_402;

architecture SYN_BEHAVIORAL of FA_402 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_401 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_401;

architecture SYN_BEHAVIORAL of FA_401 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_400 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_400;

architecture SYN_BEHAVIORAL of FA_400 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_399 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_399;

architecture SYN_BEHAVIORAL of FA_399 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_398 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_398;

architecture SYN_BEHAVIORAL of FA_398 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => A, A2 => n4, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_397 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_397;

architecture SYN_BEHAVIORAL of FA_397 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_396 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_396;

architecture SYN_BEHAVIORAL of FA_396 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_395 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_395;

architecture SYN_BEHAVIORAL of FA_395 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_394 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_394;

architecture SYN_BEHAVIORAL of FA_394 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n9, n10 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : INV_X1 port map( A => n7, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : XNOR2_X1 port map( A => n5, B => Ci, ZN => S);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n9);
   U7 : INV_X1 port map( A => n10, ZN => Co);
   U8 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n9, B2 => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_393 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_393;

architecture SYN_BEHAVIORAL of FA_393 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => A, A2 => n4, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_392 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_392;

architecture SYN_BEHAVIORAL of FA_392 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => A, A2 => n4, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_391 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_391;

architecture SYN_BEHAVIORAL of FA_391 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_390 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_390;

architecture SYN_BEHAVIORAL of FA_390 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_389 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_389;

architecture SYN_BEHAVIORAL of FA_389 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => A, A2 => n4, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_388 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_388;

architecture SYN_BEHAVIORAL of FA_388 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => A, A2 => n4, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_387 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_387;

architecture SYN_BEHAVIORAL of FA_387 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_386 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_386;

architecture SYN_BEHAVIORAL of FA_386 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n4, B2 => Ci, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_385 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_385;

architecture SYN_BEHAVIORAL of FA_385 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n8, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : CLKBUF_X1 port map( A => n8, Z => n5);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n8);
   U6 : INV_X1 port map( A => n9, ZN => Co);
   U7 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n5, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_384 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_384;

architecture SYN_BEHAVIORAL of FA_384 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => Ci, ZN => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U3 : XNOR2_X1 port map( A => n4, B => n7, ZN => S);
   U4 : XNOR2_X1 port map( A => n5, B => B, ZN => n7);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_383 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_383;

architecture SYN_BEHAVIORAL of FA_383 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_382 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_382;

architecture SYN_BEHAVIORAL of FA_382 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n4, B2 => Ci, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_381 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_381;

architecture SYN_BEHAVIORAL of FA_381 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n4, B2 => Ci, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_380 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_380;

architecture SYN_BEHAVIORAL of FA_380 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n6, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_379 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_379;

architecture SYN_BEHAVIORAL of FA_379 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_378 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_378;

architecture SYN_BEHAVIORAL of FA_378 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => A, A2 => n7, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_377 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_377;

architecture SYN_BEHAVIORAL of FA_377 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_376 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_376;

architecture SYN_BEHAVIORAL of FA_376 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_375 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_375;

architecture SYN_BEHAVIORAL of FA_375 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_374 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_374;

architecture SYN_BEHAVIORAL of FA_374 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_373 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_373;

architecture SYN_BEHAVIORAL of FA_373 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_372 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_372;

architecture SYN_BEHAVIORAL of FA_372 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_371 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_371;

architecture SYN_BEHAVIORAL of FA_371 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_370 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_370;

architecture SYN_BEHAVIORAL of FA_370 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_369 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_369;

architecture SYN_BEHAVIORAL of FA_369 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_368 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_368;

architecture SYN_BEHAVIORAL of FA_368 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_367 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_367;

architecture SYN_BEHAVIORAL of FA_367 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_366 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_366;

architecture SYN_BEHAVIORAL of FA_366 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_365 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_365;

architecture SYN_BEHAVIORAL of FA_365 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_364 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_364;

architecture SYN_BEHAVIORAL of FA_364 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_363 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_363;

architecture SYN_BEHAVIORAL of FA_363 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => A, A2 => n6, B1 => n5, B2 => Ci, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_362 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_362;

architecture SYN_BEHAVIORAL of FA_362 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_361 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_361;

architecture SYN_BEHAVIORAL of FA_361 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_360 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_360;

architecture SYN_BEHAVIORAL of FA_360 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_359 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_359;

architecture SYN_BEHAVIORAL of FA_359 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => A, A2 => n6, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_358 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_358;

architecture SYN_BEHAVIORAL of FA_358 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_357 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_357;

architecture SYN_BEHAVIORAL of FA_357 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_356 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_356;

architecture SYN_BEHAVIORAL of FA_356 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_355 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_355;

architecture SYN_BEHAVIORAL of FA_355 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_354 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_354;

architecture SYN_BEHAVIORAL of FA_354 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_353 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_353;

architecture SYN_BEHAVIORAL of FA_353 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_352 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_352;

architecture SYN_BEHAVIORAL of FA_352 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_351 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_351;

architecture SYN_BEHAVIORAL of FA_351 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : AOI21_X1 port map( B1 => n7, B2 => A, A => Ci, ZN => n5);
   U3 : NOR2_X1 port map( A1 => n7, A2 => A, ZN => n4);
   U4 : NOR2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_350 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_350;

architecture SYN_BEHAVIORAL of FA_350 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : XOR2_X1 port map( A => B, B => n8, Z => n4);
   U3 : INV_X1 port map( A => A, ZN => n8);
   U4 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n6, ZN => n5);
   U5 : INV_X1 port map( A => n5, ZN => Co);
   U6 : CLKBUF_X1 port map( A => B, Z => n7);
   U7 : XNOR2_X1 port map( A => B, B => n8, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_349 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_349;

architecture SYN_BEHAVIORAL of FA_349 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_348 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_348;

architecture SYN_BEHAVIORAL of FA_348 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_347 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_347;

architecture SYN_BEHAVIORAL of FA_347 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_346 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_346;

architecture SYN_BEHAVIORAL of FA_346 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_345 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_345;

architecture SYN_BEHAVIORAL of FA_345 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_344 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_344;

architecture SYN_BEHAVIORAL of FA_344 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n9, n10 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : INV_X1 port map( A => n7, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : XNOR2_X1 port map( A => Ci, B => n5, ZN => S);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n9);
   U7 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n9, ZN => n10);
   U8 : INV_X1 port map( A => n10, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_343 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_343;

architecture SYN_BEHAVIORAL of FA_343 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n9, n10 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : INV_X1 port map( A => n7, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : XNOR2_X1 port map( A => Ci, B => n5, ZN => S);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n9);
   U7 : INV_X1 port map( A => n10, ZN => Co);
   U8 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n9, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_342 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_342;

architecture SYN_BEHAVIORAL of FA_342 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_341 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_341;

architecture SYN_BEHAVIORAL of FA_341 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => A, A2 => n4, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_340 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_340;

architecture SYN_BEHAVIORAL of FA_340 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_339 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_339;

architecture SYN_BEHAVIORAL of FA_339 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_338 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_338;

architecture SYN_BEHAVIORAL of FA_338 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => A, A2 => n4, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_337 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_337;

architecture SYN_BEHAVIORAL of FA_337 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_336 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_336;

architecture SYN_BEHAVIORAL of FA_336 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_335 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_335;

architecture SYN_BEHAVIORAL of FA_335 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_334 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_334;

architecture SYN_BEHAVIORAL of FA_334 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_333 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_333;

architecture SYN_BEHAVIORAL of FA_333 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_332 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_332;

architecture SYN_BEHAVIORAL of FA_332 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_331 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_331;

architecture SYN_BEHAVIORAL of FA_331 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_330 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_330;

architecture SYN_BEHAVIORAL of FA_330 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_329 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_329;

architecture SYN_BEHAVIORAL of FA_329 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_328 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_328;

architecture SYN_BEHAVIORAL of FA_328 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_327 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_327;

architecture SYN_BEHAVIORAL of FA_327 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_326 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_326;

architecture SYN_BEHAVIORAL of FA_326 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_325 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_325;

architecture SYN_BEHAVIORAL of FA_325 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_324 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_324;

architecture SYN_BEHAVIORAL of FA_324 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => A, A2 => n4, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_323 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_323;

architecture SYN_BEHAVIORAL of FA_323 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_322 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_322;

architecture SYN_BEHAVIORAL of FA_322 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : XNOR2_X1 port map( A => B, B => n6, ZN => n4);
   U4 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n4, B2 => Ci, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_321 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_321;

architecture SYN_BEHAVIORAL of FA_321 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n8, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : CLKBUF_X1 port map( A => n8, Z => n5);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n8);
   U6 : INV_X1 port map( A => n9, ZN => Co);
   U7 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n5, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_320 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_320;

architecture SYN_BEHAVIORAL of FA_320 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n6, B2 => Ci, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_319 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_319;

architecture SYN_BEHAVIORAL of FA_319 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_318 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_318;

architecture SYN_BEHAVIORAL of FA_318 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n4, B2 => Ci, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_317 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_317;

architecture SYN_BEHAVIORAL of FA_317 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n4, B2 => Ci, ZN => n2);
   U4 : INV_X1 port map( A => n2, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_316 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_316;

architecture SYN_BEHAVIORAL of FA_316 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : INV_X1 port map( A => n2, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_315 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_315;

architecture SYN_BEHAVIORAL of FA_315 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_314 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_314;

architecture SYN_BEHAVIORAL of FA_314 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_313 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_313;

architecture SYN_BEHAVIORAL of FA_313 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_312 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_312;

architecture SYN_BEHAVIORAL of FA_312 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_311 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_311;

architecture SYN_BEHAVIORAL of FA_311 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_310 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_310;

architecture SYN_BEHAVIORAL of FA_310 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_309 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_309;

architecture SYN_BEHAVIORAL of FA_309 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_308 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_308;

architecture SYN_BEHAVIORAL of FA_308 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => A, A2 => n7, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_307 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_307;

architecture SYN_BEHAVIORAL of FA_307 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => A, A2 => n7, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_306 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_306;

architecture SYN_BEHAVIORAL of FA_306 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_305 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_305;

architecture SYN_BEHAVIORAL of FA_305 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n7);
   U4 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n5);
   U5 : INV_X1 port map( A => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_304 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_304;

architecture SYN_BEHAVIORAL of FA_304 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_303 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_303;

architecture SYN_BEHAVIORAL of FA_303 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_302 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_302;

architecture SYN_BEHAVIORAL of FA_302 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n5);
   U2 : NOR2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U4 : NOR2_X1 port map( A1 => B, A2 => A, ZN => n4);
   U5 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_301 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_301;

architecture SYN_BEHAVIORAL of FA_301 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_300 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_300;

architecture SYN_BEHAVIORAL of FA_300 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_299 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_299;

architecture SYN_BEHAVIORAL of FA_299 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => A, A2 => n7, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_298 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_298;

architecture SYN_BEHAVIORAL of FA_298 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_297 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_297;

architecture SYN_BEHAVIORAL of FA_297 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => A, A2 => n6, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_296 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_296;

architecture SYN_BEHAVIORAL of FA_296 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_295 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_295;

architecture SYN_BEHAVIORAL of FA_295 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_294 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_294;

architecture SYN_BEHAVIORAL of FA_294 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_293 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_293;

architecture SYN_BEHAVIORAL of FA_293 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => A, A2 => n7, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_292 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_292;

architecture SYN_BEHAVIORAL of FA_292 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : INV_X1 port map( A => n2, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_291 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_291;

architecture SYN_BEHAVIORAL of FA_291 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_290 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_290;

architecture SYN_BEHAVIORAL of FA_290 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => A, A2 => n7, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_289 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_289;

architecture SYN_BEHAVIORAL of FA_289 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_288 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_288;

architecture SYN_BEHAVIORAL of FA_288 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_287 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_287;

architecture SYN_BEHAVIORAL of FA_287 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_286 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_286;

architecture SYN_BEHAVIORAL of FA_286 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_285 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_285;

architecture SYN_BEHAVIORAL of FA_285 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_284 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_284;

architecture SYN_BEHAVIORAL of FA_284 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_283 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_283;

architecture SYN_BEHAVIORAL of FA_283 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_282 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_282;

architecture SYN_BEHAVIORAL of FA_282 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => A, A2 => n6, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_281 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_281;

architecture SYN_BEHAVIORAL of FA_281 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_280 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_280;

architecture SYN_BEHAVIORAL of FA_280 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_279 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_279;

architecture SYN_BEHAVIORAL of FA_279 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_278 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_278;

architecture SYN_BEHAVIORAL of FA_278 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_277 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_277;

architecture SYN_BEHAVIORAL of FA_277 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_276 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_276;

architecture SYN_BEHAVIORAL of FA_276 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_275 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_275;

architecture SYN_BEHAVIORAL of FA_275 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_274 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_274;

architecture SYN_BEHAVIORAL of FA_274 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_273 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_273;

architecture SYN_BEHAVIORAL of FA_273 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_272 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_272;

architecture SYN_BEHAVIORAL of FA_272 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_271 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_271;

architecture SYN_BEHAVIORAL of FA_271 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_270 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_270;

architecture SYN_BEHAVIORAL of FA_270 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_269 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_269;

architecture SYN_BEHAVIORAL of FA_269 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_268 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_268;

architecture SYN_BEHAVIORAL of FA_268 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_267 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_267;

architecture SYN_BEHAVIORAL of FA_267 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => A, A2 => n4, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_266 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_266;

architecture SYN_BEHAVIORAL of FA_266 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_265 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_265;

architecture SYN_BEHAVIORAL of FA_265 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_264 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_264;

architecture SYN_BEHAVIORAL of FA_264 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_263 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_263;

architecture SYN_BEHAVIORAL of FA_263 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_262 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_262;

architecture SYN_BEHAVIORAL of FA_262 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_261 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_261;

architecture SYN_BEHAVIORAL of FA_261 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => A, A2 => n4, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_260 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_260;

architecture SYN_BEHAVIORAL of FA_260 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_259 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_259;

architecture SYN_BEHAVIORAL of FA_259 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => A, A2 => n4, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_258 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_258;

architecture SYN_BEHAVIORAL of FA_258 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n4, B2 => Ci, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_257 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_257;

architecture SYN_BEHAVIORAL of FA_257 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n8, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : CLKBUF_X1 port map( A => n8, Z => n4);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n8);
   U6 : INV_X1 port map( A => n9, ZN => Co);
   U7 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n4, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_256 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_256;

architecture SYN_BEHAVIORAL of FA_256 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n6, B2 => Ci, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_255 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_255;

architecture SYN_BEHAVIORAL of FA_255 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_254 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_254;

architecture SYN_BEHAVIORAL of FA_254 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_253 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_253;

architecture SYN_BEHAVIORAL of FA_253 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_252 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_252;

architecture SYN_BEHAVIORAL of FA_252 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n6, B2 => Ci, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_251 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_251;

architecture SYN_BEHAVIORAL of FA_251 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_250 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_250;

architecture SYN_BEHAVIORAL of FA_250 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_249 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_249;

architecture SYN_BEHAVIORAL of FA_249 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_248 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_248;

architecture SYN_BEHAVIORAL of FA_248 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_247 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_247;

architecture SYN_BEHAVIORAL of FA_247 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_246 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_246;

architecture SYN_BEHAVIORAL of FA_246 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_245 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_245;

architecture SYN_BEHAVIORAL of FA_245 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U4 : CLKBUF_X1 port map( A => B, Z => n4);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_244 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_244;

architecture SYN_BEHAVIORAL of FA_244 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_243 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_243;

architecture SYN_BEHAVIORAL of FA_243 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_242 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_242;

architecture SYN_BEHAVIORAL of FA_242 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U3 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_241 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_241;

architecture SYN_BEHAVIORAL of FA_241 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_240 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_240;

architecture SYN_BEHAVIORAL of FA_240 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_239 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_239;

architecture SYN_BEHAVIORAL of FA_239 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_238 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_238;

architecture SYN_BEHAVIORAL of FA_238 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_237 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_237;

architecture SYN_BEHAVIORAL of FA_237 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_236 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_236;

architecture SYN_BEHAVIORAL of FA_236 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_235 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_235;

architecture SYN_BEHAVIORAL of FA_235 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_234 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_234;

architecture SYN_BEHAVIORAL of FA_234 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_233 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_233;

architecture SYN_BEHAVIORAL of FA_233 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_232 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_232;

architecture SYN_BEHAVIORAL of FA_232 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_231 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_231;

architecture SYN_BEHAVIORAL of FA_231 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n4);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_230 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_230;

architecture SYN_BEHAVIORAL of FA_230 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_229 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_229;

architecture SYN_BEHAVIORAL of FA_229 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => A, A2 => B, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_228 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_228;

architecture SYN_BEHAVIORAL of FA_228 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_227 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_227;

architecture SYN_BEHAVIORAL of FA_227 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_226 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_226;

architecture SYN_BEHAVIORAL of FA_226 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_225 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_225;

architecture SYN_BEHAVIORAL of FA_225 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_224 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_224;

architecture SYN_BEHAVIORAL of FA_224 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_223 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_223;

architecture SYN_BEHAVIORAL of FA_223 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_222 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_222;

architecture SYN_BEHAVIORAL of FA_222 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_221 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_221;

architecture SYN_BEHAVIORAL of FA_221 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_220 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_220;

architecture SYN_BEHAVIORAL of FA_220 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : XOR2_X1 port map( A => B, B => n8, Z => n4);
   U3 : CLKBUF_X1 port map( A => B, Z => n5);
   U4 : INV_X1 port map( A => A, ZN => n8);
   U5 : OAI22_X1 port map( A1 => n6, A2 => n8, B1 => n7, B2 => n4, ZN => Co);
   U6 : INV_X1 port map( A => n5, ZN => n6);
   U7 : INV_X1 port map( A => Ci, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_219 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_219;

architecture SYN_BEHAVIORAL of FA_219 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_218 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_218;

architecture SYN_BEHAVIORAL of FA_218 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : INV_X1 port map( A => n2, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_217 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_217;

architecture SYN_BEHAVIORAL of FA_217 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_216 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_216;

architecture SYN_BEHAVIORAL of FA_216 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_215 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_215;

architecture SYN_BEHAVIORAL of FA_215 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_214 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_214;

architecture SYN_BEHAVIORAL of FA_214 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_213 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_213;

architecture SYN_BEHAVIORAL of FA_213 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n6, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_212 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_212;

architecture SYN_BEHAVIORAL of FA_212 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_211 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_211;

architecture SYN_BEHAVIORAL of FA_211 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_210 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_210;

architecture SYN_BEHAVIORAL of FA_210 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => A, A2 => n4, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_209 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_209;

architecture SYN_BEHAVIORAL of FA_209 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_208 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_208;

architecture SYN_BEHAVIORAL of FA_208 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => A, A2 => n4, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_207 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_207;

architecture SYN_BEHAVIORAL of FA_207 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_206 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_206;

architecture SYN_BEHAVIORAL of FA_206 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_205 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_205;

architecture SYN_BEHAVIORAL of FA_205 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_204 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_204;

architecture SYN_BEHAVIORAL of FA_204 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_203 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_203;

architecture SYN_BEHAVIORAL of FA_203 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_202 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_202;

architecture SYN_BEHAVIORAL of FA_202 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_201 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_201;

architecture SYN_BEHAVIORAL of FA_201 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_200 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_200;

architecture SYN_BEHAVIORAL of FA_200 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_199 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_199;

architecture SYN_BEHAVIORAL of FA_199 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => A, A2 => n4, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_198 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_198;

architecture SYN_BEHAVIORAL of FA_198 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_197 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_197;

architecture SYN_BEHAVIORAL of FA_197 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => A, A2 => n4, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_196 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_196;

architecture SYN_BEHAVIORAL of FA_196 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_195 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_195;

architecture SYN_BEHAVIORAL of FA_195 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_194 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_194;

architecture SYN_BEHAVIORAL of FA_194 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_193 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_193;

architecture SYN_BEHAVIORAL of FA_193 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n9, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U4 : CLKBUF_X1 port map( A => n9, Z => n5);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n9);
   U7 : INV_X1 port map( A => n10, ZN => Co);
   U8 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n4, B2 => n5, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_192 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_192;

architecture SYN_BEHAVIORAL of FA_192 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_191 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_191;

architecture SYN_BEHAVIORAL of FA_191 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n6, B2 => Ci, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_190 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_190;

architecture SYN_BEHAVIORAL of FA_190 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n6, B2 => Ci, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_189 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_189;

architecture SYN_BEHAVIORAL of FA_189 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n6, B2 => Ci, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_188 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_188;

architecture SYN_BEHAVIORAL of FA_188 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n6, B2 => Ci, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_187 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_187;

architecture SYN_BEHAVIORAL of FA_187 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_186 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_186;

architecture SYN_BEHAVIORAL of FA_186 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n6, B2 => Ci, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_185 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_185;

architecture SYN_BEHAVIORAL of FA_185 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => A, A2 => n4, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_184 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_184;

architecture SYN_BEHAVIORAL of FA_184 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_183 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_183;

architecture SYN_BEHAVIORAL of FA_183 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_182 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_182;

architecture SYN_BEHAVIORAL of FA_182 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n7);
   U1 : BUF_X1 port map( A => Ci, Z => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_181 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_181;

architecture SYN_BEHAVIORAL of FA_181 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_180 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_180;

architecture SYN_BEHAVIORAL of FA_180 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_179 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_179;

architecture SYN_BEHAVIORAL of FA_179 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_178 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_178;

architecture SYN_BEHAVIORAL of FA_178 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_177 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_177;

architecture SYN_BEHAVIORAL of FA_177 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_176 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_176;

architecture SYN_BEHAVIORAL of FA_176 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_175 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_175;

architecture SYN_BEHAVIORAL of FA_175 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n6, B2 => Ci, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_174 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_174;

architecture SYN_BEHAVIORAL of FA_174 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_173 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_173;

architecture SYN_BEHAVIORAL of FA_173 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_172 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_172;

architecture SYN_BEHAVIORAL of FA_172 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_171 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_171;

architecture SYN_BEHAVIORAL of FA_171 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_170 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_170;

architecture SYN_BEHAVIORAL of FA_170 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_169 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_169;

architecture SYN_BEHAVIORAL of FA_169 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_168 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_168;

architecture SYN_BEHAVIORAL of FA_168 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_167 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_167;

architecture SYN_BEHAVIORAL of FA_167 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_166 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_166;

architecture SYN_BEHAVIORAL of FA_166 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_165 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_165;

architecture SYN_BEHAVIORAL of FA_165 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_164 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_164;

architecture SYN_BEHAVIORAL of FA_164 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_163 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_163;

architecture SYN_BEHAVIORAL of FA_163 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_162 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_162;

architecture SYN_BEHAVIORAL of FA_162 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => A, A2 => B, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_161 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_161;

architecture SYN_BEHAVIORAL of FA_161 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_160 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_160;

architecture SYN_BEHAVIORAL of FA_160 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_159 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_159;

architecture SYN_BEHAVIORAL of FA_159 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_158 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_158;

architecture SYN_BEHAVIORAL of FA_158 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : AOI22_X1 port map( A1 => A, A2 => B, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_157 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_157;

architecture SYN_BEHAVIORAL of FA_157 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_156 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_156;

architecture SYN_BEHAVIORAL of FA_156 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_155 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_155;

architecture SYN_BEHAVIORAL of FA_155 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_154 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_154;

architecture SYN_BEHAVIORAL of FA_154 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_153 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_153;

architecture SYN_BEHAVIORAL of FA_153 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_152 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_152;

architecture SYN_BEHAVIORAL of FA_152 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_151 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_151;

architecture SYN_BEHAVIORAL of FA_151 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_150 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_150;

architecture SYN_BEHAVIORAL of FA_150 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_149 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_149;

architecture SYN_BEHAVIORAL of FA_149 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n2);
   U5 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_148 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_148;

architecture SYN_BEHAVIORAL of FA_148 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => n6, B => B, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_147 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_147;

architecture SYN_BEHAVIORAL of FA_147 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n7);
   U4 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n5);
   U5 : INV_X1 port map( A => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_146 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_146;

architecture SYN_BEHAVIORAL of FA_146 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_145 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_145;

architecture SYN_BEHAVIORAL of FA_145 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_144 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_144;

architecture SYN_BEHAVIORAL of FA_144 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_143 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_143;

architecture SYN_BEHAVIORAL of FA_143 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_142 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_142;

architecture SYN_BEHAVIORAL of FA_142 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n6, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_141 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_141;

architecture SYN_BEHAVIORAL of FA_141 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => n4, B2 => n5, A => n7, ZN => Co);
   U2 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : AND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NOR2_X1 port map( A1 => n6, A2 => Ci, ZN => n7);
   U6 : XNOR2_X1 port map( A => B, B => A, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_140 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_140;

architecture SYN_BEHAVIORAL of FA_140 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => A, A2 => n6, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_139 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_139;

architecture SYN_BEHAVIORAL of FA_139 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n6, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_138 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_138;

architecture SYN_BEHAVIORAL of FA_138 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_137 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_137;

architecture SYN_BEHAVIORAL of FA_137 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_136 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_136;

architecture SYN_BEHAVIORAL of FA_136 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_135 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_135;

architecture SYN_BEHAVIORAL of FA_135 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => A, A2 => n4, B1 => n7, B2 => Ci, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_134 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_134;

architecture SYN_BEHAVIORAL of FA_134 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_133 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_133;

architecture SYN_BEHAVIORAL of FA_133 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_132 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_132;

architecture SYN_BEHAVIORAL of FA_132 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_131 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_131;

architecture SYN_BEHAVIORAL of FA_131 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => A, A2 => n4, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_130 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_130;

architecture SYN_BEHAVIORAL of FA_130 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U4 : AOI22_X1 port map( A1 => A, A2 => n6, B1 => n4, B2 => Ci, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_129 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_129;

architecture SYN_BEHAVIORAL of FA_129 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7, n8, n9, n10 : std_logic;

begin
   
   U1 : INV_X1 port map( A => Ci, ZN => n9);
   U2 : OR2_X1 port map( A1 => n8, A2 => n5, ZN => Co);
   U3 : AND2_X1 port map( A1 => A, A2 => n7, ZN => n5);
   U4 : CLKBUF_X1 port map( A => n10, Z => n6);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => A, ZN => n10);
   U7 : XNOR2_X1 port map( A => Ci, B => n10, ZN => S);
   U8 : NOR2_X1 port map( A1 => n9, A2 => n6, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_128 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_128;

architecture SYN_BEHAVIORAL of FA_128 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_127 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_127;

architecture SYN_BEHAVIORAL of FA_127 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_126 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_126;

architecture SYN_BEHAVIORAL of FA_126 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_125 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_125;

architecture SYN_BEHAVIORAL of FA_125 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n6, B2 => Ci, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_124 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_124;

architecture SYN_BEHAVIORAL of FA_124 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_123 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_123;

architecture SYN_BEHAVIORAL of FA_123 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n6, B2 => Ci, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_122 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_122;

architecture SYN_BEHAVIORAL of FA_122 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_121 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_121;

architecture SYN_BEHAVIORAL of FA_121 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n6, B2 => Ci, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_120 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_120;

architecture SYN_BEHAVIORAL of FA_120 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_119 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_119;

architecture SYN_BEHAVIORAL of FA_119 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_118 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_118;

architecture SYN_BEHAVIORAL of FA_118 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_117 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_117;

architecture SYN_BEHAVIORAL of FA_117 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_116 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_116;

architecture SYN_BEHAVIORAL of FA_116 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_115 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_115;

architecture SYN_BEHAVIORAL of FA_115 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_114 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_114;

architecture SYN_BEHAVIORAL of FA_114 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_113 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_113;

architecture SYN_BEHAVIORAL of FA_113 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_112 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_112;

architecture SYN_BEHAVIORAL of FA_112 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_111 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_111;

architecture SYN_BEHAVIORAL of FA_111 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_110 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_110;

architecture SYN_BEHAVIORAL of FA_110 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : BUF_X1 port map( A => Ci, Z => n5);
   U4 : XNOR2_X1 port map( A => n4, B => B, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_109 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_109;

architecture SYN_BEHAVIORAL of FA_109 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => n7, Z => S);
   U1 : XNOR2_X1 port map( A => n4, B => B, ZN => n7);
   U2 : INV_X1 port map( A => A, ZN => n4);
   U4 : CLKBUF_X1 port map( A => Ci, Z => n5);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_108 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_108;

architecture SYN_BEHAVIORAL of FA_108 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_107 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_107;

architecture SYN_BEHAVIORAL of FA_107 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_106 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_106;

architecture SYN_BEHAVIORAL of FA_106 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_105 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_105;

architecture SYN_BEHAVIORAL of FA_105 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_104 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_104;

architecture SYN_BEHAVIORAL of FA_104 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_103 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_103;

architecture SYN_BEHAVIORAL of FA_103 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : BUF_X1 port map( A => Ci, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_102 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_102;

architecture SYN_BEHAVIORAL of FA_102 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => n7, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U2 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_101 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_101;

architecture SYN_BEHAVIORAL of FA_101 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : BUF_X1 port map( A => Ci, Z => n4);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_100 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_100;

architecture SYN_BEHAVIORAL of FA_100 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_99 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_99;

architecture SYN_BEHAVIORAL of FA_99 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_98 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_98;

architecture SYN_BEHAVIORAL of FA_98 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_97 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_97;

architecture SYN_BEHAVIORAL of FA_97 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_96 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_96;

architecture SYN_BEHAVIORAL of FA_96 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_95 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_95;

architecture SYN_BEHAVIORAL of FA_95 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => n7, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U2 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_94 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_94;

architecture SYN_BEHAVIORAL of FA_94 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_93 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_93;

architecture SYN_BEHAVIORAL of FA_93 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_92 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_92;

architecture SYN_BEHAVIORAL of FA_92 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n7);
   U1 : CLKBUF_X1 port map( A => n7, Z => n4);
   U2 : CLKBUF_X1 port map( A => Ci, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_91 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_91;

architecture SYN_BEHAVIORAL of FA_91 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n7);
   U1 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U2 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_90 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_90;

architecture SYN_BEHAVIORAL of FA_90 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_89 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_89;

architecture SYN_BEHAVIORAL of FA_89 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_88 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_88;

architecture SYN_BEHAVIORAL of FA_88 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_87 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_87;

architecture SYN_BEHAVIORAL of FA_87 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_86 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_86;

architecture SYN_BEHAVIORAL of FA_86 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_85 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_85;

architecture SYN_BEHAVIORAL of FA_85 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_84 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_84;

architecture SYN_BEHAVIORAL of FA_84 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_83 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_83;

architecture SYN_BEHAVIORAL of FA_83 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => A, A2 => B, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_82 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_82;

architecture SYN_BEHAVIORAL of FA_82 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_81 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_81;

architecture SYN_BEHAVIORAL of FA_81 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_80 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_80;

architecture SYN_BEHAVIORAL of FA_80 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_79 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_79;

architecture SYN_BEHAVIORAL of FA_79 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_78 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_78;

architecture SYN_BEHAVIORAL of FA_78 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_77 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_77;

architecture SYN_BEHAVIORAL of FA_77 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n6, ZN => n5);
   U5 : INV_X1 port map( A => n5, ZN => Co);
   U6 : CLKBUF_X1 port map( A => B, Z => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_76 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_76;

architecture SYN_BEHAVIORAL of FA_76 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n2);
   U5 : INV_X1 port map( A => n2, ZN => Co);
   U6 : CLKBUF_X1 port map( A => B, Z => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_75 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_75;

architecture SYN_BEHAVIORAL of FA_75 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : INV_X1 port map( A => n2, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_74 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_74;

architecture SYN_BEHAVIORAL of FA_74 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_73 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_73;

architecture SYN_BEHAVIORAL of FA_73 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => A, A2 => n7, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_72 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_72;

architecture SYN_BEHAVIORAL of FA_72 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_71 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_71;

architecture SYN_BEHAVIORAL of FA_71 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_70 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_70;

architecture SYN_BEHAVIORAL of FA_70 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U3 : XNOR2_X1 port map( A => Ci, B => n5, ZN => S);
   U4 : INV_X1 port map( A => A, ZN => n7);
   U5 : AOI22_X1 port map( A1 => A, A2 => n8, B1 => Ci, B2 => n9, ZN => n6);
   U6 : INV_X1 port map( A => n6, ZN => Co);
   U7 : CLKBUF_X1 port map( A => B, Z => n8);
   U8 : XNOR2_X1 port map( A => B, B => n7, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_69 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_69;

architecture SYN_BEHAVIORAL of FA_69 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => n6, Z => S);
   U1 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n7);
   U4 : AOI22_X1 port map( A1 => n8, A2 => A, B1 => Ci, B2 => n6, ZN => n5);
   U5 : INV_X1 port map( A => n5, ZN => Co);
   U6 : CLKBUF_X1 port map( A => B, Z => n8);
   U7 : XNOR2_X1 port map( A => B, B => n7, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_68 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_68;

architecture SYN_BEHAVIORAL of FA_68 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => n4, Z => S);
   U1 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n7);
   U4 : AOI22_X1 port map( A1 => n8, A2 => A, B1 => Ci, B2 => n6, ZN => n5);
   U5 : INV_X1 port map( A => n5, ZN => Co);
   U6 : CLKBUF_X1 port map( A => B, Z => n8);
   U7 : XNOR2_X1 port map( A => B, B => n7, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_67 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_67;

architecture SYN_BEHAVIORAL of FA_67 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => n4, Z => S);
   U1 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n7);
   U4 : AOI22_X1 port map( A1 => n8, A2 => A, B1 => Ci, B2 => n6, ZN => n5);
   U5 : INV_X1 port map( A => n5, ZN => Co);
   U6 : CLKBUF_X1 port map( A => B, Z => n8);
   U7 : XNOR2_X1 port map( A => B, B => n7, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_66 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_66;

architecture SYN_BEHAVIORAL of FA_66 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_65 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_65;

architecture SYN_BEHAVIORAL of FA_65 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net97982, net99540, net99568, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : OR2_X1 port map( A1 => n8, A2 => n5, ZN => Co);
   U2 : AND2_X1 port map( A1 => A, A2 => n7, ZN => n5);
   U3 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);
   U4 : CLKBUF_X1 port map( A => Ci, Z => net99568);
   U5 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U6 : CLKBUF_X1 port map( A => n6, Z => net99540);
   U7 : CLKBUF_X1 port map( A => B, Z => n7);
   U8 : INV_X1 port map( A => net99568, ZN => net97982);
   U9 : NOR2_X1 port map( A1 => net97982, A2 => net99540, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_64 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_64;

architecture SYN_BEHAVIORAL of FA_64 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_63 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_63;

architecture SYN_BEHAVIORAL of FA_63 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_62 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_62;

architecture SYN_BEHAVIORAL of FA_62 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_61 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_61;

architecture SYN_BEHAVIORAL of FA_61 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_60 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_60;

architecture SYN_BEHAVIORAL of FA_60 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_59 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_59;

architecture SYN_BEHAVIORAL of FA_59 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_58 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_58;

architecture SYN_BEHAVIORAL of FA_58 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_57 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_57;

architecture SYN_BEHAVIORAL of FA_57 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_56 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_56;

architecture SYN_BEHAVIORAL of FA_56 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_55 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_55;

architecture SYN_BEHAVIORAL of FA_55 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_54 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_54;

architecture SYN_BEHAVIORAL of FA_54 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_53 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_53;

architecture SYN_BEHAVIORAL of FA_53 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_52 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_52;

architecture SYN_BEHAVIORAL of FA_52 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_51 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_51;

architecture SYN_BEHAVIORAL of FA_51 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_50 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_50;

architecture SYN_BEHAVIORAL of FA_50 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_49 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_49;

architecture SYN_BEHAVIORAL of FA_49 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_48 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_48;

architecture SYN_BEHAVIORAL of FA_48 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_47 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_47;

architecture SYN_BEHAVIORAL of FA_47 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_46 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_46;

architecture SYN_BEHAVIORAL of FA_46 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_45 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_45;

architecture SYN_BEHAVIORAL of FA_45 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_44 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_44;

architecture SYN_BEHAVIORAL of FA_44 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_43 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_43;

architecture SYN_BEHAVIORAL of FA_43 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_42 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_42;

architecture SYN_BEHAVIORAL of FA_42 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_41 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_41;

architecture SYN_BEHAVIORAL of FA_41 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_40 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_40;

architecture SYN_BEHAVIORAL of FA_40 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_39 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_39;

architecture SYN_BEHAVIORAL of FA_39 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_38 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_38;

architecture SYN_BEHAVIORAL of FA_38 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_37 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_37;

architecture SYN_BEHAVIORAL of FA_37 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_36 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_36;

architecture SYN_BEHAVIORAL of FA_36 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_35 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_35;

architecture SYN_BEHAVIORAL of FA_35 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_34 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_34;

architecture SYN_BEHAVIORAL of FA_34 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n6, B2 => Ci, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_33 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_33;

architecture SYN_BEHAVIORAL of FA_33 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_32 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_32;

architecture SYN_BEHAVIORAL of FA_32 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U2 : CLKBUF_X1 port map( A => n7, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_31 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_31;

architecture SYN_BEHAVIORAL of FA_31 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_30 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_30;

architecture SYN_BEHAVIORAL of FA_30 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : CLKBUF_X1 port map( A => n7, Z => n4);
   U2 : CLKBUF_X1 port map( A => Ci, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_29 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_29;

architecture SYN_BEHAVIORAL of FA_29 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_28 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_28;

architecture SYN_BEHAVIORAL of FA_28 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n7);
   U1 : CLKBUF_X1 port map( A => n7, Z => n4);
   U2 : CLKBUF_X1 port map( A => Ci, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_27 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_27;

architecture SYN_BEHAVIORAL of FA_27 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n7);
   U4 : CLKBUF_X1 port map( A => Ci, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_26 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_26;

architecture SYN_BEHAVIORAL of FA_26 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_25 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_25;

architecture SYN_BEHAVIORAL of FA_25 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_24 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_24;

architecture SYN_BEHAVIORAL of FA_24 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_23 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_23;

architecture SYN_BEHAVIORAL of FA_23 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_22 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_22;

architecture SYN_BEHAVIORAL of FA_22 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_21 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_21;

architecture SYN_BEHAVIORAL of FA_21 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_20 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_20;

architecture SYN_BEHAVIORAL of FA_20 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_19 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_19;

architecture SYN_BEHAVIORAL of FA_19 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_18 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_18;

architecture SYN_BEHAVIORAL of FA_18 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_17 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_17;

architecture SYN_BEHAVIORAL of FA_17 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_16 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_16;

architecture SYN_BEHAVIORAL of FA_16 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U2 : INV_X1 port map( A => n7, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_15 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_15;

architecture SYN_BEHAVIORAL of FA_15 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_14 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_14;

architecture SYN_BEHAVIORAL of FA_14 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_13 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_13;

architecture SYN_BEHAVIORAL of FA_13 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : CLKBUF_X1 port map( A => n7, Z => n4);
   U2 : CLKBUF_X1 port map( A => Ci, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_12 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_12;

architecture SYN_BEHAVIORAL of FA_12 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n7);
   U1 : CLKBUF_X1 port map( A => n7, Z => n4);
   U2 : CLKBUF_X1 port map( A => Ci, Z => n5);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U6 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_11 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_11;

architecture SYN_BEHAVIORAL of FA_11 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n8);
   U1 : CLKBUF_X1 port map( A => n8, Z => n4);
   U2 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : CLKBUF_X1 port map( A => Ci, Z => n6);
   U6 : INV_X1 port map( A => n9, ZN => Co);
   U7 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n8, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_10 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_10;

architecture SYN_BEHAVIORAL of FA_10 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => n4, Z => S);
   U1 : CLKBUF_X1 port map( A => n8, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n5);
   U4 : XNOR2_X1 port map( A => n5, B => B, ZN => n8);
   U5 : CLKBUF_X1 port map( A => Ci, Z => n6);
   U6 : INV_X1 port map( A => n9, ZN => Co);
   U7 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n8, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_9 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_9;

architecture SYN_BEHAVIORAL of FA_9 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => n8, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n8);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : CLKBUF_X1 port map( A => Ci, Z => n6);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n8, ZN => n9);
   U7 : INV_X1 port map( A => n9, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_8 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_8;

architecture SYN_BEHAVIORAL of FA_8 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => n4, Z => S);
   U1 : CLKBUF_X1 port map( A => n9, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n7);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : CLKBUF_X1 port map( A => Ci, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n9);
   U7 : INV_X1 port map( A => n10, ZN => Co);
   U8 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n9, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_7 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_7;

architecture SYN_BEHAVIORAL of FA_7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : CLKBUF_X1 port map( A => n9, Z => n5);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n9);
   U6 : CLKBUF_X1 port map( A => Ci, Z => n7);
   U7 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n9, ZN => n10);
   U8 : INV_X1 port map( A => n10, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_6 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_6;

architecture SYN_BEHAVIORAL of FA_6 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => Ci, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_5 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_5;

architecture SYN_BEHAVIORAL of FA_5 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal net91727, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => net91727, Z => S);
   U1 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U2 : NOR2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : AOI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n6);
   U5 : NOR2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U6 : CLKBUF_X1 port map( A => Ci, Z => net91727);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_4 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_4;

architecture SYN_BEHAVIORAL of FA_4 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal net90567, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => net90567, Z => S);
   U1 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U2 : NOR2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : AOI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n6);
   U5 : NOR2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U6 : CLKBUF_X1 port map( A => Ci, Z => net90567);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_3 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_3;

architecture SYN_BEHAVIORAL of FA_3 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal net94500, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => net94500, B => n4, Z => S);
   U1 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U2 : NOR2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : AOI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n6);
   U5 : NOR2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U6 : CLKBUF_X1 port map( A => Ci, Z => net94500);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_2 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2;

architecture SYN_BEHAVIORAL of FA_2 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => n4, Z => S);
   U1 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U2 : CLKBUF_X1 port map( A => Ci, Z => n5);
   U4 : AOI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n7);
   U5 : NOR2_X1 port map( A1 => n7, A2 => n6, ZN => Co);
   U6 : NOR2_X1 port map( A1 => B, A2 => A, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_1 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1;

architecture SYN_BEHAVIORAL of FA_1 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net92770, net102951, net102946, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => net92770, ZN => net102946);
   U2 : OR2_X1 port map( A1 => n8, A2 => n5, ZN => Co);
   U3 : AND2_X1 port map( A1 => A, A2 => n7, ZN => n5);
   U4 : XNOR2_X1 port map( A => n6, B => Ci, ZN => S);
   U5 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U6 : CLKBUF_X1 port map( A => n6, Z => net102951);
   U7 : CLKBUF_X1 port map( A => Ci, Z => net92770);
   U8 : CLKBUF_X1 port map( A => B, Z => n7);
   U9 : NOR2_X1 port map( A1 => net102951, A2 => net102946, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity shifter_N64_30 is

   port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
         std_logic_vector (63 downto 0));

end shifter_N64_30;

architecture SYN_beh of shifter_N64_30 is

signal X_Logic0_port : std_logic;

begin
   shiftLeftOnePos <= ( input(62), input(61), input(60), input(59), input(58), 
      input(57), input(56), input(55), input(54), input(53), input(52), 
      input(51), input(50), input(49), input(48), input(47), input(46), 
      input(45), input(44), input(43), input(42), input(41), input(40), 
      input(39), input(38), input(37), input(36), input(35), input(34), 
      input(33), input(32), input(31), input(30), input(29), input(28), 
      input(27), input(26), input(25), input(24), input(23), input(22), 
      input(21), input(20), input(19), input(18), input(17), input(16), 
      input(15), input(14), input(13), input(12), input(11), input(10), 
      input(9), input(8), input(7), input(6), input(5), input(4), input(3), 
      input(2), input(1), input(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity shifter_N64_29 is

   port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
         std_logic_vector (63 downto 0));

end shifter_N64_29;

architecture SYN_beh of shifter_N64_29 is

signal X_Logic0_port : std_logic;

begin
   shiftLeftOnePos <= ( input(62), input(61), input(60), input(59), input(58), 
      input(57), input(56), input(55), input(54), input(53), input(52), 
      input(51), input(50), input(49), input(48), input(47), input(46), 
      input(45), input(44), input(43), input(42), input(41), input(40), 
      input(39), input(38), input(37), input(36), input(35), input(34), 
      input(33), input(32), input(31), input(30), input(29), input(28), 
      input(27), input(26), input(25), input(24), input(23), input(22), 
      input(21), input(20), input(19), input(18), input(17), input(16), 
      input(15), input(14), input(13), input(12), input(11), input(10), 
      input(9), input(8), input(7), input(6), input(5), input(4), input(3), 
      input(2), input(1), input(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity shifter_N64_28 is

   port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
         std_logic_vector (63 downto 0));

end shifter_N64_28;

architecture SYN_beh of shifter_N64_28 is

signal X_Logic0_port : std_logic;

begin
   shiftLeftOnePos <= ( input(62), input(61), input(60), input(59), input(58), 
      input(57), input(56), input(55), input(54), input(53), input(52), 
      input(51), input(50), input(49), input(48), input(47), input(46), 
      input(45), input(44), input(43), input(42), input(41), input(40), 
      input(39), input(38), input(37), input(36), input(35), input(34), 
      input(33), input(32), input(31), input(30), input(29), input(28), 
      input(27), input(26), input(25), input(24), input(23), input(22), 
      input(21), input(20), input(19), input(18), input(17), input(16), 
      input(15), input(14), input(13), input(12), input(11), input(10), 
      input(9), input(8), input(7), input(6), input(5), input(4), input(3), 
      input(2), input(1), input(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity shifter_N64_27 is

   port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
         std_logic_vector (63 downto 0));

end shifter_N64_27;

architecture SYN_beh of shifter_N64_27 is

signal X_Logic0_port : std_logic;

begin
   shiftLeftOnePos <= ( input(62), input(61), input(60), input(59), input(58), 
      input(57), input(56), input(55), input(54), input(53), input(52), 
      input(51), input(50), input(49), input(48), input(47), input(46), 
      input(45), input(44), input(43), input(42), input(41), input(40), 
      input(39), input(38), input(37), input(36), input(35), input(34), 
      input(33), input(32), input(31), input(30), input(29), input(28), 
      input(27), input(26), input(25), input(24), input(23), input(22), 
      input(21), input(20), input(19), input(18), input(17), input(16), 
      input(15), input(14), input(13), input(12), input(11), input(10), 
      input(9), input(8), input(7), input(6), input(5), input(4), input(3), 
      input(2), input(1), input(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity shifter_N64_26 is

   port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
         std_logic_vector (63 downto 0));

end shifter_N64_26;

architecture SYN_beh of shifter_N64_26 is

signal X_Logic0_port : std_logic;

begin
   shiftLeftOnePos <= ( input(62), input(61), input(60), input(59), input(58), 
      input(57), input(56), input(55), input(54), input(53), input(52), 
      input(51), input(50), input(49), input(48), input(47), input(46), 
      input(45), input(44), input(43), input(42), input(41), input(40), 
      input(39), input(38), input(37), input(36), input(35), input(34), 
      input(33), input(32), input(31), input(30), input(29), input(28), 
      input(27), input(26), input(25), input(24), input(23), input(22), 
      input(21), input(20), input(19), input(18), input(17), input(16), 
      input(15), input(14), input(13), input(12), input(11), input(10), 
      input(9), input(8), input(7), input(6), input(5), input(4), input(3), 
      input(2), input(1), input(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity shifter_N64_25 is

   port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
         std_logic_vector (63 downto 0));

end shifter_N64_25;

architecture SYN_beh of shifter_N64_25 is

signal X_Logic0_port : std_logic;

begin
   shiftLeftOnePos <= ( input(62), input(61), input(60), input(59), input(58), 
      input(57), input(56), input(55), input(54), input(53), input(52), 
      input(51), input(50), input(49), input(48), input(47), input(46), 
      input(45), input(44), input(43), input(42), input(41), input(40), 
      input(39), input(38), input(37), input(36), input(35), input(34), 
      input(33), input(32), input(31), input(30), input(29), input(28), 
      input(27), input(26), input(25), input(24), input(23), input(22), 
      input(21), input(20), input(19), input(18), input(17), input(16), 
      input(15), input(14), input(13), input(12), input(11), input(10), 
      input(9), input(8), input(7), input(6), input(5), input(4), input(3), 
      input(2), input(1), input(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity shifter_N64_24 is

   port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
         std_logic_vector (63 downto 0));

end shifter_N64_24;

architecture SYN_beh of shifter_N64_24 is

signal X_Logic0_port : std_logic;

begin
   shiftLeftOnePos <= ( input(62), input(61), input(60), input(59), input(58), 
      input(57), input(56), input(55), input(54), input(53), input(52), 
      input(51), input(50), input(49), input(48), input(47), input(46), 
      input(45), input(44), input(43), input(42), input(41), input(40), 
      input(39), input(38), input(37), input(36), input(35), input(34), 
      input(33), input(32), input(31), input(30), input(29), input(28), 
      input(27), input(26), input(25), input(24), input(23), input(22), 
      input(21), input(20), input(19), input(18), input(17), input(16), 
      input(15), input(14), input(13), input(12), input(11), input(10), 
      input(9), input(8), input(7), input(6), input(5), input(4), input(3), 
      input(2), input(1), input(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity shifter_N64_23 is

   port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
         std_logic_vector (63 downto 0));

end shifter_N64_23;

architecture SYN_beh of shifter_N64_23 is

signal X_Logic0_port : std_logic;

begin
   shiftLeftOnePos <= ( input(62), input(61), input(60), input(59), input(58), 
      input(57), input(56), input(55), input(54), input(53), input(52), 
      input(51), input(50), input(49), input(48), input(47), input(46), 
      input(45), input(44), input(43), input(42), input(41), input(40), 
      input(39), input(38), input(37), input(36), input(35), input(34), 
      input(33), input(32), input(31), input(30), input(29), input(28), 
      input(27), input(26), input(25), input(24), input(23), input(22), 
      input(21), input(20), input(19), input(18), input(17), input(16), 
      input(15), input(14), input(13), input(12), input(11), input(10), 
      input(9), input(8), input(7), input(6), input(5), input(4), input(3), 
      input(2), input(1), input(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity shifter_N64_22 is

   port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
         std_logic_vector (63 downto 0));

end shifter_N64_22;

architecture SYN_beh of shifter_N64_22 is

signal X_Logic0_port : std_logic;

begin
   shiftLeftOnePos <= ( input(62), input(61), input(60), input(59), input(58), 
      input(57), input(56), input(55), input(54), input(53), input(52), 
      input(51), input(50), input(49), input(48), input(47), input(46), 
      input(45), input(44), input(43), input(42), input(41), input(40), 
      input(39), input(38), input(37), input(36), input(35), input(34), 
      input(33), input(32), input(31), input(30), input(29), input(28), 
      input(27), input(26), input(25), input(24), input(23), input(22), 
      input(21), input(20), input(19), input(18), input(17), input(16), 
      input(15), input(14), input(13), input(12), input(11), input(10), 
      input(9), input(8), input(7), input(6), input(5), input(4), input(3), 
      input(2), input(1), input(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity shifter_N64_21 is

   port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
         std_logic_vector (63 downto 0));

end shifter_N64_21;

architecture SYN_beh of shifter_N64_21 is

signal X_Logic0_port : std_logic;

begin
   shiftLeftOnePos <= ( input(62), input(61), input(60), input(59), input(58), 
      input(57), input(56), input(55), input(54), input(53), input(52), 
      input(51), input(50), input(49), input(48), input(47), input(46), 
      input(45), input(44), input(43), input(42), input(41), input(40), 
      input(39), input(38), input(37), input(36), input(35), input(34), 
      input(33), input(32), input(31), input(30), input(29), input(28), 
      input(27), input(26), input(25), input(24), input(23), input(22), 
      input(21), input(20), input(19), input(18), input(17), input(16), 
      input(15), input(14), input(13), input(12), input(11), input(10), 
      input(9), input(8), input(7), input(6), input(5), input(4), input(3), 
      input(2), input(1), input(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity shifter_N64_20 is

   port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
         std_logic_vector (63 downto 0));

end shifter_N64_20;

architecture SYN_beh of shifter_N64_20 is

signal X_Logic0_port : std_logic;

begin
   shiftLeftOnePos <= ( input(62), input(61), input(60), input(59), input(58), 
      input(57), input(56), input(55), input(54), input(53), input(52), 
      input(51), input(50), input(49), input(48), input(47), input(46), 
      input(45), input(44), input(43), input(42), input(41), input(40), 
      input(39), input(38), input(37), input(36), input(35), input(34), 
      input(33), input(32), input(31), input(30), input(29), input(28), 
      input(27), input(26), input(25), input(24), input(23), input(22), 
      input(21), input(20), input(19), input(18), input(17), input(16), 
      input(15), input(14), input(13), input(12), input(11), input(10), 
      input(9), input(8), input(7), input(6), input(5), input(4), input(3), 
      input(2), input(1), input(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity shifter_N64_19 is

   port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
         std_logic_vector (63 downto 0));

end shifter_N64_19;

architecture SYN_beh of shifter_N64_19 is

signal X_Logic0_port : std_logic;

begin
   shiftLeftOnePos <= ( input(62), input(61), input(60), input(59), input(58), 
      input(57), input(56), input(55), input(54), input(53), input(52), 
      input(51), input(50), input(49), input(48), input(47), input(46), 
      input(45), input(44), input(43), input(42), input(41), input(40), 
      input(39), input(38), input(37), input(36), input(35), input(34), 
      input(33), input(32), input(31), input(30), input(29), input(28), 
      input(27), input(26), input(25), input(24), input(23), input(22), 
      input(21), input(20), input(19), input(18), input(17), input(16), 
      input(15), input(14), input(13), input(12), input(11), input(10), 
      input(9), input(8), input(7), input(6), input(5), input(4), input(3), 
      input(2), input(1), input(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity shifter_N64_18 is

   port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
         std_logic_vector (63 downto 0));

end shifter_N64_18;

architecture SYN_beh of shifter_N64_18 is

signal X_Logic0_port : std_logic;

begin
   shiftLeftOnePos <= ( input(62), input(61), input(60), input(59), input(58), 
      input(57), input(56), input(55), input(54), input(53), input(52), 
      input(51), input(50), input(49), input(48), input(47), input(46), 
      input(45), input(44), input(43), input(42), input(41), input(40), 
      input(39), input(38), input(37), input(36), input(35), input(34), 
      input(33), input(32), input(31), input(30), input(29), input(28), 
      input(27), input(26), input(25), input(24), input(23), input(22), 
      input(21), input(20), input(19), input(18), input(17), input(16), 
      input(15), input(14), input(13), input(12), input(11), input(10), 
      input(9), input(8), input(7), input(6), input(5), input(4), input(3), 
      input(2), input(1), input(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity shifter_N64_17 is

   port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
         std_logic_vector (63 downto 0));

end shifter_N64_17;

architecture SYN_beh of shifter_N64_17 is

signal X_Logic0_port : std_logic;

begin
   shiftLeftOnePos <= ( input(62), input(61), input(60), input(59), input(58), 
      input(57), input(56), input(55), input(54), input(53), input(52), 
      input(51), input(50), input(49), input(48), input(47), input(46), 
      input(45), input(44), input(43), input(42), input(41), input(40), 
      input(39), input(38), input(37), input(36), input(35), input(34), 
      input(33), input(32), input(31), input(30), input(29), input(28), 
      input(27), input(26), input(25), input(24), input(23), input(22), 
      input(21), input(20), input(19), input(18), input(17), input(16), 
      input(15), input(14), input(13), input(12), input(11), input(10), 
      input(9), input(8), input(7), input(6), input(5), input(4), input(3), 
      input(2), input(1), input(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity shifter_N64_16 is

   port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
         std_logic_vector (63 downto 0));

end shifter_N64_16;

architecture SYN_beh of shifter_N64_16 is

signal X_Logic0_port : std_logic;

begin
   shiftLeftOnePos <= ( input(62), input(61), input(60), input(59), input(58), 
      input(57), input(56), input(55), input(54), input(53), input(52), 
      input(51), input(50), input(49), input(48), input(47), input(46), 
      input(45), input(44), input(43), input(42), input(41), input(40), 
      input(39), input(38), input(37), input(36), input(35), input(34), 
      input(33), input(32), input(31), input(30), input(29), input(28), 
      input(27), input(26), input(25), input(24), input(23), input(22), 
      input(21), input(20), input(19), input(18), input(17), input(16), 
      input(15), input(14), input(13), input(12), input(11), input(10), 
      input(9), input(8), input(7), input(6), input(5), input(4), input(3), 
      input(2), input(1), input(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity shifter_N64_15 is

   port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
         std_logic_vector (63 downto 0));

end shifter_N64_15;

architecture SYN_beh of shifter_N64_15 is

signal X_Logic0_port : std_logic;

begin
   shiftLeftOnePos <= ( input(62), input(61), input(60), input(59), input(58), 
      input(57), input(56), input(55), input(54), input(53), input(52), 
      input(51), input(50), input(49), input(48), input(47), input(46), 
      input(45), input(44), input(43), input(42), input(41), input(40), 
      input(39), input(38), input(37), input(36), input(35), input(34), 
      input(33), input(32), input(31), input(30), input(29), input(28), 
      input(27), input(26), input(25), input(24), input(23), input(22), 
      input(21), input(20), input(19), input(18), input(17), input(16), 
      input(15), input(14), input(13), input(12), input(11), input(10), 
      input(9), input(8), input(7), input(6), input(5), input(4), input(3), 
      input(2), input(1), input(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity shifter_N64_14 is

   port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
         std_logic_vector (63 downto 0));

end shifter_N64_14;

architecture SYN_beh of shifter_N64_14 is

signal X_Logic0_port : std_logic;

begin
   shiftLeftOnePos <= ( input(62), input(61), input(60), input(59), input(58), 
      input(57), input(56), input(55), input(54), input(53), input(52), 
      input(51), input(50), input(49), input(48), input(47), input(46), 
      input(45), input(44), input(43), input(42), input(41), input(40), 
      input(39), input(38), input(37), input(36), input(35), input(34), 
      input(33), input(32), input(31), input(30), input(29), input(28), 
      input(27), input(26), input(25), input(24), input(23), input(22), 
      input(21), input(20), input(19), input(18), input(17), input(16), 
      input(15), input(14), input(13), input(12), input(11), input(10), 
      input(9), input(8), input(7), input(6), input(5), input(4), input(3), 
      input(2), input(1), input(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity shifter_N64_13 is

   port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
         std_logic_vector (63 downto 0));

end shifter_N64_13;

architecture SYN_beh of shifter_N64_13 is

signal X_Logic0_port : std_logic;

begin
   shiftLeftOnePos <= ( input(62), input(61), input(60), input(59), input(58), 
      input(57), input(56), input(55), input(54), input(53), input(52), 
      input(51), input(50), input(49), input(48), input(47), input(46), 
      input(45), input(44), input(43), input(42), input(41), input(40), 
      input(39), input(38), input(37), input(36), input(35), input(34), 
      input(33), input(32), input(31), input(30), input(29), input(28), 
      input(27), input(26), input(25), input(24), input(23), input(22), 
      input(21), input(20), input(19), input(18), input(17), input(16), 
      input(15), input(14), input(13), input(12), input(11), input(10), 
      input(9), input(8), input(7), input(6), input(5), input(4), input(3), 
      input(2), input(1), input(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity shifter_N64_12 is

   port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
         std_logic_vector (63 downto 0));

end shifter_N64_12;

architecture SYN_beh of shifter_N64_12 is

signal X_Logic0_port : std_logic;

begin
   shiftLeftOnePos <= ( input(62), input(61), input(60), input(59), input(58), 
      input(57), input(56), input(55), input(54), input(53), input(52), 
      input(51), input(50), input(49), input(48), input(47), input(46), 
      input(45), input(44), input(43), input(42), input(41), input(40), 
      input(39), input(38), input(37), input(36), input(35), input(34), 
      input(33), input(32), input(31), input(30), input(29), input(28), 
      input(27), input(26), input(25), input(24), input(23), input(22), 
      input(21), input(20), input(19), input(18), input(17), input(16), 
      input(15), input(14), input(13), input(12), input(11), input(10), 
      input(9), input(8), input(7), input(6), input(5), input(4), input(3), 
      input(2), input(1), input(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity shifter_N64_11 is

   port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
         std_logic_vector (63 downto 0));

end shifter_N64_11;

architecture SYN_beh of shifter_N64_11 is

signal X_Logic0_port : std_logic;

begin
   shiftLeftOnePos <= ( input(62), input(61), input(60), input(59), input(58), 
      input(57), input(56), input(55), input(54), input(53), input(52), 
      input(51), input(50), input(49), input(48), input(47), input(46), 
      input(45), input(44), input(43), input(42), input(41), input(40), 
      input(39), input(38), input(37), input(36), input(35), input(34), 
      input(33), input(32), input(31), input(30), input(29), input(28), 
      input(27), input(26), input(25), input(24), input(23), input(22), 
      input(21), input(20), input(19), input(18), input(17), input(16), 
      input(15), input(14), input(13), input(12), input(11), input(10), 
      input(9), input(8), input(7), input(6), input(5), input(4), input(3), 
      input(2), input(1), input(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity shifter_N64_10 is

   port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
         std_logic_vector (63 downto 0));

end shifter_N64_10;

architecture SYN_beh of shifter_N64_10 is

signal X_Logic0_port : std_logic;

begin
   shiftLeftOnePos <= ( input(62), input(61), input(60), input(59), input(58), 
      input(57), input(56), input(55), input(54), input(53), input(52), 
      input(51), input(50), input(49), input(48), input(47), input(46), 
      input(45), input(44), input(43), input(42), input(41), input(40), 
      input(39), input(38), input(37), input(36), input(35), input(34), 
      input(33), input(32), input(31), input(30), input(29), input(28), 
      input(27), input(26), input(25), input(24), input(23), input(22), 
      input(21), input(20), input(19), input(18), input(17), input(16), 
      input(15), input(14), input(13), input(12), input(11), input(10), 
      input(9), input(8), input(7), input(6), input(5), input(4), input(3), 
      input(2), input(1), input(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity shifter_N64_9 is

   port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
         std_logic_vector (63 downto 0));

end shifter_N64_9;

architecture SYN_beh of shifter_N64_9 is

signal X_Logic0_port : std_logic;

begin
   shiftLeftOnePos <= ( input(62), input(61), input(60), input(59), input(58), 
      input(57), input(56), input(55), input(54), input(53), input(52), 
      input(51), input(50), input(49), input(48), input(47), input(46), 
      input(45), input(44), input(43), input(42), input(41), input(40), 
      input(39), input(38), input(37), input(36), input(35), input(34), 
      input(33), input(32), input(31), input(30), input(29), input(28), 
      input(27), input(26), input(25), input(24), input(23), input(22), 
      input(21), input(20), input(19), input(18), input(17), input(16), 
      input(15), input(14), input(13), input(12), input(11), input(10), 
      input(9), input(8), input(7), input(6), input(5), input(4), input(3), 
      input(2), input(1), input(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity shifter_N64_8 is

   port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
         std_logic_vector (63 downto 0));

end shifter_N64_8;

architecture SYN_beh of shifter_N64_8 is

signal X_Logic0_port : std_logic;

begin
   shiftLeftOnePos <= ( input(62), input(61), input(60), input(59), input(58), 
      input(57), input(56), input(55), input(54), input(53), input(52), 
      input(51), input(50), input(49), input(48), input(47), input(46), 
      input(45), input(44), input(43), input(42), input(41), input(40), 
      input(39), input(38), input(37), input(36), input(35), input(34), 
      input(33), input(32), input(31), input(30), input(29), input(28), 
      input(27), input(26), input(25), input(24), input(23), input(22), 
      input(21), input(20), input(19), input(18), input(17), input(16), 
      input(15), input(14), input(13), input(12), input(11), input(10), 
      input(9), input(8), input(7), input(6), input(5), input(4), input(3), 
      input(2), input(1), input(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity shifter_N64_7 is

   port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
         std_logic_vector (63 downto 0));

end shifter_N64_7;

architecture SYN_beh of shifter_N64_7 is

signal X_Logic0_port : std_logic;

begin
   shiftLeftOnePos <= ( input(62), input(61), input(60), input(59), input(58), 
      input(57), input(56), input(55), input(54), input(53), input(52), 
      input(51), input(50), input(49), input(48), input(47), input(46), 
      input(45), input(44), input(43), input(42), input(41), input(40), 
      input(39), input(38), input(37), input(36), input(35), input(34), 
      input(33), input(32), input(31), input(30), input(29), input(28), 
      input(27), input(26), input(25), input(24), input(23), input(22), 
      input(21), input(20), input(19), input(18), input(17), input(16), 
      input(15), input(14), input(13), input(12), input(11), input(10), 
      input(9), input(8), input(7), input(6), input(5), input(4), input(3), 
      input(2), input(1), input(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity shifter_N64_6 is

   port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
         std_logic_vector (63 downto 0));

end shifter_N64_6;

architecture SYN_beh of shifter_N64_6 is

signal X_Logic0_port : std_logic;

begin
   shiftLeftOnePos <= ( input(62), input(61), input(60), input(59), input(58), 
      input(57), input(56), input(55), input(54), input(53), input(52), 
      input(51), input(50), input(49), input(48), input(47), input(46), 
      input(45), input(44), input(43), input(42), input(41), input(40), 
      input(39), input(38), input(37), input(36), input(35), input(34), 
      input(33), input(32), input(31), input(30), input(29), input(28), 
      input(27), input(26), input(25), input(24), input(23), input(22), 
      input(21), input(20), input(19), input(18), input(17), input(16), 
      input(15), input(14), input(13), input(12), input(11), input(10), 
      input(9), input(8), input(7), input(6), input(5), input(4), input(3), 
      input(2), input(1), input(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity shifter_N64_5 is

   port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
         std_logic_vector (63 downto 0));

end shifter_N64_5;

architecture SYN_beh of shifter_N64_5 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, shiftLeftOnePos_30_port, shiftLeftOnePos_34_port, 
      shiftLeftOnePos_38_port, shiftLeftOnePos_42_port, shiftLeftOnePos_46_port
      , shiftLeftOnePos_50_port, shiftLeftOnePos_54_port : std_logic;

begin
   shiftLeftOnePos <= ( input(62), input(61), input(60), input(59), input(58), 
      input(57), input(56), input(55), input(54), shiftLeftOnePos_54_port, 
      input(52), input(51), input(50), shiftLeftOnePos_50_port, input(48), 
      input(47), input(46), shiftLeftOnePos_46_port, input(44), input(43), 
      input(42), shiftLeftOnePos_42_port, input(40), input(39), input(38), 
      shiftLeftOnePos_38_port, input(36), input(35), input(34), 
      shiftLeftOnePos_34_port, input(32), input(31), input(30), 
      shiftLeftOnePos_30_port, input(28), input(27), input(26), input(25), 
      input(24), input(23), input(22), input(21), input(20), input(19), 
      input(18), input(17), input(16), input(15), input(14), input(13), 
      input(12), input(11), input(10), input(9), input(8), input(7), input(6), 
      input(5), input(4), input(3), input(2), input(1), input(0), X_Logic0_port
      );
   
   X_Logic0_port <= '0';
   U2 : BUF_X1 port map( A => input(33), Z => shiftLeftOnePos_34_port);
   U3 : BUF_X1 port map( A => input(29), Z => shiftLeftOnePos_30_port);
   U4 : BUF_X1 port map( A => input(45), Z => shiftLeftOnePos_46_port);
   U5 : BUF_X1 port map( A => input(41), Z => shiftLeftOnePos_42_port);
   U6 : BUF_X1 port map( A => input(37), Z => shiftLeftOnePos_38_port);
   U7 : BUF_X1 port map( A => input(53), Z => shiftLeftOnePos_54_port);
   U8 : BUF_X1 port map( A => input(49), Z => shiftLeftOnePos_50_port);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity shifter_N64_4 is

   port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
         std_logic_vector (63 downto 0));

end shifter_N64_4;

architecture SYN_beh of shifter_N64_4 is

signal X_Logic0_port : std_logic;

begin
   shiftLeftOnePos <= ( input(62), input(61), input(60), input(59), input(58), 
      input(57), input(56), input(55), input(54), input(53), input(52), 
      input(51), input(50), input(49), input(48), input(47), input(46), 
      input(45), input(44), input(43), input(42), input(41), input(40), 
      input(39), input(38), input(37), input(36), input(35), input(34), 
      input(33), input(32), input(31), input(30), input(29), input(28), 
      input(27), input(26), input(25), input(24), input(23), input(22), 
      input(21), input(20), input(19), input(18), input(17), input(16), 
      input(15), input(14), input(13), input(12), input(11), input(10), 
      input(9), input(8), input(7), input(6), input(5), input(4), input(3), 
      input(2), input(1), input(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity shifter_N64_3 is

   port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
         std_logic_vector (63 downto 0));

end shifter_N64_3;

architecture SYN_beh of shifter_N64_3 is

signal X_Logic0_port : std_logic;

begin
   shiftLeftOnePos <= ( input(62), input(61), input(60), input(59), input(58), 
      input(57), input(56), input(55), input(54), input(53), input(52), 
      input(51), input(50), input(49), input(48), input(47), input(46), 
      input(45), input(44), input(43), input(42), input(41), input(40), 
      input(39), input(38), input(37), input(36), input(35), input(34), 
      input(33), input(32), input(31), input(30), input(29), input(28), 
      input(27), input(26), input(25), input(24), input(23), input(22), 
      input(21), input(20), input(19), input(18), input(17), input(16), 
      input(15), input(14), input(13), input(12), input(11), input(10), 
      input(9), input(8), input(7), input(6), input(5), input(4), input(3), 
      input(2), input(1), input(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity shifter_N64_2 is

   port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
         std_logic_vector (63 downto 0));

end shifter_N64_2;

architecture SYN_beh of shifter_N64_2 is

signal X_Logic0_port : std_logic;

begin
   shiftLeftOnePos <= ( input(62), input(61), input(60), input(59), input(58), 
      input(57), input(56), input(55), input(54), input(53), input(52), 
      input(51), input(50), input(49), input(48), input(47), input(46), 
      input(45), input(44), input(43), input(42), input(41), input(40), 
      input(39), input(38), input(37), input(36), input(35), input(34), 
      input(33), input(32), input(31), input(30), input(29), input(28), 
      input(27), input(26), input(25), input(24), input(23), input(22), 
      input(21), input(20), input(19), input(18), input(17), input(16), 
      input(15), input(14), input(13), input(12), input(11), input(10), 
      input(9), input(8), input(7), input(6), input(5), input(4), input(3), 
      input(2), input(1), input(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity shifter_N64_1 is

   port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
         std_logic_vector (63 downto 0));

end shifter_N64_1;

architecture SYN_beh of shifter_N64_1 is

signal X_Logic0_port : std_logic;

begin
   shiftLeftOnePos <= ( input(62), input(61), input(60), input(59), input(58), 
      input(57), input(56), input(55), input(54), input(53), input(52), 
      input(51), input(50), input(49), input(48), input(47), input(46), 
      input(45), input(44), input(43), input(42), input(41), input(40), 
      input(39), input(38), input(37), input(36), input(35), input(34), 
      input(33), input(32), input(31), input(30), input(29), input(28), 
      input(27), input(26), input(25), input(24), input(23), input(22), 
      input(21), input(20), input(19), input(18), input(17), input(16), 
      input(15), input(14), input(13), input(12), input(11), input(10), 
      input(9), input(8), input(7), input(6), input(5), input(4), input(3), 
      input(2), input(1), input(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity RCA_N64_14 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_N64_14;

architecture SYN_STRUCTURAL of RCA_N64_14 is

   component FA_833
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_834
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_835
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_836
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_837
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_838
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_839
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_840
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_841
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_842
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_843
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_844
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_845
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_846
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_847
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_848
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_849
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_850
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_851
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_852
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_853
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_854
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_855
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_856
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_857
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_858
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_859
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_860
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_861
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_862
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_863
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_864
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_865
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_866
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_867
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_868
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_869
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_870
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_871
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_872
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_873
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_874
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_875
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_876
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_877
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_878
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_879
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_880
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_881
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_882
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_883
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_884
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_885
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_886
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_887
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_888
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_889
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_890
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_891
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_892
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_893
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_894
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_895
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_896
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_896 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_895 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_894 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_893 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_892 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_891 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_890 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_889 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_888 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_887 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_886 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_885 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_884 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_883 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_882 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_881 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_880 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_879 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_878 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_877 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_876 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_875 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_874 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_873 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_872 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_871 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_870 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_869 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_868 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_867 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_866 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_865 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_864 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_863 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_862 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_861 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_860 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_859 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_858 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_857 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_856 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_855 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_854 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_853 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_852 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_851 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_850 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_849 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_848 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_847 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_846 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_845 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_844 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_843 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_842 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_841 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_840 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_839 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_838 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_837 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_836 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_835 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_834 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_833 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity RCA_N64_13 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_N64_13;

architecture SYN_STRUCTURAL of RCA_N64_13 is

   component FA_769
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_770
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_771
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_772
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_773
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_774
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_775
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_776
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_777
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_778
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_779
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_780
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_781
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_782
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_783
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_784
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_785
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_786
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_787
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_788
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_789
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_790
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_791
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_792
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_793
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_794
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_795
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_796
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_797
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_798
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_799
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_800
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_801
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_802
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_803
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_804
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_805
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_806
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_807
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_808
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_809
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_810
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_811
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_812
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_813
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_814
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_815
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_816
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_817
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_818
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_819
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_820
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_821
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_822
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_823
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_824
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_825
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_826
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_827
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_828
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_829
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_830
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_831
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_832
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_832 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_831 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_830 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_829 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_828 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_827 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_826 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_825 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_824 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_823 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_822 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_821 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_820 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_819 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_818 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_817 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_816 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_815 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_814 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_813 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_812 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_811 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_810 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_809 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_808 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_807 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_806 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_805 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_804 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_803 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_802 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_801 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_800 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_799 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_798 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_797 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_796 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_795 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_794 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_793 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_792 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_791 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_790 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_789 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_788 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_787 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_786 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_785 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_784 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_783 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_782 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_781 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_780 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_779 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_778 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_777 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_776 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_775 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_774 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_773 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_772 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_771 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_770 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_769 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity RCA_N64_12 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_N64_12;

architecture SYN_STRUCTURAL of RCA_N64_12 is

   component FA_705
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_706
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_707
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_708
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_709
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_710
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_711
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_712
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_713
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_714
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_715
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_716
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_717
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_718
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_719
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_720
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_721
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_722
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_723
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_724
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_725
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_726
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_727
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_728
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_729
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_730
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_731
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_732
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_733
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_734
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_735
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_736
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_737
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_738
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_739
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_740
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_741
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_742
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_743
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_744
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_745
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_746
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_747
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_748
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_749
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_750
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_751
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_752
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_753
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_754
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_755
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_756
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_757
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_758
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_759
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_760
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_761
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_762
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_763
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_764
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_765
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_766
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_767
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_768
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_768 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_767 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_766 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_765 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_764 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_763 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_762 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_761 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_760 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_759 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_758 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_757 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_756 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_755 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_754 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_753 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_752 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_751 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_750 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_749 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_748 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_747 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_746 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_745 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_744 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_743 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_742 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_741 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_740 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_739 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_738 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_737 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_736 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_735 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_734 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_733 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_732 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_731 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_730 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_729 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_728 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_727 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_726 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_725 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_724 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_723 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_722 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_721 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_720 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_719 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_718 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_717 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_716 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_715 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_714 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_713 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_712 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_711 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_710 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_709 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_708 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_707 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_706 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_705 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity RCA_N64_11 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_N64_11;

architecture SYN_STRUCTURAL of RCA_N64_11 is

   component FA_641
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_642
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_643
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_644
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_645
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_646
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_647
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_648
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_649
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_650
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_651
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_652
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_653
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_654
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_655
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_656
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_657
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_658
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_659
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_660
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_661
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_662
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_663
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_664
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_665
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_666
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_667
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_668
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_669
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_670
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_671
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_672
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_673
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_674
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_675
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_676
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_677
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_678
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_679
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_680
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_681
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_682
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_683
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_684
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_685
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_686
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_687
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_688
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_689
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_690
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_691
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_692
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_693
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_694
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_695
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_696
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_697
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_698
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_699
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_700
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_701
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_702
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_703
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_704
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_704 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_703 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_702 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_701 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_700 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_699 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_698 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_697 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_696 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_695 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_694 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_693 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_692 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_691 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_690 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_689 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_688 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_687 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_686 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_685 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_684 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_683 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_682 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_681 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_680 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_679 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_678 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_677 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_676 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_675 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_674 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_673 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_672 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_671 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_670 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_669 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_668 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_667 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_666 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_665 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_664 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_663 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_662 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_661 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_660 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_659 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_658 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_657 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_656 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_655 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_654 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_653 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_652 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_651 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_650 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_649 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_648 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_647 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_646 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_645 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_644 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_643 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_642 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_641 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity RCA_N64_10 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_N64_10;

architecture SYN_STRUCTURAL of RCA_N64_10 is

   component FA_577
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_578
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_579
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_580
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_581
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_582
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_583
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_584
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_585
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_586
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_587
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_588
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_589
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_590
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_591
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_592
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_593
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_594
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_595
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_596
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_597
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_598
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_599
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_600
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_601
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_602
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_603
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_604
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_605
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_606
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_607
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_608
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_609
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_610
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_611
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_612
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_613
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_614
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_615
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_616
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_617
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_618
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_619
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_620
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_621
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_622
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_623
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_624
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_625
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_626
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_627
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_628
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_629
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_630
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_631
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_632
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_633
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_634
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_635
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_636
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_637
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_638
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_639
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_640
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_640 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_639 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_638 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_637 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_636 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_635 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_634 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_633 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_632 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_631 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_630 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_629 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_628 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_627 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_626 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_625 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_624 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_623 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_622 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_621 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_620 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_619 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_618 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_617 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_616 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_615 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_614 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_613 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_612 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_611 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_610 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_609 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_608 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_607 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_606 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_605 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_604 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_603 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_602 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_601 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_600 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_599 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_598 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_597 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_596 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_595 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_594 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_593 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_592 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_591 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_590 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_589 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_588 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_587 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_586 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_585 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_584 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_583 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_582 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_581 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_580 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_579 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_578 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_577 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity RCA_N64_9 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_N64_9;

architecture SYN_STRUCTURAL of RCA_N64_9 is

   component FA_513
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_514
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_515
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_516
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_517
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_518
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_519
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_520
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_521
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_522
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_523
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_524
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_525
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_526
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_527
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_528
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_529
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_530
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_531
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_532
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_533
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_534
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_535
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_536
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_537
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_538
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_539
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_540
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_541
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_542
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_543
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_544
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_545
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_546
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_547
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_548
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_549
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_550
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_551
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_552
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_553
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_554
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_555
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_556
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_557
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_558
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_559
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_560
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_561
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_562
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_563
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_564
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_565
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_566
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_567
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_568
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_569
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_570
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_571
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_572
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_573
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_574
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_575
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_576
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_576 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_575 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_574 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_573 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_572 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_571 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_570 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_569 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_568 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_567 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_566 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_565 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_564 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_563 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_562 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_561 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_560 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_559 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_558 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_557 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_556 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_555 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_554 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_553 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_552 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_551 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_550 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_549 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_548 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_547 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_546 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_545 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_544 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_543 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_542 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_541 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_540 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_539 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_538 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_537 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_536 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_535 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_534 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_533 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_532 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_531 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_530 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_529 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_528 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_527 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_526 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_525 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_524 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_523 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_522 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_521 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_520 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_519 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_518 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_517 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_516 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_515 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_514 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_513 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity RCA_N64_8 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_N64_8;

architecture SYN_STRUCTURAL of RCA_N64_8 is

   component FA_449
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_450
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_451
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_452
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_453
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_454
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_455
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_456
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_457
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_458
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_459
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_460
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_461
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_462
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_463
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_464
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_465
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_466
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_467
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_468
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_469
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_470
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_471
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_472
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_473
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_474
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_475
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_476
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_477
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_478
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_479
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_480
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_481
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_482
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_483
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_484
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_485
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_486
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_487
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_488
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_489
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_490
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_491
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_492
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_493
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_494
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_495
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_496
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_497
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_498
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_499
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_500
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_501
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_502
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_503
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_504
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_505
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_506
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_507
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_508
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_509
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_510
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_511
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_512
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_512 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_511 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_510 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_509 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_508 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_507 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_506 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_505 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_504 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_503 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_502 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_501 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_500 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_499 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_498 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_497 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_496 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_495 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_494 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_493 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_492 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_491 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_490 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_489 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_488 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_487 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_486 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_485 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_484 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_483 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_482 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_481 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_480 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_479 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_478 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_477 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_476 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_475 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_474 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_473 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_472 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_471 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_470 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_469 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_468 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_467 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_466 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_465 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_464 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_463 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_462 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_461 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_460 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_459 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_458 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_457 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_456 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_455 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_454 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_453 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_452 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_451 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_450 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_449 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity RCA_N64_7 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_N64_7;

architecture SYN_STRUCTURAL of RCA_N64_7 is

   component FA_385
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_386
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_387
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_388
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_389
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_390
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_391
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_392
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_393
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_394
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_395
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_396
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_397
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_398
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_399
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_400
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_401
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_402
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_403
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_404
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_405
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_406
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_407
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_408
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_409
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_410
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_411
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_412
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_413
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_414
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_415
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_416
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_417
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_418
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_419
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_420
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_421
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_422
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_423
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_424
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_425
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_426
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_427
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_428
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_429
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_430
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_431
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_432
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_433
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_434
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_435
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_436
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_437
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_438
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_439
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_440
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_441
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_442
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_443
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_444
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_445
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_446
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_447
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_448
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_448 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_447 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_446 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_445 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_444 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_443 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_442 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_441 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_440 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_439 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_438 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_437 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_436 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_435 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_434 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_433 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_432 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_431 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_430 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_429 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_428 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_427 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_426 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_425 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_424 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_423 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_422 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_421 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_420 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_419 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_418 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_417 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_416 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_415 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_414 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_413 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_412 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_411 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_410 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_409 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_408 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_407 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_406 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_405 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_404 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_403 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_402 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_401 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_400 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_399 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_398 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_397 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_396 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_395 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_394 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_393 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_392 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_391 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_390 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_389 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_388 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_387 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_386 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_385 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity RCA_N64_6 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_N64_6;

architecture SYN_STRUCTURAL of RCA_N64_6 is

   component FA_321
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_322
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_323
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_324
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_325
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_326
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_327
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_328
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_329
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_330
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_331
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_332
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_333
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_334
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_335
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_336
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_337
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_338
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_339
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_340
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_341
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_342
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_343
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_344
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_345
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_346
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_347
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_348
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_349
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_350
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_351
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_352
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_353
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_354
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_355
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_356
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_357
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_358
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_359
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_360
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_361
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_362
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_363
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_364
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_365
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_366
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_367
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_368
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_369
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_370
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_371
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_372
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_373
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_374
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_375
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_376
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_377
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_378
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_379
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_380
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_381
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_382
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_383
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_384
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_384 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_383 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_382 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_381 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_380 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_379 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_378 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_377 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_376 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_375 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_374 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_373 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_372 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_371 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_370 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_369 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_368 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_367 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_366 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_365 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_364 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_363 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_362 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_361 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_360 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_359 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_358 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_357 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_356 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_355 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_354 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_353 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_352 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_351 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_350 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_349 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_348 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_347 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_346 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_345 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_344 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_343 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_342 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_341 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_340 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_339 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_338 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_337 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_336 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_335 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_334 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_333 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_332 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_331 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_330 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_329 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_328 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_327 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_326 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_325 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_324 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_323 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_322 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_321 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity RCA_N64_5 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_N64_5;

architecture SYN_STRUCTURAL of RCA_N64_5 is

   component FA_257
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_258
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_259
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_260
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_261
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_262
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_263
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_264
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_265
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_266
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_267
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_268
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_269
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_270
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_271
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_272
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_273
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_274
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_275
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_276
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_277
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_278
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_279
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_280
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_281
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_282
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_283
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_284
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_285
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_286
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_287
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_288
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_289
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_290
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_291
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_292
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_293
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_294
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_295
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_296
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_297
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_298
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_299
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_300
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_301
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_302
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_303
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_304
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_305
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_306
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_307
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_308
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_309
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_310
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_311
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_312
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_313
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_314
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_315
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_316
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_317
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_318
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_319
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_320
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_320 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_319 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_318 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_317 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_316 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_315 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_314 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_313 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_312 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_311 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_310 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_309 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_308 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_307 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_306 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_305 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_304 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_303 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_302 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_301 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_300 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_299 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_298 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_297 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_296 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_295 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_294 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_293 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_292 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_291 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_290 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_289 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_288 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_287 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_286 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_285 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_284 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_283 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_282 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_281 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_280 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_279 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_278 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_277 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_276 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_275 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_274 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_273 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_272 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_271 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_270 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_269 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_268 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_267 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_266 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_265 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_264 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_263 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_262 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_261 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_260 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_259 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_258 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_257 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity RCA_N64_4 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_N64_4;

architecture SYN_STRUCTURAL of RCA_N64_4 is

   component FA_193
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_194
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_195
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_196
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_197
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_198
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_199
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_200
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_201
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_202
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_203
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_204
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_205
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_206
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_207
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_208
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_209
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_210
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_211
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_212
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_213
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_214
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_215
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_216
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_217
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_218
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_219
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_220
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_221
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_222
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_223
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_224
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_225
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_226
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_227
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_228
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_229
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_230
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_231
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_232
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_233
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_234
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_235
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_236
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_237
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_238
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_239
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_240
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_241
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_242
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_243
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_244
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_245
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_246
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_247
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_248
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_249
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_250
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_251
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_252
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_253
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_254
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_255
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_256
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_256 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_255 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_254 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_253 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_252 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_251 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_250 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_249 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_248 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_247 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_246 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_245 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_244 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_243 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_242 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_241 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_240 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_239 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_238 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_237 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_236 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_235 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_234 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_233 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_232 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_231 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_230 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_229 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_228 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_227 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_226 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_225 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_224 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_223 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_222 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_221 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_220 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_219 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_218 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_217 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_216 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_215 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_214 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_213 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_212 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_211 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_210 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_209 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_208 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_207 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_206 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_205 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_204 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_203 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_202 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_201 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_200 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_199 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_198 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_197 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_196 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_195 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_194 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_193 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity RCA_N64_3 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_N64_3;

architecture SYN_STRUCTURAL of RCA_N64_3 is

   component FA_129
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_130
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_131
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_132
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_133
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_134
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_135
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_136
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_137
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_138
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_139
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_140
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_141
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_142
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_143
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_144
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_145
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_146
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_147
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_148
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_149
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_150
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_151
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_152
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_153
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_154
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_155
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_156
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_157
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_158
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_159
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_160
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_161
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_162
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_163
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_164
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_165
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_166
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_167
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_168
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_169
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_170
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_171
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_172
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_173
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_174
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_175
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_176
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_177
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_178
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_179
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_180
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_181
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_182
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_183
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_184
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_185
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_186
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_187
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_188
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_189
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_190
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_191
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_192
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_192 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_191 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_190 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_189 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_188 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_187 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_186 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_185 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_184 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_183 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_182 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_181 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_180 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_179 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_178 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_177 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_176 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_175 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_174 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_173 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_172 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_171 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_170 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_169 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_168 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_167 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_166 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_165 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_164 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_163 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_162 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_161 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_160 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_159 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_158 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_157 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_156 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_155 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_154 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_153 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_152 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_151 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_150 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_149 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_148 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_147 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_146 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_145 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_144 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_143 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_142 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_141 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_140 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_139 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_138 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_137 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_136 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_135 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_134 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_133 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_132 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_131 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_130 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_129 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity RCA_N64_2 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_N64_2;

architecture SYN_STRUCTURAL of RCA_N64_2 is

   component FA_65
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_66
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_67
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_68
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_69
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_70
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_71
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_72
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_73
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_74
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_75
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_76
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_77
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_78
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_79
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_80
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_81
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_82
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_83
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_84
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_85
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_86
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_87
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_88
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_89
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_90
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_91
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_92
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_93
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_94
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_95
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_96
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_97
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_98
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_99
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_100
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_101
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_102
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_103
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_104
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_105
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_106
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_107
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_108
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_109
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_110
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_111
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_112
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_113
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_114
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_115
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_116
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_117
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_118
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_119
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_120
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_121
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_122
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_123
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_124
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_125
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_126
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_127
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_128
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_128 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_127 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_126 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_125 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_124 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_123 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_122 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_121 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_120 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_119 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_118 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_117 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_116 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_115 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_114 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_113 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_112 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_111 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_110 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_109 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_108 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_107 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_106 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_105 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_104 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_103 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_102 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_101 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_100 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_99 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_98 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_97 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_96 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_95 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_94 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_93 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_92 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_91 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_90 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_89 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_88 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_87 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_86 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_85 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_84 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_83 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_82 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_81 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_80 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_79 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_78 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_77 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_76 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_75 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_74 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_73 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_72 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_71 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_70 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_69 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_68 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_67 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_66 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_65 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity RCA_N64_1 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_N64_1;

architecture SYN_STRUCTURAL of RCA_N64_1 is

   component FA_1
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_3
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_4
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_5
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_6
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_7
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_8
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_9
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_10
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_11
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_12
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_13
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_14
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_15
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_16
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_17
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_18
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_19
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_20
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_21
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_22
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_23
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_24
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_25
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_26
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_27
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_28
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_29
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_30
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_31
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_32
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_33
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_34
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_35
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_36
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_37
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_38
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_39
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_40
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_41
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_42
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_43
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_44
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_45
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_46
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_47
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_48
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_49
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_50
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_51
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_52
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_53
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_54
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_55
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_56
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_57
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_58
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_59
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_60
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_61
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_62
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_63
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_64
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_64 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_63 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_62 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_61 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => CTMP_4_port);
   FAI_5 : FA_60 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4), 
                           Co => CTMP_5_port);
   FAI_6 : FA_59 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5), 
                           Co => CTMP_6_port);
   FAI_7 : FA_58 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6), 
                           Co => CTMP_7_port);
   FAI_8 : FA_57 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7), 
                           Co => CTMP_8_port);
   FAI_9 : FA_56 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8), 
                           Co => CTMP_9_port);
   FAI_10 : FA_55 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9),
                           Co => CTMP_10_port);
   FAI_11 : FA_54 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_53 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_52 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_51 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_50 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_49 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_48 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_47 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_46 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_45 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_44 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_43 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_42 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_41 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_40 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_39 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_38 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_37 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_36 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_35 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_34 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_33 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_32 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_31 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_30 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_29 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_28 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_27 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_26 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_25 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_24 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_23 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_22 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_21 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_20 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_19 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_18 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_17 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_16 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_15 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_14 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_13 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_12 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_11 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_10 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_9 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_8 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_7 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_6 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_5 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_4 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_3 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_2 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_1 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity MUX_GENERIC_N64_RADIX3_15 is

   port( plusA, minusA, plus2A, minus2A : in std_logic_vector (63 downto 0);  
         SEL : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (63 
         downto 0));

end MUX_GENERIC_N64_RADIX3_15;

architecture SYN_beh of MUX_GENERIC_N64_RADIX3_15 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X8
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component TBUF_X2
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   component TBUF_X4
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   component TBUF_X1
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   signal net85116, net85117, net89097, net89095, net89093, net93069, net93945,
      net94659, net94671, n272, n273, n274, n275, n276, n277, n278, n279, n280,
      n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, 
      n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, 
      n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, 
      n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, 
      n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, 
      n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, 
      n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, 
      n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, 
      n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, 
      n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, 
      n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, 
      n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, 
      n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, 
      n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, 
      n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, 
      n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, 
      n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, 
      n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, 
      n497 : std_logic;

begin
   
   Y_tri_46_inst : TBUF_X1 port map( A => n451, EN => n280, Z => Y(46));
   Y_tri_48_inst : TBUF_X1 port map( A => n449, EN => net89095, Z => Y(48));
   Y_tri_52_inst : TBUF_X1 port map( A => n445, EN => net89095, Z => Y(52));
   Y_tri_53_inst : TBUF_X1 port map( A => n444, EN => n284, Z => Y(53));
   Y_tri_55_inst : TBUF_X1 port map( A => n442, EN => n280, Z => Y(55));
   Y_tri_57_inst : TBUF_X1 port map( A => n440, EN => n279, Z => Y(57));
   Y_tri_58_inst : TBUF_X1 port map( A => n439, EN => n284, Z => Y(58));
   Y_tri_60_inst : TBUF_X1 port map( A => n437, EN => n280, Z => Y(60));
   Y_tri_62_inst : TBUF_X1 port map( A => n435, EN => n280, Z => Y(62));
   Y_tri_63_inst : TBUF_X1 port map( A => n434, EN => n284, Z => Y(63));
   Y_tri_31_inst : TBUF_X1 port map( A => n466, EN => n284, Z => Y(31));
   Y_tri_14_inst : TBUF_X1 port map( A => n483, EN => n280, Z => Y(14));
   Y_tri_13_inst : TBUF_X1 port map( A => n484, EN => n280, Z => Y(13));
   Y_tri_15_inst : TBUF_X1 port map( A => n482, EN => net89095, Z => Y(15));
   Y_tri_16_inst : TBUF_X1 port map( A => n481, EN => n280, Z => Y(16));
   Y_tri_17_inst : TBUF_X1 port map( A => n480, EN => n280, Z => Y(17));
   Y_tri_18_inst : TBUF_X1 port map( A => n479, EN => n280, Z => Y(18));
   Y_tri_19_inst : TBUF_X1 port map( A => n478, EN => n280, Z => Y(19));
   Y_tri_20_inst : TBUF_X1 port map( A => n477, EN => n280, Z => Y(20));
   Y_tri_21_inst : TBUF_X1 port map( A => n476, EN => n280, Z => Y(21));
   Y_tri_22_inst : TBUF_X1 port map( A => n475, EN => n280, Z => Y(22));
   Y_tri_23_inst : TBUF_X1 port map( A => n474, EN => n280, Z => Y(23));
   Y_tri_24_inst : TBUF_X1 port map( A => n473, EN => n280, Z => Y(24));
   Y_tri_25_inst : TBUF_X1 port map( A => n472, EN => n280, Z => Y(25));
   Y_tri_26_inst : TBUF_X1 port map( A => n471, EN => n280, Z => Y(26));
   Y_tri_39_inst : TBUF_X1 port map( A => n458, EN => n280, Z => Y(39));
   Y_tri_27_inst : TBUF_X1 port map( A => n470, EN => n284, Z => Y(27));
   Y_tri_28_inst : TBUF_X1 port map( A => n469, EN => n280, Z => Y(28));
   Y_tri_37_inst : TBUF_X1 port map( A => n460, EN => n280, Z => Y(37));
   Y_tri_33_inst : TBUF_X1 port map( A => n464, EN => n280, Z => Y(33));
   Y_tri_29_inst : TBUF_X1 port map( A => n468, EN => n284, Z => Y(29));
   Y_tri_34_inst : TBUF_X1 port map( A => n463, EN => n284, Z => Y(34));
   Y_tri_30_inst : TBUF_X1 port map( A => n467, EN => n280, Z => Y(30));
   Y_tri_35_inst : TBUF_X1 port map( A => n462, EN => n280, Z => Y(35));
   Y_tri_41_inst : TBUF_X1 port map( A => n456, EN => n279, Z => Y(41));
   Y_tri_43_inst : TBUF_X1 port map( A => n454, EN => n284, Z => Y(43));
   Y_tri_44_inst : TBUF_X1 port map( A => n453, EN => net89095, Z => Y(44));
   Y_tri_47_inst : TBUF_X1 port map( A => n450, EN => n279, Z => Y(47));
   Y_tri_49_inst : TBUF_X1 port map( A => n448, EN => n284, Z => Y(49));
   Y_tri_50_inst : TBUF_X1 port map( A => n447, EN => n280, Z => Y(50));
   Y_tri_51_inst : TBUF_X1 port map( A => n446, EN => n279, Z => Y(51));
   Y_tri_54_inst : TBUF_X1 port map( A => n443, EN => n279, Z => Y(54));
   Y_tri_56_inst : TBUF_X1 port map( A => n441, EN => net89095, Z => Y(56));
   Y_tri_59_inst : TBUF_X1 port map( A => n438, EN => net89095, Z => Y(59));
   Y_tri_61_inst : TBUF_X1 port map( A => n436, EN => n279, Z => Y(61));
   Y_tri_36_inst : TBUF_X1 port map( A => n461, EN => n284, Z => Y(36));
   Y_tri_38_inst : TBUF_X1 port map( A => n459, EN => n284, Z => Y(38));
   Y_tri_32_inst : TBUF_X1 port map( A => n465, EN => n284, Z => Y(32));
   Y_tri_40_inst : TBUF_X1 port map( A => n457, EN => n284, Z => Y(40));
   Y_tri_42_inst : TBUF_X1 port map( A => n455, EN => n280, Z => Y(42));
   Y_tri_45_inst : TBUF_X1 port map( A => n452, EN => n284, Z => Y(45));
   Y_tri_4_inst : TBUF_X1 port map( A => n493, EN => n283, Z => Y(4));
   Y_tri_3_inst : TBUF_X1 port map( A => n494, EN => net89093, Z => Y(3));
   Y_tri_5_inst : TBUF_X1 port map( A => n492, EN => n279, Z => Y(5));
   Y_tri_6_inst : TBUF_X1 port map( A => n491, EN => net89097, Z => Y(6));
   Y_tri_7_inst : TBUF_X1 port map( A => n490, EN => net89097, Z => Y(7));
   Y_tri_8_inst : TBUF_X1 port map( A => n489, EN => net89095, Z => Y(8));
   Y_tri_1_inst : TBUF_X1 port map( A => n496, EN => net93069, Z => Y(1));
   Y_tri_12_inst : TBUF_X1 port map( A => n485, EN => n280, Z => Y(12));
   Y_tri_11_inst : TBUF_X1 port map( A => n486, EN => n280, Z => Y(11));
   Y_tri_10_inst : TBUF_X1 port map( A => n487, EN => n284, Z => Y(10));
   Y_tri_9_inst : TBUF_X1 port map( A => n488, EN => n279, Z => Y(9));
   Y_tri_2_inst : TBUF_X4 port map( A => n495, EN => net89093, Z => Y(2));
   Y_tri_0_inst : TBUF_X2 port map( A => n497, EN => net93069, Z => Y(0));
   U2 : BUF_X1 port map( A => n283, Z => n279);
   U3 : BUF_X1 port map( A => n429, Z => n282);
   U4 : BUF_X1 port map( A => n282, Z => n292);
   U5 : NOR3_X2 port map( A1 => net85117, A2 => n273, A3 => net85116, ZN => 
                           n278);
   U6 : BUF_X2 port map( A => n278, Z => n285);
   U7 : AND3_X1 port map( A1 => net93945, A2 => net94671, A3 => net85116, ZN =>
                           n430);
   U8 : INV_X1 port map( A => net93945, ZN => n272);
   U9 : AND2_X2 port map( A1 => n275, A2 => SEL(2), ZN => net93069);
   U10 : BUF_X2 port map( A => SEL(2), Z => n273);
   U11 : AND2_X2 port map( A1 => n273, A2 => n276, ZN => net89093);
   U12 : CLKBUF_X1 port map( A => SEL(0), Z => n274);
   U13 : AND2_X1 port map( A1 => net94659, A2 => n273, ZN => n431);
   U14 : INV_X1 port map( A => SEL(1), ZN => n277);
   U15 : CLKBUF_X1 port map( A => n272, Z => net85117);
   U16 : OR2_X1 port map( A1 => SEL(1), A2 => SEL(0), ZN => n275);
   U17 : INV_X1 port map( A => n275, ZN => net94659);
   U18 : INV_X1 port map( A => net94659, ZN => n276);
   U19 : CLKBUF_X3 port map( A => n431, Z => n300);
   U20 : INV_X1 port map( A => SEL(2), ZN => net94671);
   U21 : NOR2_X1 port map( A1 => net94659, A2 => net94671, ZN => n283);
   U22 : INV_X1 port map( A => n277, ZN => net93945);
   U23 : BUF_X4 port map( A => n283, Z => n280);
   U24 : BUF_X2 port map( A => net89093, Z => net89095);
   U25 : CLKBUF_X1 port map( A => n283, Z => n284);
   U26 : NOR3_X1 port map( A1 => net85117, A2 => n273, A3 => net85116, ZN => 
                           n428);
   U27 : BUF_X8 port map( A => n281, Z => n293);
   U28 : CLKBUF_X1 port map( A => net89093, Z => net89097);
   U29 : BUF_X2 port map( A => n430, Z => n281);
   U30 : CLKBUF_X1 port map( A => n281, Z => n294);
   U31 : CLKBUF_X1 port map( A => n281, Z => n295);
   U32 : CLKBUF_X1 port map( A => n281, Z => n296);
   U33 : CLKBUF_X2 port map( A => n282, Z => n290);
   U34 : CLKBUF_X1 port map( A => n431, Z => n297);
   U35 : CLKBUF_X1 port map( A => n431, Z => n298);
   U36 : CLKBUF_X1 port map( A => n278, Z => n286);
   U37 : CLKBUF_X1 port map( A => n431, Z => n299);
   U38 : CLKBUF_X1 port map( A => n278, Z => n287);
   U39 : CLKBUF_X1 port map( A => n278, Z => n288);
   U40 : NAND2_X1 port map( A1 => n319, A2 => n318, ZN => n489);
   U41 : AOI22_X1 port map( A1 => plusA(8), A2 => n292, B1 => plus2A(8), B2 => 
                           n288, ZN => n319);
   U42 : NAND2_X1 port map( A1 => n311, A2 => n310, ZN => n493);
   U43 : AOI22_X1 port map( A1 => plusA(4), A2 => n291, B1 => plus2A(4), B2 => 
                           n289, ZN => n311);
   U44 : NAND2_X1 port map( A1 => n327, A2 => n326, ZN => n485);
   U45 : AOI22_X1 port map( A1 => plusA(12), A2 => n290, B1 => plus2A(12), B2 
                           => n285, ZN => n327);
   U46 : AOI22_X1 port map( A1 => minus2A(12), A2 => n297, B1 => minusA(12), B2
                           => n293, ZN => n326);
   U47 : NAND2_X1 port map( A1 => n315, A2 => n314, ZN => n491);
   U48 : AOI22_X1 port map( A1 => plusA(6), A2 => n291, B1 => plus2A(6), B2 => 
                           n286, ZN => n315);
   U49 : NAND2_X1 port map( A1 => n323, A2 => n322, ZN => n487);
   U50 : AOI22_X1 port map( A1 => plusA(10), A2 => n290, B1 => plus2A(10), B2 
                           => n288, ZN => n323);
   U51 : NAND2_X1 port map( A1 => n308, A2 => n309, ZN => n494);
   U52 : AOI22_X1 port map( A1 => plusA(3), A2 => n282, B1 => plus2A(3), B2 => 
                           n278, ZN => n309);
   U53 : NAND2_X1 port map( A1 => n313, A2 => n312, ZN => n492);
   U54 : AOI22_X1 port map( A1 => plusA(5), A2 => n291, B1 => plus2A(5), B2 => 
                           n285, ZN => n313);
   U55 : NAND2_X1 port map( A1 => n321, A2 => n320, ZN => n488);
   U56 : AOI22_X1 port map( A1 => plusA(9), A2 => n290, B1 => plus2A(9), B2 => 
                           n288, ZN => n321);
   U57 : NAND2_X1 port map( A1 => n317, A2 => n316, ZN => n490);
   U58 : AOI22_X1 port map( A1 => plusA(7), A2 => n292, B1 => plus2A(7), B2 => 
                           n287, ZN => n317);
   U59 : NAND2_X1 port map( A1 => n325, A2 => n324, ZN => n486);
   U60 : AOI22_X1 port map( A1 => plusA(11), A2 => n290, B1 => plus2A(11), B2 
                           => n288, ZN => n325);
   U61 : INV_X1 port map( A => n274, ZN => net85116);
   U62 : NAND2_X1 port map( A1 => n369, A2 => n368, ZN => n464);
   U63 : AOI22_X1 port map( A1 => plusA(33), A2 => n292, B1 => plus2A(33), B2 
                           => n286, ZN => n369);
   U64 : AOI22_X1 port map( A1 => minus2A(33), A2 => n298, B1 => minusA(33), B2
                           => n293, ZN => n368);
   U65 : NAND2_X1 port map( A1 => n371, A2 => n370, ZN => n463);
   U66 : AOI22_X1 port map( A1 => plusA(34), A2 => n290, B1 => plus2A(34), B2 
                           => n286, ZN => n371);
   U67 : AOI22_X1 port map( A1 => minus2A(34), A2 => n298, B1 => minusA(34), B2
                           => n293, ZN => n370);
   U68 : NAND2_X1 port map( A1 => n421, A2 => n420, ZN => n438);
   U69 : AOI22_X1 port map( A1 => plusA(59), A2 => n290, B1 => plus2A(59), B2 
                           => n288, ZN => n421);
   U70 : AOI22_X1 port map( A1 => minus2A(59), A2 => n300, B1 => minusA(59), B2
                           => n293, ZN => n420);
   U71 : NAND2_X1 port map( A1 => n389, A2 => n388, ZN => n454);
   U72 : AOI22_X1 port map( A1 => plusA(43), A2 => n292, B1 => plus2A(43), B2 
                           => n287, ZN => n389);
   U73 : AOI22_X1 port map( A1 => minus2A(43), A2 => n299, B1 => minusA(43), B2
                           => n293, ZN => n388);
   U74 : NAND2_X1 port map( A1 => n381, A2 => n380, ZN => n458);
   U75 : AOI22_X1 port map( A1 => plusA(39), A2 => n292, B1 => plus2A(39), B2 
                           => n287, ZN => n381);
   U76 : AOI22_X1 port map( A1 => minus2A(39), A2 => n299, B1 => minusA(39), B2
                           => n293, ZN => n380);
   U77 : NAND2_X1 port map( A1 => n419, A2 => n418, ZN => n439);
   U78 : AOI22_X1 port map( A1 => plusA(58), A2 => n292, B1 => plus2A(58), B2 
                           => n288, ZN => n419);
   U79 : AOI22_X1 port map( A1 => minus2A(58), A2 => n300, B1 => minusA(58), B2
                           => n293, ZN => n418);
   U80 : NAND2_X1 port map( A1 => n403, A2 => n402, ZN => n447);
   U81 : AOI22_X1 port map( A1 => plusA(50), A2 => n292, B1 => plus2A(50), B2 
                           => n288, ZN => n403);
   U82 : AOI22_X1 port map( A1 => minus2A(50), A2 => n300, B1 => minusA(50), B2
                           => n296, ZN => n402);
   U83 : NAND2_X1 port map( A1 => n401, A2 => n400, ZN => n448);
   U84 : AOI22_X1 port map( A1 => plusA(49), A2 => n292, B1 => plus2A(49), B2 
                           => n288, ZN => n401);
   U85 : AOI22_X1 port map( A1 => minus2A(49), A2 => n300, B1 => minusA(49), B2
                           => n293, ZN => n400);
   U86 : NAND2_X1 port map( A1 => n335, A2 => n334, ZN => n481);
   U87 : AOI22_X1 port map( A1 => plusA(16), A2 => n290, B1 => plus2A(16), B2 
                           => n285, ZN => n335);
   U88 : AOI22_X1 port map( A1 => minus2A(16), A2 => n297, B1 => minusA(16), B2
                           => n293, ZN => n334);
   U89 : NAND2_X1 port map( A1 => n343, A2 => n342, ZN => n477);
   U90 : AOI22_X1 port map( A1 => plusA(20), A2 => n290, B1 => plus2A(20), B2 
                           => n285, ZN => n343);
   U91 : AOI22_X1 port map( A1 => minus2A(20), A2 => n297, B1 => minusA(20), B2
                           => n293, ZN => n342);
   U92 : NAND2_X1 port map( A1 => n351, A2 => n350, ZN => n473);
   U93 : AOI22_X1 port map( A1 => plusA(24), A2 => n290, B1 => plus2A(24), B2 
                           => n286, ZN => n351);
   U94 : AOI22_X1 port map( A1 => minus2A(24), A2 => n298, B1 => minusA(24), B2
                           => n293, ZN => n350);
   U95 : NAND2_X1 port map( A1 => n359, A2 => n358, ZN => n469);
   U96 : AOI22_X1 port map( A1 => plusA(28), A2 => n290, B1 => plus2A(28), B2 
                           => n286, ZN => n359);
   U97 : AOI22_X1 port map( A1 => minus2A(28), A2 => n298, B1 => minusA(28), B2
                           => n293, ZN => n358);
   U98 : NAND2_X1 port map( A1 => n367, A2 => n366, ZN => n465);
   U99 : AOI22_X1 port map( A1 => plusA(32), A2 => n290, B1 => plus2A(32), B2 
                           => n286, ZN => n367);
   U100 : AOI22_X1 port map( A1 => minus2A(32), A2 => n298, B1 => minusA(32), 
                           B2 => n293, ZN => n366);
   U101 : NAND2_X1 port map( A1 => n399, A2 => n398, ZN => n449);
   U102 : AOI22_X1 port map( A1 => plusA(48), A2 => n290, B1 => plus2A(48), B2 
                           => n288, ZN => n399);
   U103 : AOI22_X1 port map( A1 => minus2A(48), A2 => n300, B1 => minusA(48), 
                           B2 => n293, ZN => n398);
   U104 : NAND2_X1 port map( A1 => n331, A2 => n330, ZN => n483);
   U105 : AOI22_X1 port map( A1 => plusA(14), A2 => n290, B1 => plus2A(14), B2 
                           => n285, ZN => n331);
   U106 : AOI22_X1 port map( A1 => minus2A(14), A2 => n297, B1 => minusA(14), 
                           B2 => n293, ZN => n330);
   U107 : NAND2_X1 port map( A1 => n363, A2 => n362, ZN => n467);
   U108 : AOI22_X1 port map( A1 => plusA(30), A2 => n290, B1 => plus2A(30), B2 
                           => n286, ZN => n363);
   U109 : AOI22_X1 port map( A1 => minus2A(30), A2 => n298, B1 => minusA(30), 
                           B2 => n293, ZN => n362);
   U110 : NAND2_X1 port map( A1 => n339, A2 => n338, ZN => n479);
   U111 : AOI22_X1 port map( A1 => plusA(18), A2 => n290, B1 => plus2A(18), B2 
                           => n285, ZN => n339);
   U112 : AOI22_X1 port map( A1 => minus2A(18), A2 => n297, B1 => minusA(18), 
                           B2 => n293, ZN => n338);
   U113 : NAND2_X1 port map( A1 => n347, A2 => n346, ZN => n475);
   U114 : AOI22_X1 port map( A1 => plusA(22), A2 => n290, B1 => plus2A(22), B2 
                           => n285, ZN => n347);
   U115 : AOI22_X1 port map( A1 => minus2A(22), A2 => n297, B1 => minusA(22), 
                           B2 => n293, ZN => n346);
   U116 : NAND2_X1 port map( A1 => n355, A2 => n354, ZN => n471);
   U117 : AOI22_X1 port map( A1 => plusA(26), A2 => n290, B1 => plus2A(26), B2 
                           => n286, ZN => n355);
   U118 : AOI22_X1 port map( A1 => minus2A(26), A2 => n298, B1 => minusA(26), 
                           B2 => n293, ZN => n354);
   U119 : NAND2_X1 port map( A1 => n383, A2 => n382, ZN => n457);
   U120 : AOI22_X1 port map( A1 => plusA(40), A2 => n290, B1 => plus2A(40), B2 
                           => n287, ZN => n383);
   U121 : AOI22_X1 port map( A1 => minus2A(40), A2 => n299, B1 => minusA(40), 
                           B2 => n293, ZN => n382);
   U122 : NAND2_X1 port map( A1 => n379, A2 => n378, ZN => n459);
   U123 : AOI22_X1 port map( A1 => plusA(38), A2 => n290, B1 => plus2A(38), B2 
                           => n287, ZN => n379);
   U124 : AOI22_X1 port map( A1 => minus2A(38), A2 => n299, B1 => minusA(38), 
                           B2 => n293, ZN => n378);
   U125 : NAND2_X1 port map( A1 => n329, A2 => n328, ZN => n484);
   U126 : AOI22_X1 port map( A1 => plusA(13), A2 => n290, B1 => plus2A(13), B2 
                           => n285, ZN => n329);
   U127 : AOI22_X1 port map( A1 => minus2A(13), A2 => n297, B1 => minusA(13), 
                           B2 => n293, ZN => n328);
   U128 : NAND2_X1 port map( A1 => n337, A2 => n336, ZN => n480);
   U129 : AOI22_X1 port map( A1 => plusA(17), A2 => n290, B1 => plus2A(17), B2 
                           => n285, ZN => n337);
   U130 : AOI22_X1 port map( A1 => minus2A(17), A2 => n297, B1 => minusA(17), 
                           B2 => n293, ZN => n336);
   U131 : NAND2_X1 port map( A1 => n345, A2 => n344, ZN => n476);
   U132 : AOI22_X1 port map( A1 => plusA(21), A2 => n290, B1 => plus2A(21), B2 
                           => n285, ZN => n345);
   U133 : AOI22_X1 port map( A1 => minus2A(21), A2 => n297, B1 => minusA(21), 
                           B2 => n293, ZN => n344);
   U134 : NAND2_X1 port map( A1 => n353, A2 => n352, ZN => n472);
   U135 : AOI22_X1 port map( A1 => plusA(25), A2 => n290, B1 => plus2A(25), B2 
                           => n286, ZN => n353);
   U136 : AOI22_X1 port map( A1 => minus2A(25), A2 => n298, B1 => minusA(25), 
                           B2 => n293, ZN => n352);
   U137 : NAND2_X1 port map( A1 => n361, A2 => n360, ZN => n468);
   U138 : AOI22_X1 port map( A1 => plusA(29), A2 => n290, B1 => plus2A(29), B2 
                           => n286, ZN => n361);
   U139 : AOI22_X1 port map( A1 => minus2A(29), A2 => n298, B1 => minusA(29), 
                           B2 => n293, ZN => n360);
   U140 : NAND2_X1 port map( A1 => n411, A2 => n410, ZN => n443);
   U141 : AOI22_X1 port map( A1 => plusA(54), A2 => n290, B1 => plus2A(54), B2 
                           => n288, ZN => n411);
   U142 : AOI22_X1 port map( A1 => minus2A(54), A2 => n300, B1 => minusA(54), 
                           B2 => n293, ZN => n410);
   U143 : NAND2_X1 port map( A1 => n333, A2 => n332, ZN => n482);
   U144 : AOI22_X1 port map( A1 => plusA(15), A2 => n290, B1 => plus2A(15), B2 
                           => n285, ZN => n333);
   U145 : AOI22_X1 port map( A1 => minus2A(15), A2 => n297, B1 => minusA(15), 
                           B2 => n293, ZN => n332);
   U146 : NAND2_X1 port map( A1 => n341, A2 => n340, ZN => n478);
   U147 : AOI22_X1 port map( A1 => plusA(19), A2 => n290, B1 => plus2A(19), B2 
                           => n285, ZN => n341);
   U148 : AOI22_X1 port map( A1 => minus2A(19), A2 => n297, B1 => minusA(19), 
                           B2 => n293, ZN => n340);
   U149 : NAND2_X1 port map( A1 => n349, A2 => n348, ZN => n474);
   U150 : AOI22_X1 port map( A1 => plusA(23), A2 => n290, B1 => plus2A(23), B2 
                           => n285, ZN => n349);
   U151 : AOI22_X1 port map( A1 => minus2A(23), A2 => n297, B1 => minusA(23), 
                           B2 => n293, ZN => n348);
   U152 : NAND2_X1 port map( A1 => n357, A2 => n356, ZN => n470);
   U153 : AOI22_X1 port map( A1 => plusA(27), A2 => n290, B1 => plus2A(27), B2 
                           => n286, ZN => n357);
   U154 : AOI22_X1 port map( A1 => minus2A(27), A2 => n298, B1 => minusA(27), 
                           B2 => n293, ZN => n356);
   U155 : NAND2_X1 port map( A1 => n365, A2 => n364, ZN => n466);
   U156 : AOI22_X1 port map( A1 => plusA(31), A2 => n290, B1 => plus2A(31), B2 
                           => n286, ZN => n365);
   U157 : AOI22_X1 port map( A1 => minus2A(31), A2 => n298, B1 => minusA(31), 
                           B2 => n293, ZN => n364);
   U158 : NAND2_X1 port map( A1 => n391, A2 => n390, ZN => n453);
   U159 : AOI22_X1 port map( A1 => plusA(44), A2 => n290, B1 => plus2A(44), B2 
                           => n287, ZN => n391);
   U160 : AOI22_X1 port map( A1 => minus2A(44), A2 => n299, B1 => minusA(44), 
                           B2 => n293, ZN => n390);
   U161 : NAND2_X1 port map( A1 => n409, A2 => n408, ZN => n444);
   U162 : AOI22_X1 port map( A1 => plusA(53), A2 => n290, B1 => plus2A(53), B2 
                           => n288, ZN => n409);
   U163 : AOI22_X1 port map( A1 => minus2A(53), A2 => n300, B1 => minusA(53), 
                           B2 => n296, ZN => n408);
   U164 : NAND2_X1 port map( A1 => n307, A2 => n306, ZN => n495);
   U165 : AOI22_X1 port map( A1 => plusA(2), A2 => n429, B1 => plus2A(2), B2 =>
                           n428, ZN => n307);
   U166 : NAND2_X1 port map( A1 => n373, A2 => n372, ZN => n462);
   U167 : AOI22_X1 port map( A1 => plusA(35), A2 => n290, B1 => plus2A(35), B2 
                           => n286, ZN => n373);
   U168 : AOI22_X1 port map( A1 => minus2A(35), A2 => n298, B1 => minusA(35), 
                           B2 => n293, ZN => n372);
   U169 : NAND2_X1 port map( A1 => n375, A2 => n374, ZN => n461);
   U170 : AOI22_X1 port map( A1 => plusA(36), A2 => n292, B1 => plus2A(36), B2 
                           => n287, ZN => n375);
   U171 : AOI22_X1 port map( A1 => minus2A(36), A2 => n299, B1 => minusA(36), 
                           B2 => n293, ZN => n374);
   U172 : NAND2_X1 port map( A1 => n385, A2 => n384, ZN => n456);
   U173 : AOI22_X1 port map( A1 => plusA(41), A2 => n292, B1 => plus2A(41), B2 
                           => n287, ZN => n385);
   U174 : AOI22_X1 port map( A1 => minus2A(41), A2 => n299, B1 => minusA(41), 
                           B2 => n293, ZN => n384);
   U175 : NAND2_X1 port map( A1 => n433, A2 => n432, ZN => n434);
   U176 : AOI22_X1 port map( A1 => plusA(63), A2 => n292, B1 => plus2A(63), B2 
                           => n289, ZN => n433);
   U177 : AOI22_X1 port map( A1 => minus2A(63), A2 => n301, B1 => minusA(63), 
                           B2 => n293, ZN => n432);
   U178 : NAND2_X1 port map( A1 => n423, A2 => n422, ZN => n437);
   U179 : AOI22_X1 port map( A1 => plusA(60), A2 => n292, B1 => plus2A(60), B2 
                           => n289, ZN => n423);
   U180 : AOI22_X1 port map( A1 => minus2A(60), A2 => n301, B1 => minusA(60), 
                           B2 => n293, ZN => n422);
   U181 : NAND2_X1 port map( A1 => n413, A2 => n412, ZN => n442);
   U182 : AOI22_X1 port map( A1 => plusA(55), A2 => n292, B1 => plus2A(55), B2 
                           => n288, ZN => n413);
   U183 : AOI22_X1 port map( A1 => minus2A(55), A2 => n300, B1 => minusA(55), 
                           B2 => n293, ZN => n412);
   U184 : NAND2_X1 port map( A1 => n407, A2 => n406, ZN => n445);
   U185 : AOI22_X1 port map( A1 => plusA(52), A2 => n292, B1 => plus2A(52), B2 
                           => n288, ZN => n407);
   U186 : AOI22_X1 port map( A1 => minus2A(52), A2 => n300, B1 => minusA(52), 
                           B2 => n293, ZN => n406);
   U187 : NAND2_X1 port map( A1 => n405, A2 => n404, ZN => n446);
   U188 : AOI22_X1 port map( A1 => plusA(51), A2 => n292, B1 => plus2A(51), B2 
                           => n288, ZN => n405);
   U189 : AOI22_X1 port map( A1 => minus2A(51), A2 => n300, B1 => minusA(51), 
                           B2 => n293, ZN => n404);
   U190 : NAND2_X1 port map( A1 => n395, A2 => n394, ZN => n451);
   U191 : AOI22_X1 port map( A1 => plusA(46), A2 => n292, B1 => plus2A(46), B2 
                           => n287, ZN => n395);
   U192 : AOI22_X1 port map( A1 => minus2A(46), A2 => n299, B1 => minusA(46), 
                           B2 => n296, ZN => n394);
   U193 : NAND2_X1 port map( A1 => n393, A2 => n392, ZN => n452);
   U194 : AOI22_X1 port map( A1 => plusA(45), A2 => n290, B1 => plus2A(45), B2 
                           => n287, ZN => n393);
   U195 : AOI22_X1 port map( A1 => minus2A(45), A2 => n299, B1 => minusA(45), 
                           B2 => n293, ZN => n392);
   U196 : NAND2_X1 port map( A1 => n417, A2 => n416, ZN => n440);
   U197 : AOI22_X1 port map( A1 => plusA(57), A2 => n290, B1 => plus2A(57), B2 
                           => n288, ZN => n417);
   U198 : AOI22_X1 port map( A1 => minus2A(57), A2 => n300, B1 => minusA(57), 
                           B2 => n296, ZN => n416);
   U199 : NAND2_X1 port map( A1 => n387, A2 => n386, ZN => n455);
   U200 : AOI22_X1 port map( A1 => plusA(42), A2 => n290, B1 => plus2A(42), B2 
                           => n287, ZN => n387);
   U201 : AOI22_X1 port map( A1 => minus2A(42), A2 => n299, B1 => minusA(42), 
                           B2 => n296, ZN => n386);
   U202 : NAND2_X1 port map( A1 => n397, A2 => n396, ZN => n450);
   U203 : AOI22_X1 port map( A1 => plusA(47), A2 => n290, B1 => plus2A(47), B2 
                           => n287, ZN => n397);
   U204 : AOI22_X1 port map( A1 => minus2A(47), A2 => n299, B1 => minusA(47), 
                           B2 => n293, ZN => n396);
   U205 : NAND2_X1 port map( A1 => n377, A2 => n376, ZN => n460);
   U206 : AOI22_X1 port map( A1 => plusA(37), A2 => n290, B1 => plus2A(37), B2 
                           => n287, ZN => n377);
   U207 : AOI22_X1 port map( A1 => minus2A(37), A2 => n299, B1 => minusA(37), 
                           B2 => n293, ZN => n376);
   U208 : NAND2_X1 port map( A1 => n427, A2 => n426, ZN => n435);
   U209 : AOI22_X1 port map( A1 => plusA(62), A2 => n290, B1 => plus2A(62), B2 
                           => n289, ZN => n427);
   U210 : AOI22_X1 port map( A1 => minus2A(62), A2 => n301, B1 => minusA(62), 
                           B2 => n293, ZN => n426);
   U211 : NAND2_X1 port map( A1 => n425, A2 => n424, ZN => n436);
   U212 : AOI22_X1 port map( A1 => plusA(61), A2 => n290, B1 => plus2A(61), B2 
                           => n289, ZN => n425);
   U213 : AOI22_X1 port map( A1 => minus2A(61), A2 => n301, B1 => minusA(61), 
                           B2 => n296, ZN => n424);
   U214 : NAND2_X1 port map( A1 => n415, A2 => n414, ZN => n441);
   U215 : AOI22_X1 port map( A1 => plusA(56), A2 => n290, B1 => plus2A(56), B2 
                           => n288, ZN => n415);
   U216 : AOI22_X1 port map( A1 => minus2A(56), A2 => n300, B1 => minusA(56), 
                           B2 => n293, ZN => n414);
   U217 : NAND2_X1 port map( A1 => n305, A2 => n304, ZN => n496);
   U218 : AOI22_X1 port map( A1 => plusA(1), A2 => n290, B1 => plus2A(1), B2 =>
                           n288, ZN => n305);
   U219 : NAND2_X1 port map( A1 => n303, A2 => n302, ZN => n497);
   U220 : AOI22_X1 port map( A1 => plusA(0), A2 => n290, B1 => plus2A(0), B2 =>
                           n288, ZN => n303);
   U221 : NOR3_X1 port map( A1 => net85116, A2 => n273, A3 => net93945, ZN => 
                           n429);
   U222 : CLKBUF_X1 port map( A => n282, Z => n291);
   U223 : AOI22_X1 port map( A1 => minus2A(0), A2 => n297, B1 => minusA(0), B2 
                           => n293, ZN => n302);
   U224 : AOI22_X1 port map( A1 => minus2A(1), A2 => n297, B1 => minusA(1), B2 
                           => n293, ZN => n304);
   U225 : AOI22_X1 port map( A1 => minus2A(11), A2 => n297, B1 => minusA(11), 
                           B2 => n293, ZN => n324);
   U226 : AOI22_X1 port map( A1 => minus2A(10), A2 => n297, B1 => minusA(10), 
                           B2 => n293, ZN => n322);
   U227 : AOI22_X1 port map( A1 => minus2A(9), A2 => n297, B1 => minusA(9), B2 
                           => n293, ZN => n320);
   U228 : AOI22_X1 port map( A1 => minus2A(8), A2 => n297, B1 => minusA(8), B2 
                           => n296, ZN => n318);
   U229 : AOI22_X1 port map( A1 => minus2A(7), A2 => n297, B1 => minusA(7), B2 
                           => n295, ZN => n316);
   U230 : AOI22_X1 port map( A1 => minus2A(6), A2 => n298, B1 => minusA(6), B2 
                           => n295, ZN => n314);
   U231 : AOI22_X1 port map( A1 => minus2A(5), A2 => n299, B1 => minusA(5), B2 
                           => n294, ZN => n312);
   U232 : AOI22_X1 port map( A1 => minus2A(4), A2 => n300, B1 => minusA(4), B2 
                           => n294, ZN => n310);
   U233 : AOI22_X1 port map( A1 => minus2A(3), A2 => n301, B1 => minusA(3), B2 
                           => n281, ZN => n308);
   U234 : AOI22_X1 port map( A1 => minus2A(2), A2 => n431, B1 => minusA(2), B2 
                           => n430, ZN => n306);
   U235 : CLKBUF_X1 port map( A => n278, Z => n289);
   U236 : CLKBUF_X1 port map( A => n431, Z => n301);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity MUX_GENERIC_N64_RADIX3_14 is

   port( plusA, minusA, plus2A, minus2A : in std_logic_vector (63 downto 0);  
         SEL : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (63 
         downto 0));

end MUX_GENERIC_N64_RADIX3_14;

architecture SYN_beh of MUX_GENERIC_N64_RADIX3_14 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component TBUF_X4
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   component TBUF_X1
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   signal n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, 
      n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, 
      n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, 
      n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, 
      n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, 
      n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, 
      n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, 
      n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, 
      n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, 
      n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, 
      n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, 
      n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, 
      n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, 
      n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, 
      n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, 
      n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, 
      n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, 
      n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, 
      n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, 
      n499, n500, n501, n502, n503, n504 : std_logic;

begin
   
   Y_tri_60_inst : TBUF_X1 port map( A => n443, EN => n303, Z => Y(60));
   Y_tri_61_inst : TBUF_X1 port map( A => n442, EN => n303, Z => Y(61));
   Y_tri_62_inst : TBUF_X1 port map( A => n441, EN => n303, Z => Y(62));
   Y_tri_63_inst : TBUF_X1 port map( A => n440, EN => n303, Z => Y(63));
   Y_tri_38_inst : TBUF_X1 port map( A => n465, EN => n301, Z => Y(38));
   Y_tri_39_inst : TBUF_X1 port map( A => n464, EN => n301, Z => Y(39));
   Y_tri_40_inst : TBUF_X1 port map( A => n463, EN => n301, Z => Y(40));
   Y_tri_41_inst : TBUF_X1 port map( A => n462, EN => n301, Z => Y(41));
   Y_tri_42_inst : TBUF_X1 port map( A => n461, EN => n301, Z => Y(42));
   Y_tri_43_inst : TBUF_X1 port map( A => n460, EN => n301, Z => Y(43));
   Y_tri_44_inst : TBUF_X1 port map( A => n459, EN => n301, Z => Y(44));
   Y_tri_45_inst : TBUF_X1 port map( A => n458, EN => n301, Z => Y(45));
   Y_tri_46_inst : TBUF_X1 port map( A => n457, EN => n301, Z => Y(46));
   Y_tri_47_inst : TBUF_X1 port map( A => n456, EN => n301, Z => Y(47));
   Y_tri_48_inst : TBUF_X1 port map( A => n455, EN => n302, Z => Y(48));
   Y_tri_49_inst : TBUF_X1 port map( A => n454, EN => n302, Z => Y(49));
   Y_tri_50_inst : TBUF_X1 port map( A => n453, EN => n302, Z => Y(50));
   Y_tri_51_inst : TBUF_X1 port map( A => n452, EN => n302, Z => Y(51));
   Y_tri_52_inst : TBUF_X1 port map( A => n451, EN => n302, Z => Y(52));
   Y_tri_53_inst : TBUF_X1 port map( A => n450, EN => n302, Z => Y(53));
   Y_tri_54_inst : TBUF_X1 port map( A => n449, EN => n302, Z => Y(54));
   Y_tri_55_inst : TBUF_X1 port map( A => n448, EN => n302, Z => Y(55));
   Y_tri_56_inst : TBUF_X1 port map( A => n447, EN => n302, Z => Y(56));
   Y_tri_57_inst : TBUF_X1 port map( A => n446, EN => n302, Z => Y(57));
   Y_tri_58_inst : TBUF_X1 port map( A => n445, EN => n302, Z => Y(58));
   Y_tri_59_inst : TBUF_X1 port map( A => n444, EN => n302, Z => Y(59));
   Y_tri_32_inst : TBUF_X1 port map( A => n471, EN => n300, Z => Y(32));
   Y_tri_30_inst : TBUF_X1 port map( A => n473, EN => n300, Z => Y(30));
   Y_tri_29_inst : TBUF_X1 port map( A => n474, EN => n300, Z => Y(29));
   Y_tri_28_inst : TBUF_X1 port map( A => n475, EN => n300, Z => Y(28));
   Y_tri_27_inst : TBUF_X1 port map( A => n476, EN => n300, Z => Y(27));
   Y_tri_26_inst : TBUF_X1 port map( A => n477, EN => n300, Z => Y(26));
   Y_tri_25_inst : TBUF_X1 port map( A => n478, EN => n300, Z => Y(25));
   Y_tri_24_inst : TBUF_X1 port map( A => n479, EN => n300, Z => Y(24));
   Y_tri_23_inst : TBUF_X1 port map( A => n480, EN => n299, Z => Y(23));
   Y_tri_22_inst : TBUF_X1 port map( A => n481, EN => n299, Z => Y(22));
   Y_tri_21_inst : TBUF_X1 port map( A => n482, EN => n299, Z => Y(21));
   Y_tri_20_inst : TBUF_X1 port map( A => n483, EN => n299, Z => Y(20));
   Y_tri_19_inst : TBUF_X1 port map( A => n484, EN => n299, Z => Y(19));
   Y_tri_18_inst : TBUF_X1 port map( A => n485, EN => n299, Z => Y(18));
   Y_tri_17_inst : TBUF_X1 port map( A => n486, EN => n299, Z => Y(17));
   Y_tri_16_inst : TBUF_X1 port map( A => n487, EN => n299, Z => Y(16));
   Y_tri_15_inst : TBUF_X1 port map( A => n488, EN => n299, Z => Y(15));
   Y_tri_14_inst : TBUF_X1 port map( A => n489, EN => n299, Z => Y(14));
   Y_tri_33_inst : TBUF_X1 port map( A => n470, EN => n300, Z => Y(33));
   Y_tri_13_inst : TBUF_X1 port map( A => n490, EN => n299, Z => Y(13));
   Y_tri_12_inst : TBUF_X1 port map( A => n491, EN => n299, Z => Y(12));
   Y_tri_34_inst : TBUF_X1 port map( A => n469, EN => n300, Z => Y(34));
   Y_tri_35_inst : TBUF_X1 port map( A => n468, EN => n300, Z => Y(35));
   Y_tri_36_inst : TBUF_X1 port map( A => n467, EN => n301, Z => Y(36));
   Y_tri_37_inst : TBUF_X1 port map( A => n466, EN => n301, Z => Y(37));
   Y_tri_7_inst : TBUF_X1 port map( A => n497, EN => n298, Z => Y(7));
   Y_tri_8_inst : TBUF_X1 port map( A => n496, EN => n298, Z => Y(8));
   Y_tri_9_inst : TBUF_X1 port map( A => n494, EN => n298, Z => Y(9));
   Y_tri_11_inst : TBUF_X1 port map( A => n492, EN => n298, Z => Y(11));
   Y_tri_10_inst : TBUF_X1 port map( A => n493, EN => n298, Z => Y(10));
   Y_tri_31_inst : TBUF_X1 port map( A => n472, EN => n300, Z => Y(31));
   Y_tri_5_inst : TBUF_X1 port map( A => n499, EN => n298, Z => Y(5));
   Y_tri_3_inst : TBUF_X1 port map( A => n501, EN => n298, Z => Y(3));
   Y_tri_4_inst : TBUF_X1 port map( A => n500, EN => n298, Z => Y(4));
   Y_tri_2_inst : TBUF_X1 port map( A => n502, EN => n298, Z => Y(2));
   Y_tri_6_inst : TBUF_X1 port map( A => n498, EN => n298, Z => Y(6));
   Y_tri_1_inst : TBUF_X1 port map( A => n503, EN => n298, Z => Y(1));
   Y_tri_0_inst : TBUF_X4 port map( A => n504, EN => n298, Z => Y(0));
   U2 : CLKBUF_X3 port map( A => n495, Z => n298);
   U3 : NOR2_X2 port map( A1 => n325, A2 => n306, ZN => n495);
   U4 : BUF_X1 port map( A => SEL(1), Z => n272);
   U5 : NOR3_X1 port map( A1 => n273, A2 => SEL(2), A3 => n304, ZN => n436);
   U6 : NOR3_X1 port map( A1 => n304, A2 => SEL(2), A3 => n305, ZN => n434);
   U7 : NOR3_X1 port map( A1 => n272, A2 => SEL(2), A3 => n305, ZN => n435);
   U8 : INV_X1 port map( A => n305, ZN => n273);
   U9 : CLKBUF_X1 port map( A => n495, Z => n299);
   U10 : CLKBUF_X1 port map( A => n495, Z => n300);
   U11 : CLKBUF_X1 port map( A => n437, Z => n294);
   U12 : CLKBUF_X1 port map( A => n437, Z => n293);
   U13 : CLKBUF_X1 port map( A => n495, Z => n301);
   U14 : CLKBUF_X1 port map( A => n437, Z => n295);
   U15 : CLKBUF_X1 port map( A => n495, Z => n302);
   U16 : CLKBUF_X1 port map( A => n437, Z => n296);
   U17 : BUF_X1 port map( A => n435, Z => n280);
   U18 : BUF_X1 port map( A => n436, Z => n286);
   U19 : BUF_X1 port map( A => n434, Z => n274);
   U20 : BUF_X1 port map( A => n437, Z => n292);
   U21 : CLKBUF_X1 port map( A => n435, Z => n281);
   U22 : CLKBUF_X1 port map( A => n435, Z => n282);
   U23 : CLKBUF_X1 port map( A => n436, Z => n287);
   U24 : CLKBUF_X1 port map( A => n434, Z => n275);
   U25 : CLKBUF_X1 port map( A => n436, Z => n288);
   U26 : CLKBUF_X1 port map( A => n434, Z => n276);
   U27 : CLKBUF_X1 port map( A => n435, Z => n283);
   U28 : CLKBUF_X1 port map( A => n436, Z => n289);
   U29 : CLKBUF_X1 port map( A => n434, Z => n277);
   U30 : CLKBUF_X1 port map( A => n435, Z => n284);
   U31 : CLKBUF_X1 port map( A => n436, Z => n290);
   U32 : CLKBUF_X1 port map( A => n434, Z => n278);
   U33 : INV_X1 port map( A => SEL(2), ZN => n306);
   U34 : AND2_X1 port map( A1 => SEL(2), A2 => n325, ZN => n437);
   U35 : NOR2_X1 port map( A1 => SEL(1), A2 => SEL(0), ZN => n325);
   U36 : INV_X1 port map( A => n272, ZN => n304);
   U37 : INV_X1 port map( A => SEL(0), ZN => n305);
   U38 : NAND2_X1 port map( A1 => n320, A2 => n319, ZN => n498);
   U39 : AOI22_X1 port map( A1 => plusA(6), A2 => n280, B1 => plus2A(6), B2 => 
                           n274, ZN => n320);
   U40 : AOI22_X1 port map( A1 => minus2A(6), A2 => n292, B1 => minusA(6), B2 
                           => n286, ZN => n319);
   U41 : NAND2_X1 port map( A1 => n318, A2 => n317, ZN => n499);
   U42 : AOI22_X1 port map( A1 => plusA(5), A2 => n280, B1 => plus2A(5), B2 => 
                           n274, ZN => n318);
   U43 : AOI22_X1 port map( A1 => minus2A(5), A2 => n292, B1 => minusA(5), B2 
                           => n286, ZN => n317);
   U44 : NAND2_X1 port map( A1 => n322, A2 => n321, ZN => n497);
   U45 : AOI22_X1 port map( A1 => plusA(7), A2 => n280, B1 => plus2A(7), B2 => 
                           n274, ZN => n322);
   U46 : AOI22_X1 port map( A1 => minus2A(7), A2 => n292, B1 => minusA(7), B2 
                           => n286, ZN => n321);
   U47 : NAND2_X1 port map( A1 => n427, A2 => n426, ZN => n444);
   U48 : AOI22_X1 port map( A1 => plusA(59), A2 => n284, B1 => plus2A(59), B2 
                           => n278, ZN => n427);
   U49 : AOI22_X1 port map( A1 => minus2A(59), A2 => n296, B1 => minusA(59), B2
                           => n290, ZN => n426);
   U50 : NAND2_X1 port map( A1 => n425, A2 => n424, ZN => n445);
   U51 : AOI22_X1 port map( A1 => plusA(58), A2 => n284, B1 => plus2A(58), B2 
                           => n278, ZN => n425);
   U52 : AOI22_X1 port map( A1 => minus2A(58), A2 => n296, B1 => minusA(58), B2
                           => n290, ZN => n424);
   U53 : NAND2_X1 port map( A1 => n423, A2 => n422, ZN => n446);
   U54 : AOI22_X1 port map( A1 => plusA(57), A2 => n284, B1 => plus2A(57), B2 
                           => n278, ZN => n423);
   U55 : AOI22_X1 port map( A1 => minus2A(57), A2 => n296, B1 => minusA(57), B2
                           => n290, ZN => n422);
   U56 : NAND2_X1 port map( A1 => n329, A2 => n328, ZN => n493);
   U57 : AOI22_X1 port map( A1 => plusA(10), A2 => n280, B1 => plus2A(10), B2 
                           => n274, ZN => n329);
   U58 : AOI22_X1 port map( A1 => minus2A(10), A2 => n292, B1 => minusA(10), B2
                           => n286, ZN => n328);
   U59 : NAND2_X1 port map( A1 => n337, A2 => n336, ZN => n489);
   U60 : AOI22_X1 port map( A1 => plusA(14), A2 => n281, B1 => plus2A(14), B2 
                           => n275, ZN => n337);
   U61 : AOI22_X1 port map( A1 => minus2A(14), A2 => n293, B1 => minusA(14), B2
                           => n287, ZN => n336);
   U62 : NAND2_X1 port map( A1 => n345, A2 => n344, ZN => n485);
   U63 : AOI22_X1 port map( A1 => plusA(18), A2 => n281, B1 => plus2A(18), B2 
                           => n275, ZN => n345);
   U64 : AOI22_X1 port map( A1 => minus2A(18), A2 => n293, B1 => minusA(18), B2
                           => n287, ZN => n344);
   U65 : NAND2_X1 port map( A1 => n353, A2 => n352, ZN => n481);
   U66 : AOI22_X1 port map( A1 => plusA(22), A2 => n281, B1 => plus2A(22), B2 
                           => n275, ZN => n353);
   U67 : AOI22_X1 port map( A1 => minus2A(22), A2 => n293, B1 => minusA(22), B2
                           => n287, ZN => n352);
   U68 : NAND2_X1 port map( A1 => n377, A2 => n376, ZN => n469);
   U69 : AOI22_X1 port map( A1 => plusA(34), A2 => n282, B1 => plus2A(34), B2 
                           => n276, ZN => n377);
   U70 : AOI22_X1 port map( A1 => minus2A(34), A2 => n294, B1 => minusA(34), B2
                           => n288, ZN => n376);
   U71 : NAND2_X1 port map( A1 => n361, A2 => n360, ZN => n477);
   U72 : AOI22_X1 port map( A1 => plusA(26), A2 => n282, B1 => plus2A(26), B2 
                           => n276, ZN => n361);
   U73 : AOI22_X1 port map( A1 => minus2A(26), A2 => n294, B1 => minusA(26), B2
                           => n288, ZN => n360);
   U74 : NAND2_X1 port map( A1 => n369, A2 => n368, ZN => n473);
   U75 : AOI22_X1 port map( A1 => plusA(30), A2 => n282, B1 => plus2A(30), B2 
                           => n276, ZN => n369);
   U76 : AOI22_X1 port map( A1 => minus2A(30), A2 => n294, B1 => minusA(30), B2
                           => n288, ZN => n368);
   U77 : NAND2_X1 port map( A1 => n409, A2 => n408, ZN => n453);
   U78 : AOI22_X1 port map( A1 => plusA(50), A2 => n284, B1 => plus2A(50), B2 
                           => n278, ZN => n409);
   U79 : AOI22_X1 port map( A1 => minus2A(50), A2 => n296, B1 => minusA(50), B2
                           => n290, ZN => n408);
   U80 : NAND2_X1 port map( A1 => n405, A2 => n404, ZN => n455);
   U81 : AOI22_X1 port map( A1 => plusA(48), A2 => n284, B1 => plus2A(48), B2 
                           => n278, ZN => n405);
   U82 : AOI22_X1 port map( A1 => minus2A(48), A2 => n296, B1 => minusA(48), B2
                           => n290, ZN => n404);
   U83 : NAND2_X1 port map( A1 => n395, A2 => n394, ZN => n460);
   U84 : AOI22_X1 port map( A1 => plusA(43), A2 => n283, B1 => plus2A(43), B2 
                           => n277, ZN => n395);
   U85 : AOI22_X1 port map( A1 => minus2A(43), A2 => n295, B1 => minusA(43), B2
                           => n289, ZN => n394);
   U86 : NAND2_X1 port map( A1 => n379, A2 => n378, ZN => n468);
   U87 : AOI22_X1 port map( A1 => plusA(35), A2 => n282, B1 => plus2A(35), B2 
                           => n276, ZN => n379);
   U88 : AOI22_X1 port map( A1 => minus2A(35), A2 => n294, B1 => minusA(35), B2
                           => n288, ZN => n378);
   U89 : NAND2_X1 port map( A1 => n403, A2 => n402, ZN => n456);
   U90 : AOI22_X1 port map( A1 => plusA(47), A2 => n283, B1 => plus2A(47), B2 
                           => n277, ZN => n403);
   U91 : AOI22_X1 port map( A1 => minus2A(47), A2 => n295, B1 => minusA(47), B2
                           => n289, ZN => n402);
   U92 : NAND2_X1 port map( A1 => n399, A2 => n398, ZN => n458);
   U93 : AOI22_X1 port map( A1 => plusA(45), A2 => n283, B1 => plus2A(45), B2 
                           => n277, ZN => n399);
   U94 : AOI22_X1 port map( A1 => minus2A(45), A2 => n295, B1 => minusA(45), B2
                           => n289, ZN => n398);
   U95 : NAND2_X1 port map( A1 => n324, A2 => n323, ZN => n496);
   U96 : AOI22_X1 port map( A1 => plusA(8), A2 => n280, B1 => plus2A(8), B2 => 
                           n274, ZN => n324);
   U97 : AOI22_X1 port map( A1 => minus2A(8), A2 => n292, B1 => minusA(8), B2 
                           => n286, ZN => n323);
   U98 : NAND2_X1 port map( A1 => n333, A2 => n332, ZN => n491);
   U99 : AOI22_X1 port map( A1 => plusA(12), A2 => n281, B1 => plus2A(12), B2 
                           => n275, ZN => n333);
   U100 : AOI22_X1 port map( A1 => minus2A(12), A2 => n293, B1 => minusA(12), 
                           B2 => n287, ZN => n332);
   U101 : NAND2_X1 port map( A1 => n341, A2 => n340, ZN => n487);
   U102 : AOI22_X1 port map( A1 => plusA(16), A2 => n281, B1 => plus2A(16), B2 
                           => n275, ZN => n341);
   U103 : AOI22_X1 port map( A1 => minus2A(16), A2 => n293, B1 => minusA(16), 
                           B2 => n287, ZN => n340);
   U104 : NAND2_X1 port map( A1 => n349, A2 => n348, ZN => n483);
   U105 : AOI22_X1 port map( A1 => plusA(20), A2 => n281, B1 => plus2A(20), B2 
                           => n275, ZN => n349);
   U106 : AOI22_X1 port map( A1 => minus2A(20), A2 => n293, B1 => minusA(20), 
                           B2 => n287, ZN => n348);
   U107 : NAND2_X1 port map( A1 => n357, A2 => n356, ZN => n479);
   U108 : AOI22_X1 port map( A1 => plusA(24), A2 => n282, B1 => plus2A(24), B2 
                           => n276, ZN => n357);
   U109 : AOI22_X1 port map( A1 => minus2A(24), A2 => n294, B1 => minusA(24), 
                           B2 => n288, ZN => n356);
   U110 : NAND2_X1 port map( A1 => n365, A2 => n364, ZN => n475);
   U111 : AOI22_X1 port map( A1 => plusA(28), A2 => n282, B1 => plus2A(28), B2 
                           => n276, ZN => n365);
   U112 : AOI22_X1 port map( A1 => minus2A(28), A2 => n294, B1 => minusA(28), 
                           B2 => n288, ZN => n364);
   U113 : NAND2_X1 port map( A1 => n373, A2 => n372, ZN => n471);
   U114 : AOI22_X1 port map( A1 => plusA(32), A2 => n282, B1 => plus2A(32), B2 
                           => n276, ZN => n373);
   U115 : AOI22_X1 port map( A1 => minus2A(32), A2 => n294, B1 => minusA(32), 
                           B2 => n288, ZN => n372);
   U116 : NAND2_X1 port map( A1 => n389, A2 => n388, ZN => n463);
   U117 : AOI22_X1 port map( A1 => plusA(40), A2 => n283, B1 => plus2A(40), B2 
                           => n277, ZN => n389);
   U118 : AOI22_X1 port map( A1 => minus2A(40), A2 => n295, B1 => minusA(40), 
                           B2 => n289, ZN => n388);
   U119 : NAND2_X1 port map( A1 => n385, A2 => n384, ZN => n465);
   U120 : AOI22_X1 port map( A1 => plusA(38), A2 => n283, B1 => plus2A(38), B2 
                           => n277, ZN => n385);
   U121 : AOI22_X1 port map( A1 => minus2A(38), A2 => n295, B1 => minusA(38), 
                           B2 => n289, ZN => n384);
   U122 : NAND2_X1 port map( A1 => n383, A2 => n382, ZN => n466);
   U123 : AOI22_X1 port map( A1 => plusA(37), A2 => n283, B1 => plus2A(37), B2 
                           => n277, ZN => n383);
   U124 : AOI22_X1 port map( A1 => minus2A(37), A2 => n295, B1 => minusA(37), 
                           B2 => n289, ZN => n382);
   U125 : NAND2_X1 port map( A1 => n331, A2 => n330, ZN => n492);
   U126 : AOI22_X1 port map( A1 => plusA(11), A2 => n280, B1 => plus2A(11), B2 
                           => n274, ZN => n331);
   U127 : AOI22_X1 port map( A1 => minus2A(11), A2 => n292, B1 => minusA(11), 
                           B2 => n286, ZN => n330);
   U128 : NAND2_X1 port map( A1 => n339, A2 => n338, ZN => n488);
   U129 : AOI22_X1 port map( A1 => plusA(15), A2 => n281, B1 => plus2A(15), B2 
                           => n275, ZN => n339);
   U130 : AOI22_X1 port map( A1 => minus2A(15), A2 => n293, B1 => minusA(15), 
                           B2 => n287, ZN => n338);
   U131 : NAND2_X1 port map( A1 => n347, A2 => n346, ZN => n484);
   U132 : AOI22_X1 port map( A1 => plusA(19), A2 => n281, B1 => plus2A(19), B2 
                           => n275, ZN => n347);
   U133 : AOI22_X1 port map( A1 => minus2A(19), A2 => n293, B1 => minusA(19), 
                           B2 => n287, ZN => n346);
   U134 : NAND2_X1 port map( A1 => n355, A2 => n354, ZN => n480);
   U135 : AOI22_X1 port map( A1 => plusA(23), A2 => n281, B1 => plus2A(23), B2 
                           => n275, ZN => n355);
   U136 : AOI22_X1 port map( A1 => minus2A(23), A2 => n293, B1 => minusA(23), 
                           B2 => n287, ZN => n354);
   U137 : NAND2_X1 port map( A1 => n363, A2 => n362, ZN => n476);
   U138 : AOI22_X1 port map( A1 => plusA(27), A2 => n282, B1 => plus2A(27), B2 
                           => n276, ZN => n363);
   U139 : AOI22_X1 port map( A1 => minus2A(27), A2 => n294, B1 => minusA(27), 
                           B2 => n288, ZN => n362);
   U140 : NAND2_X1 port map( A1 => n371, A2 => n370, ZN => n472);
   U141 : AOI22_X1 port map( A1 => plusA(31), A2 => n282, B1 => plus2A(31), B2 
                           => n276, ZN => n371);
   U142 : AOI22_X1 port map( A1 => minus2A(31), A2 => n294, B1 => minusA(31), 
                           B2 => n288, ZN => n370);
   U143 : NAND2_X1 port map( A1 => n411, A2 => n410, ZN => n452);
   U144 : AOI22_X1 port map( A1 => plusA(51), A2 => n284, B1 => plus2A(51), B2 
                           => n278, ZN => n411);
   U145 : AOI22_X1 port map( A1 => minus2A(51), A2 => n296, B1 => minusA(51), 
                           B2 => n290, ZN => n410);
   U146 : NAND2_X1 port map( A1 => n407, A2 => n406, ZN => n454);
   U147 : AOI22_X1 port map( A1 => plusA(49), A2 => n284, B1 => plus2A(49), B2 
                           => n278, ZN => n407);
   U148 : AOI22_X1 port map( A1 => minus2A(49), A2 => n296, B1 => minusA(49), 
                           B2 => n290, ZN => n406);
   U149 : NAND2_X1 port map( A1 => n413, A2 => n412, ZN => n451);
   U150 : AOI22_X1 port map( A1 => plusA(52), A2 => n284, B1 => plus2A(52), B2 
                           => n278, ZN => n413);
   U151 : AOI22_X1 port map( A1 => minus2A(52), A2 => n296, B1 => minusA(52), 
                           B2 => n290, ZN => n412);
   U152 : NAND2_X1 port map( A1 => n381, A2 => n380, ZN => n467);
   U153 : AOI22_X1 port map( A1 => plusA(36), A2 => n283, B1 => plus2A(36), B2 
                           => n277, ZN => n381);
   U154 : AOI22_X1 port map( A1 => minus2A(36), A2 => n295, B1 => minusA(36), 
                           B2 => n289, ZN => n380);
   U155 : NAND2_X1 port map( A1 => n421, A2 => n420, ZN => n447);
   U156 : AOI22_X1 port map( A1 => plusA(56), A2 => n284, B1 => plus2A(56), B2 
                           => n278, ZN => n421);
   U157 : AOI22_X1 port map( A1 => minus2A(56), A2 => n296, B1 => minusA(56), 
                           B2 => n290, ZN => n420);
   U158 : NAND2_X1 port map( A1 => n417, A2 => n416, ZN => n449);
   U159 : AOI22_X1 port map( A1 => plusA(54), A2 => n284, B1 => plus2A(54), B2 
                           => n278, ZN => n417);
   U160 : AOI22_X1 port map( A1 => minus2A(54), A2 => n296, B1 => minusA(54), 
                           B2 => n290, ZN => n416);
   U161 : NAND2_X1 port map( A1 => n327, A2 => n326, ZN => n494);
   U162 : AOI22_X1 port map( A1 => plusA(9), A2 => n280, B1 => plus2A(9), B2 =>
                           n274, ZN => n327);
   U163 : AOI22_X1 port map( A1 => minus2A(9), A2 => n292, B1 => minusA(9), B2 
                           => n286, ZN => n326);
   U164 : NAND2_X1 port map( A1 => n335, A2 => n334, ZN => n490);
   U165 : AOI22_X1 port map( A1 => plusA(13), A2 => n281, B1 => plus2A(13), B2 
                           => n275, ZN => n335);
   U166 : AOI22_X1 port map( A1 => minus2A(13), A2 => n293, B1 => minusA(13), 
                           B2 => n287, ZN => n334);
   U167 : NAND2_X1 port map( A1 => n343, A2 => n342, ZN => n486);
   U168 : AOI22_X1 port map( A1 => plusA(17), A2 => n281, B1 => plus2A(17), B2 
                           => n275, ZN => n343);
   U169 : AOI22_X1 port map( A1 => minus2A(17), A2 => n293, B1 => minusA(17), 
                           B2 => n287, ZN => n342);
   U170 : NAND2_X1 port map( A1 => n351, A2 => n350, ZN => n482);
   U171 : AOI22_X1 port map( A1 => plusA(21), A2 => n281, B1 => plus2A(21), B2 
                           => n275, ZN => n351);
   U172 : AOI22_X1 port map( A1 => minus2A(21), A2 => n293, B1 => minusA(21), 
                           B2 => n287, ZN => n350);
   U173 : NAND2_X1 port map( A1 => n375, A2 => n374, ZN => n470);
   U174 : AOI22_X1 port map( A1 => plusA(33), A2 => n282, B1 => plus2A(33), B2 
                           => n276, ZN => n375);
   U175 : AOI22_X1 port map( A1 => minus2A(33), A2 => n294, B1 => minusA(33), 
                           B2 => n288, ZN => n374);
   U176 : NAND2_X1 port map( A1 => n359, A2 => n358, ZN => n478);
   U177 : AOI22_X1 port map( A1 => plusA(25), A2 => n282, B1 => plus2A(25), B2 
                           => n276, ZN => n359);
   U178 : AOI22_X1 port map( A1 => minus2A(25), A2 => n294, B1 => minusA(25), 
                           B2 => n288, ZN => n358);
   U179 : NAND2_X1 port map( A1 => n367, A2 => n366, ZN => n474);
   U180 : AOI22_X1 port map( A1 => plusA(29), A2 => n282, B1 => plus2A(29), B2 
                           => n276, ZN => n367);
   U181 : AOI22_X1 port map( A1 => minus2A(29), A2 => n294, B1 => minusA(29), 
                           B2 => n288, ZN => n366);
   U182 : NAND2_X1 port map( A1 => n391, A2 => n390, ZN => n462);
   U183 : AOI22_X1 port map( A1 => plusA(41), A2 => n283, B1 => plus2A(41), B2 
                           => n277, ZN => n391);
   U184 : AOI22_X1 port map( A1 => minus2A(41), A2 => n295, B1 => minusA(41), 
                           B2 => n289, ZN => n390);
   U185 : NAND2_X1 port map( A1 => n387, A2 => n386, ZN => n464);
   U186 : AOI22_X1 port map( A1 => plusA(39), A2 => n283, B1 => plus2A(39), B2 
                           => n277, ZN => n387);
   U187 : AOI22_X1 port map( A1 => minus2A(39), A2 => n295, B1 => minusA(39), 
                           B2 => n289, ZN => n386);
   U188 : NAND2_X1 port map( A1 => n393, A2 => n392, ZN => n461);
   U189 : AOI22_X1 port map( A1 => plusA(42), A2 => n283, B1 => plus2A(42), B2 
                           => n277, ZN => n393);
   U190 : AOI22_X1 port map( A1 => minus2A(42), A2 => n295, B1 => minusA(42), 
                           B2 => n289, ZN => n392);
   U191 : NAND2_X1 port map( A1 => n401, A2 => n400, ZN => n457);
   U192 : AOI22_X1 port map( A1 => plusA(46), A2 => n283, B1 => plus2A(46), B2 
                           => n277, ZN => n401);
   U193 : AOI22_X1 port map( A1 => minus2A(46), A2 => n295, B1 => minusA(46), 
                           B2 => n289, ZN => n400);
   U194 : NAND2_X1 port map( A1 => n397, A2 => n396, ZN => n459);
   U195 : AOI22_X1 port map( A1 => plusA(44), A2 => n283, B1 => plus2A(44), B2 
                           => n277, ZN => n397);
   U196 : AOI22_X1 port map( A1 => minus2A(44), A2 => n295, B1 => minusA(44), 
                           B2 => n289, ZN => n396);
   U197 : NAND2_X1 port map( A1 => n415, A2 => n414, ZN => n450);
   U198 : AOI22_X1 port map( A1 => plusA(53), A2 => n284, B1 => plus2A(53), B2 
                           => n278, ZN => n415);
   U199 : AOI22_X1 port map( A1 => minus2A(53), A2 => n296, B1 => minusA(53), 
                           B2 => n290, ZN => n414);
   U200 : NAND2_X1 port map( A1 => n419, A2 => n418, ZN => n448);
   U201 : AOI22_X1 port map( A1 => plusA(55), A2 => n284, B1 => plus2A(55), B2 
                           => n278, ZN => n419);
   U202 : AOI22_X1 port map( A1 => minus2A(55), A2 => n296, B1 => minusA(55), 
                           B2 => n290, ZN => n418);
   U203 : NAND2_X1 port map( A1 => n431, A2 => n430, ZN => n442);
   U204 : AOI22_X1 port map( A1 => plusA(61), A2 => n285, B1 => plus2A(61), B2 
                           => n279, ZN => n431);
   U205 : AOI22_X1 port map( A1 => minus2A(61), A2 => n297, B1 => minusA(61), 
                           B2 => n291, ZN => n430);
   U206 : NAND2_X1 port map( A1 => n429, A2 => n428, ZN => n443);
   U207 : AOI22_X1 port map( A1 => plusA(60), A2 => n285, B1 => plus2A(60), B2 
                           => n279, ZN => n429);
   U208 : AOI22_X1 port map( A1 => minus2A(60), A2 => n297, B1 => minusA(60), 
                           B2 => n291, ZN => n428);
   U209 : NAND2_X1 port map( A1 => n316, A2 => n315, ZN => n500);
   U210 : AOI22_X1 port map( A1 => plusA(4), A2 => n280, B1 => plus2A(4), B2 =>
                           n274, ZN => n316);
   U211 : AOI22_X1 port map( A1 => minus2A(4), A2 => n292, B1 => minusA(4), B2 
                           => n286, ZN => n315);
   U212 : NAND2_X1 port map( A1 => n439, A2 => n438, ZN => n440);
   U213 : AOI22_X1 port map( A1 => plusA(63), A2 => n285, B1 => plus2A(63), B2 
                           => n279, ZN => n439);
   U214 : AOI22_X1 port map( A1 => minus2A(63), A2 => n297, B1 => minusA(63), 
                           B2 => n291, ZN => n438);
   U215 : NAND2_X1 port map( A1 => n433, A2 => n432, ZN => n441);
   U216 : AOI22_X1 port map( A1 => plusA(62), A2 => n285, B1 => plus2A(62), B2 
                           => n279, ZN => n433);
   U217 : AOI22_X1 port map( A1 => minus2A(62), A2 => n297, B1 => minusA(62), 
                           B2 => n291, ZN => n432);
   U218 : NAND2_X1 port map( A1 => n314, A2 => n313, ZN => n501);
   U219 : AOI22_X1 port map( A1 => plusA(3), A2 => n280, B1 => plus2A(3), B2 =>
                           n274, ZN => n314);
   U220 : AOI22_X1 port map( A1 => minus2A(3), A2 => n292, B1 => minusA(3), B2 
                           => n286, ZN => n313);
   U221 : NAND2_X1 port map( A1 => n312, A2 => n311, ZN => n502);
   U222 : AOI22_X1 port map( A1 => plusA(2), A2 => n280, B1 => plus2A(2), B2 =>
                           n274, ZN => n312);
   U223 : AOI22_X1 port map( A1 => minus2A(2), A2 => n292, B1 => minusA(2), B2 
                           => n286, ZN => n311);
   U224 : NAND2_X1 port map( A1 => n310, A2 => n309, ZN => n503);
   U225 : AOI22_X1 port map( A1 => plusA(1), A2 => n280, B1 => plus2A(1), B2 =>
                           n274, ZN => n310);
   U226 : AOI22_X1 port map( A1 => minus2A(1), A2 => n292, B1 => minusA(1), B2 
                           => n286, ZN => n309);
   U227 : NAND2_X1 port map( A1 => n308, A2 => n307, ZN => n504);
   U228 : AOI22_X1 port map( A1 => plusA(0), A2 => n280, B1 => plus2A(0), B2 =>
                           n274, ZN => n308);
   U229 : AOI22_X1 port map( A1 => minus2A(0), A2 => n292, B1 => minusA(0), B2 
                           => n286, ZN => n307);
   U230 : CLKBUF_X1 port map( A => n434, Z => n279);
   U231 : CLKBUF_X1 port map( A => n435, Z => n285);
   U232 : CLKBUF_X1 port map( A => n436, Z => n291);
   U233 : CLKBUF_X1 port map( A => n437, Z => n297);
   U234 : CLKBUF_X1 port map( A => n495, Z => n303);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity MUX_GENERIC_N64_RADIX3_13 is

   port( plusA, minusA, plus2A, minus2A : in std_logic_vector (63 downto 0);  
         SEL : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (63 
         downto 0));

end MUX_GENERIC_N64_RADIX3_13;

architecture SYN_beh of MUX_GENERIC_N64_RADIX3_13 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component TBUF_X1
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   component TBUF_X4
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, 
      n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, 
      n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, 
      n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, 
      n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, 
      n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, 
      n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, 
      n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, 
      n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, 
      n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, 
      n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, 
      n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, 
      n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, 
      n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, 
      n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, 
      n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, 
      n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, 
      n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, 
      n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, 
      n499, n500, n501, n502 : std_logic;

begin
   
   U194 : NOR3_X2 port map( A1 => SEL(0), A2 => SEL(2), A3 => n302, ZN => n434)
                           ;
   U198 : NOR3_X2 port map( A1 => n302, A2 => SEL(2), A3 => n303, ZN => n432);
   U199 : NOR3_X2 port map( A1 => SEL(1), A2 => SEL(2), A3 => n303, ZN => n433)
                           ;
   Y_tri_60_inst : TBUF_X1 port map( A => n441, EN => n301, Z => Y(60));
   Y_tri_61_inst : TBUF_X1 port map( A => n440, EN => n301, Z => Y(61));
   Y_tri_62_inst : TBUF_X1 port map( A => n439, EN => n301, Z => Y(62));
   Y_tri_63_inst : TBUF_X1 port map( A => n438, EN => n301, Z => Y(63));
   Y_tri_53_inst : TBUF_X1 port map( A => n448, EN => n300, Z => Y(53));
   Y_tri_54_inst : TBUF_X1 port map( A => n447, EN => n300, Z => Y(54));
   Y_tri_55_inst : TBUF_X1 port map( A => n446, EN => n300, Z => Y(55));
   Y_tri_56_inst : TBUF_X1 port map( A => n445, EN => n300, Z => Y(56));
   Y_tri_57_inst : TBUF_X1 port map( A => n444, EN => n300, Z => Y(57));
   Y_tri_59_inst : TBUF_X1 port map( A => n442, EN => n300, Z => Y(59));
   Y_tri_58_inst : TBUF_X1 port map( A => n443, EN => n300, Z => Y(58));
   Y_tri_32_inst : TBUF_X1 port map( A => n469, EN => n298, Z => Y(32));
   Y_tri_33_inst : TBUF_X1 port map( A => n468, EN => n298, Z => Y(33));
   Y_tri_34_inst : TBUF_X1 port map( A => n467, EN => n298, Z => Y(34));
   Y_tri_35_inst : TBUF_X1 port map( A => n466, EN => n298, Z => Y(35));
   Y_tri_37_inst : TBUF_X1 port map( A => n464, EN => n299, Z => Y(37));
   Y_tri_38_inst : TBUF_X1 port map( A => n463, EN => n299, Z => Y(38));
   Y_tri_39_inst : TBUF_X1 port map( A => n462, EN => n299, Z => Y(39));
   Y_tri_40_inst : TBUF_X1 port map( A => n461, EN => n299, Z => Y(40));
   Y_tri_41_inst : TBUF_X1 port map( A => n460, EN => n299, Z => Y(41));
   Y_tri_42_inst : TBUF_X1 port map( A => n459, EN => n299, Z => Y(42));
   Y_tri_43_inst : TBUF_X1 port map( A => n458, EN => n299, Z => Y(43));
   Y_tri_44_inst : TBUF_X1 port map( A => n457, EN => n299, Z => Y(44));
   Y_tri_45_inst : TBUF_X1 port map( A => n456, EN => n299, Z => Y(45));
   Y_tri_46_inst : TBUF_X1 port map( A => n455, EN => n299, Z => Y(46));
   Y_tri_47_inst : TBUF_X1 port map( A => n454, EN => n299, Z => Y(47));
   Y_tri_48_inst : TBUF_X1 port map( A => n453, EN => n300, Z => Y(48));
   Y_tri_49_inst : TBUF_X1 port map( A => n452, EN => n300, Z => Y(49));
   Y_tri_50_inst : TBUF_X1 port map( A => n451, EN => n300, Z => Y(50));
   Y_tri_51_inst : TBUF_X1 port map( A => n450, EN => n300, Z => Y(51));
   Y_tri_52_inst : TBUF_X1 port map( A => n449, EN => n300, Z => Y(52));
   Y_tri_25_inst : TBUF_X1 port map( A => n476, EN => n298, Z => Y(25));
   Y_tri_24_inst : TBUF_X1 port map( A => n477, EN => n298, Z => Y(24));
   Y_tri_23_inst : TBUF_X1 port map( A => n478, EN => n297, Z => Y(23));
   Y_tri_22_inst : TBUF_X1 port map( A => n479, EN => n297, Z => Y(22));
   Y_tri_21_inst : TBUF_X1 port map( A => n480, EN => n297, Z => Y(21));
   Y_tri_20_inst : TBUF_X1 port map( A => n481, EN => n297, Z => Y(20));
   Y_tri_19_inst : TBUF_X1 port map( A => n482, EN => n297, Z => Y(19));
   Y_tri_18_inst : TBUF_X1 port map( A => n483, EN => n297, Z => Y(18));
   Y_tri_26_inst : TBUF_X1 port map( A => n475, EN => n298, Z => Y(26));
   Y_tri_17_inst : TBUF_X1 port map( A => n484, EN => n297, Z => Y(17));
   Y_tri_27_inst : TBUF_X1 port map( A => n474, EN => n298, Z => Y(27));
   Y_tri_28_inst : TBUF_X1 port map( A => n473, EN => n298, Z => Y(28));
   Y_tri_30_inst : TBUF_X1 port map( A => n471, EN => n298, Z => Y(30));
   Y_tri_16_inst : TBUF_X1 port map( A => n485, EN => n297, Z => Y(16));
   Y_tri_31_inst : TBUF_X1 port map( A => n470, EN => n298, Z => Y(31));
   Y_tri_15_inst : TBUF_X1 port map( A => n486, EN => n297, Z => Y(15));
   Y_tri_14_inst : TBUF_X1 port map( A => n487, EN => n297, Z => Y(14));
   Y_tri_13_inst : TBUF_X1 port map( A => n488, EN => n297, Z => Y(13));
   Y_tri_12_inst : TBUF_X1 port map( A => n489, EN => n297, Z => Y(12));
   Y_tri_6_inst : TBUF_X1 port map( A => n496, EN => n296, Z => Y(6));
   Y_tri_7_inst : TBUF_X1 port map( A => n495, EN => n296, Z => Y(7));
   Y_tri_8_inst : TBUF_X1 port map( A => n494, EN => n296, Z => Y(8));
   Y_tri_9_inst : TBUF_X1 port map( A => n492, EN => n296, Z => Y(9));
   Y_tri_10_inst : TBUF_X1 port map( A => n491, EN => n296, Z => Y(10));
   Y_tri_11_inst : TBUF_X1 port map( A => n490, EN => n296, Z => Y(11));
   Y_tri_36_inst : TBUF_X1 port map( A => n465, EN => n299, Z => Y(36));
   Y_tri_4_inst : TBUF_X1 port map( A => n498, EN => n296, Z => Y(4));
   Y_tri_3_inst : TBUF_X1 port map( A => n499, EN => n296, Z => Y(3));
   Y_tri_1_inst : TBUF_X1 port map( A => n501, EN => n296, Z => Y(1));
   Y_tri_2_inst : TBUF_X1 port map( A => n500, EN => n296, Z => Y(2));
   Y_tri_0_inst : TBUF_X1 port map( A => n502, EN => n296, Z => Y(0));
   Y_tri_5_inst : TBUF_X4 port map( A => n497, EN => n296, Z => Y(5));
   Y_tri_29_inst : TBUF_X1 port map( A => n472, EN => n298, Z => Y(29));
   U2 : CLKBUF_X3 port map( A => n493, Z => n296);
   U3 : CLKBUF_X1 port map( A => n435, Z => n292);
   U4 : CLKBUF_X1 port map( A => n435, Z => n293);
   U5 : CLKBUF_X1 port map( A => n435, Z => n294);
   U6 : CLKBUF_X1 port map( A => n493, Z => n298);
   U7 : CLKBUF_X1 port map( A => n493, Z => n297);
   U8 : CLKBUF_X1 port map( A => n435, Z => n291);
   U9 : CLKBUF_X1 port map( A => n493, Z => n299);
   U10 : CLKBUF_X1 port map( A => n493, Z => n300);
   U11 : BUF_X1 port map( A => n433, Z => n278);
   U12 : CLKBUF_X1 port map( A => n433, Z => n279);
   U13 : CLKBUF_X1 port map( A => n433, Z => n280);
   U14 : BUF_X1 port map( A => n434, Z => n284);
   U15 : BUF_X1 port map( A => n432, Z => n272);
   U16 : CLKBUF_X1 port map( A => n434, Z => n285);
   U17 : CLKBUF_X1 port map( A => n432, Z => n273);
   U18 : CLKBUF_X1 port map( A => n434, Z => n286);
   U19 : CLKBUF_X1 port map( A => n432, Z => n274);
   U20 : BUF_X1 port map( A => n435, Z => n290);
   U21 : NAND2_X1 port map( A1 => n403, A2 => n402, ZN => n453);
   U22 : AOI22_X1 port map( A1 => plusA(48), A2 => n282, B1 => plus2A(48), B2 
                           => n276, ZN => n403);
   U23 : AOI22_X1 port map( A1 => minus2A(48), A2 => n294, B1 => minusA(48), B2
                           => n288, ZN => n402);
   U24 : NAND2_X1 port map( A1 => n393, A2 => n392, ZN => n458);
   U25 : AOI22_X1 port map( A1 => plusA(43), A2 => n281, B1 => plus2A(43), B2 
                           => n275, ZN => n393);
   U26 : AOI22_X1 port map( A1 => minus2A(43), A2 => n293, B1 => minusA(43), B2
                           => n287, ZN => n392);
   U27 : NAND2_X1 port map( A1 => n383, A2 => n382, ZN => n463);
   U28 : AOI22_X1 port map( A1 => plusA(38), A2 => n281, B1 => plus2A(38), B2 
                           => n275, ZN => n383);
   U29 : AOI22_X1 port map( A1 => minus2A(38), A2 => n293, B1 => minusA(38), B2
                           => n287, ZN => n382);
   U30 : NAND2_X1 port map( A1 => n381, A2 => n380, ZN => n464);
   U31 : AOI22_X1 port map( A1 => plusA(37), A2 => n281, B1 => plus2A(37), B2 
                           => n275, ZN => n381);
   U32 : AOI22_X1 port map( A1 => minus2A(37), A2 => n293, B1 => minusA(37), B2
                           => n287, ZN => n380);
   U33 : NAND2_X1 port map( A1 => n379, A2 => n378, ZN => n465);
   U34 : AOI22_X1 port map( A1 => plusA(36), A2 => n281, B1 => plus2A(36), B2 
                           => n275, ZN => n379);
   U35 : AOI22_X1 port map( A1 => minus2A(36), A2 => n293, B1 => minusA(36), B2
                           => n287, ZN => n378);
   U36 : NAND2_X1 port map( A1 => n395, A2 => n394, ZN => n457);
   U37 : AOI22_X1 port map( A1 => plusA(44), A2 => n281, B1 => plus2A(44), B2 
                           => n275, ZN => n395);
   U38 : AOI22_X1 port map( A1 => minus2A(44), A2 => n293, B1 => minusA(44), B2
                           => n287, ZN => n394);
   U39 : CLKBUF_X1 port map( A => n433, Z => n281);
   U40 : CLKBUF_X1 port map( A => n434, Z => n287);
   U41 : CLKBUF_X1 port map( A => n432, Z => n275);
   U42 : NAND2_X1 port map( A1 => n423, A2 => n422, ZN => n443);
   U43 : AOI22_X1 port map( A1 => plusA(58), A2 => n282, B1 => plus2A(58), B2 
                           => n276, ZN => n423);
   U44 : AOI22_X1 port map( A1 => minus2A(58), A2 => n294, B1 => minusA(58), B2
                           => n288, ZN => n422);
   U45 : NAND2_X1 port map( A1 => n421, A2 => n420, ZN => n444);
   U46 : AOI22_X1 port map( A1 => plusA(57), A2 => n282, B1 => plus2A(57), B2 
                           => n276, ZN => n421);
   U47 : AOI22_X1 port map( A1 => minus2A(57), A2 => n294, B1 => minusA(57), B2
                           => n288, ZN => n420);
   U48 : NAND2_X1 port map( A1 => n415, A2 => n414, ZN => n447);
   U49 : AOI22_X1 port map( A1 => plusA(54), A2 => n282, B1 => plus2A(54), B2 
                           => n276, ZN => n415);
   U50 : AOI22_X1 port map( A1 => minus2A(54), A2 => n294, B1 => minusA(54), B2
                           => n288, ZN => n414);
   U51 : NAND2_X1 port map( A1 => n413, A2 => n412, ZN => n448);
   U52 : AOI22_X1 port map( A1 => plusA(53), A2 => n282, B1 => plus2A(53), B2 
                           => n276, ZN => n413);
   U53 : AOI22_X1 port map( A1 => minus2A(53), A2 => n294, B1 => minusA(53), B2
                           => n288, ZN => n412);
   U54 : CLKBUF_X1 port map( A => n433, Z => n282);
   U55 : CLKBUF_X1 port map( A => n434, Z => n288);
   U56 : CLKBUF_X1 port map( A => n432, Z => n276);
   U57 : NOR2_X1 port map( A1 => n323, A2 => n304, ZN => n493);
   U58 : INV_X1 port map( A => SEL(2), ZN => n304);
   U59 : NOR2_X1 port map( A1 => SEL(1), A2 => SEL(0), ZN => n323);
   U60 : AND2_X1 port map( A1 => SEL(2), A2 => n323, ZN => n435);
   U61 : NAND2_X1 port map( A1 => n322, A2 => n321, ZN => n494);
   U62 : AOI22_X1 port map( A1 => plusA(8), A2 => n278, B1 => plus2A(8), B2 => 
                           n272, ZN => n322);
   U63 : AOI22_X1 port map( A1 => minus2A(8), A2 => n290, B1 => minusA(8), B2 
                           => n284, ZN => n321);
   U64 : INV_X1 port map( A => SEL(1), ZN => n302);
   U65 : INV_X1 port map( A => SEL(0), ZN => n303);
   U66 : NAND2_X1 port map( A1 => n407, A2 => n406, ZN => n451);
   U67 : AOI22_X1 port map( A1 => plusA(50), A2 => n282, B1 => plus2A(50), B2 
                           => n276, ZN => n407);
   U68 : AOI22_X1 port map( A1 => minus2A(50), A2 => n294, B1 => minusA(50), B2
                           => n288, ZN => n406);
   U69 : NAND2_X1 port map( A1 => n320, A2 => n319, ZN => n495);
   U70 : AOI22_X1 port map( A1 => plusA(7), A2 => n278, B1 => plus2A(7), B2 => 
                           n272, ZN => n320);
   U71 : AOI22_X1 port map( A1 => minus2A(7), A2 => n290, B1 => minusA(7), B2 
                           => n284, ZN => n319);
   U72 : NAND2_X1 port map( A1 => n329, A2 => n328, ZN => n490);
   U73 : AOI22_X1 port map( A1 => plusA(11), A2 => n278, B1 => plus2A(11), B2 
                           => n272, ZN => n329);
   U74 : AOI22_X1 port map( A1 => minus2A(11), A2 => n290, B1 => minusA(11), B2
                           => n284, ZN => n328);
   U75 : NAND2_X1 port map( A1 => n337, A2 => n336, ZN => n486);
   U76 : AOI22_X1 port map( A1 => plusA(15), A2 => n279, B1 => plus2A(15), B2 
                           => n273, ZN => n337);
   U77 : AOI22_X1 port map( A1 => minus2A(15), A2 => n291, B1 => minusA(15), B2
                           => n285, ZN => n336);
   U78 : NAND2_X1 port map( A1 => n369, A2 => n368, ZN => n470);
   U79 : AOI22_X1 port map( A1 => plusA(31), A2 => n280, B1 => plus2A(31), B2 
                           => n274, ZN => n369);
   U80 : AOI22_X1 port map( A1 => minus2A(31), A2 => n292, B1 => minusA(31), B2
                           => n286, ZN => n368);
   U81 : NAND2_X1 port map( A1 => n361, A2 => n360, ZN => n474);
   U82 : AOI22_X1 port map( A1 => plusA(27), A2 => n280, B1 => plus2A(27), B2 
                           => n274, ZN => n361);
   U83 : AOI22_X1 port map( A1 => minus2A(27), A2 => n292, B1 => minusA(27), B2
                           => n286, ZN => n360);
   U84 : NAND2_X1 port map( A1 => n345, A2 => n344, ZN => n482);
   U85 : AOI22_X1 port map( A1 => plusA(19), A2 => n279, B1 => plus2A(19), B2 
                           => n273, ZN => n345);
   U86 : AOI22_X1 port map( A1 => minus2A(19), A2 => n291, B1 => minusA(19), B2
                           => n285, ZN => n344);
   U87 : NAND2_X1 port map( A1 => n353, A2 => n352, ZN => n478);
   U88 : AOI22_X1 port map( A1 => plusA(23), A2 => n279, B1 => plus2A(23), B2 
                           => n273, ZN => n353);
   U89 : AOI22_X1 port map( A1 => minus2A(23), A2 => n291, B1 => minusA(23), B2
                           => n285, ZN => n352);
   U90 : NAND2_X1 port map( A1 => n397, A2 => n396, ZN => n456);
   U91 : AOI22_X1 port map( A1 => plusA(45), A2 => n281, B1 => plus2A(45), B2 
                           => n275, ZN => n397);
   U92 : AOI22_X1 port map( A1 => minus2A(45), A2 => n293, B1 => minusA(45), B2
                           => n287, ZN => n396);
   U93 : NAND2_X1 port map( A1 => n377, A2 => n376, ZN => n466);
   U94 : AOI22_X1 port map( A1 => plusA(35), A2 => n280, B1 => plus2A(35), B2 
                           => n274, ZN => n377);
   U95 : AOI22_X1 port map( A1 => minus2A(35), A2 => n292, B1 => minusA(35), B2
                           => n286, ZN => n376);
   U96 : NAND2_X1 port map( A1 => n401, A2 => n400, ZN => n454);
   U97 : AOI22_X1 port map( A1 => plusA(47), A2 => n281, B1 => plus2A(47), B2 
                           => n275, ZN => n401);
   U98 : AOI22_X1 port map( A1 => minus2A(47), A2 => n293, B1 => minusA(47), B2
                           => n287, ZN => n400);
   U99 : NAND2_X1 port map( A1 => n387, A2 => n386, ZN => n461);
   U100 : AOI22_X1 port map( A1 => plusA(40), A2 => n281, B1 => plus2A(40), B2 
                           => n275, ZN => n387);
   U101 : AOI22_X1 port map( A1 => minus2A(40), A2 => n293, B1 => minusA(40), 
                           B2 => n287, ZN => n386);
   U102 : NAND2_X1 port map( A1 => n325, A2 => n324, ZN => n492);
   U103 : AOI22_X1 port map( A1 => plusA(9), A2 => n278, B1 => plus2A(9), B2 =>
                           n272, ZN => n325);
   U104 : AOI22_X1 port map( A1 => minus2A(9), A2 => n290, B1 => minusA(9), B2 
                           => n284, ZN => n324);
   U105 : NAND2_X1 port map( A1 => n333, A2 => n332, ZN => n488);
   U106 : AOI22_X1 port map( A1 => plusA(13), A2 => n279, B1 => plus2A(13), B2 
                           => n273, ZN => n333);
   U107 : AOI22_X1 port map( A1 => minus2A(13), A2 => n291, B1 => minusA(13), 
                           B2 => n285, ZN => n332);
   U108 : NAND2_X1 port map( A1 => n341, A2 => n340, ZN => n484);
   U109 : AOI22_X1 port map( A1 => plusA(17), A2 => n279, B1 => plus2A(17), B2 
                           => n273, ZN => n341);
   U110 : AOI22_X1 port map( A1 => minus2A(17), A2 => n291, B1 => minusA(17), 
                           B2 => n285, ZN => n340);
   U111 : NAND2_X1 port map( A1 => n365, A2 => n364, ZN => n472);
   U112 : AOI22_X1 port map( A1 => plusA(29), A2 => n280, B1 => plus2A(29), B2 
                           => n274, ZN => n365);
   U113 : AOI22_X1 port map( A1 => minus2A(29), A2 => n292, B1 => minusA(29), 
                           B2 => n286, ZN => n364);
   U114 : NAND2_X1 port map( A1 => n349, A2 => n348, ZN => n480);
   U115 : AOI22_X1 port map( A1 => plusA(21), A2 => n279, B1 => plus2A(21), B2 
                           => n273, ZN => n349);
   U116 : AOI22_X1 port map( A1 => minus2A(21), A2 => n291, B1 => minusA(21), 
                           B2 => n285, ZN => n348);
   U117 : NAND2_X1 port map( A1 => n357, A2 => n356, ZN => n476);
   U118 : AOI22_X1 port map( A1 => plusA(25), A2 => n280, B1 => plus2A(25), B2 
                           => n274, ZN => n357);
   U119 : AOI22_X1 port map( A1 => minus2A(25), A2 => n292, B1 => minusA(25), 
                           B2 => n286, ZN => n356);
   U120 : NAND2_X1 port map( A1 => n373, A2 => n372, ZN => n468);
   U121 : AOI22_X1 port map( A1 => plusA(33), A2 => n280, B1 => plus2A(33), B2 
                           => n274, ZN => n373);
   U122 : AOI22_X1 port map( A1 => minus2A(33), A2 => n292, B1 => minusA(33), 
                           B2 => n286, ZN => n372);
   U123 : NAND2_X1 port map( A1 => n405, A2 => n404, ZN => n452);
   U124 : AOI22_X1 port map( A1 => plusA(49), A2 => n282, B1 => plus2A(49), B2 
                           => n276, ZN => n405);
   U125 : AOI22_X1 port map( A1 => minus2A(49), A2 => n294, B1 => minusA(49), 
                           B2 => n288, ZN => n404);
   U126 : NAND2_X1 port map( A1 => n409, A2 => n408, ZN => n450);
   U127 : AOI22_X1 port map( A1 => plusA(51), A2 => n282, B1 => plus2A(51), B2 
                           => n276, ZN => n409);
   U128 : AOI22_X1 port map( A1 => minus2A(51), A2 => n294, B1 => minusA(51), 
                           B2 => n288, ZN => n408);
   U129 : NAND2_X1 port map( A1 => n331, A2 => n330, ZN => n489);
   U130 : AOI22_X1 port map( A1 => plusA(12), A2 => n279, B1 => plus2A(12), B2 
                           => n273, ZN => n331);
   U131 : AOI22_X1 port map( A1 => minus2A(12), A2 => n291, B1 => minusA(12), 
                           B2 => n285, ZN => n330);
   U132 : NAND2_X1 port map( A1 => n339, A2 => n338, ZN => n485);
   U133 : AOI22_X1 port map( A1 => plusA(16), A2 => n279, B1 => plus2A(16), B2 
                           => n273, ZN => n339);
   U134 : AOI22_X1 port map( A1 => minus2A(16), A2 => n291, B1 => minusA(16), 
                           B2 => n285, ZN => n338);
   U135 : NAND2_X1 port map( A1 => n363, A2 => n362, ZN => n473);
   U136 : AOI22_X1 port map( A1 => plusA(28), A2 => n280, B1 => plus2A(28), B2 
                           => n274, ZN => n363);
   U137 : AOI22_X1 port map( A1 => minus2A(28), A2 => n292, B1 => minusA(28), 
                           B2 => n286, ZN => n362);
   U138 : NAND2_X1 port map( A1 => n347, A2 => n346, ZN => n481);
   U139 : AOI22_X1 port map( A1 => plusA(20), A2 => n279, B1 => plus2A(20), B2 
                           => n273, ZN => n347);
   U140 : AOI22_X1 port map( A1 => minus2A(20), A2 => n291, B1 => minusA(20), 
                           B2 => n285, ZN => n346);
   U141 : NAND2_X1 port map( A1 => n355, A2 => n354, ZN => n477);
   U142 : AOI22_X1 port map( A1 => plusA(24), A2 => n280, B1 => plus2A(24), B2 
                           => n274, ZN => n355);
   U143 : AOI22_X1 port map( A1 => minus2A(24), A2 => n292, B1 => minusA(24), 
                           B2 => n286, ZN => n354);
   U144 : NAND2_X1 port map( A1 => n411, A2 => n410, ZN => n449);
   U145 : AOI22_X1 port map( A1 => plusA(52), A2 => n282, B1 => plus2A(52), B2 
                           => n276, ZN => n411);
   U146 : AOI22_X1 port map( A1 => minus2A(52), A2 => n294, B1 => minusA(52), 
                           B2 => n288, ZN => n410);
   U147 : NAND2_X1 port map( A1 => n371, A2 => n370, ZN => n469);
   U148 : AOI22_X1 port map( A1 => plusA(32), A2 => n280, B1 => plus2A(32), B2 
                           => n274, ZN => n371);
   U149 : AOI22_X1 port map( A1 => minus2A(32), A2 => n292, B1 => minusA(32), 
                           B2 => n286, ZN => n370);
   U150 : NAND2_X1 port map( A1 => n385, A2 => n384, ZN => n462);
   U151 : AOI22_X1 port map( A1 => plusA(39), A2 => n281, B1 => plus2A(39), B2 
                           => n275, ZN => n385);
   U152 : AOI22_X1 port map( A1 => minus2A(39), A2 => n293, B1 => minusA(39), 
                           B2 => n287, ZN => n384);
   U153 : NAND2_X1 port map( A1 => n389, A2 => n388, ZN => n460);
   U154 : AOI22_X1 port map( A1 => plusA(41), A2 => n281, B1 => plus2A(41), B2 
                           => n275, ZN => n389);
   U155 : AOI22_X1 port map( A1 => minus2A(41), A2 => n293, B1 => minusA(41), 
                           B2 => n287, ZN => n388);
   U156 : NAND2_X1 port map( A1 => n327, A2 => n326, ZN => n491);
   U157 : AOI22_X1 port map( A1 => plusA(10), A2 => n278, B1 => plus2A(10), B2 
                           => n272, ZN => n327);
   U158 : AOI22_X1 port map( A1 => minus2A(10), A2 => n290, B1 => minusA(10), 
                           B2 => n284, ZN => n326);
   U159 : NAND2_X1 port map( A1 => n335, A2 => n334, ZN => n487);
   U160 : AOI22_X1 port map( A1 => plusA(14), A2 => n279, B1 => plus2A(14), B2 
                           => n273, ZN => n335);
   U161 : AOI22_X1 port map( A1 => minus2A(14), A2 => n291, B1 => minusA(14), 
                           B2 => n285, ZN => n334);
   U162 : NAND2_X1 port map( A1 => n367, A2 => n366, ZN => n471);
   U163 : AOI22_X1 port map( A1 => plusA(30), A2 => n280, B1 => plus2A(30), B2 
                           => n274, ZN => n367);
   U164 : AOI22_X1 port map( A1 => minus2A(30), A2 => n292, B1 => minusA(30), 
                           B2 => n286, ZN => n366);
   U165 : NAND2_X1 port map( A1 => n359, A2 => n358, ZN => n475);
   U166 : AOI22_X1 port map( A1 => plusA(26), A2 => n280, B1 => plus2A(26), B2 
                           => n274, ZN => n359);
   U167 : AOI22_X1 port map( A1 => minus2A(26), A2 => n292, B1 => minusA(26), 
                           B2 => n286, ZN => n358);
   U168 : NAND2_X1 port map( A1 => n343, A2 => n342, ZN => n483);
   U169 : AOI22_X1 port map( A1 => plusA(18), A2 => n279, B1 => plus2A(18), B2 
                           => n273, ZN => n343);
   U170 : AOI22_X1 port map( A1 => minus2A(18), A2 => n291, B1 => minusA(18), 
                           B2 => n285, ZN => n342);
   U171 : NAND2_X1 port map( A1 => n351, A2 => n350, ZN => n479);
   U172 : AOI22_X1 port map( A1 => plusA(22), A2 => n279, B1 => plus2A(22), B2 
                           => n273, ZN => n351);
   U173 : AOI22_X1 port map( A1 => minus2A(22), A2 => n291, B1 => minusA(22), 
                           B2 => n285, ZN => n350);
   U174 : NAND2_X1 port map( A1 => n391, A2 => n390, ZN => n459);
   U175 : AOI22_X1 port map( A1 => plusA(42), A2 => n281, B1 => plus2A(42), B2 
                           => n275, ZN => n391);
   U176 : AOI22_X1 port map( A1 => minus2A(42), A2 => n293, B1 => minusA(42), 
                           B2 => n287, ZN => n390);
   U177 : NAND2_X1 port map( A1 => n375, A2 => n374, ZN => n467);
   U178 : AOI22_X1 port map( A1 => plusA(34), A2 => n280, B1 => plus2A(34), B2 
                           => n274, ZN => n375);
   U179 : AOI22_X1 port map( A1 => minus2A(34), A2 => n292, B1 => minusA(34), 
                           B2 => n286, ZN => n374);
   U180 : NAND2_X1 port map( A1 => n399, A2 => n398, ZN => n455);
   U181 : AOI22_X1 port map( A1 => plusA(46), A2 => n281, B1 => plus2A(46), B2 
                           => n275, ZN => n399);
   U182 : AOI22_X1 port map( A1 => minus2A(46), A2 => n293, B1 => minusA(46), 
                           B2 => n287, ZN => n398);
   U183 : NAND2_X1 port map( A1 => n437, A2 => n436, ZN => n438);
   U184 : AOI22_X1 port map( A1 => plusA(63), A2 => n283, B1 => plus2A(63), B2 
                           => n277, ZN => n437);
   U185 : AOI22_X1 port map( A1 => minus2A(63), A2 => n295, B1 => minusA(63), 
                           B2 => n289, ZN => n436);
   U186 : NAND2_X1 port map( A1 => n431, A2 => n430, ZN => n439);
   U187 : AOI22_X1 port map( A1 => plusA(62), A2 => n283, B1 => plus2A(62), B2 
                           => n277, ZN => n431);
   U188 : AOI22_X1 port map( A1 => minus2A(62), A2 => n295, B1 => minusA(62), 
                           B2 => n289, ZN => n430);
   U189 : NAND2_X1 port map( A1 => n429, A2 => n428, ZN => n440);
   U190 : AOI22_X1 port map( A1 => plusA(61), A2 => n283, B1 => plus2A(61), B2 
                           => n277, ZN => n429);
   U191 : AOI22_X1 port map( A1 => minus2A(61), A2 => n295, B1 => minusA(61), 
                           B2 => n289, ZN => n428);
   U192 : NAND2_X1 port map( A1 => n427, A2 => n426, ZN => n441);
   U193 : AOI22_X1 port map( A1 => plusA(60), A2 => n283, B1 => plus2A(60), B2 
                           => n277, ZN => n427);
   U195 : AOI22_X1 port map( A1 => minus2A(60), A2 => n295, B1 => minusA(60), 
                           B2 => n289, ZN => n426);
   U196 : NAND2_X1 port map( A1 => n425, A2 => n424, ZN => n442);
   U197 : AOI22_X1 port map( A1 => plusA(59), A2 => n282, B1 => plus2A(59), B2 
                           => n276, ZN => n425);
   U200 : AOI22_X1 port map( A1 => minus2A(59), A2 => n294, B1 => minusA(59), 
                           B2 => n288, ZN => n424);
   U201 : NAND2_X1 port map( A1 => n419, A2 => n418, ZN => n445);
   U202 : AOI22_X1 port map( A1 => plusA(56), A2 => n282, B1 => plus2A(56), B2 
                           => n276, ZN => n419);
   U203 : AOI22_X1 port map( A1 => minus2A(56), A2 => n294, B1 => minusA(56), 
                           B2 => n288, ZN => n418);
   U204 : NAND2_X1 port map( A1 => n417, A2 => n416, ZN => n446);
   U205 : AOI22_X1 port map( A1 => plusA(55), A2 => n282, B1 => plus2A(55), B2 
                           => n276, ZN => n417);
   U206 : AOI22_X1 port map( A1 => minus2A(55), A2 => n294, B1 => minusA(55), 
                           B2 => n288, ZN => n416);
   U207 : NAND2_X1 port map( A1 => n318, A2 => n317, ZN => n496);
   U208 : AOI22_X1 port map( A1 => plusA(6), A2 => n278, B1 => plus2A(6), B2 =>
                           n272, ZN => n318);
   U209 : AOI22_X1 port map( A1 => minus2A(6), A2 => n290, B1 => minusA(6), B2 
                           => n284, ZN => n317);
   U210 : NAND2_X1 port map( A1 => n316, A2 => n315, ZN => n497);
   U211 : AOI22_X1 port map( A1 => plusA(5), A2 => n278, B1 => plus2A(5), B2 =>
                           n272, ZN => n316);
   U212 : AOI22_X1 port map( A1 => minus2A(5), A2 => n290, B1 => minusA(5), B2 
                           => n284, ZN => n315);
   U213 : NAND2_X1 port map( A1 => n312, A2 => n311, ZN => n499);
   U214 : AOI22_X1 port map( A1 => plusA(3), A2 => n278, B1 => plus2A(3), B2 =>
                           n272, ZN => n312);
   U215 : AOI22_X1 port map( A1 => minus2A(3), A2 => n290, B1 => minusA(3), B2 
                           => n284, ZN => n311);
   U216 : NAND2_X1 port map( A1 => n314, A2 => n313, ZN => n498);
   U217 : AOI22_X1 port map( A1 => plusA(4), A2 => n278, B1 => plus2A(4), B2 =>
                           n272, ZN => n314);
   U218 : AOI22_X1 port map( A1 => minus2A(4), A2 => n290, B1 => minusA(4), B2 
                           => n284, ZN => n313);
   U219 : NAND2_X1 port map( A1 => n310, A2 => n309, ZN => n500);
   U220 : AOI22_X1 port map( A1 => plusA(2), A2 => n278, B1 => plus2A(2), B2 =>
                           n272, ZN => n310);
   U221 : AOI22_X1 port map( A1 => minus2A(2), A2 => n290, B1 => minusA(2), B2 
                           => n284, ZN => n309);
   U222 : NAND2_X1 port map( A1 => n308, A2 => n307, ZN => n501);
   U223 : AOI22_X1 port map( A1 => plusA(1), A2 => n278, B1 => plus2A(1), B2 =>
                           n272, ZN => n308);
   U224 : AOI22_X1 port map( A1 => minus2A(1), A2 => n290, B1 => minusA(1), B2 
                           => n284, ZN => n307);
   U225 : NAND2_X1 port map( A1 => n306, A2 => n305, ZN => n502);
   U226 : AOI22_X1 port map( A1 => plusA(0), A2 => n278, B1 => plus2A(0), B2 =>
                           n272, ZN => n306);
   U227 : AOI22_X1 port map( A1 => minus2A(0), A2 => n290, B1 => minusA(0), B2 
                           => n284, ZN => n305);
   U228 : CLKBUF_X1 port map( A => n432, Z => n277);
   U229 : CLKBUF_X1 port map( A => n433, Z => n283);
   U230 : CLKBUF_X1 port map( A => n434, Z => n289);
   U231 : CLKBUF_X1 port map( A => n435, Z => n295);
   U232 : CLKBUF_X1 port map( A => n493, Z => n301);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity MUX_GENERIC_N64_RADIX3_11 is

   port( plusA, minusA, plus2A, minus2A : in std_logic_vector (63 downto 0);  
         SEL : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (63 
         downto 0));

end MUX_GENERIC_N64_RADIX3_11;

architecture SYN_beh of MUX_GENERIC_N64_RADIX3_11 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component TBUF_X1
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   component TBUF_X4
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   signal n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, 
      n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, 
      n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, 
      n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, 
      n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, 
      n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, 
      n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, 
      n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, 
      n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, 
      n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, 
      n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, 
      n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, 
      n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, 
      n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, 
      n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, 
      n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, 
      n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, 
      n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, 
      n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, 
      n499, n500, n501, n502 : std_logic;

begin
   
   Y_tri_60_inst : TBUF_X1 port map( A => n441, EN => n301, Z => Y(60));
   Y_tri_61_inst : TBUF_X1 port map( A => n440, EN => n301, Z => Y(61));
   Y_tri_62_inst : TBUF_X1 port map( A => n439, EN => n301, Z => Y(62));
   Y_tri_63_inst : TBUF_X1 port map( A => n438, EN => n301, Z => Y(63));
   Y_tri_40_inst : TBUF_X1 port map( A => n461, EN => n299, Z => Y(40));
   Y_tri_41_inst : TBUF_X1 port map( A => n460, EN => n299, Z => Y(41));
   Y_tri_42_inst : TBUF_X1 port map( A => n459, EN => n299, Z => Y(42));
   Y_tri_43_inst : TBUF_X1 port map( A => n458, EN => n299, Z => Y(43));
   Y_tri_44_inst : TBUF_X1 port map( A => n457, EN => n299, Z => Y(44));
   Y_tri_45_inst : TBUF_X1 port map( A => n456, EN => n299, Z => Y(45));
   Y_tri_46_inst : TBUF_X1 port map( A => n455, EN => n299, Z => Y(46));
   Y_tri_47_inst : TBUF_X1 port map( A => n454, EN => n299, Z => Y(47));
   Y_tri_48_inst : TBUF_X1 port map( A => n453, EN => n300, Z => Y(48));
   Y_tri_49_inst : TBUF_X1 port map( A => n452, EN => n300, Z => Y(49));
   Y_tri_50_inst : TBUF_X1 port map( A => n451, EN => n300, Z => Y(50));
   Y_tri_51_inst : TBUF_X1 port map( A => n450, EN => n300, Z => Y(51));
   Y_tri_52_inst : TBUF_X1 port map( A => n449, EN => n300, Z => Y(52));
   Y_tri_53_inst : TBUF_X1 port map( A => n448, EN => n300, Z => Y(53));
   Y_tri_54_inst : TBUF_X1 port map( A => n447, EN => n300, Z => Y(54));
   Y_tri_55_inst : TBUF_X1 port map( A => n446, EN => n300, Z => Y(55));
   Y_tri_56_inst : TBUF_X1 port map( A => n445, EN => n300, Z => Y(56));
   Y_tri_57_inst : TBUF_X1 port map( A => n444, EN => n300, Z => Y(57));
   Y_tri_58_inst : TBUF_X1 port map( A => n443, EN => n300, Z => Y(58));
   Y_tri_59_inst : TBUF_X1 port map( A => n442, EN => n300, Z => Y(59));
   Y_tri_19_inst : TBUF_X1 port map( A => n482, EN => n297, Z => Y(19));
   Y_tri_20_inst : TBUF_X1 port map( A => n481, EN => n297, Z => Y(20));
   Y_tri_21_inst : TBUF_X1 port map( A => n480, EN => n297, Z => Y(21));
   Y_tri_22_inst : TBUF_X1 port map( A => n479, EN => n297, Z => Y(22));
   Y_tri_23_inst : TBUF_X1 port map( A => n478, EN => n297, Z => Y(23));
   Y_tri_24_inst : TBUF_X1 port map( A => n477, EN => n298, Z => Y(24));
   Y_tri_25_inst : TBUF_X1 port map( A => n476, EN => n298, Z => Y(25));
   Y_tri_26_inst : TBUF_X1 port map( A => n475, EN => n298, Z => Y(26));
   Y_tri_27_inst : TBUF_X1 port map( A => n474, EN => n298, Z => Y(27));
   Y_tri_28_inst : TBUF_X1 port map( A => n473, EN => n298, Z => Y(28));
   Y_tri_29_inst : TBUF_X1 port map( A => n472, EN => n298, Z => Y(29));
   Y_tri_30_inst : TBUF_X1 port map( A => n471, EN => n298, Z => Y(30));
   Y_tri_31_inst : TBUF_X1 port map( A => n470, EN => n298, Z => Y(31));
   Y_tri_32_inst : TBUF_X1 port map( A => n469, EN => n298, Z => Y(32));
   Y_tri_33_inst : TBUF_X1 port map( A => n468, EN => n298, Z => Y(33));
   Y_tri_34_inst : TBUF_X1 port map( A => n467, EN => n298, Z => Y(34));
   Y_tri_35_inst : TBUF_X1 port map( A => n466, EN => n298, Z => Y(35));
   Y_tri_36_inst : TBUF_X1 port map( A => n465, EN => n299, Z => Y(36));
   Y_tri_37_inst : TBUF_X1 port map( A => n464, EN => n299, Z => Y(37));
   Y_tri_38_inst : TBUF_X1 port map( A => n463, EN => n299, Z => Y(38));
   Y_tri_13_inst : TBUF_X1 port map( A => n488, EN => n297, Z => Y(13));
   Y_tri_12_inst : TBUF_X1 port map( A => n489, EN => n297, Z => Y(12));
   Y_tri_11_inst : TBUF_X1 port map( A => n490, EN => n296, Z => Y(11));
   Y_tri_10_inst : TBUF_X1 port map( A => n491, EN => n296, Z => Y(10));
   Y_tri_9_inst : TBUF_X1 port map( A => n492, EN => n296, Z => Y(9));
   Y_tri_14_inst : TBUF_X1 port map( A => n487, EN => n297, Z => Y(14));
   Y_tri_8_inst : TBUF_X1 port map( A => n494, EN => n296, Z => Y(8));
   Y_tri_15_inst : TBUF_X1 port map( A => n486, EN => n297, Z => Y(15));
   Y_tri_16_inst : TBUF_X1 port map( A => n485, EN => n297, Z => Y(16));
   Y_tri_17_inst : TBUF_X1 port map( A => n484, EN => n297, Z => Y(17));
   Y_tri_18_inst : TBUF_X1 port map( A => n483, EN => n297, Z => Y(18));
   Y_tri_7_inst : TBUF_X1 port map( A => n495, EN => n296, Z => Y(7));
   Y_tri_6_inst : TBUF_X1 port map( A => n496, EN => n296, Z => Y(6));
   Y_tri_5_inst : TBUF_X1 port map( A => n497, EN => n296, Z => Y(5));
   Y_tri_4_inst : TBUF_X1 port map( A => n498, EN => n296, Z => Y(4));
   Y_tri_3_inst : TBUF_X1 port map( A => n499, EN => n296, Z => Y(3));
   Y_tri_2_inst : TBUF_X1 port map( A => n500, EN => n296, Z => Y(2));
   Y_tri_1_inst : TBUF_X1 port map( A => n501, EN => n296, Z => Y(1));
   Y_tri_0_inst : TBUF_X4 port map( A => n502, EN => n296, Z => Y(0));
   Y_tri_39_inst : TBUF_X1 port map( A => n462, EN => n299, Z => Y(39));
   U2 : NOR3_X1 port map( A1 => SEL(0), A2 => SEL(2), A3 => n302, ZN => n434);
   U3 : NOR3_X1 port map( A1 => n302, A2 => SEL(2), A3 => n303, ZN => n432);
   U4 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n303, ZN => n433);
   U5 : CLKBUF_X3 port map( A => n493, Z => n296);
   U6 : CLKBUF_X1 port map( A => n493, Z => n297);
   U7 : CLKBUF_X1 port map( A => n493, Z => n298);
   U8 : CLKBUF_X1 port map( A => n493, Z => n299);
   U9 : CLKBUF_X1 port map( A => n493, Z => n300);
   U10 : NAND2_X1 port map( A1 => n423, A2 => n422, ZN => n443);
   U11 : AOI22_X1 port map( A1 => plusA(58), A2 => n282, B1 => plus2A(58), B2 
                           => n276, ZN => n423);
   U12 : AOI22_X1 port map( A1 => minus2A(58), A2 => n294, B1 => minusA(58), B2
                           => n288, ZN => n422);
   U13 : NAND2_X1 port map( A1 => n403, A2 => n402, ZN => n453);
   U14 : AOI22_X1 port map( A1 => plusA(48), A2 => n282, B1 => plus2A(48), B2 
                           => n276, ZN => n403);
   U15 : AOI22_X1 port map( A1 => minus2A(48), A2 => n294, B1 => minusA(48), B2
                           => n288, ZN => n402);
   U16 : BUF_X1 port map( A => n433, Z => n278);
   U17 : CLKBUF_X1 port map( A => n433, Z => n279);
   U18 : BUF_X1 port map( A => n434, Z => n284);
   U19 : BUF_X1 port map( A => n432, Z => n272);
   U20 : CLKBUF_X1 port map( A => n434, Z => n285);
   U21 : CLKBUF_X1 port map( A => n432, Z => n273);
   U22 : BUF_X1 port map( A => n435, Z => n291);
   U23 : BUF_X1 port map( A => n435, Z => n290);
   U24 : NAND2_X1 port map( A1 => n337, A2 => n336, ZN => n486);
   U25 : AOI22_X1 port map( A1 => plusA(15), A2 => n279, B1 => plus2A(15), B2 
                           => n273, ZN => n337);
   U26 : AOI22_X1 port map( A1 => minus2A(15), A2 => n291, B1 => minusA(15), B2
                           => n285, ZN => n336);
   U27 : NAND2_X1 port map( A1 => n385, A2 => n384, ZN => n462);
   U28 : AOI22_X1 port map( A1 => plusA(39), A2 => n281, B1 => plus2A(39), B2 
                           => n275, ZN => n385);
   U29 : AOI22_X1 port map( A1 => minus2A(39), A2 => n293, B1 => minusA(39), B2
                           => n287, ZN => n384);
   U30 : NAND2_X1 port map( A1 => n377, A2 => n376, ZN => n466);
   U31 : AOI22_X1 port map( A1 => plusA(35), A2 => n280, B1 => plus2A(35), B2 
                           => n274, ZN => n377);
   U32 : AOI22_X1 port map( A1 => minus2A(35), A2 => n292, B1 => minusA(35), B2
                           => n286, ZN => n376);
   U33 : NAND2_X1 port map( A1 => n369, A2 => n368, ZN => n470);
   U34 : AOI22_X1 port map( A1 => plusA(31), A2 => n280, B1 => plus2A(31), B2 
                           => n274, ZN => n369);
   U35 : AOI22_X1 port map( A1 => minus2A(31), A2 => n292, B1 => minusA(31), B2
                           => n286, ZN => n368);
   U36 : NAND2_X1 port map( A1 => n361, A2 => n360, ZN => n474);
   U37 : AOI22_X1 port map( A1 => plusA(27), A2 => n280, B1 => plus2A(27), B2 
                           => n274, ZN => n361);
   U38 : AOI22_X1 port map( A1 => minus2A(27), A2 => n292, B1 => minusA(27), B2
                           => n286, ZN => n360);
   U39 : NAND2_X1 port map( A1 => n353, A2 => n352, ZN => n478);
   U40 : AOI22_X1 port map( A1 => plusA(23), A2 => n279, B1 => plus2A(23), B2 
                           => n273, ZN => n353);
   U41 : AOI22_X1 port map( A1 => minus2A(23), A2 => n291, B1 => minusA(23), B2
                           => n285, ZN => n352);
   U42 : NAND2_X1 port map( A1 => n345, A2 => n344, ZN => n482);
   U43 : AOI22_X1 port map( A1 => plusA(19), A2 => n279, B1 => plus2A(19), B2 
                           => n273, ZN => n345);
   U44 : AOI22_X1 port map( A1 => minus2A(19), A2 => n291, B1 => minusA(19), B2
                           => n285, ZN => n344);
   U45 : NAND2_X1 port map( A1 => n341, A2 => n340, ZN => n484);
   U46 : AOI22_X1 port map( A1 => plusA(17), A2 => n279, B1 => plus2A(17), B2 
                           => n273, ZN => n341);
   U47 : AOI22_X1 port map( A1 => minus2A(17), A2 => n291, B1 => minusA(17), B2
                           => n285, ZN => n340);
   U48 : NAND2_X1 port map( A1 => n333, A2 => n332, ZN => n488);
   U49 : AOI22_X1 port map( A1 => plusA(13), A2 => n279, B1 => plus2A(13), B2 
                           => n273, ZN => n333);
   U50 : AOI22_X1 port map( A1 => minus2A(13), A2 => n291, B1 => minusA(13), B2
                           => n285, ZN => n332);
   U51 : NAND2_X1 port map( A1 => n381, A2 => n380, ZN => n464);
   U52 : AOI22_X1 port map( A1 => plusA(37), A2 => n281, B1 => plus2A(37), B2 
                           => n275, ZN => n381);
   U53 : AOI22_X1 port map( A1 => minus2A(37), A2 => n293, B1 => minusA(37), B2
                           => n287, ZN => n380);
   U54 : NAND2_X1 port map( A1 => n373, A2 => n372, ZN => n468);
   U55 : AOI22_X1 port map( A1 => plusA(33), A2 => n280, B1 => plus2A(33), B2 
                           => n274, ZN => n373);
   U56 : AOI22_X1 port map( A1 => minus2A(33), A2 => n292, B1 => minusA(33), B2
                           => n286, ZN => n372);
   U57 : NAND2_X1 port map( A1 => n365, A2 => n364, ZN => n472);
   U58 : AOI22_X1 port map( A1 => plusA(29), A2 => n280, B1 => plus2A(29), B2 
                           => n274, ZN => n365);
   U59 : AOI22_X1 port map( A1 => minus2A(29), A2 => n292, B1 => minusA(29), B2
                           => n286, ZN => n364);
   U60 : NAND2_X1 port map( A1 => n357, A2 => n356, ZN => n476);
   U61 : AOI22_X1 port map( A1 => plusA(25), A2 => n280, B1 => plus2A(25), B2 
                           => n274, ZN => n357);
   U62 : AOI22_X1 port map( A1 => minus2A(25), A2 => n292, B1 => minusA(25), B2
                           => n286, ZN => n356);
   U63 : NAND2_X1 port map( A1 => n349, A2 => n348, ZN => n480);
   U64 : AOI22_X1 port map( A1 => plusA(21), A2 => n279, B1 => plus2A(21), B2 
                           => n273, ZN => n349);
   U65 : AOI22_X1 port map( A1 => minus2A(21), A2 => n291, B1 => minusA(21), B2
                           => n285, ZN => n348);
   U66 : NAND2_X1 port map( A1 => n339, A2 => n338, ZN => n485);
   U67 : AOI22_X1 port map( A1 => plusA(16), A2 => n279, B1 => plus2A(16), B2 
                           => n273, ZN => n339);
   U68 : AOI22_X1 port map( A1 => minus2A(16), A2 => n291, B1 => minusA(16), B2
                           => n285, ZN => n338);
   U69 : NAND2_X1 port map( A1 => n331, A2 => n330, ZN => n489);
   U70 : AOI22_X1 port map( A1 => plusA(12), A2 => n279, B1 => plus2A(12), B2 
                           => n273, ZN => n331);
   U71 : AOI22_X1 port map( A1 => minus2A(12), A2 => n291, B1 => minusA(12), B2
                           => n285, ZN => n330);
   U72 : NAND2_X1 port map( A1 => n379, A2 => n378, ZN => n465);
   U73 : AOI22_X1 port map( A1 => plusA(36), A2 => n281, B1 => plus2A(36), B2 
                           => n275, ZN => n379);
   U74 : AOI22_X1 port map( A1 => minus2A(36), A2 => n293, B1 => minusA(36), B2
                           => n287, ZN => n378);
   U75 : NAND2_X1 port map( A1 => n371, A2 => n370, ZN => n469);
   U76 : AOI22_X1 port map( A1 => plusA(32), A2 => n280, B1 => plus2A(32), B2 
                           => n274, ZN => n371);
   U77 : AOI22_X1 port map( A1 => minus2A(32), A2 => n292, B1 => minusA(32), B2
                           => n286, ZN => n370);
   U78 : NAND2_X1 port map( A1 => n363, A2 => n362, ZN => n473);
   U79 : AOI22_X1 port map( A1 => plusA(28), A2 => n280, B1 => plus2A(28), B2 
                           => n274, ZN => n363);
   U80 : AOI22_X1 port map( A1 => minus2A(28), A2 => n292, B1 => minusA(28), B2
                           => n286, ZN => n362);
   U81 : NAND2_X1 port map( A1 => n355, A2 => n354, ZN => n477);
   U82 : AOI22_X1 port map( A1 => plusA(24), A2 => n280, B1 => plus2A(24), B2 
                           => n274, ZN => n355);
   U83 : AOI22_X1 port map( A1 => minus2A(24), A2 => n292, B1 => minusA(24), B2
                           => n286, ZN => n354);
   U84 : NAND2_X1 port map( A1 => n347, A2 => n346, ZN => n481);
   U85 : AOI22_X1 port map( A1 => plusA(20), A2 => n279, B1 => plus2A(20), B2 
                           => n273, ZN => n347);
   U86 : AOI22_X1 port map( A1 => minus2A(20), A2 => n291, B1 => minusA(20), B2
                           => n285, ZN => n346);
   U87 : NAND2_X1 port map( A1 => n343, A2 => n342, ZN => n483);
   U88 : AOI22_X1 port map( A1 => plusA(18), A2 => n279, B1 => plus2A(18), B2 
                           => n273, ZN => n343);
   U89 : AOI22_X1 port map( A1 => minus2A(18), A2 => n291, B1 => minusA(18), B2
                           => n285, ZN => n342);
   U90 : NAND2_X1 port map( A1 => n335, A2 => n334, ZN => n487);
   U91 : AOI22_X1 port map( A1 => plusA(14), A2 => n279, B1 => plus2A(14), B2 
                           => n273, ZN => n335);
   U92 : AOI22_X1 port map( A1 => minus2A(14), A2 => n291, B1 => minusA(14), B2
                           => n285, ZN => n334);
   U93 : NAND2_X1 port map( A1 => n383, A2 => n382, ZN => n463);
   U94 : AOI22_X1 port map( A1 => plusA(38), A2 => n281, B1 => plus2A(38), B2 
                           => n275, ZN => n383);
   U95 : AOI22_X1 port map( A1 => minus2A(38), A2 => n293, B1 => minusA(38), B2
                           => n287, ZN => n382);
   U96 : NAND2_X1 port map( A1 => n375, A2 => n374, ZN => n467);
   U97 : AOI22_X1 port map( A1 => plusA(34), A2 => n280, B1 => plus2A(34), B2 
                           => n274, ZN => n375);
   U98 : AOI22_X1 port map( A1 => minus2A(34), A2 => n292, B1 => minusA(34), B2
                           => n286, ZN => n374);
   U99 : NAND2_X1 port map( A1 => n367, A2 => n366, ZN => n471);
   U100 : AOI22_X1 port map( A1 => plusA(30), A2 => n280, B1 => plus2A(30), B2 
                           => n274, ZN => n367);
   U101 : AOI22_X1 port map( A1 => minus2A(30), A2 => n292, B1 => minusA(30), 
                           B2 => n286, ZN => n366);
   U102 : NAND2_X1 port map( A1 => n359, A2 => n358, ZN => n475);
   U103 : AOI22_X1 port map( A1 => plusA(26), A2 => n280, B1 => plus2A(26), B2 
                           => n274, ZN => n359);
   U104 : AOI22_X1 port map( A1 => minus2A(26), A2 => n292, B1 => minusA(26), 
                           B2 => n286, ZN => n358);
   U105 : NAND2_X1 port map( A1 => n351, A2 => n350, ZN => n479);
   U106 : AOI22_X1 port map( A1 => plusA(22), A2 => n279, B1 => plus2A(22), B2 
                           => n273, ZN => n351);
   U107 : AOI22_X1 port map( A1 => minus2A(22), A2 => n291, B1 => minusA(22), 
                           B2 => n285, ZN => n350);
   U108 : CLKBUF_X1 port map( A => n433, Z => n280);
   U109 : CLKBUF_X1 port map( A => n434, Z => n286);
   U110 : CLKBUF_X1 port map( A => n432, Z => n274);
   U111 : BUF_X1 port map( A => n435, Z => n292);
   U112 : NAND2_X1 port map( A1 => n431, A2 => n430, ZN => n439);
   U113 : AOI22_X1 port map( A1 => plusA(62), A2 => n283, B1 => plus2A(62), B2 
                           => n277, ZN => n431);
   U114 : AOI22_X1 port map( A1 => minus2A(62), A2 => n295, B1 => minusA(62), 
                           B2 => n289, ZN => n430);
   U115 : NAND2_X1 port map( A1 => n429, A2 => n428, ZN => n440);
   U116 : AOI22_X1 port map( A1 => plusA(61), A2 => n283, B1 => plus2A(61), B2 
                           => n277, ZN => n429);
   U117 : AOI22_X1 port map( A1 => minus2A(61), A2 => n295, B1 => minusA(61), 
                           B2 => n289, ZN => n428);
   U118 : NAND2_X1 port map( A1 => n427, A2 => n426, ZN => n441);
   U119 : AOI22_X1 port map( A1 => plusA(60), A2 => n283, B1 => plus2A(60), B2 
                           => n277, ZN => n427);
   U120 : AOI22_X1 port map( A1 => minus2A(60), A2 => n295, B1 => minusA(60), 
                           B2 => n289, ZN => n426);
   U121 : NAND2_X1 port map( A1 => n425, A2 => n424, ZN => n442);
   U122 : AOI22_X1 port map( A1 => plusA(59), A2 => n282, B1 => plus2A(59), B2 
                           => n276, ZN => n425);
   U123 : AOI22_X1 port map( A1 => minus2A(59), A2 => n294, B1 => minusA(59), 
                           B2 => n288, ZN => n424);
   U124 : NAND2_X1 port map( A1 => n421, A2 => n420, ZN => n444);
   U125 : AOI22_X1 port map( A1 => plusA(57), A2 => n282, B1 => plus2A(57), B2 
                           => n276, ZN => n421);
   U126 : AOI22_X1 port map( A1 => minus2A(57), A2 => n294, B1 => minusA(57), 
                           B2 => n288, ZN => n420);
   U127 : NAND2_X1 port map( A1 => n417, A2 => n416, ZN => n446);
   U128 : AOI22_X1 port map( A1 => plusA(55), A2 => n282, B1 => plus2A(55), B2 
                           => n276, ZN => n417);
   U129 : AOI22_X1 port map( A1 => minus2A(55), A2 => n294, B1 => minusA(55), 
                           B2 => n288, ZN => n416);
   U130 : NAND2_X1 port map( A1 => n415, A2 => n414, ZN => n447);
   U131 : AOI22_X1 port map( A1 => plusA(54), A2 => n282, B1 => plus2A(54), B2 
                           => n276, ZN => n415);
   U132 : AOI22_X1 port map( A1 => minus2A(54), A2 => n294, B1 => minusA(54), 
                           B2 => n288, ZN => n414);
   U133 : NAND2_X1 port map( A1 => n413, A2 => n412, ZN => n448);
   U134 : AOI22_X1 port map( A1 => plusA(53), A2 => n282, B1 => plus2A(53), B2 
                           => n276, ZN => n413);
   U135 : AOI22_X1 port map( A1 => minus2A(53), A2 => n294, B1 => minusA(53), 
                           B2 => n288, ZN => n412);
   U136 : NAND2_X1 port map( A1 => n411, A2 => n410, ZN => n449);
   U137 : AOI22_X1 port map( A1 => plusA(52), A2 => n282, B1 => plus2A(52), B2 
                           => n276, ZN => n411);
   U138 : AOI22_X1 port map( A1 => minus2A(52), A2 => n294, B1 => minusA(52), 
                           B2 => n288, ZN => n410);
   U139 : NAND2_X1 port map( A1 => n409, A2 => n408, ZN => n450);
   U140 : AOI22_X1 port map( A1 => plusA(51), A2 => n282, B1 => plus2A(51), B2 
                           => n276, ZN => n409);
   U141 : AOI22_X1 port map( A1 => minus2A(51), A2 => n294, B1 => minusA(51), 
                           B2 => n288, ZN => n408);
   U142 : NAND2_X1 port map( A1 => n407, A2 => n406, ZN => n451);
   U143 : AOI22_X1 port map( A1 => plusA(50), A2 => n282, B1 => plus2A(50), B2 
                           => n276, ZN => n407);
   U144 : AOI22_X1 port map( A1 => minus2A(50), A2 => n294, B1 => minusA(50), 
                           B2 => n288, ZN => n406);
   U145 : NAND2_X1 port map( A1 => n401, A2 => n400, ZN => n454);
   U146 : AOI22_X1 port map( A1 => plusA(47), A2 => n281, B1 => plus2A(47), B2 
                           => n275, ZN => n401);
   U147 : AOI22_X1 port map( A1 => minus2A(47), A2 => n293, B1 => minusA(47), 
                           B2 => n287, ZN => n400);
   U148 : NAND2_X1 port map( A1 => n397, A2 => n396, ZN => n456);
   U149 : AOI22_X1 port map( A1 => plusA(45), A2 => n281, B1 => plus2A(45), B2 
                           => n275, ZN => n397);
   U150 : AOI22_X1 port map( A1 => minus2A(45), A2 => n293, B1 => minusA(45), 
                           B2 => n287, ZN => n396);
   U151 : NAND2_X1 port map( A1 => n393, A2 => n392, ZN => n458);
   U152 : AOI22_X1 port map( A1 => plusA(43), A2 => n281, B1 => plus2A(43), B2 
                           => n275, ZN => n393);
   U153 : AOI22_X1 port map( A1 => minus2A(43), A2 => n293, B1 => minusA(43), 
                           B2 => n287, ZN => n392);
   U154 : NAND2_X1 port map( A1 => n389, A2 => n388, ZN => n460);
   U155 : AOI22_X1 port map( A1 => plusA(41), A2 => n281, B1 => plus2A(41), B2 
                           => n275, ZN => n389);
   U156 : AOI22_X1 port map( A1 => minus2A(41), A2 => n293, B1 => minusA(41), 
                           B2 => n287, ZN => n388);
   U157 : NAND2_X1 port map( A1 => n405, A2 => n404, ZN => n452);
   U158 : AOI22_X1 port map( A1 => plusA(49), A2 => n282, B1 => plus2A(49), B2 
                           => n276, ZN => n405);
   U159 : AOI22_X1 port map( A1 => minus2A(49), A2 => n294, B1 => minusA(49), 
                           B2 => n288, ZN => n404);
   U160 : NAND2_X1 port map( A1 => n419, A2 => n418, ZN => n445);
   U161 : AOI22_X1 port map( A1 => plusA(56), A2 => n282, B1 => plus2A(56), B2 
                           => n276, ZN => n419);
   U162 : AOI22_X1 port map( A1 => minus2A(56), A2 => n294, B1 => minusA(56), 
                           B2 => n288, ZN => n418);
   U163 : NAND2_X1 port map( A1 => n387, A2 => n386, ZN => n461);
   U164 : AOI22_X1 port map( A1 => plusA(40), A2 => n281, B1 => plus2A(40), B2 
                           => n275, ZN => n387);
   U165 : AOI22_X1 port map( A1 => minus2A(40), A2 => n293, B1 => minusA(40), 
                           B2 => n287, ZN => n386);
   U166 : NAND2_X1 port map( A1 => n399, A2 => n398, ZN => n455);
   U167 : AOI22_X1 port map( A1 => plusA(46), A2 => n281, B1 => plus2A(46), B2 
                           => n275, ZN => n399);
   U168 : AOI22_X1 port map( A1 => minus2A(46), A2 => n293, B1 => minusA(46), 
                           B2 => n287, ZN => n398);
   U169 : NAND2_X1 port map( A1 => n395, A2 => n394, ZN => n457);
   U170 : AOI22_X1 port map( A1 => plusA(44), A2 => n281, B1 => plus2A(44), B2 
                           => n275, ZN => n395);
   U171 : AOI22_X1 port map( A1 => minus2A(44), A2 => n293, B1 => minusA(44), 
                           B2 => n287, ZN => n394);
   U172 : NAND2_X1 port map( A1 => n391, A2 => n390, ZN => n459);
   U173 : AOI22_X1 port map( A1 => plusA(42), A2 => n281, B1 => plus2A(42), B2 
                           => n275, ZN => n391);
   U174 : AOI22_X1 port map( A1 => minus2A(42), A2 => n293, B1 => minusA(42), 
                           B2 => n287, ZN => n390);
   U175 : CLKBUF_X1 port map( A => n433, Z => n281);
   U176 : CLKBUF_X1 port map( A => n434, Z => n287);
   U177 : CLKBUF_X1 port map( A => n432, Z => n275);
   U178 : BUF_X1 port map( A => n435, Z => n293);
   U179 : CLKBUF_X1 port map( A => n433, Z => n282);
   U180 : CLKBUF_X1 port map( A => n434, Z => n288);
   U181 : CLKBUF_X1 port map( A => n432, Z => n276);
   U182 : BUF_X1 port map( A => n435, Z => n294);
   U183 : NOR2_X1 port map( A1 => n323, A2 => n304, ZN => n493);
   U184 : INV_X1 port map( A => SEL(2), ZN => n304);
   U185 : AND2_X1 port map( A1 => SEL(2), A2 => n323, ZN => n435);
   U186 : NOR2_X1 port map( A1 => SEL(1), A2 => SEL(0), ZN => n323);
   U187 : INV_X1 port map( A => SEL(1), ZN => n302);
   U188 : INV_X1 port map( A => SEL(0), ZN => n303);
   U189 : NAND2_X1 port map( A1 => n329, A2 => n328, ZN => n490);
   U190 : AOI22_X1 port map( A1 => plusA(11), A2 => n278, B1 => plus2A(11), B2 
                           => n272, ZN => n329);
   U191 : AOI22_X1 port map( A1 => minus2A(11), A2 => n290, B1 => minusA(11), 
                           B2 => n284, ZN => n328);
   U192 : NAND2_X1 port map( A1 => n437, A2 => n436, ZN => n438);
   U193 : AOI22_X1 port map( A1 => plusA(63), A2 => n283, B1 => plus2A(63), B2 
                           => n277, ZN => n437);
   U194 : AOI22_X1 port map( A1 => minus2A(63), A2 => n295, B1 => minusA(63), 
                           B2 => n289, ZN => n436);
   U195 : NAND2_X1 port map( A1 => n327, A2 => n326, ZN => n491);
   U196 : AOI22_X1 port map( A1 => plusA(10), A2 => n278, B1 => plus2A(10), B2 
                           => n272, ZN => n327);
   U197 : AOI22_X1 port map( A1 => minus2A(10), A2 => n290, B1 => minusA(10), 
                           B2 => n284, ZN => n326);
   U198 : NAND2_X1 port map( A1 => n325, A2 => n324, ZN => n492);
   U199 : AOI22_X1 port map( A1 => plusA(9), A2 => n278, B1 => plus2A(9), B2 =>
                           n272, ZN => n325);
   U200 : AOI22_X1 port map( A1 => minus2A(9), A2 => n290, B1 => minusA(9), B2 
                           => n284, ZN => n324);
   U201 : NAND2_X1 port map( A1 => n320, A2 => n319, ZN => n495);
   U202 : AOI22_X1 port map( A1 => plusA(7), A2 => n278, B1 => plus2A(7), B2 =>
                           n272, ZN => n320);
   U203 : AOI22_X1 port map( A1 => minus2A(7), A2 => n290, B1 => minusA(7), B2 
                           => n284, ZN => n319);
   U204 : NAND2_X1 port map( A1 => n318, A2 => n317, ZN => n496);
   U205 : AOI22_X1 port map( A1 => plusA(6), A2 => n278, B1 => plus2A(6), B2 =>
                           n272, ZN => n318);
   U206 : AOI22_X1 port map( A1 => minus2A(6), A2 => n290, B1 => minusA(6), B2 
                           => n284, ZN => n317);
   U207 : NAND2_X1 port map( A1 => n316, A2 => n315, ZN => n497);
   U208 : AOI22_X1 port map( A1 => plusA(5), A2 => n278, B1 => plus2A(5), B2 =>
                           n272, ZN => n316);
   U209 : AOI22_X1 port map( A1 => minus2A(5), A2 => n290, B1 => minusA(5), B2 
                           => n284, ZN => n315);
   U210 : NAND2_X1 port map( A1 => n312, A2 => n311, ZN => n499);
   U211 : AOI22_X1 port map( A1 => plusA(3), A2 => n278, B1 => plus2A(3), B2 =>
                           n272, ZN => n312);
   U212 : AOI22_X1 port map( A1 => minus2A(3), A2 => n290, B1 => minusA(3), B2 
                           => n284, ZN => n311);
   U213 : NAND2_X1 port map( A1 => n322, A2 => n321, ZN => n494);
   U214 : AOI22_X1 port map( A1 => plusA(8), A2 => n278, B1 => plus2A(8), B2 =>
                           n272, ZN => n322);
   U215 : AOI22_X1 port map( A1 => minus2A(8), A2 => n290, B1 => minusA(8), B2 
                           => n284, ZN => n321);
   U216 : NAND2_X1 port map( A1 => n314, A2 => n313, ZN => n498);
   U217 : AOI22_X1 port map( A1 => plusA(4), A2 => n278, B1 => plus2A(4), B2 =>
                           n272, ZN => n314);
   U218 : AOI22_X1 port map( A1 => minus2A(4), A2 => n290, B1 => minusA(4), B2 
                           => n284, ZN => n313);
   U219 : NAND2_X1 port map( A1 => n310, A2 => n309, ZN => n500);
   U220 : AOI22_X1 port map( A1 => plusA(2), A2 => n278, B1 => plus2A(2), B2 =>
                           n272, ZN => n310);
   U221 : AOI22_X1 port map( A1 => minus2A(2), A2 => n290, B1 => minusA(2), B2 
                           => n284, ZN => n309);
   U222 : NAND2_X1 port map( A1 => n308, A2 => n307, ZN => n501);
   U223 : AOI22_X1 port map( A1 => plusA(1), A2 => n278, B1 => plus2A(1), B2 =>
                           n272, ZN => n308);
   U224 : AOI22_X1 port map( A1 => minus2A(1), A2 => n290, B1 => minusA(1), B2 
                           => n284, ZN => n307);
   U225 : NAND2_X1 port map( A1 => n306, A2 => n305, ZN => n502);
   U226 : AOI22_X1 port map( A1 => plusA(0), A2 => n278, B1 => plus2A(0), B2 =>
                           n272, ZN => n306);
   U227 : AOI22_X1 port map( A1 => minus2A(0), A2 => n290, B1 => minusA(0), B2 
                           => n284, ZN => n305);
   U228 : CLKBUF_X1 port map( A => n432, Z => n277);
   U229 : CLKBUF_X1 port map( A => n433, Z => n283);
   U230 : CLKBUF_X1 port map( A => n434, Z => n289);
   U231 : CLKBUF_X1 port map( A => n435, Z => n295);
   U232 : CLKBUF_X1 port map( A => n493, Z => n301);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity MUX_GENERIC_N64_RADIX3_10 is

   port( plusA, minusA, plus2A, minus2A : in std_logic_vector (63 downto 0);  
         SEL : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (63 
         downto 0));

end MUX_GENERIC_N64_RADIX3_10;

architecture SYN_beh of MUX_GENERIC_N64_RADIX3_10 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component TBUF_X4
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   component TBUF_X1
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   signal n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, 
      n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, 
      n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, 
      n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, 
      n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, 
      n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, 
      n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, 
      n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, 
      n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, 
      n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, 
      n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, 
      n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, 
      n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, 
      n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, 
      n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, 
      n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, 
      n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, 
      n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, 
      n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, 
      n499, n500, n501, n502 : std_logic;

begin
   
   Y_tri_60_inst : TBUF_X1 port map( A => n441, EN => n301, Z => Y(60));
   Y_tri_61_inst : TBUF_X1 port map( A => n440, EN => n301, Z => Y(61));
   Y_tri_62_inst : TBUF_X1 port map( A => n439, EN => n301, Z => Y(62));
   Y_tri_63_inst : TBUF_X1 port map( A => n438, EN => n301, Z => Y(63));
   Y_tri_37_inst : TBUF_X1 port map( A => n464, EN => n299, Z => Y(37));
   Y_tri_38_inst : TBUF_X1 port map( A => n463, EN => n299, Z => Y(38));
   Y_tri_39_inst : TBUF_X1 port map( A => n462, EN => n299, Z => Y(39));
   Y_tri_40_inst : TBUF_X1 port map( A => n461, EN => n299, Z => Y(40));
   Y_tri_41_inst : TBUF_X1 port map( A => n460, EN => n299, Z => Y(41));
   Y_tri_42_inst : TBUF_X1 port map( A => n459, EN => n299, Z => Y(42));
   Y_tri_43_inst : TBUF_X1 port map( A => n458, EN => n299, Z => Y(43));
   Y_tri_44_inst : TBUF_X1 port map( A => n457, EN => n299, Z => Y(44));
   Y_tri_45_inst : TBUF_X1 port map( A => n456, EN => n299, Z => Y(45));
   Y_tri_46_inst : TBUF_X1 port map( A => n455, EN => n299, Z => Y(46));
   Y_tri_47_inst : TBUF_X1 port map( A => n454, EN => n299, Z => Y(47));
   Y_tri_48_inst : TBUF_X1 port map( A => n453, EN => n300, Z => Y(48));
   Y_tri_49_inst : TBUF_X1 port map( A => n452, EN => n300, Z => Y(49));
   Y_tri_50_inst : TBUF_X1 port map( A => n451, EN => n300, Z => Y(50));
   Y_tri_51_inst : TBUF_X1 port map( A => n450, EN => n300, Z => Y(51));
   Y_tri_52_inst : TBUF_X1 port map( A => n449, EN => n300, Z => Y(52));
   Y_tri_53_inst : TBUF_X1 port map( A => n448, EN => n300, Z => Y(53));
   Y_tri_54_inst : TBUF_X1 port map( A => n447, EN => n300, Z => Y(54));
   Y_tri_55_inst : TBUF_X1 port map( A => n446, EN => n300, Z => Y(55));
   Y_tri_56_inst : TBUF_X1 port map( A => n445, EN => n300, Z => Y(56));
   Y_tri_58_inst : TBUF_X1 port map( A => n443, EN => n300, Z => Y(58));
   Y_tri_59_inst : TBUF_X1 port map( A => n442, EN => n300, Z => Y(59));
   Y_tri_57_inst : TBUF_X1 port map( A => n444, EN => n300, Z => Y(57));
   Y_tri_15_inst : TBUF_X1 port map( A => n486, EN => n297, Z => Y(15));
   Y_tri_16_inst : TBUF_X1 port map( A => n485, EN => n297, Z => Y(16));
   Y_tri_17_inst : TBUF_X1 port map( A => n484, EN => n297, Z => Y(17));
   Y_tri_18_inst : TBUF_X1 port map( A => n483, EN => n297, Z => Y(18));
   Y_tri_19_inst : TBUF_X1 port map( A => n482, EN => n297, Z => Y(19));
   Y_tri_20_inst : TBUF_X1 port map( A => n481, EN => n297, Z => Y(20));
   Y_tri_21_inst : TBUF_X1 port map( A => n480, EN => n297, Z => Y(21));
   Y_tri_22_inst : TBUF_X1 port map( A => n479, EN => n297, Z => Y(22));
   Y_tri_23_inst : TBUF_X1 port map( A => n478, EN => n297, Z => Y(23));
   Y_tri_24_inst : TBUF_X1 port map( A => n477, EN => n298, Z => Y(24));
   Y_tri_25_inst : TBUF_X1 port map( A => n476, EN => n298, Z => Y(25));
   Y_tri_26_inst : TBUF_X1 port map( A => n475, EN => n298, Z => Y(26));
   Y_tri_27_inst : TBUF_X1 port map( A => n474, EN => n298, Z => Y(27));
   Y_tri_28_inst : TBUF_X1 port map( A => n473, EN => n298, Z => Y(28));
   Y_tri_29_inst : TBUF_X1 port map( A => n472, EN => n298, Z => Y(29));
   Y_tri_30_inst : TBUF_X1 port map( A => n471, EN => n298, Z => Y(30));
   Y_tri_31_inst : TBUF_X1 port map( A => n470, EN => n298, Z => Y(31));
   Y_tri_32_inst : TBUF_X1 port map( A => n469, EN => n298, Z => Y(32));
   Y_tri_33_inst : TBUF_X1 port map( A => n468, EN => n298, Z => Y(33));
   Y_tri_34_inst : TBUF_X1 port map( A => n467, EN => n298, Z => Y(34));
   Y_tri_35_inst : TBUF_X1 port map( A => n466, EN => n298, Z => Y(35));
   Y_tri_36_inst : TBUF_X1 port map( A => n465, EN => n299, Z => Y(36));
   Y_tri_8_inst : TBUF_X1 port map( A => n494, EN => n296, Z => Y(8));
   Y_tri_7_inst : TBUF_X1 port map( A => n495, EN => n296, Z => Y(7));
   Y_tri_6_inst : TBUF_X1 port map( A => n496, EN => n296, Z => Y(6));
   Y_tri_13_inst : TBUF_X1 port map( A => n488, EN => n297, Z => Y(13));
   Y_tri_14_inst : TBUF_X1 port map( A => n487, EN => n297, Z => Y(14));
   Y_tri_12_inst : TBUF_X1 port map( A => n489, EN => n297, Z => Y(12));
   Y_tri_10_inst : TBUF_X1 port map( A => n491, EN => n296, Z => Y(10));
   Y_tri_11_inst : TBUF_X1 port map( A => n490, EN => n296, Z => Y(11));
   Y_tri_5_inst : TBUF_X1 port map( A => n497, EN => n296, Z => Y(5));
   Y_tri_4_inst : TBUF_X1 port map( A => n498, EN => n296, Z => Y(4));
   Y_tri_3_inst : TBUF_X1 port map( A => n499, EN => n296, Z => Y(3));
   Y_tri_2_inst : TBUF_X1 port map( A => n500, EN => n296, Z => Y(2));
   Y_tri_1_inst : TBUF_X1 port map( A => n501, EN => n296, Z => Y(1));
   Y_tri_0_inst : TBUF_X1 port map( A => n502, EN => n296, Z => Y(0));
   Y_tri_9_inst : TBUF_X4 port map( A => n492, EN => n296, Z => Y(9));
   U2 : NOR3_X1 port map( A1 => SEL(0), A2 => SEL(2), A3 => n302, ZN => n434);
   U3 : NOR3_X1 port map( A1 => n302, A2 => SEL(2), A3 => n303, ZN => n432);
   U4 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n303, ZN => n433);
   U5 : CLKBUF_X3 port map( A => n493, Z => n296);
   U6 : CLKBUF_X1 port map( A => n493, Z => n297);
   U7 : CLKBUF_X1 port map( A => n493, Z => n298);
   U8 : CLKBUF_X1 port map( A => n493, Z => n299);
   U9 : CLKBUF_X1 port map( A => n493, Z => n300);
   U10 : NAND2_X1 port map( A1 => n379, A2 => n378, ZN => n465);
   U11 : AOI22_X1 port map( A1 => plusA(36), A2 => n281, B1 => plus2A(36), B2 
                           => n275, ZN => n379);
   U12 : AOI22_X1 port map( A1 => minus2A(36), A2 => n293, B1 => minusA(36), B2
                           => n287, ZN => n378);
   U13 : NAND2_X1 port map( A1 => n371, A2 => n370, ZN => n469);
   U14 : AOI22_X1 port map( A1 => plusA(32), A2 => n280, B1 => plus2A(32), B2 
                           => n274, ZN => n371);
   U15 : AOI22_X1 port map( A1 => minus2A(32), A2 => n292, B1 => minusA(32), B2
                           => n286, ZN => n370);
   U16 : NAND2_X1 port map( A1 => n363, A2 => n362, ZN => n473);
   U17 : AOI22_X1 port map( A1 => plusA(28), A2 => n280, B1 => plus2A(28), B2 
                           => n274, ZN => n363);
   U18 : AOI22_X1 port map( A1 => minus2A(28), A2 => n292, B1 => minusA(28), B2
                           => n286, ZN => n362);
   U19 : NAND2_X1 port map( A1 => n355, A2 => n354, ZN => n477);
   U20 : AOI22_X1 port map( A1 => plusA(24), A2 => n280, B1 => plus2A(24), B2 
                           => n274, ZN => n355);
   U21 : AOI22_X1 port map( A1 => minus2A(24), A2 => n292, B1 => minusA(24), B2
                           => n286, ZN => n354);
   U22 : NAND2_X1 port map( A1 => n347, A2 => n346, ZN => n481);
   U23 : AOI22_X1 port map( A1 => plusA(20), A2 => n279, B1 => plus2A(20), B2 
                           => n273, ZN => n347);
   U24 : AOI22_X1 port map( A1 => minus2A(20), A2 => n291, B1 => minusA(20), B2
                           => n285, ZN => n346);
   U25 : NAND2_X1 port map( A1 => n339, A2 => n338, ZN => n485);
   U26 : AOI22_X1 port map( A1 => plusA(16), A2 => n279, B1 => plus2A(16), B2 
                           => n273, ZN => n339);
   U27 : AOI22_X1 port map( A1 => minus2A(16), A2 => n291, B1 => minusA(16), B2
                           => n285, ZN => n338);
   U28 : NAND2_X1 port map( A1 => n375, A2 => n374, ZN => n467);
   U29 : AOI22_X1 port map( A1 => plusA(34), A2 => n280, B1 => plus2A(34), B2 
                           => n274, ZN => n375);
   U30 : AOI22_X1 port map( A1 => minus2A(34), A2 => n292, B1 => minusA(34), B2
                           => n286, ZN => n374);
   U31 : NAND2_X1 port map( A1 => n367, A2 => n366, ZN => n471);
   U32 : AOI22_X1 port map( A1 => plusA(30), A2 => n280, B1 => plus2A(30), B2 
                           => n274, ZN => n367);
   U33 : AOI22_X1 port map( A1 => minus2A(30), A2 => n292, B1 => minusA(30), B2
                           => n286, ZN => n366);
   U34 : NAND2_X1 port map( A1 => n359, A2 => n358, ZN => n475);
   U35 : AOI22_X1 port map( A1 => plusA(26), A2 => n280, B1 => plus2A(26), B2 
                           => n274, ZN => n359);
   U36 : AOI22_X1 port map( A1 => minus2A(26), A2 => n292, B1 => minusA(26), B2
                           => n286, ZN => n358);
   U37 : NAND2_X1 port map( A1 => n351, A2 => n350, ZN => n479);
   U38 : AOI22_X1 port map( A1 => plusA(22), A2 => n279, B1 => plus2A(22), B2 
                           => n273, ZN => n351);
   U39 : AOI22_X1 port map( A1 => minus2A(22), A2 => n291, B1 => minusA(22), B2
                           => n285, ZN => n350);
   U40 : NAND2_X1 port map( A1 => n343, A2 => n342, ZN => n483);
   U41 : AOI22_X1 port map( A1 => plusA(18), A2 => n279, B1 => plus2A(18), B2 
                           => n273, ZN => n343);
   U42 : AOI22_X1 port map( A1 => minus2A(18), A2 => n291, B1 => minusA(18), B2
                           => n285, ZN => n342);
   U43 : NAND2_X1 port map( A1 => n373, A2 => n372, ZN => n468);
   U44 : AOI22_X1 port map( A1 => plusA(33), A2 => n280, B1 => plus2A(33), B2 
                           => n274, ZN => n373);
   U45 : AOI22_X1 port map( A1 => minus2A(33), A2 => n292, B1 => minusA(33), B2
                           => n286, ZN => n372);
   U46 : NAND2_X1 port map( A1 => n365, A2 => n364, ZN => n472);
   U47 : AOI22_X1 port map( A1 => plusA(29), A2 => n280, B1 => plus2A(29), B2 
                           => n274, ZN => n365);
   U48 : AOI22_X1 port map( A1 => minus2A(29), A2 => n292, B1 => minusA(29), B2
                           => n286, ZN => n364);
   U49 : NAND2_X1 port map( A1 => n357, A2 => n356, ZN => n476);
   U50 : AOI22_X1 port map( A1 => plusA(25), A2 => n280, B1 => plus2A(25), B2 
                           => n274, ZN => n357);
   U51 : AOI22_X1 port map( A1 => minus2A(25), A2 => n292, B1 => minusA(25), B2
                           => n286, ZN => n356);
   U52 : NAND2_X1 port map( A1 => n349, A2 => n348, ZN => n480);
   U53 : AOI22_X1 port map( A1 => plusA(21), A2 => n279, B1 => plus2A(21), B2 
                           => n273, ZN => n349);
   U54 : AOI22_X1 port map( A1 => minus2A(21), A2 => n291, B1 => minusA(21), B2
                           => n285, ZN => n348);
   U55 : NAND2_X1 port map( A1 => n341, A2 => n340, ZN => n484);
   U56 : AOI22_X1 port map( A1 => plusA(17), A2 => n279, B1 => plus2A(17), B2 
                           => n273, ZN => n341);
   U57 : AOI22_X1 port map( A1 => minus2A(17), A2 => n291, B1 => minusA(17), B2
                           => n285, ZN => n340);
   U58 : NAND2_X1 port map( A1 => n377, A2 => n376, ZN => n466);
   U59 : AOI22_X1 port map( A1 => plusA(35), A2 => n280, B1 => plus2A(35), B2 
                           => n274, ZN => n377);
   U60 : AOI22_X1 port map( A1 => minus2A(35), A2 => n292, B1 => minusA(35), B2
                           => n286, ZN => n376);
   U61 : NAND2_X1 port map( A1 => n369, A2 => n368, ZN => n470);
   U62 : AOI22_X1 port map( A1 => plusA(31), A2 => n280, B1 => plus2A(31), B2 
                           => n274, ZN => n369);
   U63 : AOI22_X1 port map( A1 => minus2A(31), A2 => n292, B1 => minusA(31), B2
                           => n286, ZN => n368);
   U64 : NAND2_X1 port map( A1 => n361, A2 => n360, ZN => n474);
   U65 : AOI22_X1 port map( A1 => plusA(27), A2 => n280, B1 => plus2A(27), B2 
                           => n274, ZN => n361);
   U66 : AOI22_X1 port map( A1 => minus2A(27), A2 => n292, B1 => minusA(27), B2
                           => n286, ZN => n360);
   U67 : NAND2_X1 port map( A1 => n353, A2 => n352, ZN => n478);
   U68 : AOI22_X1 port map( A1 => plusA(23), A2 => n279, B1 => plus2A(23), B2 
                           => n273, ZN => n353);
   U69 : AOI22_X1 port map( A1 => minus2A(23), A2 => n291, B1 => minusA(23), B2
                           => n285, ZN => n352);
   U70 : NAND2_X1 port map( A1 => n345, A2 => n344, ZN => n482);
   U71 : AOI22_X1 port map( A1 => plusA(19), A2 => n279, B1 => plus2A(19), B2 
                           => n273, ZN => n345);
   U72 : AOI22_X1 port map( A1 => minus2A(19), A2 => n291, B1 => minusA(19), B2
                           => n285, ZN => n344);
   U73 : NAND2_X1 port map( A1 => n427, A2 => n426, ZN => n441);
   U74 : AOI22_X1 port map( A1 => plusA(60), A2 => n283, B1 => plus2A(60), B2 
                           => n277, ZN => n427);
   U75 : AOI22_X1 port map( A1 => minus2A(60), A2 => n295, B1 => minusA(60), B2
                           => n289, ZN => n426);
   U76 : NAND2_X1 port map( A1 => n425, A2 => n424, ZN => n442);
   U77 : AOI22_X1 port map( A1 => plusA(59), A2 => n282, B1 => plus2A(59), B2 
                           => n276, ZN => n425);
   U78 : AOI22_X1 port map( A1 => minus2A(59), A2 => n294, B1 => minusA(59), B2
                           => n288, ZN => n424);
   U79 : NAND2_X1 port map( A1 => n423, A2 => n422, ZN => n443);
   U80 : AOI22_X1 port map( A1 => plusA(58), A2 => n282, B1 => plus2A(58), B2 
                           => n276, ZN => n423);
   U81 : AOI22_X1 port map( A1 => minus2A(58), A2 => n294, B1 => minusA(58), B2
                           => n288, ZN => n422);
   U82 : NAND2_X1 port map( A1 => n415, A2 => n414, ZN => n447);
   U83 : AOI22_X1 port map( A1 => plusA(54), A2 => n282, B1 => plus2A(54), B2 
                           => n276, ZN => n415);
   U84 : AOI22_X1 port map( A1 => minus2A(54), A2 => n294, B1 => minusA(54), B2
                           => n288, ZN => n414);
   U85 : NAND2_X1 port map( A1 => n413, A2 => n412, ZN => n448);
   U86 : AOI22_X1 port map( A1 => plusA(53), A2 => n282, B1 => plus2A(53), B2 
                           => n276, ZN => n413);
   U87 : AOI22_X1 port map( A1 => minus2A(53), A2 => n294, B1 => minusA(53), B2
                           => n288, ZN => n412);
   U88 : NAND2_X1 port map( A1 => n407, A2 => n406, ZN => n451);
   U89 : AOI22_X1 port map( A1 => plusA(50), A2 => n282, B1 => plus2A(50), B2 
                           => n276, ZN => n407);
   U90 : AOI22_X1 port map( A1 => minus2A(50), A2 => n294, B1 => minusA(50), B2
                           => n288, ZN => n406);
   U91 : NAND2_X1 port map( A1 => n405, A2 => n404, ZN => n452);
   U92 : AOI22_X1 port map( A1 => plusA(49), A2 => n282, B1 => plus2A(49), B2 
                           => n276, ZN => n405);
   U93 : AOI22_X1 port map( A1 => minus2A(49), A2 => n294, B1 => minusA(49), B2
                           => n288, ZN => n404);
   U94 : NAND2_X1 port map( A1 => n403, A2 => n402, ZN => n453);
   U95 : AOI22_X1 port map( A1 => plusA(48), A2 => n282, B1 => plus2A(48), B2 
                           => n276, ZN => n403);
   U96 : AOI22_X1 port map( A1 => minus2A(48), A2 => n294, B1 => minusA(48), B2
                           => n288, ZN => n402);
   U97 : NAND2_X1 port map( A1 => n387, A2 => n386, ZN => n461);
   U98 : AOI22_X1 port map( A1 => plusA(40), A2 => n281, B1 => plus2A(40), B2 
                           => n275, ZN => n387);
   U99 : AOI22_X1 port map( A1 => minus2A(40), A2 => n293, B1 => minusA(40), B2
                           => n287, ZN => n386);
   U100 : NAND2_X1 port map( A1 => n391, A2 => n390, ZN => n459);
   U101 : AOI22_X1 port map( A1 => plusA(42), A2 => n281, B1 => plus2A(42), B2 
                           => n275, ZN => n391);
   U102 : AOI22_X1 port map( A1 => minus2A(42), A2 => n293, B1 => minusA(42), 
                           B2 => n287, ZN => n390);
   U103 : NAND2_X1 port map( A1 => n383, A2 => n382, ZN => n463);
   U104 : AOI22_X1 port map( A1 => plusA(38), A2 => n281, B1 => plus2A(38), B2 
                           => n275, ZN => n383);
   U105 : AOI22_X1 port map( A1 => minus2A(38), A2 => n293, B1 => minusA(38), 
                           B2 => n287, ZN => n382);
   U106 : NAND2_X1 port map( A1 => n393, A2 => n392, ZN => n458);
   U107 : AOI22_X1 port map( A1 => plusA(43), A2 => n281, B1 => plus2A(43), B2 
                           => n275, ZN => n393);
   U108 : AOI22_X1 port map( A1 => minus2A(43), A2 => n293, B1 => minusA(43), 
                           B2 => n287, ZN => n392);
   U109 : NAND2_X1 port map( A1 => n389, A2 => n388, ZN => n460);
   U110 : AOI22_X1 port map( A1 => plusA(41), A2 => n281, B1 => plus2A(41), B2 
                           => n275, ZN => n389);
   U111 : AOI22_X1 port map( A1 => minus2A(41), A2 => n293, B1 => minusA(41), 
                           B2 => n287, ZN => n388);
   U112 : NAND2_X1 port map( A1 => n381, A2 => n380, ZN => n464);
   U113 : AOI22_X1 port map( A1 => plusA(37), A2 => n281, B1 => plus2A(37), B2 
                           => n275, ZN => n381);
   U114 : AOI22_X1 port map( A1 => minus2A(37), A2 => n293, B1 => minusA(37), 
                           B2 => n287, ZN => n380);
   U115 : NAND2_X1 port map( A1 => n385, A2 => n384, ZN => n462);
   U116 : AOI22_X1 port map( A1 => plusA(39), A2 => n281, B1 => plus2A(39), B2 
                           => n275, ZN => n385);
   U117 : AOI22_X1 port map( A1 => minus2A(39), A2 => n293, B1 => minusA(39), 
                           B2 => n287, ZN => n384);
   U118 : NAND2_X1 port map( A1 => n395, A2 => n394, ZN => n457);
   U119 : AOI22_X1 port map( A1 => plusA(44), A2 => n281, B1 => plus2A(44), B2 
                           => n275, ZN => n395);
   U120 : AOI22_X1 port map( A1 => minus2A(44), A2 => n293, B1 => minusA(44), 
                           B2 => n287, ZN => n394);
   U121 : BUF_X1 port map( A => n433, Z => n279);
   U122 : BUF_X1 port map( A => n434, Z => n285);
   U123 : BUF_X1 port map( A => n432, Z => n273);
   U124 : BUF_X1 port map( A => n435, Z => n291);
   U125 : NAND2_X1 port map( A1 => n335, A2 => n334, ZN => n487);
   U126 : AOI22_X1 port map( A1 => plusA(14), A2 => n279, B1 => plus2A(14), B2 
                           => n273, ZN => n335);
   U127 : AOI22_X1 port map( A1 => minus2A(14), A2 => n291, B1 => minusA(14), 
                           B2 => n285, ZN => n334);
   U128 : NAND2_X1 port map( A1 => n337, A2 => n336, ZN => n486);
   U129 : AOI22_X1 port map( A1 => plusA(15), A2 => n279, B1 => plus2A(15), B2 
                           => n273, ZN => n337);
   U130 : AOI22_X1 port map( A1 => minus2A(15), A2 => n291, B1 => minusA(15), 
                           B2 => n285, ZN => n336);
   U131 : BUF_X1 port map( A => n433, Z => n280);
   U132 : BUF_X1 port map( A => n434, Z => n286);
   U133 : BUF_X1 port map( A => n432, Z => n274);
   U134 : BUF_X1 port map( A => n435, Z => n292);
   U135 : NAND2_X1 port map( A1 => n437, A2 => n436, ZN => n438);
   U136 : AOI22_X1 port map( A1 => plusA(63), A2 => n283, B1 => plus2A(63), B2 
                           => n277, ZN => n437);
   U137 : AOI22_X1 port map( A1 => minus2A(63), A2 => n295, B1 => minusA(63), 
                           B2 => n289, ZN => n436);
   U138 : NAND2_X1 port map( A1 => n431, A2 => n430, ZN => n439);
   U139 : AOI22_X1 port map( A1 => plusA(62), A2 => n283, B1 => plus2A(62), B2 
                           => n277, ZN => n431);
   U140 : AOI22_X1 port map( A1 => minus2A(62), A2 => n295, B1 => minusA(62), 
                           B2 => n289, ZN => n430);
   U141 : NAND2_X1 port map( A1 => n429, A2 => n428, ZN => n440);
   U142 : AOI22_X1 port map( A1 => plusA(61), A2 => n283, B1 => plus2A(61), B2 
                           => n277, ZN => n429);
   U143 : AOI22_X1 port map( A1 => minus2A(61), A2 => n295, B1 => minusA(61), 
                           B2 => n289, ZN => n428);
   U144 : NAND2_X1 port map( A1 => n421, A2 => n420, ZN => n444);
   U145 : AOI22_X1 port map( A1 => plusA(57), A2 => n282, B1 => plus2A(57), B2 
                           => n276, ZN => n421);
   U146 : AOI22_X1 port map( A1 => minus2A(57), A2 => n294, B1 => minusA(57), 
                           B2 => n288, ZN => n420);
   U147 : NAND2_X1 port map( A1 => n417, A2 => n416, ZN => n446);
   U148 : AOI22_X1 port map( A1 => plusA(55), A2 => n282, B1 => plus2A(55), B2 
                           => n276, ZN => n417);
   U149 : AOI22_X1 port map( A1 => minus2A(55), A2 => n294, B1 => minusA(55), 
                           B2 => n288, ZN => n416);
   U150 : NAND2_X1 port map( A1 => n411, A2 => n410, ZN => n449);
   U151 : AOI22_X1 port map( A1 => plusA(52), A2 => n282, B1 => plus2A(52), B2 
                           => n276, ZN => n411);
   U152 : AOI22_X1 port map( A1 => minus2A(52), A2 => n294, B1 => minusA(52), 
                           B2 => n288, ZN => n410);
   U153 : NAND2_X1 port map( A1 => n409, A2 => n408, ZN => n450);
   U154 : AOI22_X1 port map( A1 => plusA(51), A2 => n282, B1 => plus2A(51), B2 
                           => n276, ZN => n409);
   U155 : AOI22_X1 port map( A1 => minus2A(51), A2 => n294, B1 => minusA(51), 
                           B2 => n288, ZN => n408);
   U156 : NAND2_X1 port map( A1 => n401, A2 => n400, ZN => n454);
   U157 : AOI22_X1 port map( A1 => plusA(47), A2 => n281, B1 => plus2A(47), B2 
                           => n275, ZN => n401);
   U158 : AOI22_X1 port map( A1 => minus2A(47), A2 => n293, B1 => minusA(47), 
                           B2 => n287, ZN => n400);
   U159 : NAND2_X1 port map( A1 => n397, A2 => n396, ZN => n456);
   U160 : AOI22_X1 port map( A1 => plusA(45), A2 => n281, B1 => plus2A(45), B2 
                           => n275, ZN => n397);
   U161 : AOI22_X1 port map( A1 => minus2A(45), A2 => n293, B1 => minusA(45), 
                           B2 => n287, ZN => n396);
   U162 : NAND2_X1 port map( A1 => n419, A2 => n418, ZN => n445);
   U163 : AOI22_X1 port map( A1 => plusA(56), A2 => n282, B1 => plus2A(56), B2 
                           => n276, ZN => n419);
   U164 : AOI22_X1 port map( A1 => minus2A(56), A2 => n294, B1 => minusA(56), 
                           B2 => n288, ZN => n418);
   U165 : NAND2_X1 port map( A1 => n399, A2 => n398, ZN => n455);
   U166 : AOI22_X1 port map( A1 => plusA(46), A2 => n281, B1 => plus2A(46), B2 
                           => n275, ZN => n399);
   U167 : AOI22_X1 port map( A1 => minus2A(46), A2 => n293, B1 => minusA(46), 
                           B2 => n287, ZN => n398);
   U168 : BUF_X1 port map( A => n433, Z => n281);
   U169 : BUF_X1 port map( A => n434, Z => n287);
   U170 : BUF_X1 port map( A => n432, Z => n275);
   U171 : BUF_X1 port map( A => n435, Z => n293);
   U172 : BUF_X1 port map( A => n433, Z => n282);
   U173 : BUF_X1 port map( A => n434, Z => n288);
   U174 : BUF_X1 port map( A => n432, Z => n276);
   U175 : BUF_X1 port map( A => n435, Z => n294);
   U176 : BUF_X1 port map( A => n433, Z => n278);
   U177 : BUF_X1 port map( A => n434, Z => n284);
   U178 : BUF_X1 port map( A => n432, Z => n272);
   U179 : BUF_X1 port map( A => n435, Z => n290);
   U180 : NOR2_X1 port map( A1 => n323, A2 => n304, ZN => n493);
   U181 : INV_X1 port map( A => SEL(2), ZN => n304);
   U182 : AND2_X1 port map( A1 => SEL(2), A2 => n323, ZN => n435);
   U183 : NOR2_X1 port map( A1 => SEL(1), A2 => SEL(0), ZN => n323);
   U184 : INV_X1 port map( A => SEL(1), ZN => n302);
   U185 : INV_X1 port map( A => SEL(0), ZN => n303);
   U186 : NAND2_X1 port map( A1 => n333, A2 => n332, ZN => n488);
   U187 : AOI22_X1 port map( A1 => plusA(13), A2 => n279, B1 => plus2A(13), B2 
                           => n273, ZN => n333);
   U188 : AOI22_X1 port map( A1 => minus2A(13), A2 => n291, B1 => minusA(13), 
                           B2 => n285, ZN => n332);
   U189 : NAND2_X1 port map( A1 => n331, A2 => n330, ZN => n489);
   U190 : AOI22_X1 port map( A1 => plusA(12), A2 => n279, B1 => plus2A(12), B2 
                           => n273, ZN => n331);
   U191 : AOI22_X1 port map( A1 => minus2A(12), A2 => n291, B1 => minusA(12), 
                           B2 => n285, ZN => n330);
   U192 : NAND2_X1 port map( A1 => n329, A2 => n328, ZN => n490);
   U193 : AOI22_X1 port map( A1 => plusA(11), A2 => n278, B1 => plus2A(11), B2 
                           => n272, ZN => n329);
   U194 : AOI22_X1 port map( A1 => minus2A(11), A2 => n290, B1 => minusA(11), 
                           B2 => n284, ZN => n328);
   U195 : NAND2_X1 port map( A1 => n327, A2 => n326, ZN => n491);
   U196 : AOI22_X1 port map( A1 => plusA(10), A2 => n278, B1 => plus2A(10), B2 
                           => n272, ZN => n327);
   U197 : AOI22_X1 port map( A1 => minus2A(10), A2 => n290, B1 => minusA(10), 
                           B2 => n284, ZN => n326);
   U198 : NAND2_X1 port map( A1 => n325, A2 => n324, ZN => n492);
   U199 : AOI22_X1 port map( A1 => plusA(9), A2 => n278, B1 => plus2A(9), B2 =>
                           n272, ZN => n325);
   U200 : AOI22_X1 port map( A1 => minus2A(9), A2 => n290, B1 => minusA(9), B2 
                           => n284, ZN => n324);
   U201 : NAND2_X1 port map( A1 => n320, A2 => n319, ZN => n495);
   U202 : AOI22_X1 port map( A1 => plusA(7), A2 => n278, B1 => plus2A(7), B2 =>
                           n272, ZN => n320);
   U203 : AOI22_X1 port map( A1 => minus2A(7), A2 => n290, B1 => minusA(7), B2 
                           => n284, ZN => n319);
   U204 : NAND2_X1 port map( A1 => n318, A2 => n317, ZN => n496);
   U205 : AOI22_X1 port map( A1 => plusA(6), A2 => n278, B1 => plus2A(6), B2 =>
                           n272, ZN => n318);
   U206 : AOI22_X1 port map( A1 => minus2A(6), A2 => n290, B1 => minusA(6), B2 
                           => n284, ZN => n317);
   U207 : NAND2_X1 port map( A1 => n316, A2 => n315, ZN => n497);
   U208 : AOI22_X1 port map( A1 => plusA(5), A2 => n278, B1 => plus2A(5), B2 =>
                           n272, ZN => n316);
   U209 : AOI22_X1 port map( A1 => minus2A(5), A2 => n290, B1 => minusA(5), B2 
                           => n284, ZN => n315);
   U210 : NAND2_X1 port map( A1 => n312, A2 => n311, ZN => n499);
   U211 : AOI22_X1 port map( A1 => plusA(3), A2 => n278, B1 => plus2A(3), B2 =>
                           n272, ZN => n312);
   U212 : AOI22_X1 port map( A1 => minus2A(3), A2 => n290, B1 => minusA(3), B2 
                           => n284, ZN => n311);
   U213 : NAND2_X1 port map( A1 => n322, A2 => n321, ZN => n494);
   U214 : AOI22_X1 port map( A1 => plusA(8), A2 => n278, B1 => plus2A(8), B2 =>
                           n272, ZN => n322);
   U215 : AOI22_X1 port map( A1 => minus2A(8), A2 => n290, B1 => minusA(8), B2 
                           => n284, ZN => n321);
   U216 : NAND2_X1 port map( A1 => n314, A2 => n313, ZN => n498);
   U217 : AOI22_X1 port map( A1 => plusA(4), A2 => n278, B1 => plus2A(4), B2 =>
                           n272, ZN => n314);
   U218 : AOI22_X1 port map( A1 => minus2A(4), A2 => n290, B1 => minusA(4), B2 
                           => n284, ZN => n313);
   U219 : NAND2_X1 port map( A1 => n310, A2 => n309, ZN => n500);
   U220 : AOI22_X1 port map( A1 => plusA(2), A2 => n278, B1 => plus2A(2), B2 =>
                           n272, ZN => n310);
   U221 : AOI22_X1 port map( A1 => minus2A(2), A2 => n290, B1 => minusA(2), B2 
                           => n284, ZN => n309);
   U222 : NAND2_X1 port map( A1 => n308, A2 => n307, ZN => n501);
   U223 : AOI22_X1 port map( A1 => plusA(1), A2 => n278, B1 => plus2A(1), B2 =>
                           n272, ZN => n308);
   U224 : AOI22_X1 port map( A1 => minus2A(1), A2 => n290, B1 => minusA(1), B2 
                           => n284, ZN => n307);
   U225 : NAND2_X1 port map( A1 => n306, A2 => n305, ZN => n502);
   U226 : AOI22_X1 port map( A1 => plusA(0), A2 => n278, B1 => plus2A(0), B2 =>
                           n272, ZN => n306);
   U227 : AOI22_X1 port map( A1 => minus2A(0), A2 => n290, B1 => minusA(0), B2 
                           => n284, ZN => n305);
   U228 : CLKBUF_X1 port map( A => n432, Z => n277);
   U229 : CLKBUF_X1 port map( A => n433, Z => n283);
   U230 : CLKBUF_X1 port map( A => n434, Z => n289);
   U231 : CLKBUF_X1 port map( A => n435, Z => n295);
   U232 : CLKBUF_X1 port map( A => n493, Z => n301);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity MUX_GENERIC_N64_RADIX3_9 is

   port( plusA, minusA, plus2A, minus2A : in std_logic_vector (63 downto 0);  
         SEL : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (63 
         downto 0));

end MUX_GENERIC_N64_RADIX3_9;

architecture SYN_beh of MUX_GENERIC_N64_RADIX3_9 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component TBUF_X1
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   component TBUF_X4
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   signal n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, 
      n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, 
      n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, 
      n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, 
      n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, 
      n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, 
      n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, 
      n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, 
      n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, 
      n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, 
      n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, 
      n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, 
      n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, 
      n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, 
      n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, 
      n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, 
      n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, 
      n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, 
      n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, 
      n499, n500, n501, n502 : std_logic;

begin
   
   Y_tri_60_inst : TBUF_X1 port map( A => n441, EN => n301, Z => Y(60));
   Y_tri_61_inst : TBUF_X1 port map( A => n440, EN => n301, Z => Y(61));
   Y_tri_62_inst : TBUF_X1 port map( A => n439, EN => n301, Z => Y(62));
   Y_tri_63_inst : TBUF_X1 port map( A => n438, EN => n301, Z => Y(63));
   Y_tri_57_inst : TBUF_X1 port map( A => n444, EN => n300, Z => Y(57));
   Y_tri_58_inst : TBUF_X1 port map( A => n443, EN => n300, Z => Y(58));
   Y_tri_59_inst : TBUF_X1 port map( A => n442, EN => n300, Z => Y(59));
   Y_tri_56_inst : TBUF_X1 port map( A => n445, EN => n300, Z => Y(56));
   Y_tri_30_inst : TBUF_X1 port map( A => n471, EN => n298, Z => Y(30));
   Y_tri_31_inst : TBUF_X1 port map( A => n470, EN => n298, Z => Y(31));
   Y_tri_32_inst : TBUF_X1 port map( A => n469, EN => n298, Z => Y(32));
   Y_tri_33_inst : TBUF_X1 port map( A => n468, EN => n298, Z => Y(33));
   Y_tri_35_inst : TBUF_X1 port map( A => n466, EN => n298, Z => Y(35));
   Y_tri_36_inst : TBUF_X1 port map( A => n465, EN => n299, Z => Y(36));
   Y_tri_37_inst : TBUF_X1 port map( A => n464, EN => n299, Z => Y(37));
   Y_tri_38_inst : TBUF_X1 port map( A => n463, EN => n299, Z => Y(38));
   Y_tri_39_inst : TBUF_X1 port map( A => n462, EN => n299, Z => Y(39));
   Y_tri_40_inst : TBUF_X1 port map( A => n461, EN => n299, Z => Y(40));
   Y_tri_41_inst : TBUF_X1 port map( A => n460, EN => n299, Z => Y(41));
   Y_tri_42_inst : TBUF_X1 port map( A => n459, EN => n299, Z => Y(42));
   Y_tri_43_inst : TBUF_X1 port map( A => n458, EN => n299, Z => Y(43));
   Y_tri_44_inst : TBUF_X1 port map( A => n457, EN => n299, Z => Y(44));
   Y_tri_45_inst : TBUF_X1 port map( A => n456, EN => n299, Z => Y(45));
   Y_tri_46_inst : TBUF_X1 port map( A => n455, EN => n299, Z => Y(46));
   Y_tri_47_inst : TBUF_X1 port map( A => n454, EN => n299, Z => Y(47));
   Y_tri_48_inst : TBUF_X1 port map( A => n453, EN => n300, Z => Y(48));
   Y_tri_49_inst : TBUF_X1 port map( A => n452, EN => n300, Z => Y(49));
   Y_tri_52_inst : TBUF_X1 port map( A => n449, EN => n300, Z => Y(52));
   Y_tri_53_inst : TBUF_X1 port map( A => n448, EN => n300, Z => Y(53));
   Y_tri_54_inst : TBUF_X1 port map( A => n447, EN => n300, Z => Y(54));
   Y_tri_55_inst : TBUF_X1 port map( A => n446, EN => n300, Z => Y(55));
   Y_tri_34_inst : TBUF_X1 port map( A => n467, EN => n298, Z => Y(34));
   Y_tri_51_inst : TBUF_X1 port map( A => n450, EN => n300, Z => Y(51));
   Y_tri_11_inst : TBUF_X1 port map( A => n490, EN => n296, Z => Y(11));
   Y_tri_12_inst : TBUF_X1 port map( A => n489, EN => n297, Z => Y(12));
   Y_tri_13_inst : TBUF_X1 port map( A => n488, EN => n297, Z => Y(13));
   Y_tri_14_inst : TBUF_X1 port map( A => n487, EN => n297, Z => Y(14));
   Y_tri_15_inst : TBUF_X1 port map( A => n486, EN => n297, Z => Y(15));
   Y_tri_16_inst : TBUF_X1 port map( A => n485, EN => n297, Z => Y(16));
   Y_tri_17_inst : TBUF_X1 port map( A => n484, EN => n297, Z => Y(17));
   Y_tri_18_inst : TBUF_X1 port map( A => n483, EN => n297, Z => Y(18));
   Y_tri_19_inst : TBUF_X1 port map( A => n482, EN => n297, Z => Y(19));
   Y_tri_20_inst : TBUF_X1 port map( A => n481, EN => n297, Z => Y(20));
   Y_tri_21_inst : TBUF_X1 port map( A => n480, EN => n297, Z => Y(21));
   Y_tri_22_inst : TBUF_X1 port map( A => n479, EN => n297, Z => Y(22));
   Y_tri_23_inst : TBUF_X1 port map( A => n478, EN => n297, Z => Y(23));
   Y_tri_24_inst : TBUF_X1 port map( A => n477, EN => n298, Z => Y(24));
   Y_tri_25_inst : TBUF_X1 port map( A => n476, EN => n298, Z => Y(25));
   Y_tri_26_inst : TBUF_X1 port map( A => n475, EN => n298, Z => Y(26));
   Y_tri_27_inst : TBUF_X1 port map( A => n474, EN => n298, Z => Y(27));
   Y_tri_28_inst : TBUF_X1 port map( A => n473, EN => n298, Z => Y(28));
   Y_tri_29_inst : TBUF_X1 port map( A => n472, EN => n298, Z => Y(29));
   Y_tri_7_inst : TBUF_X1 port map( A => n495, EN => n296, Z => Y(7));
   Y_tri_6_inst : TBUF_X1 port map( A => n496, EN => n296, Z => Y(6));
   Y_tri_5_inst : TBUF_X1 port map( A => n497, EN => n296, Z => Y(5));
   Y_tri_8_inst : TBUF_X1 port map( A => n494, EN => n296, Z => Y(8));
   Y_tri_9_inst : TBUF_X1 port map( A => n492, EN => n296, Z => Y(9));
   Y_tri_4_inst : TBUF_X1 port map( A => n498, EN => n296, Z => Y(4));
   Y_tri_3_inst : TBUF_X1 port map( A => n499, EN => n296, Z => Y(3));
   Y_tri_2_inst : TBUF_X1 port map( A => n500, EN => n296, Z => Y(2));
   Y_tri_1_inst : TBUF_X1 port map( A => n501, EN => n296, Z => Y(1));
   Y_tri_0_inst : TBUF_X1 port map( A => n502, EN => n296, Z => Y(0));
   Y_tri_10_inst : TBUF_X4 port map( A => n491, EN => n296, Z => Y(10));
   Y_tri_50_inst : TBUF_X1 port map( A => n451, EN => n300, Z => Y(50));
   U2 : NOR3_X1 port map( A1 => SEL(0), A2 => SEL(2), A3 => n302, ZN => n434);
   U3 : NOR3_X1 port map( A1 => n302, A2 => SEL(2), A3 => n303, ZN => n432);
   U4 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n303, ZN => n433);
   U5 : CLKBUF_X3 port map( A => n493, Z => n296);
   U6 : CLKBUF_X1 port map( A => n493, Z => n297);
   U7 : CLKBUF_X1 port map( A => n493, Z => n298);
   U8 : CLKBUF_X1 port map( A => n493, Z => n299);
   U9 : CLKBUF_X1 port map( A => n493, Z => n300);
   U10 : NAND2_X1 port map( A1 => n359, A2 => n358, ZN => n475);
   U11 : AOI22_X1 port map( A1 => plusA(26), A2 => n280, B1 => plus2A(26), B2 
                           => n274, ZN => n359);
   U12 : AOI22_X1 port map( A1 => minus2A(26), A2 => n292, B1 => minusA(26), B2
                           => n286, ZN => n358);
   U13 : NAND2_X1 port map( A1 => n351, A2 => n350, ZN => n479);
   U14 : AOI22_X1 port map( A1 => plusA(22), A2 => n279, B1 => plus2A(22), B2 
                           => n273, ZN => n351);
   U15 : AOI22_X1 port map( A1 => minus2A(22), A2 => n291, B1 => minusA(22), B2
                           => n285, ZN => n350);
   U16 : NAND2_X1 port map( A1 => n343, A2 => n342, ZN => n483);
   U17 : AOI22_X1 port map( A1 => plusA(18), A2 => n279, B1 => plus2A(18), B2 
                           => n273, ZN => n343);
   U18 : AOI22_X1 port map( A1 => minus2A(18), A2 => n291, B1 => minusA(18), B2
                           => n285, ZN => n342);
   U19 : NAND2_X1 port map( A1 => n363, A2 => n362, ZN => n473);
   U20 : AOI22_X1 port map( A1 => plusA(28), A2 => n280, B1 => plus2A(28), B2 
                           => n274, ZN => n363);
   U21 : AOI22_X1 port map( A1 => minus2A(28), A2 => n292, B1 => minusA(28), B2
                           => n286, ZN => n362);
   U22 : NAND2_X1 port map( A1 => n355, A2 => n354, ZN => n477);
   U23 : AOI22_X1 port map( A1 => plusA(24), A2 => n280, B1 => plus2A(24), B2 
                           => n274, ZN => n355);
   U24 : AOI22_X1 port map( A1 => minus2A(24), A2 => n292, B1 => minusA(24), B2
                           => n286, ZN => n354);
   U25 : NAND2_X1 port map( A1 => n347, A2 => n346, ZN => n481);
   U26 : AOI22_X1 port map( A1 => plusA(20), A2 => n279, B1 => plus2A(20), B2 
                           => n273, ZN => n347);
   U27 : AOI22_X1 port map( A1 => minus2A(20), A2 => n291, B1 => minusA(20), B2
                           => n285, ZN => n346);
   U28 : NAND2_X1 port map( A1 => n361, A2 => n360, ZN => n474);
   U29 : AOI22_X1 port map( A1 => plusA(27), A2 => n280, B1 => plus2A(27), B2 
                           => n274, ZN => n361);
   U30 : AOI22_X1 port map( A1 => minus2A(27), A2 => n292, B1 => minusA(27), B2
                           => n286, ZN => n360);
   U31 : NAND2_X1 port map( A1 => n353, A2 => n352, ZN => n478);
   U32 : AOI22_X1 port map( A1 => plusA(23), A2 => n279, B1 => plus2A(23), B2 
                           => n273, ZN => n353);
   U33 : AOI22_X1 port map( A1 => minus2A(23), A2 => n291, B1 => minusA(23), B2
                           => n285, ZN => n352);
   U34 : NAND2_X1 port map( A1 => n345, A2 => n344, ZN => n482);
   U35 : AOI22_X1 port map( A1 => plusA(19), A2 => n279, B1 => plus2A(19), B2 
                           => n273, ZN => n345);
   U36 : AOI22_X1 port map( A1 => minus2A(19), A2 => n291, B1 => minusA(19), B2
                           => n285, ZN => n344);
   U37 : NAND2_X1 port map( A1 => n365, A2 => n364, ZN => n472);
   U38 : AOI22_X1 port map( A1 => plusA(29), A2 => n280, B1 => plus2A(29), B2 
                           => n274, ZN => n365);
   U39 : AOI22_X1 port map( A1 => minus2A(29), A2 => n292, B1 => minusA(29), B2
                           => n286, ZN => n364);
   U40 : NAND2_X1 port map( A1 => n357, A2 => n356, ZN => n476);
   U41 : AOI22_X1 port map( A1 => plusA(25), A2 => n280, B1 => plus2A(25), B2 
                           => n274, ZN => n357);
   U42 : AOI22_X1 port map( A1 => minus2A(25), A2 => n292, B1 => minusA(25), B2
                           => n286, ZN => n356);
   U43 : NAND2_X1 port map( A1 => n349, A2 => n348, ZN => n480);
   U44 : AOI22_X1 port map( A1 => plusA(21), A2 => n279, B1 => plus2A(21), B2 
                           => n273, ZN => n349);
   U45 : AOI22_X1 port map( A1 => minus2A(21), A2 => n291, B1 => minusA(21), B2
                           => n285, ZN => n348);
   U46 : NAND2_X1 port map( A1 => n417, A2 => n416, ZN => n446);
   U47 : AOI22_X1 port map( A1 => plusA(55), A2 => n282, B1 => plus2A(55), B2 
                           => n276, ZN => n417);
   U48 : AOI22_X1 port map( A1 => minus2A(55), A2 => n294, B1 => minusA(55), B2
                           => n288, ZN => n416);
   U49 : NAND2_X1 port map( A1 => n415, A2 => n414, ZN => n447);
   U50 : AOI22_X1 port map( A1 => plusA(54), A2 => n282, B1 => plus2A(54), B2 
                           => n276, ZN => n415);
   U51 : AOI22_X1 port map( A1 => minus2A(54), A2 => n294, B1 => minusA(54), B2
                           => n288, ZN => n414);
   U52 : NAND2_X1 port map( A1 => n413, A2 => n412, ZN => n448);
   U53 : AOI22_X1 port map( A1 => plusA(53), A2 => n282, B1 => plus2A(53), B2 
                           => n276, ZN => n413);
   U54 : AOI22_X1 port map( A1 => minus2A(53), A2 => n294, B1 => minusA(53), B2
                           => n288, ZN => n412);
   U55 : NAND2_X1 port map( A1 => n411, A2 => n410, ZN => n449);
   U56 : AOI22_X1 port map( A1 => plusA(52), A2 => n282, B1 => plus2A(52), B2 
                           => n276, ZN => n411);
   U57 : AOI22_X1 port map( A1 => minus2A(52), A2 => n294, B1 => minusA(52), B2
                           => n288, ZN => n410);
   U58 : NAND2_X1 port map( A1 => n409, A2 => n408, ZN => n450);
   U59 : AOI22_X1 port map( A1 => plusA(51), A2 => n282, B1 => plus2A(51), B2 
                           => n276, ZN => n409);
   U60 : AOI22_X1 port map( A1 => minus2A(51), A2 => n294, B1 => minusA(51), B2
                           => n288, ZN => n408);
   U61 : NAND2_X1 port map( A1 => n407, A2 => n406, ZN => n451);
   U62 : AOI22_X1 port map( A1 => plusA(50), A2 => n282, B1 => plus2A(50), B2 
                           => n276, ZN => n407);
   U63 : AOI22_X1 port map( A1 => minus2A(50), A2 => n294, B1 => minusA(50), B2
                           => n288, ZN => n406);
   U64 : NAND2_X1 port map( A1 => n405, A2 => n404, ZN => n452);
   U65 : AOI22_X1 port map( A1 => plusA(49), A2 => n282, B1 => plus2A(49), B2 
                           => n276, ZN => n405);
   U66 : AOI22_X1 port map( A1 => minus2A(49), A2 => n294, B1 => minusA(49), B2
                           => n288, ZN => n404);
   U67 : NAND2_X1 port map( A1 => n403, A2 => n402, ZN => n453);
   U68 : AOI22_X1 port map( A1 => plusA(48), A2 => n282, B1 => plus2A(48), B2 
                           => n276, ZN => n403);
   U69 : AOI22_X1 port map( A1 => minus2A(48), A2 => n294, B1 => minusA(48), B2
                           => n288, ZN => n402);
   U70 : NAND2_X1 port map( A1 => n401, A2 => n400, ZN => n454);
   U71 : AOI22_X1 port map( A1 => plusA(47), A2 => n281, B1 => plus2A(47), B2 
                           => n275, ZN => n401);
   U72 : AOI22_X1 port map( A1 => minus2A(47), A2 => n293, B1 => minusA(47), B2
                           => n287, ZN => n400);
   U73 : NAND2_X1 port map( A1 => n391, A2 => n390, ZN => n459);
   U74 : AOI22_X1 port map( A1 => plusA(42), A2 => n281, B1 => plus2A(42), B2 
                           => n275, ZN => n391);
   U75 : AOI22_X1 port map( A1 => minus2A(42), A2 => n293, B1 => minusA(42), B2
                           => n287, ZN => n390);
   U76 : NAND2_X1 port map( A1 => n383, A2 => n382, ZN => n463);
   U77 : AOI22_X1 port map( A1 => plusA(38), A2 => n281, B1 => plus2A(38), B2 
                           => n275, ZN => n383);
   U78 : AOI22_X1 port map( A1 => minus2A(38), A2 => n293, B1 => minusA(38), B2
                           => n287, ZN => n382);
   U79 : NAND2_X1 port map( A1 => n375, A2 => n374, ZN => n467);
   U80 : AOI22_X1 port map( A1 => plusA(34), A2 => n280, B1 => plus2A(34), B2 
                           => n274, ZN => n375);
   U81 : AOI22_X1 port map( A1 => minus2A(34), A2 => n292, B1 => minusA(34), B2
                           => n286, ZN => n374);
   U82 : NAND2_X1 port map( A1 => n367, A2 => n366, ZN => n471);
   U83 : AOI22_X1 port map( A1 => plusA(30), A2 => n280, B1 => plus2A(30), B2 
                           => n274, ZN => n367);
   U84 : AOI22_X1 port map( A1 => minus2A(30), A2 => n292, B1 => minusA(30), B2
                           => n286, ZN => n366);
   U85 : NAND2_X1 port map( A1 => n395, A2 => n394, ZN => n457);
   U86 : AOI22_X1 port map( A1 => plusA(44), A2 => n281, B1 => plus2A(44), B2 
                           => n275, ZN => n395);
   U87 : AOI22_X1 port map( A1 => minus2A(44), A2 => n293, B1 => minusA(44), B2
                           => n287, ZN => n394);
   U88 : NAND2_X1 port map( A1 => n387, A2 => n386, ZN => n461);
   U89 : AOI22_X1 port map( A1 => plusA(40), A2 => n281, B1 => plus2A(40), B2 
                           => n275, ZN => n387);
   U90 : AOI22_X1 port map( A1 => minus2A(40), A2 => n293, B1 => minusA(40), B2
                           => n287, ZN => n386);
   U91 : NAND2_X1 port map( A1 => n379, A2 => n378, ZN => n465);
   U92 : AOI22_X1 port map( A1 => plusA(36), A2 => n281, B1 => plus2A(36), B2 
                           => n275, ZN => n379);
   U93 : AOI22_X1 port map( A1 => minus2A(36), A2 => n293, B1 => minusA(36), B2
                           => n287, ZN => n378);
   U94 : NAND2_X1 port map( A1 => n371, A2 => n370, ZN => n469);
   U95 : AOI22_X1 port map( A1 => plusA(32), A2 => n280, B1 => plus2A(32), B2 
                           => n274, ZN => n371);
   U96 : AOI22_X1 port map( A1 => minus2A(32), A2 => n292, B1 => minusA(32), B2
                           => n286, ZN => n370);
   U97 : NAND2_X1 port map( A1 => n397, A2 => n396, ZN => n456);
   U98 : AOI22_X1 port map( A1 => plusA(45), A2 => n281, B1 => plus2A(45), B2 
                           => n275, ZN => n397);
   U99 : AOI22_X1 port map( A1 => minus2A(45), A2 => n293, B1 => minusA(45), B2
                           => n287, ZN => n396);
   U100 : NAND2_X1 port map( A1 => n393, A2 => n392, ZN => n458);
   U101 : AOI22_X1 port map( A1 => plusA(43), A2 => n281, B1 => plus2A(43), B2 
                           => n275, ZN => n393);
   U102 : AOI22_X1 port map( A1 => minus2A(43), A2 => n293, B1 => minusA(43), 
                           B2 => n287, ZN => n392);
   U103 : NAND2_X1 port map( A1 => n385, A2 => n384, ZN => n462);
   U104 : AOI22_X1 port map( A1 => plusA(39), A2 => n281, B1 => plus2A(39), B2 
                           => n275, ZN => n385);
   U105 : AOI22_X1 port map( A1 => minus2A(39), A2 => n293, B1 => minusA(39), 
                           B2 => n287, ZN => n384);
   U106 : NAND2_X1 port map( A1 => n377, A2 => n376, ZN => n466);
   U107 : AOI22_X1 port map( A1 => plusA(35), A2 => n280, B1 => plus2A(35), B2 
                           => n274, ZN => n377);
   U108 : AOI22_X1 port map( A1 => minus2A(35), A2 => n292, B1 => minusA(35), 
                           B2 => n286, ZN => n376);
   U109 : NAND2_X1 port map( A1 => n369, A2 => n368, ZN => n470);
   U110 : AOI22_X1 port map( A1 => plusA(31), A2 => n280, B1 => plus2A(31), B2 
                           => n274, ZN => n369);
   U111 : AOI22_X1 port map( A1 => minus2A(31), A2 => n292, B1 => minusA(31), 
                           B2 => n286, ZN => n368);
   U112 : NAND2_X1 port map( A1 => n389, A2 => n388, ZN => n460);
   U113 : AOI22_X1 port map( A1 => plusA(41), A2 => n281, B1 => plus2A(41), B2 
                           => n275, ZN => n389);
   U114 : AOI22_X1 port map( A1 => minus2A(41), A2 => n293, B1 => minusA(41), 
                           B2 => n287, ZN => n388);
   U115 : NAND2_X1 port map( A1 => n381, A2 => n380, ZN => n464);
   U116 : AOI22_X1 port map( A1 => plusA(37), A2 => n281, B1 => plus2A(37), B2 
                           => n275, ZN => n381);
   U117 : AOI22_X1 port map( A1 => minus2A(37), A2 => n293, B1 => minusA(37), 
                           B2 => n287, ZN => n380);
   U118 : NAND2_X1 port map( A1 => n373, A2 => n372, ZN => n468);
   U119 : AOI22_X1 port map( A1 => plusA(33), A2 => n280, B1 => plus2A(33), B2 
                           => n274, ZN => n373);
   U120 : AOI22_X1 port map( A1 => minus2A(33), A2 => n292, B1 => minusA(33), 
                           B2 => n286, ZN => n372);
   U121 : NAND2_X1 port map( A1 => n399, A2 => n398, ZN => n455);
   U122 : AOI22_X1 port map( A1 => plusA(46), A2 => n281, B1 => plus2A(46), B2 
                           => n275, ZN => n399);
   U123 : AOI22_X1 port map( A1 => minus2A(46), A2 => n293, B1 => minusA(46), 
                           B2 => n287, ZN => n398);
   U124 : NAND2_X1 port map( A1 => n431, A2 => n430, ZN => n439);
   U125 : AOI22_X1 port map( A1 => plusA(62), A2 => n283, B1 => plus2A(62), B2 
                           => n277, ZN => n431);
   U126 : AOI22_X1 port map( A1 => minus2A(62), A2 => n295, B1 => minusA(62), 
                           B2 => n289, ZN => n430);
   U127 : NAND2_X1 port map( A1 => n429, A2 => n428, ZN => n440);
   U128 : AOI22_X1 port map( A1 => plusA(61), A2 => n283, B1 => plus2A(61), B2 
                           => n277, ZN => n429);
   U129 : AOI22_X1 port map( A1 => minus2A(61), A2 => n295, B1 => minusA(61), 
                           B2 => n289, ZN => n428);
   U130 : NAND2_X1 port map( A1 => n427, A2 => n426, ZN => n441);
   U131 : AOI22_X1 port map( A1 => plusA(60), A2 => n283, B1 => plus2A(60), B2 
                           => n277, ZN => n427);
   U132 : AOI22_X1 port map( A1 => minus2A(60), A2 => n295, B1 => minusA(60), 
                           B2 => n289, ZN => n426);
   U133 : NAND2_X1 port map( A1 => n425, A2 => n424, ZN => n442);
   U134 : AOI22_X1 port map( A1 => plusA(59), A2 => n282, B1 => plus2A(59), B2 
                           => n276, ZN => n425);
   U135 : AOI22_X1 port map( A1 => minus2A(59), A2 => n294, B1 => minusA(59), 
                           B2 => n288, ZN => n424);
   U136 : NAND2_X1 port map( A1 => n423, A2 => n422, ZN => n443);
   U137 : AOI22_X1 port map( A1 => plusA(58), A2 => n282, B1 => plus2A(58), B2 
                           => n276, ZN => n423);
   U138 : AOI22_X1 port map( A1 => minus2A(58), A2 => n294, B1 => minusA(58), 
                           B2 => n288, ZN => n422);
   U139 : NAND2_X1 port map( A1 => n421, A2 => n420, ZN => n444);
   U140 : AOI22_X1 port map( A1 => plusA(57), A2 => n282, B1 => plus2A(57), B2 
                           => n276, ZN => n421);
   U141 : AOI22_X1 port map( A1 => minus2A(57), A2 => n294, B1 => minusA(57), 
                           B2 => n288, ZN => n420);
   U142 : NAND2_X1 port map( A1 => n419, A2 => n418, ZN => n445);
   U143 : AOI22_X1 port map( A1 => plusA(56), A2 => n282, B1 => plus2A(56), B2 
                           => n276, ZN => n419);
   U144 : AOI22_X1 port map( A1 => minus2A(56), A2 => n294, B1 => minusA(56), 
                           B2 => n288, ZN => n418);
   U145 : BUF_X1 port map( A => n433, Z => n279);
   U146 : BUF_X1 port map( A => n434, Z => n285);
   U147 : BUF_X1 port map( A => n432, Z => n273);
   U148 : BUF_X1 port map( A => n435, Z => n291);
   U149 : NAND2_X1 port map( A1 => n339, A2 => n338, ZN => n485);
   U150 : AOI22_X1 port map( A1 => plusA(16), A2 => n279, B1 => plus2A(16), B2 
                           => n273, ZN => n339);
   U151 : AOI22_X1 port map( A1 => minus2A(16), A2 => n291, B1 => minusA(16), 
                           B2 => n285, ZN => n338);
   U152 : NAND2_X1 port map( A1 => n341, A2 => n340, ZN => n484);
   U153 : AOI22_X1 port map( A1 => plusA(17), A2 => n279, B1 => plus2A(17), B2 
                           => n273, ZN => n341);
   U154 : AOI22_X1 port map( A1 => minus2A(17), A2 => n291, B1 => minusA(17), 
                           B2 => n285, ZN => n340);
   U155 : BUF_X1 port map( A => n433, Z => n280);
   U156 : BUF_X1 port map( A => n434, Z => n286);
   U157 : BUF_X1 port map( A => n432, Z => n274);
   U158 : BUF_X1 port map( A => n435, Z => n292);
   U159 : BUF_X1 port map( A => n433, Z => n281);
   U160 : BUF_X1 port map( A => n434, Z => n287);
   U161 : BUF_X1 port map( A => n432, Z => n275);
   U162 : BUF_X1 port map( A => n435, Z => n293);
   U163 : NAND2_X1 port map( A1 => n437, A2 => n436, ZN => n438);
   U164 : AOI22_X1 port map( A1 => plusA(63), A2 => n283, B1 => plus2A(63), B2 
                           => n277, ZN => n437);
   U165 : AOI22_X1 port map( A1 => minus2A(63), A2 => n295, B1 => minusA(63), 
                           B2 => n289, ZN => n436);
   U166 : BUF_X1 port map( A => n433, Z => n282);
   U167 : BUF_X1 port map( A => n434, Z => n288);
   U168 : BUF_X1 port map( A => n432, Z => n276);
   U169 : BUF_X1 port map( A => n435, Z => n294);
   U170 : BUF_X1 port map( A => n433, Z => n278);
   U171 : BUF_X1 port map( A => n434, Z => n284);
   U172 : BUF_X1 port map( A => n432, Z => n272);
   U173 : BUF_X1 port map( A => n435, Z => n290);
   U174 : NOR2_X1 port map( A1 => n323, A2 => n304, ZN => n493);
   U175 : INV_X1 port map( A => SEL(2), ZN => n304);
   U176 : AND2_X1 port map( A1 => SEL(2), A2 => n323, ZN => n435);
   U177 : NOR2_X1 port map( A1 => SEL(1), A2 => SEL(0), ZN => n323);
   U178 : INV_X1 port map( A => SEL(1), ZN => n302);
   U179 : INV_X1 port map( A => SEL(0), ZN => n303);
   U180 : NAND2_X1 port map( A1 => n337, A2 => n336, ZN => n486);
   U181 : AOI22_X1 port map( A1 => plusA(15), A2 => n279, B1 => plus2A(15), B2 
                           => n273, ZN => n337);
   U182 : AOI22_X1 port map( A1 => minus2A(15), A2 => n291, B1 => minusA(15), 
                           B2 => n285, ZN => n336);
   U183 : NAND2_X1 port map( A1 => n335, A2 => n334, ZN => n487);
   U184 : AOI22_X1 port map( A1 => plusA(14), A2 => n279, B1 => plus2A(14), B2 
                           => n273, ZN => n335);
   U185 : AOI22_X1 port map( A1 => minus2A(14), A2 => n291, B1 => minusA(14), 
                           B2 => n285, ZN => n334);
   U186 : NAND2_X1 port map( A1 => n333, A2 => n332, ZN => n488);
   U187 : AOI22_X1 port map( A1 => plusA(13), A2 => n279, B1 => plus2A(13), B2 
                           => n273, ZN => n333);
   U188 : AOI22_X1 port map( A1 => minus2A(13), A2 => n291, B1 => minusA(13), 
                           B2 => n285, ZN => n332);
   U189 : NAND2_X1 port map( A1 => n329, A2 => n328, ZN => n490);
   U190 : AOI22_X1 port map( A1 => plusA(11), A2 => n278, B1 => plus2A(11), B2 
                           => n272, ZN => n329);
   U191 : AOI22_X1 port map( A1 => minus2A(11), A2 => n290, B1 => minusA(11), 
                           B2 => n284, ZN => n328);
   U192 : NAND2_X1 port map( A1 => n327, A2 => n326, ZN => n491);
   U193 : AOI22_X1 port map( A1 => plusA(10), A2 => n278, B1 => plus2A(10), B2 
                           => n272, ZN => n327);
   U194 : AOI22_X1 port map( A1 => minus2A(10), A2 => n290, B1 => minusA(10), 
                           B2 => n284, ZN => n326);
   U195 : NAND2_X1 port map( A1 => n325, A2 => n324, ZN => n492);
   U196 : AOI22_X1 port map( A1 => plusA(9), A2 => n278, B1 => plus2A(9), B2 =>
                           n272, ZN => n325);
   U197 : AOI22_X1 port map( A1 => minus2A(9), A2 => n290, B1 => minusA(9), B2 
                           => n284, ZN => n324);
   U198 : NAND2_X1 port map( A1 => n320, A2 => n319, ZN => n495);
   U199 : AOI22_X1 port map( A1 => plusA(7), A2 => n278, B1 => plus2A(7), B2 =>
                           n272, ZN => n320);
   U200 : AOI22_X1 port map( A1 => minus2A(7), A2 => n290, B1 => minusA(7), B2 
                           => n284, ZN => n319);
   U201 : NAND2_X1 port map( A1 => n318, A2 => n317, ZN => n496);
   U202 : AOI22_X1 port map( A1 => plusA(6), A2 => n278, B1 => plus2A(6), B2 =>
                           n272, ZN => n318);
   U203 : AOI22_X1 port map( A1 => minus2A(6), A2 => n290, B1 => minusA(6), B2 
                           => n284, ZN => n317);
   U204 : NAND2_X1 port map( A1 => n316, A2 => n315, ZN => n497);
   U205 : AOI22_X1 port map( A1 => plusA(5), A2 => n278, B1 => plus2A(5), B2 =>
                           n272, ZN => n316);
   U206 : AOI22_X1 port map( A1 => minus2A(5), A2 => n290, B1 => minusA(5), B2 
                           => n284, ZN => n315);
   U207 : NAND2_X1 port map( A1 => n312, A2 => n311, ZN => n499);
   U208 : AOI22_X1 port map( A1 => plusA(3), A2 => n278, B1 => plus2A(3), B2 =>
                           n272, ZN => n312);
   U209 : AOI22_X1 port map( A1 => minus2A(3), A2 => n290, B1 => minusA(3), B2 
                           => n284, ZN => n311);
   U210 : NAND2_X1 port map( A1 => n331, A2 => n330, ZN => n489);
   U211 : AOI22_X1 port map( A1 => plusA(12), A2 => n279, B1 => plus2A(12), B2 
                           => n273, ZN => n331);
   U212 : AOI22_X1 port map( A1 => minus2A(12), A2 => n291, B1 => minusA(12), 
                           B2 => n285, ZN => n330);
   U213 : NAND2_X1 port map( A1 => n322, A2 => n321, ZN => n494);
   U214 : AOI22_X1 port map( A1 => plusA(8), A2 => n278, B1 => plus2A(8), B2 =>
                           n272, ZN => n322);
   U215 : AOI22_X1 port map( A1 => minus2A(8), A2 => n290, B1 => minusA(8), B2 
                           => n284, ZN => n321);
   U216 : NAND2_X1 port map( A1 => n314, A2 => n313, ZN => n498);
   U217 : AOI22_X1 port map( A1 => plusA(4), A2 => n278, B1 => plus2A(4), B2 =>
                           n272, ZN => n314);
   U218 : AOI22_X1 port map( A1 => minus2A(4), A2 => n290, B1 => minusA(4), B2 
                           => n284, ZN => n313);
   U219 : NAND2_X1 port map( A1 => n310, A2 => n309, ZN => n500);
   U220 : AOI22_X1 port map( A1 => plusA(2), A2 => n278, B1 => plus2A(2), B2 =>
                           n272, ZN => n310);
   U221 : AOI22_X1 port map( A1 => minus2A(2), A2 => n290, B1 => minusA(2), B2 
                           => n284, ZN => n309);
   U222 : NAND2_X1 port map( A1 => n308, A2 => n307, ZN => n501);
   U223 : AOI22_X1 port map( A1 => plusA(1), A2 => n278, B1 => plus2A(1), B2 =>
                           n272, ZN => n308);
   U224 : AOI22_X1 port map( A1 => minus2A(1), A2 => n290, B1 => minusA(1), B2 
                           => n284, ZN => n307);
   U225 : NAND2_X1 port map( A1 => n306, A2 => n305, ZN => n502);
   U226 : AOI22_X1 port map( A1 => plusA(0), A2 => n278, B1 => plus2A(0), B2 =>
                           n272, ZN => n306);
   U227 : AOI22_X1 port map( A1 => minus2A(0), A2 => n290, B1 => minusA(0), B2 
                           => n284, ZN => n305);
   U228 : CLKBUF_X1 port map( A => n432, Z => n277);
   U229 : CLKBUF_X1 port map( A => n433, Z => n283);
   U230 : CLKBUF_X1 port map( A => n434, Z => n289);
   U231 : CLKBUF_X1 port map( A => n435, Z => n295);
   U232 : CLKBUF_X1 port map( A => n493, Z => n301);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity MUX_GENERIC_N64_RADIX3_8 is

   port( plusA, minusA, plus2A, minus2A : in std_logic_vector (63 downto 0);  
         SEL : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (63 
         downto 0));

end MUX_GENERIC_N64_RADIX3_8;

architecture SYN_beh of MUX_GENERIC_N64_RADIX3_8 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component TBUF_X2
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   component TBUF_X1
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   signal n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, 
      n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, 
      n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, 
      n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, 
      n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, 
      n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, 
      n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, 
      n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, 
      n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, 
      n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, 
      n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, 
      n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, 
      n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, 
      n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, 
      n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, 
      n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, 
      n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, 
      n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, 
      n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, 
      n499, n500, n501, n502 : std_logic;

begin
   
   Y_tri_60_inst : TBUF_X1 port map( A => n441, EN => n301, Z => Y(60));
   Y_tri_61_inst : TBUF_X1 port map( A => n440, EN => n301, Z => Y(61));
   Y_tri_62_inst : TBUF_X1 port map( A => n439, EN => n301, Z => Y(62));
   Y_tri_63_inst : TBUF_X1 port map( A => n438, EN => n301, Z => Y(63));
   Y_tri_50_inst : TBUF_X1 port map( A => n451, EN => n300, Z => Y(50));
   Y_tri_51_inst : TBUF_X1 port map( A => n450, EN => n300, Z => Y(51));
   Y_tri_52_inst : TBUF_X1 port map( A => n449, EN => n300, Z => Y(52));
   Y_tri_53_inst : TBUF_X1 port map( A => n448, EN => n300, Z => Y(53));
   Y_tri_54_inst : TBUF_X1 port map( A => n447, EN => n300, Z => Y(54));
   Y_tri_55_inst : TBUF_X1 port map( A => n446, EN => n300, Z => Y(55));
   Y_tri_56_inst : TBUF_X1 port map( A => n445, EN => n300, Z => Y(56));
   Y_tri_57_inst : TBUF_X1 port map( A => n444, EN => n300, Z => Y(57));
   Y_tri_58_inst : TBUF_X1 port map( A => n443, EN => n300, Z => Y(58));
   Y_tri_59_inst : TBUF_X1 port map( A => n442, EN => n300, Z => Y(59));
   Y_tri_23_inst : TBUF_X1 port map( A => n478, EN => n297, Z => Y(23));
   Y_tri_24_inst : TBUF_X1 port map( A => n477, EN => n298, Z => Y(24));
   Y_tri_25_inst : TBUF_X1 port map( A => n476, EN => n298, Z => Y(25));
   Y_tri_26_inst : TBUF_X1 port map( A => n475, EN => n298, Z => Y(26));
   Y_tri_27_inst : TBUF_X1 port map( A => n474, EN => n298, Z => Y(27));
   Y_tri_28_inst : TBUF_X1 port map( A => n473, EN => n298, Z => Y(28));
   Y_tri_29_inst : TBUF_X1 port map( A => n472, EN => n298, Z => Y(29));
   Y_tri_30_inst : TBUF_X1 port map( A => n471, EN => n298, Z => Y(30));
   Y_tri_31_inst : TBUF_X1 port map( A => n470, EN => n298, Z => Y(31));
   Y_tri_32_inst : TBUF_X1 port map( A => n469, EN => n298, Z => Y(32));
   Y_tri_33_inst : TBUF_X1 port map( A => n468, EN => n298, Z => Y(33));
   Y_tri_34_inst : TBUF_X1 port map( A => n467, EN => n298, Z => Y(34));
   Y_tri_35_inst : TBUF_X1 port map( A => n466, EN => n298, Z => Y(35));
   Y_tri_36_inst : TBUF_X1 port map( A => n465, EN => n299, Z => Y(36));
   Y_tri_37_inst : TBUF_X1 port map( A => n464, EN => n299, Z => Y(37));
   Y_tri_38_inst : TBUF_X1 port map( A => n463, EN => n299, Z => Y(38));
   Y_tri_39_inst : TBUF_X1 port map( A => n462, EN => n299, Z => Y(39));
   Y_tri_40_inst : TBUF_X1 port map( A => n461, EN => n299, Z => Y(40));
   Y_tri_41_inst : TBUF_X1 port map( A => n460, EN => n299, Z => Y(41));
   Y_tri_42_inst : TBUF_X1 port map( A => n459, EN => n299, Z => Y(42));
   Y_tri_43_inst : TBUF_X1 port map( A => n458, EN => n299, Z => Y(43));
   Y_tri_45_inst : TBUF_X1 port map( A => n456, EN => n299, Z => Y(45));
   Y_tri_46_inst : TBUF_X1 port map( A => n455, EN => n299, Z => Y(46));
   Y_tri_47_inst : TBUF_X1 port map( A => n454, EN => n299, Z => Y(47));
   Y_tri_48_inst : TBUF_X1 port map( A => n453, EN => n300, Z => Y(48));
   Y_tri_49_inst : TBUF_X1 port map( A => n452, EN => n300, Z => Y(49));
   Y_tri_44_inst : TBUF_X1 port map( A => n457, EN => n299, Z => Y(44));
   Y_tri_10_inst : TBUF_X1 port map( A => n491, EN => n296, Z => Y(10));
   Y_tri_11_inst : TBUF_X1 port map( A => n490, EN => n296, Z => Y(11));
   Y_tri_12_inst : TBUF_X1 port map( A => n489, EN => n297, Z => Y(12));
   Y_tri_13_inst : TBUF_X1 port map( A => n488, EN => n297, Z => Y(13));
   Y_tri_14_inst : TBUF_X1 port map( A => n487, EN => n297, Z => Y(14));
   Y_tri_15_inst : TBUF_X1 port map( A => n486, EN => n297, Z => Y(15));
   Y_tri_16_inst : TBUF_X1 port map( A => n485, EN => n297, Z => Y(16));
   Y_tri_17_inst : TBUF_X1 port map( A => n484, EN => n297, Z => Y(17));
   Y_tri_18_inst : TBUF_X1 port map( A => n483, EN => n297, Z => Y(18));
   Y_tri_19_inst : TBUF_X1 port map( A => n482, EN => n297, Z => Y(19));
   Y_tri_20_inst : TBUF_X1 port map( A => n481, EN => n297, Z => Y(20));
   Y_tri_21_inst : TBUF_X1 port map( A => n480, EN => n297, Z => Y(21));
   Y_tri_22_inst : TBUF_X1 port map( A => n479, EN => n297, Z => Y(22));
   Y_tri_5_inst : TBUF_X1 port map( A => n497, EN => n296, Z => Y(5));
   Y_tri_4_inst : TBUF_X1 port map( A => n498, EN => n296, Z => Y(4));
   Y_tri_3_inst : TBUF_X1 port map( A => n499, EN => n296, Z => Y(3));
   Y_tri_6_inst : TBUF_X1 port map( A => n496, EN => n296, Z => Y(6));
   Y_tri_7_inst : TBUF_X1 port map( A => n495, EN => n296, Z => Y(7));
   Y_tri_8_inst : TBUF_X1 port map( A => n494, EN => n296, Z => Y(8));
   Y_tri_2_inst : TBUF_X1 port map( A => n500, EN => n296, Z => Y(2));
   Y_tri_1_inst : TBUF_X1 port map( A => n501, EN => n296, Z => Y(1));
   Y_tri_0_inst : TBUF_X1 port map( A => n502, EN => n296, Z => Y(0));
   Y_tri_9_inst : TBUF_X2 port map( A => n492, EN => n296, Z => Y(9));
   U2 : NOR3_X1 port map( A1 => SEL(0), A2 => SEL(2), A3 => n302, ZN => n434);
   U3 : NOR3_X1 port map( A1 => n302, A2 => SEL(2), A3 => n303, ZN => n432);
   U4 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n303, ZN => n433);
   U5 : CLKBUF_X3 port map( A => n493, Z => n296);
   U6 : CLKBUF_X1 port map( A => n493, Z => n297);
   U7 : CLKBUF_X1 port map( A => n493, Z => n298);
   U8 : CLKBUF_X1 port map( A => n493, Z => n299);
   U9 : CLKBUF_X1 port map( A => n493, Z => n300);
   U10 : NAND2_X1 port map( A1 => n349, A2 => n348, ZN => n480);
   U11 : AOI22_X1 port map( A1 => plusA(21), A2 => n279, B1 => plus2A(21), B2 
                           => n273, ZN => n349);
   U12 : AOI22_X1 port map( A1 => minus2A(21), A2 => n291, B1 => minusA(21), B2
                           => n285, ZN => n348);
   U13 : NAND2_X1 port map( A1 => n347, A2 => n346, ZN => n481);
   U14 : AOI22_X1 port map( A1 => plusA(20), A2 => n279, B1 => plus2A(20), B2 
                           => n273, ZN => n347);
   U15 : AOI22_X1 port map( A1 => minus2A(20), A2 => n291, B1 => minusA(20), B2
                           => n285, ZN => n346);
   U16 : NAND2_X1 port map( A1 => n351, A2 => n350, ZN => n479);
   U17 : AOI22_X1 port map( A1 => plusA(22), A2 => n279, B1 => plus2A(22), B2 
                           => n273, ZN => n351);
   U18 : AOI22_X1 port map( A1 => minus2A(22), A2 => n291, B1 => minusA(22), B2
                           => n285, ZN => n350);
   U19 : NAND2_X1 port map( A1 => n405, A2 => n404, ZN => n452);
   U20 : AOI22_X1 port map( A1 => plusA(49), A2 => n282, B1 => plus2A(49), B2 
                           => n276, ZN => n405);
   U21 : AOI22_X1 port map( A1 => minus2A(49), A2 => n294, B1 => minusA(49), B2
                           => n288, ZN => n404);
   U22 : NAND2_X1 port map( A1 => n403, A2 => n402, ZN => n453);
   U23 : AOI22_X1 port map( A1 => plusA(48), A2 => n282, B1 => plus2A(48), B2 
                           => n276, ZN => n403);
   U24 : AOI22_X1 port map( A1 => minus2A(48), A2 => n294, B1 => minusA(48), B2
                           => n288, ZN => n402);
   U25 : NAND2_X1 port map( A1 => n401, A2 => n400, ZN => n454);
   U26 : AOI22_X1 port map( A1 => plusA(47), A2 => n281, B1 => plus2A(47), B2 
                           => n275, ZN => n401);
   U27 : AOI22_X1 port map( A1 => minus2A(47), A2 => n293, B1 => minusA(47), B2
                           => n287, ZN => n400);
   U28 : NAND2_X1 port map( A1 => n399, A2 => n398, ZN => n455);
   U29 : AOI22_X1 port map( A1 => plusA(46), A2 => n281, B1 => plus2A(46), B2 
                           => n275, ZN => n399);
   U30 : AOI22_X1 port map( A1 => minus2A(46), A2 => n293, B1 => minusA(46), B2
                           => n287, ZN => n398);
   U31 : NAND2_X1 port map( A1 => n397, A2 => n396, ZN => n456);
   U32 : AOI22_X1 port map( A1 => plusA(45), A2 => n281, B1 => plus2A(45), B2 
                           => n275, ZN => n397);
   U33 : AOI22_X1 port map( A1 => minus2A(45), A2 => n293, B1 => minusA(45), B2
                           => n287, ZN => n396);
   U34 : NAND2_X1 port map( A1 => n393, A2 => n392, ZN => n458);
   U35 : AOI22_X1 port map( A1 => plusA(43), A2 => n281, B1 => plus2A(43), B2 
                           => n275, ZN => n393);
   U36 : AOI22_X1 port map( A1 => minus2A(43), A2 => n293, B1 => minusA(43), B2
                           => n287, ZN => n392);
   U37 : NAND2_X1 port map( A1 => n385, A2 => n384, ZN => n462);
   U38 : AOI22_X1 port map( A1 => plusA(39), A2 => n281, B1 => plus2A(39), B2 
                           => n275, ZN => n385);
   U39 : AOI22_X1 port map( A1 => minus2A(39), A2 => n293, B1 => minusA(39), B2
                           => n287, ZN => n384);
   U40 : NAND2_X1 port map( A1 => n377, A2 => n376, ZN => n466);
   U41 : AOI22_X1 port map( A1 => plusA(35), A2 => n280, B1 => plus2A(35), B2 
                           => n274, ZN => n377);
   U42 : AOI22_X1 port map( A1 => minus2A(35), A2 => n292, B1 => minusA(35), B2
                           => n286, ZN => n376);
   U43 : NAND2_X1 port map( A1 => n369, A2 => n368, ZN => n470);
   U44 : AOI22_X1 port map( A1 => plusA(31), A2 => n280, B1 => plus2A(31), B2 
                           => n274, ZN => n369);
   U45 : AOI22_X1 port map( A1 => minus2A(31), A2 => n292, B1 => minusA(31), B2
                           => n286, ZN => n368);
   U46 : NAND2_X1 port map( A1 => n361, A2 => n360, ZN => n474);
   U47 : AOI22_X1 port map( A1 => plusA(27), A2 => n280, B1 => plus2A(27), B2 
                           => n274, ZN => n361);
   U48 : AOI22_X1 port map( A1 => minus2A(27), A2 => n292, B1 => minusA(27), B2
                           => n286, ZN => n360);
   U49 : NAND2_X1 port map( A1 => n353, A2 => n352, ZN => n478);
   U50 : AOI22_X1 port map( A1 => plusA(23), A2 => n279, B1 => plus2A(23), B2 
                           => n273, ZN => n353);
   U51 : AOI22_X1 port map( A1 => minus2A(23), A2 => n291, B1 => minusA(23), B2
                           => n285, ZN => n352);
   U52 : NAND2_X1 port map( A1 => n389, A2 => n388, ZN => n460);
   U53 : AOI22_X1 port map( A1 => plusA(41), A2 => n281, B1 => plus2A(41), B2 
                           => n275, ZN => n389);
   U54 : AOI22_X1 port map( A1 => minus2A(41), A2 => n293, B1 => minusA(41), B2
                           => n287, ZN => n388);
   U55 : NAND2_X1 port map( A1 => n381, A2 => n380, ZN => n464);
   U56 : AOI22_X1 port map( A1 => plusA(37), A2 => n281, B1 => plus2A(37), B2 
                           => n275, ZN => n381);
   U57 : AOI22_X1 port map( A1 => minus2A(37), A2 => n293, B1 => minusA(37), B2
                           => n287, ZN => n380);
   U58 : NAND2_X1 port map( A1 => n373, A2 => n372, ZN => n468);
   U59 : AOI22_X1 port map( A1 => plusA(33), A2 => n280, B1 => plus2A(33), B2 
                           => n274, ZN => n373);
   U60 : AOI22_X1 port map( A1 => minus2A(33), A2 => n292, B1 => minusA(33), B2
                           => n286, ZN => n372);
   U61 : NAND2_X1 port map( A1 => n365, A2 => n364, ZN => n472);
   U62 : AOI22_X1 port map( A1 => plusA(29), A2 => n280, B1 => plus2A(29), B2 
                           => n274, ZN => n365);
   U63 : AOI22_X1 port map( A1 => minus2A(29), A2 => n292, B1 => minusA(29), B2
                           => n286, ZN => n364);
   U64 : NAND2_X1 port map( A1 => n357, A2 => n356, ZN => n476);
   U65 : AOI22_X1 port map( A1 => plusA(25), A2 => n280, B1 => plus2A(25), B2 
                           => n274, ZN => n357);
   U66 : AOI22_X1 port map( A1 => minus2A(25), A2 => n292, B1 => minusA(25), B2
                           => n286, ZN => n356);
   U67 : NAND2_X1 port map( A1 => n395, A2 => n394, ZN => n457);
   U68 : AOI22_X1 port map( A1 => plusA(44), A2 => n281, B1 => plus2A(44), B2 
                           => n275, ZN => n395);
   U69 : AOI22_X1 port map( A1 => minus2A(44), A2 => n293, B1 => minusA(44), B2
                           => n287, ZN => n394);
   U70 : NAND2_X1 port map( A1 => n387, A2 => n386, ZN => n461);
   U71 : AOI22_X1 port map( A1 => plusA(40), A2 => n281, B1 => plus2A(40), B2 
                           => n275, ZN => n387);
   U72 : AOI22_X1 port map( A1 => minus2A(40), A2 => n293, B1 => minusA(40), B2
                           => n287, ZN => n386);
   U73 : NAND2_X1 port map( A1 => n379, A2 => n378, ZN => n465);
   U74 : AOI22_X1 port map( A1 => plusA(36), A2 => n281, B1 => plus2A(36), B2 
                           => n275, ZN => n379);
   U75 : AOI22_X1 port map( A1 => minus2A(36), A2 => n293, B1 => minusA(36), B2
                           => n287, ZN => n378);
   U76 : NAND2_X1 port map( A1 => n371, A2 => n370, ZN => n469);
   U77 : AOI22_X1 port map( A1 => plusA(32), A2 => n280, B1 => plus2A(32), B2 
                           => n274, ZN => n371);
   U78 : AOI22_X1 port map( A1 => minus2A(32), A2 => n292, B1 => minusA(32), B2
                           => n286, ZN => n370);
   U79 : NAND2_X1 port map( A1 => n363, A2 => n362, ZN => n473);
   U80 : AOI22_X1 port map( A1 => plusA(28), A2 => n280, B1 => plus2A(28), B2 
                           => n274, ZN => n363);
   U81 : AOI22_X1 port map( A1 => minus2A(28), A2 => n292, B1 => minusA(28), B2
                           => n286, ZN => n362);
   U82 : NAND2_X1 port map( A1 => n355, A2 => n354, ZN => n477);
   U83 : AOI22_X1 port map( A1 => plusA(24), A2 => n280, B1 => plus2A(24), B2 
                           => n274, ZN => n355);
   U84 : AOI22_X1 port map( A1 => minus2A(24), A2 => n292, B1 => minusA(24), B2
                           => n286, ZN => n354);
   U85 : NAND2_X1 port map( A1 => n391, A2 => n390, ZN => n459);
   U86 : AOI22_X1 port map( A1 => plusA(42), A2 => n281, B1 => plus2A(42), B2 
                           => n275, ZN => n391);
   U87 : AOI22_X1 port map( A1 => minus2A(42), A2 => n293, B1 => minusA(42), B2
                           => n287, ZN => n390);
   U88 : NAND2_X1 port map( A1 => n383, A2 => n382, ZN => n463);
   U89 : AOI22_X1 port map( A1 => plusA(38), A2 => n281, B1 => plus2A(38), B2 
                           => n275, ZN => n383);
   U90 : AOI22_X1 port map( A1 => minus2A(38), A2 => n293, B1 => minusA(38), B2
                           => n287, ZN => n382);
   U91 : NAND2_X1 port map( A1 => n375, A2 => n374, ZN => n467);
   U92 : AOI22_X1 port map( A1 => plusA(34), A2 => n280, B1 => plus2A(34), B2 
                           => n274, ZN => n375);
   U93 : AOI22_X1 port map( A1 => minus2A(34), A2 => n292, B1 => minusA(34), B2
                           => n286, ZN => n374);
   U94 : NAND2_X1 port map( A1 => n367, A2 => n366, ZN => n471);
   U95 : AOI22_X1 port map( A1 => plusA(30), A2 => n280, B1 => plus2A(30), B2 
                           => n274, ZN => n367);
   U96 : AOI22_X1 port map( A1 => minus2A(30), A2 => n292, B1 => minusA(30), B2
                           => n286, ZN => n366);
   U97 : NAND2_X1 port map( A1 => n359, A2 => n358, ZN => n475);
   U98 : AOI22_X1 port map( A1 => plusA(26), A2 => n280, B1 => plus2A(26), B2 
                           => n274, ZN => n359);
   U99 : AOI22_X1 port map( A1 => minus2A(26), A2 => n292, B1 => minusA(26), B2
                           => n286, ZN => n358);
   U100 : NAND2_X1 port map( A1 => n437, A2 => n436, ZN => n438);
   U101 : AOI22_X1 port map( A1 => plusA(63), A2 => n283, B1 => plus2A(63), B2 
                           => n277, ZN => n437);
   U102 : AOI22_X1 port map( A1 => minus2A(63), A2 => n295, B1 => minusA(63), 
                           B2 => n289, ZN => n436);
   U103 : NAND2_X1 port map( A1 => n431, A2 => n430, ZN => n439);
   U104 : AOI22_X1 port map( A1 => plusA(62), A2 => n283, B1 => plus2A(62), B2 
                           => n277, ZN => n431);
   U105 : AOI22_X1 port map( A1 => minus2A(62), A2 => n295, B1 => minusA(62), 
                           B2 => n289, ZN => n430);
   U106 : NAND2_X1 port map( A1 => n429, A2 => n428, ZN => n440);
   U107 : AOI22_X1 port map( A1 => plusA(61), A2 => n283, B1 => plus2A(61), B2 
                           => n277, ZN => n429);
   U108 : AOI22_X1 port map( A1 => minus2A(61), A2 => n295, B1 => minusA(61), 
                           B2 => n289, ZN => n428);
   U109 : NAND2_X1 port map( A1 => n427, A2 => n426, ZN => n441);
   U110 : AOI22_X1 port map( A1 => plusA(60), A2 => n283, B1 => plus2A(60), B2 
                           => n277, ZN => n427);
   U111 : AOI22_X1 port map( A1 => minus2A(60), A2 => n295, B1 => minusA(60), 
                           B2 => n289, ZN => n426);
   U112 : NAND2_X1 port map( A1 => n425, A2 => n424, ZN => n442);
   U113 : AOI22_X1 port map( A1 => plusA(59), A2 => n282, B1 => plus2A(59), B2 
                           => n276, ZN => n425);
   U114 : AOI22_X1 port map( A1 => minus2A(59), A2 => n294, B1 => minusA(59), 
                           B2 => n288, ZN => n424);
   U115 : NAND2_X1 port map( A1 => n423, A2 => n422, ZN => n443);
   U116 : AOI22_X1 port map( A1 => plusA(58), A2 => n282, B1 => plus2A(58), B2 
                           => n276, ZN => n423);
   U117 : AOI22_X1 port map( A1 => minus2A(58), A2 => n294, B1 => minusA(58), 
                           B2 => n288, ZN => n422);
   U118 : NAND2_X1 port map( A1 => n421, A2 => n420, ZN => n444);
   U119 : AOI22_X1 port map( A1 => plusA(57), A2 => n282, B1 => plus2A(57), B2 
                           => n276, ZN => n421);
   U120 : AOI22_X1 port map( A1 => minus2A(57), A2 => n294, B1 => minusA(57), 
                           B2 => n288, ZN => n420);
   U121 : NAND2_X1 port map( A1 => n419, A2 => n418, ZN => n445);
   U122 : AOI22_X1 port map( A1 => plusA(56), A2 => n282, B1 => plus2A(56), B2 
                           => n276, ZN => n419);
   U123 : AOI22_X1 port map( A1 => minus2A(56), A2 => n294, B1 => minusA(56), 
                           B2 => n288, ZN => n418);
   U124 : NAND2_X1 port map( A1 => n417, A2 => n416, ZN => n446);
   U125 : AOI22_X1 port map( A1 => plusA(55), A2 => n282, B1 => plus2A(55), B2 
                           => n276, ZN => n417);
   U126 : AOI22_X1 port map( A1 => minus2A(55), A2 => n294, B1 => minusA(55), 
                           B2 => n288, ZN => n416);
   U127 : NAND2_X1 port map( A1 => n415, A2 => n414, ZN => n447);
   U128 : AOI22_X1 port map( A1 => plusA(54), A2 => n282, B1 => plus2A(54), B2 
                           => n276, ZN => n415);
   U129 : AOI22_X1 port map( A1 => minus2A(54), A2 => n294, B1 => minusA(54), 
                           B2 => n288, ZN => n414);
   U130 : NAND2_X1 port map( A1 => n413, A2 => n412, ZN => n448);
   U131 : AOI22_X1 port map( A1 => plusA(53), A2 => n282, B1 => plus2A(53), B2 
                           => n276, ZN => n413);
   U132 : AOI22_X1 port map( A1 => minus2A(53), A2 => n294, B1 => minusA(53), 
                           B2 => n288, ZN => n412);
   U133 : NAND2_X1 port map( A1 => n411, A2 => n410, ZN => n449);
   U134 : AOI22_X1 port map( A1 => plusA(52), A2 => n282, B1 => plus2A(52), B2 
                           => n276, ZN => n411);
   U135 : AOI22_X1 port map( A1 => minus2A(52), A2 => n294, B1 => minusA(52), 
                           B2 => n288, ZN => n410);
   U136 : NAND2_X1 port map( A1 => n409, A2 => n408, ZN => n450);
   U137 : AOI22_X1 port map( A1 => plusA(51), A2 => n282, B1 => plus2A(51), B2 
                           => n276, ZN => n409);
   U138 : AOI22_X1 port map( A1 => minus2A(51), A2 => n294, B1 => minusA(51), 
                           B2 => n288, ZN => n408);
   U139 : NAND2_X1 port map( A1 => n407, A2 => n406, ZN => n451);
   U140 : AOI22_X1 port map( A1 => plusA(50), A2 => n282, B1 => plus2A(50), B2 
                           => n276, ZN => n407);
   U141 : AOI22_X1 port map( A1 => minus2A(50), A2 => n294, B1 => minusA(50), 
                           B2 => n288, ZN => n406);
   U142 : BUF_X1 port map( A => n433, Z => n279);
   U143 : BUF_X1 port map( A => n434, Z => n285);
   U144 : BUF_X1 port map( A => n432, Z => n273);
   U145 : NAND2_X1 port map( A1 => n345, A2 => n344, ZN => n482);
   U146 : AOI22_X1 port map( A1 => plusA(19), A2 => n279, B1 => plus2A(19), B2 
                           => n273, ZN => n345);
   U147 : AOI22_X1 port map( A1 => minus2A(19), A2 => n291, B1 => minusA(19), 
                           B2 => n285, ZN => n344);
   U148 : NAND2_X1 port map( A1 => n343, A2 => n342, ZN => n483);
   U149 : AOI22_X1 port map( A1 => plusA(18), A2 => n279, B1 => plus2A(18), B2 
                           => n273, ZN => n343);
   U150 : AOI22_X1 port map( A1 => minus2A(18), A2 => n291, B1 => minusA(18), 
                           B2 => n285, ZN => n342);
   U151 : BUF_X1 port map( A => n433, Z => n280);
   U152 : BUF_X1 port map( A => n434, Z => n286);
   U153 : BUF_X1 port map( A => n432, Z => n274);
   U154 : BUF_X1 port map( A => n435, Z => n292);
   U155 : BUF_X1 port map( A => n435, Z => n291);
   U156 : BUF_X1 port map( A => n433, Z => n281);
   U157 : BUF_X1 port map( A => n434, Z => n287);
   U158 : BUF_X1 port map( A => n432, Z => n275);
   U159 : BUF_X1 port map( A => n435, Z => n293);
   U160 : BUF_X1 port map( A => n433, Z => n282);
   U161 : BUF_X1 port map( A => n434, Z => n288);
   U162 : BUF_X1 port map( A => n432, Z => n276);
   U163 : BUF_X1 port map( A => n435, Z => n294);
   U164 : BUF_X1 port map( A => n433, Z => n278);
   U165 : BUF_X1 port map( A => n434, Z => n284);
   U166 : BUF_X1 port map( A => n432, Z => n272);
   U167 : BUF_X1 port map( A => n435, Z => n290);
   U168 : NOR2_X1 port map( A1 => n323, A2 => n304, ZN => n493);
   U169 : INV_X1 port map( A => SEL(2), ZN => n304);
   U170 : NOR2_X1 port map( A1 => SEL(1), A2 => SEL(0), ZN => n323);
   U171 : INV_X1 port map( A => SEL(1), ZN => n302);
   U172 : INV_X1 port map( A => SEL(0), ZN => n303);
   U173 : NAND2_X1 port map( A1 => n341, A2 => n340, ZN => n484);
   U174 : AOI22_X1 port map( A1 => plusA(17), A2 => n279, B1 => plus2A(17), B2 
                           => n273, ZN => n341);
   U175 : AOI22_X1 port map( A1 => minus2A(17), A2 => n291, B1 => minusA(17), 
                           B2 => n285, ZN => n340);
   U176 : AND2_X1 port map( A1 => SEL(2), A2 => n323, ZN => n435);
   U177 : NAND2_X1 port map( A1 => n339, A2 => n338, ZN => n485);
   U178 : AOI22_X1 port map( A1 => plusA(16), A2 => n279, B1 => plus2A(16), B2 
                           => n273, ZN => n339);
   U179 : AOI22_X1 port map( A1 => minus2A(16), A2 => n291, B1 => minusA(16), 
                           B2 => n285, ZN => n338);
   U180 : NAND2_X1 port map( A1 => n337, A2 => n336, ZN => n486);
   U181 : AOI22_X1 port map( A1 => plusA(15), A2 => n279, B1 => plus2A(15), B2 
                           => n273, ZN => n337);
   U182 : AOI22_X1 port map( A1 => minus2A(15), A2 => n291, B1 => minusA(15), 
                           B2 => n285, ZN => n336);
   U183 : NAND2_X1 port map( A1 => n335, A2 => n334, ZN => n487);
   U184 : AOI22_X1 port map( A1 => plusA(14), A2 => n279, B1 => plus2A(14), B2 
                           => n273, ZN => n335);
   U185 : AOI22_X1 port map( A1 => minus2A(14), A2 => n291, B1 => minusA(14), 
                           B2 => n285, ZN => n334);
   U186 : NAND2_X1 port map( A1 => n333, A2 => n332, ZN => n488);
   U187 : AOI22_X1 port map( A1 => plusA(13), A2 => n279, B1 => plus2A(13), B2 
                           => n273, ZN => n333);
   U188 : AOI22_X1 port map( A1 => minus2A(13), A2 => n291, B1 => minusA(13), 
                           B2 => n285, ZN => n332);
   U189 : NAND2_X1 port map( A1 => n329, A2 => n328, ZN => n490);
   U190 : AOI22_X1 port map( A1 => plusA(11), A2 => n278, B1 => plus2A(11), B2 
                           => n272, ZN => n329);
   U191 : AOI22_X1 port map( A1 => minus2A(11), A2 => n290, B1 => minusA(11), 
                           B2 => n284, ZN => n328);
   U192 : NAND2_X1 port map( A1 => n327, A2 => n326, ZN => n491);
   U193 : AOI22_X1 port map( A1 => plusA(10), A2 => n278, B1 => plus2A(10), B2 
                           => n272, ZN => n327);
   U194 : AOI22_X1 port map( A1 => minus2A(10), A2 => n290, B1 => minusA(10), 
                           B2 => n284, ZN => n326);
   U195 : NAND2_X1 port map( A1 => n325, A2 => n324, ZN => n492);
   U196 : AOI22_X1 port map( A1 => plusA(9), A2 => n278, B1 => plus2A(9), B2 =>
                           n272, ZN => n325);
   U197 : AOI22_X1 port map( A1 => minus2A(9), A2 => n290, B1 => minusA(9), B2 
                           => n284, ZN => n324);
   U198 : NAND2_X1 port map( A1 => n320, A2 => n319, ZN => n495);
   U199 : AOI22_X1 port map( A1 => plusA(7), A2 => n278, B1 => plus2A(7), B2 =>
                           n272, ZN => n320);
   U200 : AOI22_X1 port map( A1 => minus2A(7), A2 => n290, B1 => minusA(7), B2 
                           => n284, ZN => n319);
   U201 : NAND2_X1 port map( A1 => n318, A2 => n317, ZN => n496);
   U202 : AOI22_X1 port map( A1 => plusA(6), A2 => n278, B1 => plus2A(6), B2 =>
                           n272, ZN => n318);
   U203 : AOI22_X1 port map( A1 => minus2A(6), A2 => n290, B1 => minusA(6), B2 
                           => n284, ZN => n317);
   U204 : NAND2_X1 port map( A1 => n316, A2 => n315, ZN => n497);
   U205 : AOI22_X1 port map( A1 => plusA(5), A2 => n278, B1 => plus2A(5), B2 =>
                           n272, ZN => n316);
   U206 : AOI22_X1 port map( A1 => minus2A(5), A2 => n290, B1 => minusA(5), B2 
                           => n284, ZN => n315);
   U207 : NAND2_X1 port map( A1 => n312, A2 => n311, ZN => n499);
   U208 : AOI22_X1 port map( A1 => plusA(3), A2 => n278, B1 => plus2A(3), B2 =>
                           n272, ZN => n312);
   U209 : AOI22_X1 port map( A1 => minus2A(3), A2 => n290, B1 => minusA(3), B2 
                           => n284, ZN => n311);
   U210 : NAND2_X1 port map( A1 => n331, A2 => n330, ZN => n489);
   U211 : AOI22_X1 port map( A1 => plusA(12), A2 => n279, B1 => plus2A(12), B2 
                           => n273, ZN => n331);
   U212 : AOI22_X1 port map( A1 => minus2A(12), A2 => n291, B1 => minusA(12), 
                           B2 => n285, ZN => n330);
   U213 : NAND2_X1 port map( A1 => n322, A2 => n321, ZN => n494);
   U214 : AOI22_X1 port map( A1 => plusA(8), A2 => n278, B1 => plus2A(8), B2 =>
                           n272, ZN => n322);
   U215 : AOI22_X1 port map( A1 => minus2A(8), A2 => n290, B1 => minusA(8), B2 
                           => n284, ZN => n321);
   U216 : NAND2_X1 port map( A1 => n314, A2 => n313, ZN => n498);
   U217 : AOI22_X1 port map( A1 => plusA(4), A2 => n278, B1 => plus2A(4), B2 =>
                           n272, ZN => n314);
   U218 : AOI22_X1 port map( A1 => minus2A(4), A2 => n290, B1 => minusA(4), B2 
                           => n284, ZN => n313);
   U219 : NAND2_X1 port map( A1 => n310, A2 => n309, ZN => n500);
   U220 : AOI22_X1 port map( A1 => plusA(2), A2 => n278, B1 => plus2A(2), B2 =>
                           n272, ZN => n310);
   U221 : AOI22_X1 port map( A1 => minus2A(2), A2 => n290, B1 => minusA(2), B2 
                           => n284, ZN => n309);
   U222 : NAND2_X1 port map( A1 => n308, A2 => n307, ZN => n501);
   U223 : AOI22_X1 port map( A1 => plusA(1), A2 => n278, B1 => plus2A(1), B2 =>
                           n272, ZN => n308);
   U224 : AOI22_X1 port map( A1 => minus2A(1), A2 => n290, B1 => minusA(1), B2 
                           => n284, ZN => n307);
   U225 : NAND2_X1 port map( A1 => n306, A2 => n305, ZN => n502);
   U226 : AOI22_X1 port map( A1 => plusA(0), A2 => n278, B1 => plus2A(0), B2 =>
                           n272, ZN => n306);
   U227 : AOI22_X1 port map( A1 => minus2A(0), A2 => n290, B1 => minusA(0), B2 
                           => n284, ZN => n305);
   U228 : CLKBUF_X1 port map( A => n432, Z => n277);
   U229 : CLKBUF_X1 port map( A => n433, Z => n283);
   U230 : CLKBUF_X1 port map( A => n434, Z => n289);
   U231 : CLKBUF_X1 port map( A => n435, Z => n295);
   U232 : CLKBUF_X1 port map( A => n493, Z => n301);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity MUX_GENERIC_N64_RADIX3_7 is

   port( plusA, minusA, plus2A, minus2A : in std_logic_vector (63 downto 0);  
         SEL : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (63 
         downto 0));

end MUX_GENERIC_N64_RADIX3_7;

architecture SYN_beh of MUX_GENERIC_N64_RADIX3_7 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component TBUF_X2
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   component TBUF_X1
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   signal n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, 
      n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, 
      n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, 
      n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, 
      n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, 
      n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, 
      n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, 
      n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, 
      n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, 
      n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, 
      n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, 
      n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, 
      n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, 
      n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, 
      n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, 
      n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, 
      n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, 
      n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, 
      n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, 
      n499, n500, n501, n502 : std_logic;

begin
   
   Y_tri_60_inst : TBUF_X1 port map( A => n441, EN => n301, Z => Y(60));
   Y_tri_61_inst : TBUF_X1 port map( A => n440, EN => n301, Z => Y(61));
   Y_tri_62_inst : TBUF_X1 port map( A => n439, EN => n301, Z => Y(62));
   Y_tri_63_inst : TBUF_X1 port map( A => n438, EN => n301, Z => Y(63));
   Y_tri_45_inst : TBUF_X1 port map( A => n456, EN => n299, Z => Y(45));
   Y_tri_46_inst : TBUF_X1 port map( A => n455, EN => n299, Z => Y(46));
   Y_tri_47_inst : TBUF_X1 port map( A => n454, EN => n299, Z => Y(47));
   Y_tri_48_inst : TBUF_X1 port map( A => n453, EN => n300, Z => Y(48));
   Y_tri_49_inst : TBUF_X1 port map( A => n452, EN => n300, Z => Y(49));
   Y_tri_50_inst : TBUF_X1 port map( A => n451, EN => n300, Z => Y(50));
   Y_tri_51_inst : TBUF_X1 port map( A => n450, EN => n300, Z => Y(51));
   Y_tri_52_inst : TBUF_X1 port map( A => n449, EN => n300, Z => Y(52));
   Y_tri_53_inst : TBUF_X1 port map( A => n448, EN => n300, Z => Y(53));
   Y_tri_55_inst : TBUF_X1 port map( A => n446, EN => n300, Z => Y(55));
   Y_tri_56_inst : TBUF_X1 port map( A => n445, EN => n300, Z => Y(56));
   Y_tri_57_inst : TBUF_X1 port map( A => n444, EN => n300, Z => Y(57));
   Y_tri_58_inst : TBUF_X1 port map( A => n443, EN => n300, Z => Y(58));
   Y_tri_59_inst : TBUF_X1 port map( A => n442, EN => n300, Z => Y(59));
   Y_tri_16_inst : TBUF_X1 port map( A => n485, EN => n297, Z => Y(16));
   Y_tri_17_inst : TBUF_X1 port map( A => n484, EN => n297, Z => Y(17));
   Y_tri_18_inst : TBUF_X1 port map( A => n483, EN => n297, Z => Y(18));
   Y_tri_19_inst : TBUF_X1 port map( A => n482, EN => n297, Z => Y(19));
   Y_tri_20_inst : TBUF_X1 port map( A => n481, EN => n297, Z => Y(20));
   Y_tri_21_inst : TBUF_X1 port map( A => n480, EN => n297, Z => Y(21));
   Y_tri_22_inst : TBUF_X1 port map( A => n479, EN => n297, Z => Y(22));
   Y_tri_24_inst : TBUF_X1 port map( A => n477, EN => n298, Z => Y(24));
   Y_tri_25_inst : TBUF_X1 port map( A => n476, EN => n298, Z => Y(25));
   Y_tri_26_inst : TBUF_X1 port map( A => n475, EN => n298, Z => Y(26));
   Y_tri_27_inst : TBUF_X1 port map( A => n474, EN => n298, Z => Y(27));
   Y_tri_28_inst : TBUF_X1 port map( A => n473, EN => n298, Z => Y(28));
   Y_tri_29_inst : TBUF_X1 port map( A => n472, EN => n298, Z => Y(29));
   Y_tri_30_inst : TBUF_X1 port map( A => n471, EN => n298, Z => Y(30));
   Y_tri_31_inst : TBUF_X1 port map( A => n470, EN => n298, Z => Y(31));
   Y_tri_32_inst : TBUF_X1 port map( A => n469, EN => n298, Z => Y(32));
   Y_tri_34_inst : TBUF_X1 port map( A => n467, EN => n298, Z => Y(34));
   Y_tri_35_inst : TBUF_X1 port map( A => n466, EN => n298, Z => Y(35));
   Y_tri_36_inst : TBUF_X1 port map( A => n465, EN => n299, Z => Y(36));
   Y_tri_38_inst : TBUF_X1 port map( A => n463, EN => n299, Z => Y(38));
   Y_tri_39_inst : TBUF_X1 port map( A => n462, EN => n299, Z => Y(39));
   Y_tri_40_inst : TBUF_X1 port map( A => n461, EN => n299, Z => Y(40));
   Y_tri_41_inst : TBUF_X1 port map( A => n460, EN => n299, Z => Y(41));
   Y_tri_42_inst : TBUF_X1 port map( A => n459, EN => n299, Z => Y(42));
   Y_tri_43_inst : TBUF_X1 port map( A => n458, EN => n299, Z => Y(43));
   Y_tri_44_inst : TBUF_X1 port map( A => n457, EN => n299, Z => Y(44));
   Y_tri_23_inst : TBUF_X1 port map( A => n478, EN => n297, Z => Y(23));
   Y_tri_33_inst : TBUF_X1 port map( A => n468, EN => n298, Z => Y(33));
   Y_tri_8_inst : TBUF_X1 port map( A => n494, EN => n296, Z => Y(8));
   Y_tri_9_inst : TBUF_X1 port map( A => n492, EN => n296, Z => Y(9));
   Y_tri_10_inst : TBUF_X1 port map( A => n491, EN => n296, Z => Y(10));
   Y_tri_11_inst : TBUF_X1 port map( A => n490, EN => n296, Z => Y(11));
   Y_tri_12_inst : TBUF_X1 port map( A => n489, EN => n297, Z => Y(12));
   Y_tri_13_inst : TBUF_X1 port map( A => n488, EN => n297, Z => Y(13));
   Y_tri_14_inst : TBUF_X1 port map( A => n487, EN => n297, Z => Y(14));
   Y_tri_15_inst : TBUF_X1 port map( A => n486, EN => n297, Z => Y(15));
   Y_tri_4_inst : TBUF_X1 port map( A => n498, EN => n296, Z => Y(4));
   Y_tri_3_inst : TBUF_X1 port map( A => n499, EN => n296, Z => Y(3));
   Y_tri_2_inst : TBUF_X1 port map( A => n500, EN => n296, Z => Y(2));
   Y_tri_1_inst : TBUF_X1 port map( A => n501, EN => n296, Z => Y(1));
   Y_tri_5_inst : TBUF_X1 port map( A => n497, EN => n296, Z => Y(5));
   Y_tri_6_inst : TBUF_X1 port map( A => n496, EN => n296, Z => Y(6));
   Y_tri_0_inst : TBUF_X1 port map( A => n502, EN => n296, Z => Y(0));
   Y_tri_54_inst : TBUF_X1 port map( A => n447, EN => n300, Z => Y(54));
   Y_tri_37_inst : TBUF_X1 port map( A => n464, EN => n299, Z => Y(37));
   Y_tri_7_inst : TBUF_X2 port map( A => n495, EN => n296, Z => Y(7));
   U2 : NOR3_X1 port map( A1 => SEL(0), A2 => SEL(2), A3 => n302, ZN => n434);
   U3 : NOR3_X1 port map( A1 => n302, A2 => SEL(2), A3 => n303, ZN => n432);
   U4 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n303, ZN => n433);
   U5 : BUF_X2 port map( A => n493, Z => n296);
   U6 : CLKBUF_X1 port map( A => n493, Z => n297);
   U7 : CLKBUF_X1 port map( A => n493, Z => n298);
   U8 : CLKBUF_X1 port map( A => n493, Z => n299);
   U9 : CLKBUF_X1 port map( A => n493, Z => n300);
   U10 : NAND2_X1 port map( A1 => n395, A2 => n394, ZN => n457);
   U11 : AOI22_X1 port map( A1 => plusA(44), A2 => n281, B1 => plus2A(44), B2 
                           => n275, ZN => n395);
   U12 : AOI22_X1 port map( A1 => minus2A(44), A2 => n293, B1 => minusA(44), B2
                           => n287, ZN => n394);
   U13 : NAND2_X1 port map( A1 => n393, A2 => n392, ZN => n458);
   U14 : AOI22_X1 port map( A1 => plusA(43), A2 => n281, B1 => plus2A(43), B2 
                           => n275, ZN => n393);
   U15 : AOI22_X1 port map( A1 => minus2A(43), A2 => n293, B1 => minusA(43), B2
                           => n287, ZN => n392);
   U16 : NAND2_X1 port map( A1 => n389, A2 => n388, ZN => n460);
   U17 : AOI22_X1 port map( A1 => plusA(41), A2 => n281, B1 => plus2A(41), B2 
                           => n275, ZN => n389);
   U18 : AOI22_X1 port map( A1 => minus2A(41), A2 => n293, B1 => minusA(41), B2
                           => n287, ZN => n388);
   U19 : NAND2_X1 port map( A1 => n381, A2 => n380, ZN => n464);
   U20 : AOI22_X1 port map( A1 => plusA(37), A2 => n281, B1 => plus2A(37), B2 
                           => n275, ZN => n381);
   U21 : AOI22_X1 port map( A1 => minus2A(37), A2 => n293, B1 => minusA(37), B2
                           => n287, ZN => n380);
   U22 : NAND2_X1 port map( A1 => n373, A2 => n372, ZN => n468);
   U23 : AOI22_X1 port map( A1 => plusA(33), A2 => n280, B1 => plus2A(33), B2 
                           => n274, ZN => n373);
   U24 : AOI22_X1 port map( A1 => minus2A(33), A2 => n292, B1 => minusA(33), B2
                           => n286, ZN => n372);
   U25 : NAND2_X1 port map( A1 => n365, A2 => n364, ZN => n472);
   U26 : AOI22_X1 port map( A1 => plusA(29), A2 => n280, B1 => plus2A(29), B2 
                           => n274, ZN => n365);
   U27 : AOI22_X1 port map( A1 => minus2A(29), A2 => n292, B1 => minusA(29), B2
                           => n286, ZN => n364);
   U28 : NAND2_X1 port map( A1 => n357, A2 => n356, ZN => n476);
   U29 : AOI22_X1 port map( A1 => plusA(25), A2 => n280, B1 => plus2A(25), B2 
                           => n274, ZN => n357);
   U30 : AOI22_X1 port map( A1 => minus2A(25), A2 => n292, B1 => minusA(25), B2
                           => n286, ZN => n356);
   U31 : NAND2_X1 port map( A1 => n385, A2 => n384, ZN => n462);
   U32 : AOI22_X1 port map( A1 => plusA(39), A2 => n281, B1 => plus2A(39), B2 
                           => n275, ZN => n385);
   U33 : AOI22_X1 port map( A1 => minus2A(39), A2 => n293, B1 => minusA(39), B2
                           => n287, ZN => n384);
   U34 : NAND2_X1 port map( A1 => n377, A2 => n376, ZN => n466);
   U35 : AOI22_X1 port map( A1 => plusA(35), A2 => n280, B1 => plus2A(35), B2 
                           => n274, ZN => n377);
   U36 : AOI22_X1 port map( A1 => minus2A(35), A2 => n292, B1 => minusA(35), B2
                           => n286, ZN => n376);
   U37 : NAND2_X1 port map( A1 => n369, A2 => n368, ZN => n470);
   U38 : AOI22_X1 port map( A1 => plusA(31), A2 => n280, B1 => plus2A(31), B2 
                           => n274, ZN => n369);
   U39 : AOI22_X1 port map( A1 => minus2A(31), A2 => n292, B1 => minusA(31), B2
                           => n286, ZN => n368);
   U40 : NAND2_X1 port map( A1 => n361, A2 => n360, ZN => n474);
   U41 : AOI22_X1 port map( A1 => plusA(27), A2 => n280, B1 => plus2A(27), B2 
                           => n274, ZN => n361);
   U42 : AOI22_X1 port map( A1 => minus2A(27), A2 => n292, B1 => minusA(27), B2
                           => n286, ZN => n360);
   U43 : NAND2_X1 port map( A1 => n353, A2 => n352, ZN => n478);
   U44 : AOI22_X1 port map( A1 => plusA(23), A2 => n279, B1 => plus2A(23), B2 
                           => n273, ZN => n353);
   U45 : AOI22_X1 port map( A1 => minus2A(23), A2 => n291, B1 => minusA(23), B2
                           => n285, ZN => n352);
   U46 : NAND2_X1 port map( A1 => n391, A2 => n390, ZN => n459);
   U47 : AOI22_X1 port map( A1 => plusA(42), A2 => n281, B1 => plus2A(42), B2 
                           => n275, ZN => n391);
   U48 : AOI22_X1 port map( A1 => minus2A(42), A2 => n293, B1 => minusA(42), B2
                           => n287, ZN => n390);
   U49 : NAND2_X1 port map( A1 => n383, A2 => n382, ZN => n463);
   U50 : AOI22_X1 port map( A1 => plusA(38), A2 => n281, B1 => plus2A(38), B2 
                           => n275, ZN => n383);
   U51 : AOI22_X1 port map( A1 => minus2A(38), A2 => n293, B1 => minusA(38), B2
                           => n287, ZN => n382);
   U52 : NAND2_X1 port map( A1 => n375, A2 => n374, ZN => n467);
   U53 : AOI22_X1 port map( A1 => plusA(34), A2 => n280, B1 => plus2A(34), B2 
                           => n274, ZN => n375);
   U54 : AOI22_X1 port map( A1 => minus2A(34), A2 => n292, B1 => minusA(34), B2
                           => n286, ZN => n374);
   U55 : NAND2_X1 port map( A1 => n367, A2 => n366, ZN => n471);
   U56 : AOI22_X1 port map( A1 => plusA(30), A2 => n280, B1 => plus2A(30), B2 
                           => n274, ZN => n367);
   U57 : AOI22_X1 port map( A1 => minus2A(30), A2 => n292, B1 => minusA(30), B2
                           => n286, ZN => n366);
   U58 : NAND2_X1 port map( A1 => n359, A2 => n358, ZN => n475);
   U59 : AOI22_X1 port map( A1 => plusA(26), A2 => n280, B1 => plus2A(26), B2 
                           => n274, ZN => n359);
   U60 : AOI22_X1 port map( A1 => minus2A(26), A2 => n292, B1 => minusA(26), B2
                           => n286, ZN => n358);
   U61 : NAND2_X1 port map( A1 => n351, A2 => n350, ZN => n479);
   U62 : AOI22_X1 port map( A1 => plusA(22), A2 => n279, B1 => plus2A(22), B2 
                           => n273, ZN => n351);
   U63 : AOI22_X1 port map( A1 => minus2A(22), A2 => n291, B1 => minusA(22), B2
                           => n285, ZN => n350);
   U64 : NAND2_X1 port map( A1 => n387, A2 => n386, ZN => n461);
   U65 : AOI22_X1 port map( A1 => plusA(40), A2 => n281, B1 => plus2A(40), B2 
                           => n275, ZN => n387);
   U66 : AOI22_X1 port map( A1 => minus2A(40), A2 => n293, B1 => minusA(40), B2
                           => n287, ZN => n386);
   U67 : NAND2_X1 port map( A1 => n379, A2 => n378, ZN => n465);
   U68 : AOI22_X1 port map( A1 => plusA(36), A2 => n281, B1 => plus2A(36), B2 
                           => n275, ZN => n379);
   U69 : AOI22_X1 port map( A1 => minus2A(36), A2 => n293, B1 => minusA(36), B2
                           => n287, ZN => n378);
   U70 : NAND2_X1 port map( A1 => n371, A2 => n370, ZN => n469);
   U71 : AOI22_X1 port map( A1 => plusA(32), A2 => n280, B1 => plus2A(32), B2 
                           => n274, ZN => n371);
   U72 : AOI22_X1 port map( A1 => minus2A(32), A2 => n292, B1 => minusA(32), B2
                           => n286, ZN => n370);
   U73 : NAND2_X1 port map( A1 => n363, A2 => n362, ZN => n473);
   U74 : AOI22_X1 port map( A1 => plusA(28), A2 => n280, B1 => plus2A(28), B2 
                           => n274, ZN => n363);
   U75 : AOI22_X1 port map( A1 => minus2A(28), A2 => n292, B1 => minusA(28), B2
                           => n286, ZN => n362);
   U76 : NAND2_X1 port map( A1 => n355, A2 => n354, ZN => n477);
   U77 : AOI22_X1 port map( A1 => plusA(24), A2 => n280, B1 => plus2A(24), B2 
                           => n274, ZN => n355);
   U78 : AOI22_X1 port map( A1 => minus2A(24), A2 => n292, B1 => minusA(24), B2
                           => n286, ZN => n354);
   U79 : NAND2_X1 port map( A1 => n437, A2 => n436, ZN => n438);
   U80 : AOI22_X1 port map( A1 => plusA(63), A2 => n283, B1 => plus2A(63), B2 
                           => n277, ZN => n437);
   U81 : AOI22_X1 port map( A1 => minus2A(63), A2 => n295, B1 => minusA(63), B2
                           => n289, ZN => n436);
   U82 : NAND2_X1 port map( A1 => n431, A2 => n430, ZN => n439);
   U83 : AOI22_X1 port map( A1 => plusA(62), A2 => n283, B1 => plus2A(62), B2 
                           => n277, ZN => n431);
   U84 : AOI22_X1 port map( A1 => minus2A(62), A2 => n295, B1 => minusA(62), B2
                           => n289, ZN => n430);
   U85 : NAND2_X1 port map( A1 => n429, A2 => n428, ZN => n440);
   U86 : AOI22_X1 port map( A1 => plusA(61), A2 => n283, B1 => plus2A(61), B2 
                           => n277, ZN => n429);
   U87 : AOI22_X1 port map( A1 => minus2A(61), A2 => n295, B1 => minusA(61), B2
                           => n289, ZN => n428);
   U88 : NAND2_X1 port map( A1 => n427, A2 => n426, ZN => n441);
   U89 : AOI22_X1 port map( A1 => plusA(60), A2 => n283, B1 => plus2A(60), B2 
                           => n277, ZN => n427);
   U90 : AOI22_X1 port map( A1 => minus2A(60), A2 => n295, B1 => minusA(60), B2
                           => n289, ZN => n426);
   U91 : NAND2_X1 port map( A1 => n425, A2 => n424, ZN => n442);
   U92 : AOI22_X1 port map( A1 => plusA(59), A2 => n282, B1 => plus2A(59), B2 
                           => n276, ZN => n425);
   U93 : AOI22_X1 port map( A1 => minus2A(59), A2 => n294, B1 => minusA(59), B2
                           => n288, ZN => n424);
   U94 : NAND2_X1 port map( A1 => n423, A2 => n422, ZN => n443);
   U95 : AOI22_X1 port map( A1 => plusA(58), A2 => n282, B1 => plus2A(58), B2 
                           => n276, ZN => n423);
   U96 : AOI22_X1 port map( A1 => minus2A(58), A2 => n294, B1 => minusA(58), B2
                           => n288, ZN => n422);
   U97 : NAND2_X1 port map( A1 => n421, A2 => n420, ZN => n444);
   U98 : AOI22_X1 port map( A1 => plusA(57), A2 => n282, B1 => plus2A(57), B2 
                           => n276, ZN => n421);
   U99 : AOI22_X1 port map( A1 => minus2A(57), A2 => n294, B1 => minusA(57), B2
                           => n288, ZN => n420);
   U100 : NAND2_X1 port map( A1 => n419, A2 => n418, ZN => n445);
   U101 : AOI22_X1 port map( A1 => plusA(56), A2 => n282, B1 => plus2A(56), B2 
                           => n276, ZN => n419);
   U102 : AOI22_X1 port map( A1 => minus2A(56), A2 => n294, B1 => minusA(56), 
                           B2 => n288, ZN => n418);
   U103 : NAND2_X1 port map( A1 => n417, A2 => n416, ZN => n446);
   U104 : AOI22_X1 port map( A1 => plusA(55), A2 => n282, B1 => plus2A(55), B2 
                           => n276, ZN => n417);
   U105 : AOI22_X1 port map( A1 => minus2A(55), A2 => n294, B1 => minusA(55), 
                           B2 => n288, ZN => n416);
   U106 : NAND2_X1 port map( A1 => n415, A2 => n414, ZN => n447);
   U107 : AOI22_X1 port map( A1 => plusA(54), A2 => n282, B1 => plus2A(54), B2 
                           => n276, ZN => n415);
   U108 : AOI22_X1 port map( A1 => minus2A(54), A2 => n294, B1 => minusA(54), 
                           B2 => n288, ZN => n414);
   U109 : NAND2_X1 port map( A1 => n413, A2 => n412, ZN => n448);
   U110 : AOI22_X1 port map( A1 => plusA(53), A2 => n282, B1 => plus2A(53), B2 
                           => n276, ZN => n413);
   U111 : AOI22_X1 port map( A1 => minus2A(53), A2 => n294, B1 => minusA(53), 
                           B2 => n288, ZN => n412);
   U112 : NAND2_X1 port map( A1 => n411, A2 => n410, ZN => n449);
   U113 : AOI22_X1 port map( A1 => plusA(52), A2 => n282, B1 => plus2A(52), B2 
                           => n276, ZN => n411);
   U114 : AOI22_X1 port map( A1 => minus2A(52), A2 => n294, B1 => minusA(52), 
                           B2 => n288, ZN => n410);
   U115 : NAND2_X1 port map( A1 => n409, A2 => n408, ZN => n450);
   U116 : AOI22_X1 port map( A1 => plusA(51), A2 => n282, B1 => plus2A(51), B2 
                           => n276, ZN => n409);
   U117 : AOI22_X1 port map( A1 => minus2A(51), A2 => n294, B1 => minusA(51), 
                           B2 => n288, ZN => n408);
   U118 : NAND2_X1 port map( A1 => n407, A2 => n406, ZN => n451);
   U119 : AOI22_X1 port map( A1 => plusA(50), A2 => n282, B1 => plus2A(50), B2 
                           => n276, ZN => n407);
   U120 : AOI22_X1 port map( A1 => minus2A(50), A2 => n294, B1 => minusA(50), 
                           B2 => n288, ZN => n406);
   U121 : NAND2_X1 port map( A1 => n405, A2 => n404, ZN => n452);
   U122 : AOI22_X1 port map( A1 => plusA(49), A2 => n282, B1 => plus2A(49), B2 
                           => n276, ZN => n405);
   U123 : AOI22_X1 port map( A1 => minus2A(49), A2 => n294, B1 => minusA(49), 
                           B2 => n288, ZN => n404);
   U124 : NAND2_X1 port map( A1 => n403, A2 => n402, ZN => n453);
   U125 : AOI22_X1 port map( A1 => plusA(48), A2 => n282, B1 => plus2A(48), B2 
                           => n276, ZN => n403);
   U126 : AOI22_X1 port map( A1 => minus2A(48), A2 => n294, B1 => minusA(48), 
                           B2 => n288, ZN => n402);
   U127 : NAND2_X1 port map( A1 => n401, A2 => n400, ZN => n454);
   U128 : AOI22_X1 port map( A1 => plusA(47), A2 => n281, B1 => plus2A(47), B2 
                           => n275, ZN => n401);
   U129 : AOI22_X1 port map( A1 => minus2A(47), A2 => n293, B1 => minusA(47), 
                           B2 => n287, ZN => n400);
   U130 : NAND2_X1 port map( A1 => n399, A2 => n398, ZN => n455);
   U131 : AOI22_X1 port map( A1 => plusA(46), A2 => n281, B1 => plus2A(46), B2 
                           => n275, ZN => n399);
   U132 : AOI22_X1 port map( A1 => minus2A(46), A2 => n293, B1 => minusA(46), 
                           B2 => n287, ZN => n398);
   U133 : NAND2_X1 port map( A1 => n397, A2 => n396, ZN => n456);
   U134 : AOI22_X1 port map( A1 => plusA(45), A2 => n281, B1 => plus2A(45), B2 
                           => n275, ZN => n397);
   U135 : AOI22_X1 port map( A1 => minus2A(45), A2 => n293, B1 => minusA(45), 
                           B2 => n287, ZN => n396);
   U136 : BUF_X1 port map( A => n433, Z => n280);
   U137 : BUF_X1 port map( A => n433, Z => n279);
   U138 : BUF_X1 port map( A => n434, Z => n286);
   U139 : BUF_X1 port map( A => n432, Z => n274);
   U140 : BUF_X1 port map( A => n434, Z => n285);
   U141 : BUF_X1 port map( A => n432, Z => n273);
   U142 : BUF_X1 port map( A => n435, Z => n292);
   U143 : BUF_X1 port map( A => n435, Z => n291);
   U144 : NAND2_X1 port map( A1 => n349, A2 => n348, ZN => n480);
   U145 : AOI22_X1 port map( A1 => plusA(21), A2 => n279, B1 => plus2A(21), B2 
                           => n273, ZN => n349);
   U146 : AOI22_X1 port map( A1 => minus2A(21), A2 => n291, B1 => minusA(21), 
                           B2 => n285, ZN => n348);
   U147 : NAND2_X1 port map( A1 => n347, A2 => n346, ZN => n481);
   U148 : AOI22_X1 port map( A1 => plusA(20), A2 => n279, B1 => plus2A(20), B2 
                           => n273, ZN => n347);
   U149 : AOI22_X1 port map( A1 => minus2A(20), A2 => n291, B1 => minusA(20), 
                           B2 => n285, ZN => n346);
   U150 : BUF_X1 port map( A => n433, Z => n281);
   U151 : BUF_X1 port map( A => n434, Z => n287);
   U152 : BUF_X1 port map( A => n432, Z => n275);
   U153 : BUF_X1 port map( A => n435, Z => n293);
   U154 : BUF_X1 port map( A => n433, Z => n282);
   U155 : BUF_X1 port map( A => n434, Z => n288);
   U156 : BUF_X1 port map( A => n432, Z => n276);
   U157 : BUF_X1 port map( A => n435, Z => n294);
   U158 : BUF_X1 port map( A => n433, Z => n278);
   U159 : BUF_X1 port map( A => n434, Z => n284);
   U160 : BUF_X1 port map( A => n432, Z => n272);
   U161 : BUF_X1 port map( A => n435, Z => n290);
   U162 : NOR2_X1 port map( A1 => n323, A2 => n304, ZN => n493);
   U163 : INV_X1 port map( A => SEL(2), ZN => n304);
   U164 : NOR2_X1 port map( A1 => SEL(1), A2 => SEL(0), ZN => n323);
   U165 : AND2_X1 port map( A1 => SEL(2), A2 => n323, ZN => n435);
   U166 : INV_X1 port map( A => SEL(1), ZN => n302);
   U167 : INV_X1 port map( A => SEL(0), ZN => n303);
   U168 : NAND2_X1 port map( A1 => n345, A2 => n344, ZN => n482);
   U169 : AOI22_X1 port map( A1 => plusA(19), A2 => n279, B1 => plus2A(19), B2 
                           => n273, ZN => n345);
   U170 : AOI22_X1 port map( A1 => minus2A(19), A2 => n291, B1 => minusA(19), 
                           B2 => n285, ZN => n344);
   U171 : NAND2_X1 port map( A1 => n343, A2 => n342, ZN => n483);
   U172 : AOI22_X1 port map( A1 => plusA(18), A2 => n279, B1 => plus2A(18), B2 
                           => n273, ZN => n343);
   U173 : AOI22_X1 port map( A1 => minus2A(18), A2 => n291, B1 => minusA(18), 
                           B2 => n285, ZN => n342);
   U174 : NAND2_X1 port map( A1 => n341, A2 => n340, ZN => n484);
   U175 : AOI22_X1 port map( A1 => plusA(17), A2 => n279, B1 => plus2A(17), B2 
                           => n273, ZN => n341);
   U176 : AOI22_X1 port map( A1 => minus2A(17), A2 => n291, B1 => minusA(17), 
                           B2 => n285, ZN => n340);
   U177 : NAND2_X1 port map( A1 => n337, A2 => n336, ZN => n486);
   U178 : AOI22_X1 port map( A1 => plusA(15), A2 => n279, B1 => plus2A(15), B2 
                           => n273, ZN => n337);
   U179 : AOI22_X1 port map( A1 => minus2A(15), A2 => n291, B1 => minusA(15), 
                           B2 => n285, ZN => n336);
   U180 : NAND2_X1 port map( A1 => n335, A2 => n334, ZN => n487);
   U181 : AOI22_X1 port map( A1 => plusA(14), A2 => n279, B1 => plus2A(14), B2 
                           => n273, ZN => n335);
   U182 : AOI22_X1 port map( A1 => minus2A(14), A2 => n291, B1 => minusA(14), 
                           B2 => n285, ZN => n334);
   U183 : NAND2_X1 port map( A1 => n333, A2 => n332, ZN => n488);
   U184 : AOI22_X1 port map( A1 => plusA(13), A2 => n279, B1 => plus2A(13), B2 
                           => n273, ZN => n333);
   U185 : AOI22_X1 port map( A1 => minus2A(13), A2 => n291, B1 => minusA(13), 
                           B2 => n285, ZN => n332);
   U186 : NAND2_X1 port map( A1 => n329, A2 => n328, ZN => n490);
   U187 : AOI22_X1 port map( A1 => plusA(11), A2 => n278, B1 => plus2A(11), B2 
                           => n272, ZN => n329);
   U188 : AOI22_X1 port map( A1 => minus2A(11), A2 => n290, B1 => minusA(11), 
                           B2 => n284, ZN => n328);
   U189 : NAND2_X1 port map( A1 => n327, A2 => n326, ZN => n491);
   U190 : AOI22_X1 port map( A1 => plusA(10), A2 => n278, B1 => plus2A(10), B2 
                           => n272, ZN => n327);
   U191 : AOI22_X1 port map( A1 => minus2A(10), A2 => n290, B1 => minusA(10), 
                           B2 => n284, ZN => n326);
   U192 : NAND2_X1 port map( A1 => n325, A2 => n324, ZN => n492);
   U193 : AOI22_X1 port map( A1 => plusA(9), A2 => n278, B1 => plus2A(9), B2 =>
                           n272, ZN => n325);
   U194 : AOI22_X1 port map( A1 => minus2A(9), A2 => n290, B1 => minusA(9), B2 
                           => n284, ZN => n324);
   U195 : NAND2_X1 port map( A1 => n320, A2 => n319, ZN => n495);
   U196 : AOI22_X1 port map( A1 => plusA(7), A2 => n278, B1 => plus2A(7), B2 =>
                           n272, ZN => n320);
   U197 : AOI22_X1 port map( A1 => minus2A(7), A2 => n290, B1 => minusA(7), B2 
                           => n284, ZN => n319);
   U198 : NAND2_X1 port map( A1 => n318, A2 => n317, ZN => n496);
   U199 : AOI22_X1 port map( A1 => plusA(6), A2 => n278, B1 => plus2A(6), B2 =>
                           n272, ZN => n318);
   U200 : AOI22_X1 port map( A1 => minus2A(6), A2 => n290, B1 => minusA(6), B2 
                           => n284, ZN => n317);
   U201 : NAND2_X1 port map( A1 => n316, A2 => n315, ZN => n497);
   U202 : AOI22_X1 port map( A1 => plusA(5), A2 => n278, B1 => plus2A(5), B2 =>
                           n272, ZN => n316);
   U203 : AOI22_X1 port map( A1 => minus2A(5), A2 => n290, B1 => minusA(5), B2 
                           => n284, ZN => n315);
   U204 : NAND2_X1 port map( A1 => n312, A2 => n311, ZN => n499);
   U205 : AOI22_X1 port map( A1 => plusA(3), A2 => n278, B1 => plus2A(3), B2 =>
                           n272, ZN => n312);
   U206 : AOI22_X1 port map( A1 => minus2A(3), A2 => n290, B1 => minusA(3), B2 
                           => n284, ZN => n311);
   U207 : NAND2_X1 port map( A1 => n339, A2 => n338, ZN => n485);
   U208 : AOI22_X1 port map( A1 => plusA(16), A2 => n279, B1 => plus2A(16), B2 
                           => n273, ZN => n339);
   U209 : AOI22_X1 port map( A1 => minus2A(16), A2 => n291, B1 => minusA(16), 
                           B2 => n285, ZN => n338);
   U210 : NAND2_X1 port map( A1 => n331, A2 => n330, ZN => n489);
   U211 : AOI22_X1 port map( A1 => plusA(12), A2 => n279, B1 => plus2A(12), B2 
                           => n273, ZN => n331);
   U212 : AOI22_X1 port map( A1 => minus2A(12), A2 => n291, B1 => minusA(12), 
                           B2 => n285, ZN => n330);
   U213 : NAND2_X1 port map( A1 => n322, A2 => n321, ZN => n494);
   U214 : AOI22_X1 port map( A1 => plusA(8), A2 => n278, B1 => plus2A(8), B2 =>
                           n272, ZN => n322);
   U215 : AOI22_X1 port map( A1 => minus2A(8), A2 => n290, B1 => minusA(8), B2 
                           => n284, ZN => n321);
   U216 : NAND2_X1 port map( A1 => n314, A2 => n313, ZN => n498);
   U217 : AOI22_X1 port map( A1 => plusA(4), A2 => n278, B1 => plus2A(4), B2 =>
                           n272, ZN => n314);
   U218 : AOI22_X1 port map( A1 => minus2A(4), A2 => n290, B1 => minusA(4), B2 
                           => n284, ZN => n313);
   U219 : NAND2_X1 port map( A1 => n310, A2 => n309, ZN => n500);
   U220 : AOI22_X1 port map( A1 => plusA(2), A2 => n278, B1 => plus2A(2), B2 =>
                           n272, ZN => n310);
   U221 : AOI22_X1 port map( A1 => minus2A(2), A2 => n290, B1 => minusA(2), B2 
                           => n284, ZN => n309);
   U222 : NAND2_X1 port map( A1 => n308, A2 => n307, ZN => n501);
   U223 : AOI22_X1 port map( A1 => plusA(1), A2 => n278, B1 => plus2A(1), B2 =>
                           n272, ZN => n308);
   U224 : AOI22_X1 port map( A1 => minus2A(1), A2 => n290, B1 => minusA(1), B2 
                           => n284, ZN => n307);
   U225 : NAND2_X1 port map( A1 => n306, A2 => n305, ZN => n502);
   U226 : AOI22_X1 port map( A1 => plusA(0), A2 => n278, B1 => plus2A(0), B2 =>
                           n272, ZN => n306);
   U227 : AOI22_X1 port map( A1 => minus2A(0), A2 => n290, B1 => minusA(0), B2 
                           => n284, ZN => n305);
   U228 : CLKBUF_X1 port map( A => n432, Z => n277);
   U229 : CLKBUF_X1 port map( A => n433, Z => n283);
   U230 : CLKBUF_X1 port map( A => n434, Z => n289);
   U231 : CLKBUF_X1 port map( A => n435, Z => n295);
   U232 : CLKBUF_X1 port map( A => n493, Z => n301);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity MUX_GENERIC_N64_RADIX3_6 is

   port( plusA, minusA, plus2A, minus2A : in std_logic_vector (63 downto 0);  
         SEL : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (63 
         downto 0));

end MUX_GENERIC_N64_RADIX3_6;

architecture SYN_beh of MUX_GENERIC_N64_RADIX3_6 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component TBUF_X2
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   component TBUF_X1
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   signal n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, 
      n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, 
      n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, 
      n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, 
      n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, 
      n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, 
      n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, 
      n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, 
      n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, 
      n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, 
      n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, 
      n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, 
      n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, 
      n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, 
      n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, 
      n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, 
      n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, 
      n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, 
      n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, 
      n499, n500, n501, n502 : std_logic;

begin
   
   Y_tri_60_inst : TBUF_X1 port map( A => n441, EN => n301, Z => Y(60));
   Y_tri_61_inst : TBUF_X1 port map( A => n440, EN => n301, Z => Y(61));
   Y_tri_62_inst : TBUF_X1 port map( A => n439, EN => n301, Z => Y(62));
   Y_tri_63_inst : TBUF_X1 port map( A => n438, EN => n301, Z => Y(63));
   Y_tri_38_inst : TBUF_X1 port map( A => n463, EN => n299, Z => Y(38));
   Y_tri_39_inst : TBUF_X1 port map( A => n462, EN => n299, Z => Y(39));
   Y_tri_42_inst : TBUF_X1 port map( A => n459, EN => n299, Z => Y(42));
   Y_tri_43_inst : TBUF_X1 port map( A => n458, EN => n299, Z => Y(43));
   Y_tri_44_inst : TBUF_X1 port map( A => n457, EN => n299, Z => Y(44));
   Y_tri_45_inst : TBUF_X1 port map( A => n456, EN => n299, Z => Y(45));
   Y_tri_46_inst : TBUF_X1 port map( A => n455, EN => n299, Z => Y(46));
   Y_tri_47_inst : TBUF_X1 port map( A => n454, EN => n299, Z => Y(47));
   Y_tri_48_inst : TBUF_X1 port map( A => n453, EN => n300, Z => Y(48));
   Y_tri_49_inst : TBUF_X1 port map( A => n452, EN => n300, Z => Y(49));
   Y_tri_51_inst : TBUF_X1 port map( A => n450, EN => n300, Z => Y(51));
   Y_tri_52_inst : TBUF_X1 port map( A => n449, EN => n300, Z => Y(52));
   Y_tri_53_inst : TBUF_X1 port map( A => n448, EN => n300, Z => Y(53));
   Y_tri_54_inst : TBUF_X1 port map( A => n447, EN => n300, Z => Y(54));
   Y_tri_55_inst : TBUF_X1 port map( A => n446, EN => n300, Z => Y(55));
   Y_tri_56_inst : TBUF_X1 port map( A => n445, EN => n300, Z => Y(56));
   Y_tri_57_inst : TBUF_X1 port map( A => n444, EN => n300, Z => Y(57));
   Y_tri_58_inst : TBUF_X1 port map( A => n443, EN => n300, Z => Y(58));
   Y_tri_59_inst : TBUF_X1 port map( A => n442, EN => n300, Z => Y(59));
   Y_tri_50_inst : TBUF_X1 port map( A => n451, EN => n300, Z => Y(50));
   Y_tri_14_inst : TBUF_X1 port map( A => n487, EN => n297, Z => Y(14));
   Y_tri_15_inst : TBUF_X1 port map( A => n486, EN => n297, Z => Y(15));
   Y_tri_16_inst : TBUF_X1 port map( A => n485, EN => n297, Z => Y(16));
   Y_tri_17_inst : TBUF_X1 port map( A => n484, EN => n297, Z => Y(17));
   Y_tri_18_inst : TBUF_X1 port map( A => n483, EN => n297, Z => Y(18));
   Y_tri_19_inst : TBUF_X1 port map( A => n482, EN => n297, Z => Y(19));
   Y_tri_21_inst : TBUF_X1 port map( A => n480, EN => n297, Z => Y(21));
   Y_tri_22_inst : TBUF_X1 port map( A => n479, EN => n297, Z => Y(22));
   Y_tri_23_inst : TBUF_X1 port map( A => n478, EN => n297, Z => Y(23));
   Y_tri_24_inst : TBUF_X1 port map( A => n477, EN => n298, Z => Y(24));
   Y_tri_25_inst : TBUF_X1 port map( A => n476, EN => n298, Z => Y(25));
   Y_tri_26_inst : TBUF_X1 port map( A => n475, EN => n298, Z => Y(26));
   Y_tri_27_inst : TBUF_X1 port map( A => n474, EN => n298, Z => Y(27));
   Y_tri_28_inst : TBUF_X1 port map( A => n473, EN => n298, Z => Y(28));
   Y_tri_29_inst : TBUF_X1 port map( A => n472, EN => n298, Z => Y(29));
   Y_tri_31_inst : TBUF_X1 port map( A => n470, EN => n298, Z => Y(31));
   Y_tri_32_inst : TBUF_X1 port map( A => n469, EN => n298, Z => Y(32));
   Y_tri_33_inst : TBUF_X1 port map( A => n468, EN => n298, Z => Y(33));
   Y_tri_34_inst : TBUF_X1 port map( A => n467, EN => n298, Z => Y(34));
   Y_tri_35_inst : TBUF_X1 port map( A => n466, EN => n298, Z => Y(35));
   Y_tri_36_inst : TBUF_X1 port map( A => n465, EN => n299, Z => Y(36));
   Y_tri_37_inst : TBUF_X1 port map( A => n464, EN => n299, Z => Y(37));
   Y_tri_20_inst : TBUF_X1 port map( A => n481, EN => n297, Z => Y(20));
   Y_tri_30_inst : TBUF_X1 port map( A => n471, EN => n298, Z => Y(30));
   Y_tri_6_inst : TBUF_X1 port map( A => n496, EN => n296, Z => Y(6));
   Y_tri_7_inst : TBUF_X1 port map( A => n495, EN => n296, Z => Y(7));
   Y_tri_8_inst : TBUF_X1 port map( A => n494, EN => n296, Z => Y(8));
   Y_tri_9_inst : TBUF_X1 port map( A => n492, EN => n296, Z => Y(9));
   Y_tri_10_inst : TBUF_X1 port map( A => n491, EN => n296, Z => Y(10));
   Y_tri_11_inst : TBUF_X1 port map( A => n490, EN => n296, Z => Y(11));
   Y_tri_12_inst : TBUF_X1 port map( A => n489, EN => n297, Z => Y(12));
   Y_tri_13_inst : TBUF_X1 port map( A => n488, EN => n297, Z => Y(13));
   Y_tri_2_inst : TBUF_X1 port map( A => n500, EN => n296, Z => Y(2));
   Y_tri_1_inst : TBUF_X1 port map( A => n501, EN => n296, Z => Y(1));
   Y_tri_3_inst : TBUF_X1 port map( A => n499, EN => n296, Z => Y(3));
   Y_tri_4_inst : TBUF_X1 port map( A => n498, EN => n296, Z => Y(4));
   Y_tri_0_inst : TBUF_X1 port map( A => n502, EN => n296, Z => Y(0));
   Y_tri_40_inst : TBUF_X1 port map( A => n461, EN => n299, Z => Y(40));
   Y_tri_41_inst : TBUF_X1 port map( A => n460, EN => n299, Z => Y(41));
   Y_tri_5_inst : TBUF_X2 port map( A => n497, EN => n296, Z => Y(5));
   U2 : NOR3_X1 port map( A1 => SEL(0), A2 => SEL(2), A3 => n302, ZN => n434);
   U3 : NOR3_X1 port map( A1 => n302, A2 => SEL(2), A3 => n303, ZN => n432);
   U4 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n303, ZN => n433);
   U5 : BUF_X1 port map( A => n493, Z => n296);
   U6 : CLKBUF_X1 port map( A => n493, Z => n297);
   U7 : CLKBUF_X1 port map( A => n493, Z => n298);
   U8 : CLKBUF_X1 port map( A => n493, Z => n299);
   U9 : CLKBUF_X1 port map( A => n493, Z => n300);
   U10 : NAND2_X1 port map( A1 => n377, A2 => n376, ZN => n466);
   U11 : AOI22_X1 port map( A1 => plusA(35), A2 => n280, B1 => plus2A(35), B2 
                           => n274, ZN => n377);
   U12 : AOI22_X1 port map( A1 => minus2A(35), A2 => n292, B1 => minusA(35), B2
                           => n286, ZN => n376);
   U13 : NAND2_X1 port map( A1 => n369, A2 => n368, ZN => n470);
   U14 : AOI22_X1 port map( A1 => plusA(31), A2 => n280, B1 => plus2A(31), B2 
                           => n274, ZN => n369);
   U15 : AOI22_X1 port map( A1 => minus2A(31), A2 => n292, B1 => minusA(31), B2
                           => n286, ZN => n368);
   U16 : NAND2_X1 port map( A1 => n361, A2 => n360, ZN => n474);
   U17 : AOI22_X1 port map( A1 => plusA(27), A2 => n280, B1 => plus2A(27), B2 
                           => n274, ZN => n361);
   U18 : AOI22_X1 port map( A1 => minus2A(27), A2 => n292, B1 => minusA(27), B2
                           => n286, ZN => n360);
   U19 : NAND2_X1 port map( A1 => n381, A2 => n380, ZN => n464);
   U20 : AOI22_X1 port map( A1 => plusA(37), A2 => n281, B1 => plus2A(37), B2 
                           => n275, ZN => n381);
   U21 : AOI22_X1 port map( A1 => minus2A(37), A2 => n293, B1 => minusA(37), B2
                           => n287, ZN => n380);
   U22 : NAND2_X1 port map( A1 => n373, A2 => n372, ZN => n468);
   U23 : AOI22_X1 port map( A1 => plusA(33), A2 => n280, B1 => plus2A(33), B2 
                           => n274, ZN => n373);
   U24 : AOI22_X1 port map( A1 => minus2A(33), A2 => n292, B1 => minusA(33), B2
                           => n286, ZN => n372);
   U25 : NAND2_X1 port map( A1 => n365, A2 => n364, ZN => n472);
   U26 : AOI22_X1 port map( A1 => plusA(29), A2 => n280, B1 => plus2A(29), B2 
                           => n274, ZN => n365);
   U27 : AOI22_X1 port map( A1 => minus2A(29), A2 => n292, B1 => minusA(29), B2
                           => n286, ZN => n364);
   U28 : NAND2_X1 port map( A1 => n357, A2 => n356, ZN => n476);
   U29 : AOI22_X1 port map( A1 => plusA(25), A2 => n280, B1 => plus2A(25), B2 
                           => n274, ZN => n357);
   U30 : AOI22_X1 port map( A1 => minus2A(25), A2 => n292, B1 => minusA(25), B2
                           => n286, ZN => n356);
   U31 : NAND2_X1 port map( A1 => n379, A2 => n378, ZN => n465);
   U32 : AOI22_X1 port map( A1 => plusA(36), A2 => n281, B1 => plus2A(36), B2 
                           => n275, ZN => n379);
   U33 : AOI22_X1 port map( A1 => minus2A(36), A2 => n293, B1 => minusA(36), B2
                           => n287, ZN => n378);
   U34 : NAND2_X1 port map( A1 => n371, A2 => n370, ZN => n469);
   U35 : AOI22_X1 port map( A1 => plusA(32), A2 => n280, B1 => plus2A(32), B2 
                           => n274, ZN => n371);
   U36 : AOI22_X1 port map( A1 => minus2A(32), A2 => n292, B1 => minusA(32), B2
                           => n286, ZN => n370);
   U37 : NAND2_X1 port map( A1 => n363, A2 => n362, ZN => n473);
   U38 : AOI22_X1 port map( A1 => plusA(28), A2 => n280, B1 => plus2A(28), B2 
                           => n274, ZN => n363);
   U39 : AOI22_X1 port map( A1 => minus2A(28), A2 => n292, B1 => minusA(28), B2
                           => n286, ZN => n362);
   U40 : NAND2_X1 port map( A1 => n355, A2 => n354, ZN => n477);
   U41 : AOI22_X1 port map( A1 => plusA(24), A2 => n280, B1 => plus2A(24), B2 
                           => n274, ZN => n355);
   U42 : AOI22_X1 port map( A1 => minus2A(24), A2 => n292, B1 => minusA(24), B2
                           => n286, ZN => n354);
   U43 : NAND2_X1 port map( A1 => n375, A2 => n374, ZN => n467);
   U44 : AOI22_X1 port map( A1 => plusA(34), A2 => n280, B1 => plus2A(34), B2 
                           => n274, ZN => n375);
   U45 : AOI22_X1 port map( A1 => minus2A(34), A2 => n292, B1 => minusA(34), B2
                           => n286, ZN => n374);
   U46 : NAND2_X1 port map( A1 => n367, A2 => n366, ZN => n471);
   U47 : AOI22_X1 port map( A1 => plusA(30), A2 => n280, B1 => plus2A(30), B2 
                           => n274, ZN => n367);
   U48 : AOI22_X1 port map( A1 => minus2A(30), A2 => n292, B1 => minusA(30), B2
                           => n286, ZN => n366);
   U49 : NAND2_X1 port map( A1 => n359, A2 => n358, ZN => n475);
   U50 : AOI22_X1 port map( A1 => plusA(26), A2 => n280, B1 => plus2A(26), B2 
                           => n274, ZN => n359);
   U51 : AOI22_X1 port map( A1 => minus2A(26), A2 => n292, B1 => minusA(26), B2
                           => n286, ZN => n358);
   U52 : NAND2_X1 port map( A1 => n437, A2 => n436, ZN => n438);
   U53 : AOI22_X1 port map( A1 => plusA(63), A2 => n283, B1 => plus2A(63), B2 
                           => n277, ZN => n437);
   U54 : AOI22_X1 port map( A1 => minus2A(63), A2 => n295, B1 => minusA(63), B2
                           => n289, ZN => n436);
   U55 : NAND2_X1 port map( A1 => n431, A2 => n430, ZN => n439);
   U56 : AOI22_X1 port map( A1 => plusA(62), A2 => n283, B1 => plus2A(62), B2 
                           => n277, ZN => n431);
   U57 : AOI22_X1 port map( A1 => minus2A(62), A2 => n295, B1 => minusA(62), B2
                           => n289, ZN => n430);
   U58 : NAND2_X1 port map( A1 => n429, A2 => n428, ZN => n440);
   U59 : AOI22_X1 port map( A1 => plusA(61), A2 => n283, B1 => plus2A(61), B2 
                           => n277, ZN => n429);
   U60 : AOI22_X1 port map( A1 => minus2A(61), A2 => n295, B1 => minusA(61), B2
                           => n289, ZN => n428);
   U61 : NAND2_X1 port map( A1 => n427, A2 => n426, ZN => n441);
   U62 : AOI22_X1 port map( A1 => plusA(60), A2 => n283, B1 => plus2A(60), B2 
                           => n277, ZN => n427);
   U63 : AOI22_X1 port map( A1 => minus2A(60), A2 => n295, B1 => minusA(60), B2
                           => n289, ZN => n426);
   U64 : NAND2_X1 port map( A1 => n425, A2 => n424, ZN => n442);
   U65 : AOI22_X1 port map( A1 => plusA(59), A2 => n282, B1 => plus2A(59), B2 
                           => n276, ZN => n425);
   U66 : AOI22_X1 port map( A1 => minus2A(59), A2 => n294, B1 => minusA(59), B2
                           => n288, ZN => n424);
   U67 : NAND2_X1 port map( A1 => n423, A2 => n422, ZN => n443);
   U68 : AOI22_X1 port map( A1 => plusA(58), A2 => n282, B1 => plus2A(58), B2 
                           => n276, ZN => n423);
   U69 : AOI22_X1 port map( A1 => minus2A(58), A2 => n294, B1 => minusA(58), B2
                           => n288, ZN => n422);
   U70 : NAND2_X1 port map( A1 => n421, A2 => n420, ZN => n444);
   U71 : AOI22_X1 port map( A1 => plusA(57), A2 => n282, B1 => plus2A(57), B2 
                           => n276, ZN => n421);
   U72 : AOI22_X1 port map( A1 => minus2A(57), A2 => n294, B1 => minusA(57), B2
                           => n288, ZN => n420);
   U73 : NAND2_X1 port map( A1 => n419, A2 => n418, ZN => n445);
   U74 : AOI22_X1 port map( A1 => plusA(56), A2 => n282, B1 => plus2A(56), B2 
                           => n276, ZN => n419);
   U75 : AOI22_X1 port map( A1 => minus2A(56), A2 => n294, B1 => minusA(56), B2
                           => n288, ZN => n418);
   U76 : NAND2_X1 port map( A1 => n417, A2 => n416, ZN => n446);
   U77 : AOI22_X1 port map( A1 => plusA(55), A2 => n282, B1 => plus2A(55), B2 
                           => n276, ZN => n417);
   U78 : AOI22_X1 port map( A1 => minus2A(55), A2 => n294, B1 => minusA(55), B2
                           => n288, ZN => n416);
   U79 : NAND2_X1 port map( A1 => n415, A2 => n414, ZN => n447);
   U80 : AOI22_X1 port map( A1 => plusA(54), A2 => n282, B1 => plus2A(54), B2 
                           => n276, ZN => n415);
   U81 : AOI22_X1 port map( A1 => minus2A(54), A2 => n294, B1 => minusA(54), B2
                           => n288, ZN => n414);
   U82 : NAND2_X1 port map( A1 => n413, A2 => n412, ZN => n448);
   U83 : AOI22_X1 port map( A1 => plusA(53), A2 => n282, B1 => plus2A(53), B2 
                           => n276, ZN => n413);
   U84 : AOI22_X1 port map( A1 => minus2A(53), A2 => n294, B1 => minusA(53), B2
                           => n288, ZN => n412);
   U85 : NAND2_X1 port map( A1 => n411, A2 => n410, ZN => n449);
   U86 : AOI22_X1 port map( A1 => plusA(52), A2 => n282, B1 => plus2A(52), B2 
                           => n276, ZN => n411);
   U87 : AOI22_X1 port map( A1 => minus2A(52), A2 => n294, B1 => minusA(52), B2
                           => n288, ZN => n410);
   U88 : NAND2_X1 port map( A1 => n409, A2 => n408, ZN => n450);
   U89 : AOI22_X1 port map( A1 => plusA(51), A2 => n282, B1 => plus2A(51), B2 
                           => n276, ZN => n409);
   U90 : AOI22_X1 port map( A1 => minus2A(51), A2 => n294, B1 => minusA(51), B2
                           => n288, ZN => n408);
   U91 : NAND2_X1 port map( A1 => n407, A2 => n406, ZN => n451);
   U92 : AOI22_X1 port map( A1 => plusA(50), A2 => n282, B1 => plus2A(50), B2 
                           => n276, ZN => n407);
   U93 : AOI22_X1 port map( A1 => minus2A(50), A2 => n294, B1 => minusA(50), B2
                           => n288, ZN => n406);
   U94 : NAND2_X1 port map( A1 => n405, A2 => n404, ZN => n452);
   U95 : AOI22_X1 port map( A1 => plusA(49), A2 => n282, B1 => plus2A(49), B2 
                           => n276, ZN => n405);
   U96 : AOI22_X1 port map( A1 => minus2A(49), A2 => n294, B1 => minusA(49), B2
                           => n288, ZN => n404);
   U97 : NAND2_X1 port map( A1 => n403, A2 => n402, ZN => n453);
   U98 : AOI22_X1 port map( A1 => plusA(48), A2 => n282, B1 => plus2A(48), B2 
                           => n276, ZN => n403);
   U99 : AOI22_X1 port map( A1 => minus2A(48), A2 => n294, B1 => minusA(48), B2
                           => n288, ZN => n402);
   U100 : NAND2_X1 port map( A1 => n401, A2 => n400, ZN => n454);
   U101 : AOI22_X1 port map( A1 => plusA(47), A2 => n281, B1 => plus2A(47), B2 
                           => n275, ZN => n401);
   U102 : AOI22_X1 port map( A1 => minus2A(47), A2 => n293, B1 => minusA(47), 
                           B2 => n287, ZN => n400);
   U103 : NAND2_X1 port map( A1 => n399, A2 => n398, ZN => n455);
   U104 : AOI22_X1 port map( A1 => plusA(46), A2 => n281, B1 => plus2A(46), B2 
                           => n275, ZN => n399);
   U105 : AOI22_X1 port map( A1 => minus2A(46), A2 => n293, B1 => minusA(46), 
                           B2 => n287, ZN => n398);
   U106 : NAND2_X1 port map( A1 => n397, A2 => n396, ZN => n456);
   U107 : AOI22_X1 port map( A1 => plusA(45), A2 => n281, B1 => plus2A(45), B2 
                           => n275, ZN => n397);
   U108 : AOI22_X1 port map( A1 => minus2A(45), A2 => n293, B1 => minusA(45), 
                           B2 => n287, ZN => n396);
   U109 : NAND2_X1 port map( A1 => n395, A2 => n394, ZN => n457);
   U110 : AOI22_X1 port map( A1 => plusA(44), A2 => n281, B1 => plus2A(44), B2 
                           => n275, ZN => n395);
   U111 : AOI22_X1 port map( A1 => minus2A(44), A2 => n293, B1 => minusA(44), 
                           B2 => n287, ZN => n394);
   U112 : NAND2_X1 port map( A1 => n391, A2 => n390, ZN => n459);
   U113 : AOI22_X1 port map( A1 => plusA(42), A2 => n281, B1 => plus2A(42), B2 
                           => n275, ZN => n391);
   U114 : AOI22_X1 port map( A1 => minus2A(42), A2 => n293, B1 => minusA(42), 
                           B2 => n287, ZN => n390);
   U115 : NAND2_X1 port map( A1 => n393, A2 => n392, ZN => n458);
   U116 : AOI22_X1 port map( A1 => plusA(43), A2 => n281, B1 => plus2A(43), B2 
                           => n275, ZN => n393);
   U117 : AOI22_X1 port map( A1 => minus2A(43), A2 => n293, B1 => minusA(43), 
                           B2 => n287, ZN => n392);
   U118 : NAND2_X1 port map( A1 => n385, A2 => n384, ZN => n462);
   U119 : AOI22_X1 port map( A1 => plusA(39), A2 => n281, B1 => plus2A(39), B2 
                           => n275, ZN => n385);
   U120 : AOI22_X1 port map( A1 => minus2A(39), A2 => n293, B1 => minusA(39), 
                           B2 => n287, ZN => n384);
   U121 : NAND2_X1 port map( A1 => n389, A2 => n388, ZN => n460);
   U122 : AOI22_X1 port map( A1 => plusA(41), A2 => n281, B1 => plus2A(41), B2 
                           => n275, ZN => n389);
   U123 : AOI22_X1 port map( A1 => minus2A(41), A2 => n293, B1 => minusA(41), 
                           B2 => n287, ZN => n388);
   U124 : NAND2_X1 port map( A1 => n387, A2 => n386, ZN => n461);
   U125 : AOI22_X1 port map( A1 => plusA(40), A2 => n281, B1 => plus2A(40), B2 
                           => n275, ZN => n387);
   U126 : AOI22_X1 port map( A1 => minus2A(40), A2 => n293, B1 => minusA(40), 
                           B2 => n287, ZN => n386);
   U127 : NAND2_X1 port map( A1 => n383, A2 => n382, ZN => n463);
   U128 : AOI22_X1 port map( A1 => plusA(38), A2 => n281, B1 => plus2A(38), B2 
                           => n275, ZN => n383);
   U129 : AOI22_X1 port map( A1 => minus2A(38), A2 => n293, B1 => minusA(38), 
                           B2 => n287, ZN => n382);
   U130 : BUF_X1 port map( A => n433, Z => n280);
   U131 : BUF_X1 port map( A => n433, Z => n279);
   U132 : BUF_X1 port map( A => n434, Z => n286);
   U133 : BUF_X1 port map( A => n432, Z => n274);
   U134 : BUF_X1 port map( A => n434, Z => n285);
   U135 : BUF_X1 port map( A => n432, Z => n273);
   U136 : BUF_X1 port map( A => n435, Z => n292);
   U137 : BUF_X1 port map( A => n435, Z => n291);
   U138 : NAND2_X1 port map( A1 => n353, A2 => n352, ZN => n478);
   U139 : AOI22_X1 port map( A1 => plusA(23), A2 => n279, B1 => plus2A(23), B2 
                           => n273, ZN => n353);
   U140 : AOI22_X1 port map( A1 => minus2A(23), A2 => n291, B1 => minusA(23), 
                           B2 => n285, ZN => n352);
   U141 : NAND2_X1 port map( A1 => n351, A2 => n350, ZN => n479);
   U142 : AOI22_X1 port map( A1 => plusA(22), A2 => n279, B1 => plus2A(22), B2 
                           => n273, ZN => n351);
   U143 : AOI22_X1 port map( A1 => minus2A(22), A2 => n291, B1 => minusA(22), 
                           B2 => n285, ZN => n350);
   U144 : BUF_X1 port map( A => n434, Z => n287);
   U145 : BUF_X1 port map( A => n433, Z => n281);
   U146 : BUF_X1 port map( A => n432, Z => n275);
   U147 : BUF_X1 port map( A => n435, Z => n293);
   U148 : BUF_X1 port map( A => n433, Z => n282);
   U149 : BUF_X1 port map( A => n434, Z => n288);
   U150 : BUF_X1 port map( A => n432, Z => n276);
   U151 : BUF_X1 port map( A => n435, Z => n294);
   U152 : BUF_X1 port map( A => n433, Z => n278);
   U153 : BUF_X1 port map( A => n434, Z => n284);
   U154 : BUF_X1 port map( A => n432, Z => n272);
   U155 : BUF_X1 port map( A => n435, Z => n290);
   U156 : NOR2_X1 port map( A1 => n323, A2 => n304, ZN => n493);
   U157 : INV_X1 port map( A => SEL(2), ZN => n304);
   U158 : NOR2_X1 port map( A1 => SEL(1), A2 => SEL(0), ZN => n323);
   U159 : AND2_X1 port map( A1 => SEL(2), A2 => n323, ZN => n435);
   U160 : INV_X1 port map( A => SEL(1), ZN => n302);
   U161 : INV_X1 port map( A => SEL(0), ZN => n303);
   U162 : NAND2_X1 port map( A1 => n349, A2 => n348, ZN => n480);
   U163 : AOI22_X1 port map( A1 => plusA(21), A2 => n279, B1 => plus2A(21), B2 
                           => n273, ZN => n349);
   U164 : AOI22_X1 port map( A1 => minus2A(21), A2 => n291, B1 => minusA(21), 
                           B2 => n285, ZN => n348);
   U165 : NAND2_X1 port map( A1 => n347, A2 => n346, ZN => n481);
   U166 : AOI22_X1 port map( A1 => plusA(20), A2 => n279, B1 => plus2A(20), B2 
                           => n273, ZN => n347);
   U167 : AOI22_X1 port map( A1 => minus2A(20), A2 => n291, B1 => minusA(20), 
                           B2 => n285, ZN => n346);
   U168 : NAND2_X1 port map( A1 => n345, A2 => n344, ZN => n482);
   U169 : AOI22_X1 port map( A1 => plusA(19), A2 => n279, B1 => plus2A(19), B2 
                           => n273, ZN => n345);
   U170 : AOI22_X1 port map( A1 => minus2A(19), A2 => n291, B1 => minusA(19), 
                           B2 => n285, ZN => n344);
   U171 : NAND2_X1 port map( A1 => n343, A2 => n342, ZN => n483);
   U172 : AOI22_X1 port map( A1 => plusA(18), A2 => n279, B1 => plus2A(18), B2 
                           => n273, ZN => n343);
   U173 : AOI22_X1 port map( A1 => minus2A(18), A2 => n291, B1 => minusA(18), 
                           B2 => n285, ZN => n342);
   U174 : NAND2_X1 port map( A1 => n341, A2 => n340, ZN => n484);
   U175 : AOI22_X1 port map( A1 => plusA(17), A2 => n279, B1 => plus2A(17), B2 
                           => n273, ZN => n341);
   U176 : AOI22_X1 port map( A1 => minus2A(17), A2 => n291, B1 => minusA(17), 
                           B2 => n285, ZN => n340);
   U177 : NAND2_X1 port map( A1 => n337, A2 => n336, ZN => n486);
   U178 : AOI22_X1 port map( A1 => plusA(15), A2 => n279, B1 => plus2A(15), B2 
                           => n273, ZN => n337);
   U179 : AOI22_X1 port map( A1 => minus2A(15), A2 => n291, B1 => minusA(15), 
                           B2 => n285, ZN => n336);
   U180 : NAND2_X1 port map( A1 => n335, A2 => n334, ZN => n487);
   U181 : AOI22_X1 port map( A1 => plusA(14), A2 => n279, B1 => plus2A(14), B2 
                           => n273, ZN => n335);
   U182 : AOI22_X1 port map( A1 => minus2A(14), A2 => n291, B1 => minusA(14), 
                           B2 => n285, ZN => n334);
   U183 : NAND2_X1 port map( A1 => n333, A2 => n332, ZN => n488);
   U184 : AOI22_X1 port map( A1 => plusA(13), A2 => n279, B1 => plus2A(13), B2 
                           => n273, ZN => n333);
   U185 : AOI22_X1 port map( A1 => minus2A(13), A2 => n291, B1 => minusA(13), 
                           B2 => n285, ZN => n332);
   U186 : NAND2_X1 port map( A1 => n329, A2 => n328, ZN => n490);
   U187 : AOI22_X1 port map( A1 => plusA(11), A2 => n278, B1 => plus2A(11), B2 
                           => n272, ZN => n329);
   U188 : AOI22_X1 port map( A1 => minus2A(11), A2 => n290, B1 => minusA(11), 
                           B2 => n284, ZN => n328);
   U189 : NAND2_X1 port map( A1 => n327, A2 => n326, ZN => n491);
   U190 : AOI22_X1 port map( A1 => plusA(10), A2 => n278, B1 => plus2A(10), B2 
                           => n272, ZN => n327);
   U191 : AOI22_X1 port map( A1 => minus2A(10), A2 => n290, B1 => minusA(10), 
                           B2 => n284, ZN => n326);
   U192 : NAND2_X1 port map( A1 => n325, A2 => n324, ZN => n492);
   U193 : AOI22_X1 port map( A1 => plusA(9), A2 => n278, B1 => plus2A(9), B2 =>
                           n272, ZN => n325);
   U194 : AOI22_X1 port map( A1 => minus2A(9), A2 => n290, B1 => minusA(9), B2 
                           => n284, ZN => n324);
   U195 : NAND2_X1 port map( A1 => n320, A2 => n319, ZN => n495);
   U196 : AOI22_X1 port map( A1 => plusA(7), A2 => n278, B1 => plus2A(7), B2 =>
                           n272, ZN => n320);
   U197 : AOI22_X1 port map( A1 => minus2A(7), A2 => n290, B1 => minusA(7), B2 
                           => n284, ZN => n319);
   U198 : NAND2_X1 port map( A1 => n318, A2 => n317, ZN => n496);
   U199 : AOI22_X1 port map( A1 => plusA(6), A2 => n278, B1 => plus2A(6), B2 =>
                           n272, ZN => n318);
   U200 : AOI22_X1 port map( A1 => minus2A(6), A2 => n290, B1 => minusA(6), B2 
                           => n284, ZN => n317);
   U201 : NAND2_X1 port map( A1 => n316, A2 => n315, ZN => n497);
   U202 : AOI22_X1 port map( A1 => plusA(5), A2 => n278, B1 => plus2A(5), B2 =>
                           n272, ZN => n316);
   U203 : AOI22_X1 port map( A1 => minus2A(5), A2 => n290, B1 => minusA(5), B2 
                           => n284, ZN => n315);
   U204 : NAND2_X1 port map( A1 => n312, A2 => n311, ZN => n499);
   U205 : AOI22_X1 port map( A1 => plusA(3), A2 => n278, B1 => plus2A(3), B2 =>
                           n272, ZN => n312);
   U206 : AOI22_X1 port map( A1 => minus2A(3), A2 => n290, B1 => minusA(3), B2 
                           => n284, ZN => n311);
   U207 : NAND2_X1 port map( A1 => n339, A2 => n338, ZN => n485);
   U208 : AOI22_X1 port map( A1 => plusA(16), A2 => n279, B1 => plus2A(16), B2 
                           => n273, ZN => n339);
   U209 : AOI22_X1 port map( A1 => minus2A(16), A2 => n291, B1 => minusA(16), 
                           B2 => n285, ZN => n338);
   U210 : NAND2_X1 port map( A1 => n331, A2 => n330, ZN => n489);
   U211 : AOI22_X1 port map( A1 => plusA(12), A2 => n279, B1 => plus2A(12), B2 
                           => n273, ZN => n331);
   U212 : AOI22_X1 port map( A1 => minus2A(12), A2 => n291, B1 => minusA(12), 
                           B2 => n285, ZN => n330);
   U213 : NAND2_X1 port map( A1 => n322, A2 => n321, ZN => n494);
   U214 : AOI22_X1 port map( A1 => plusA(8), A2 => n278, B1 => plus2A(8), B2 =>
                           n272, ZN => n322);
   U215 : AOI22_X1 port map( A1 => minus2A(8), A2 => n290, B1 => minusA(8), B2 
                           => n284, ZN => n321);
   U216 : NAND2_X1 port map( A1 => n314, A2 => n313, ZN => n498);
   U217 : AOI22_X1 port map( A1 => plusA(4), A2 => n278, B1 => plus2A(4), B2 =>
                           n272, ZN => n314);
   U218 : AOI22_X1 port map( A1 => minus2A(4), A2 => n290, B1 => minusA(4), B2 
                           => n284, ZN => n313);
   U219 : NAND2_X1 port map( A1 => n310, A2 => n309, ZN => n500);
   U220 : AOI22_X1 port map( A1 => plusA(2), A2 => n278, B1 => plus2A(2), B2 =>
                           n272, ZN => n310);
   U221 : AOI22_X1 port map( A1 => minus2A(2), A2 => n290, B1 => minusA(2), B2 
                           => n284, ZN => n309);
   U222 : NAND2_X1 port map( A1 => n308, A2 => n307, ZN => n501);
   U223 : AOI22_X1 port map( A1 => plusA(1), A2 => n278, B1 => plus2A(1), B2 =>
                           n272, ZN => n308);
   U224 : AOI22_X1 port map( A1 => minus2A(1), A2 => n290, B1 => minusA(1), B2 
                           => n284, ZN => n307);
   U225 : NAND2_X1 port map( A1 => n306, A2 => n305, ZN => n502);
   U226 : AOI22_X1 port map( A1 => plusA(0), A2 => n278, B1 => plus2A(0), B2 =>
                           n272, ZN => n306);
   U227 : AOI22_X1 port map( A1 => minus2A(0), A2 => n290, B1 => minusA(0), B2 
                           => n284, ZN => n305);
   U228 : CLKBUF_X1 port map( A => n432, Z => n277);
   U229 : CLKBUF_X1 port map( A => n433, Z => n283);
   U230 : CLKBUF_X1 port map( A => n434, Z => n289);
   U231 : CLKBUF_X1 port map( A => n435, Z => n295);
   U232 : CLKBUF_X1 port map( A => n493, Z => n301);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity MUX_GENERIC_N64_RADIX3_5 is

   port( plusA, minusA, plus2A, minus2A : in std_logic_vector (63 downto 0);  
         SEL : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (63 
         downto 0));

end MUX_GENERIC_N64_RADIX3_5;

architecture SYN_beh of MUX_GENERIC_N64_RADIX3_5 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component TBUF_X1
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   signal n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, 
      n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, 
      n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, 
      n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, 
      n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, 
      n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, 
      n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, 
      n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, 
      n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, 
      n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, 
      n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, 
      n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, 
      n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, 
      n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, 
      n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, 
      n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, 
      n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, 
      n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, 
      n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, 
      n499, n500, n501, n502 : std_logic;

begin
   
   Y_tri_60_inst : TBUF_X1 port map( A => n441, EN => n301, Z => Y(60));
   Y_tri_61_inst : TBUF_X1 port map( A => n440, EN => n301, Z => Y(61));
   Y_tri_62_inst : TBUF_X1 port map( A => n439, EN => n301, Z => Y(62));
   Y_tri_63_inst : TBUF_X1 port map( A => n438, EN => n301, Z => Y(63));
   Y_tri_34_inst : TBUF_X1 port map( A => n467, EN => n298, Z => Y(34));
   Y_tri_35_inst : TBUF_X1 port map( A => n466, EN => n298, Z => Y(35));
   Y_tri_36_inst : TBUF_X1 port map( A => n465, EN => n299, Z => Y(36));
   Y_tri_37_inst : TBUF_X1 port map( A => n464, EN => n299, Z => Y(37));
   Y_tri_38_inst : TBUF_X1 port map( A => n463, EN => n299, Z => Y(38));
   Y_tri_39_inst : TBUF_X1 port map( A => n462, EN => n299, Z => Y(39));
   Y_tri_40_inst : TBUF_X1 port map( A => n461, EN => n299, Z => Y(40));
   Y_tri_41_inst : TBUF_X1 port map( A => n460, EN => n299, Z => Y(41));
   Y_tri_42_inst : TBUF_X1 port map( A => n459, EN => n299, Z => Y(42));
   Y_tri_43_inst : TBUF_X1 port map( A => n458, EN => n299, Z => Y(43));
   Y_tri_44_inst : TBUF_X1 port map( A => n457, EN => n299, Z => Y(44));
   Y_tri_45_inst : TBUF_X1 port map( A => n456, EN => n299, Z => Y(45));
   Y_tri_46_inst : TBUF_X1 port map( A => n455, EN => n299, Z => Y(46));
   Y_tri_47_inst : TBUF_X1 port map( A => n454, EN => n299, Z => Y(47));
   Y_tri_48_inst : TBUF_X1 port map( A => n453, EN => n300, Z => Y(48));
   Y_tri_49_inst : TBUF_X1 port map( A => n452, EN => n300, Z => Y(49));
   Y_tri_50_inst : TBUF_X1 port map( A => n451, EN => n300, Z => Y(50));
   Y_tri_51_inst : TBUF_X1 port map( A => n450, EN => n300, Z => Y(51));
   Y_tri_52_inst : TBUF_X1 port map( A => n449, EN => n300, Z => Y(52));
   Y_tri_53_inst : TBUF_X1 port map( A => n448, EN => n300, Z => Y(53));
   Y_tri_54_inst : TBUF_X1 port map( A => n447, EN => n300, Z => Y(54));
   Y_tri_55_inst : TBUF_X1 port map( A => n446, EN => n300, Z => Y(55));
   Y_tri_56_inst : TBUF_X1 port map( A => n445, EN => n300, Z => Y(56));
   Y_tri_57_inst : TBUF_X1 port map( A => n444, EN => n300, Z => Y(57));
   Y_tri_58_inst : TBUF_X1 port map( A => n443, EN => n300, Z => Y(58));
   Y_tri_59_inst : TBUF_X1 port map( A => n442, EN => n300, Z => Y(59));
   Y_tri_12_inst : TBUF_X1 port map( A => n489, EN => n297, Z => Y(12));
   Y_tri_13_inst : TBUF_X1 port map( A => n488, EN => n297, Z => Y(13));
   Y_tri_14_inst : TBUF_X1 port map( A => n487, EN => n297, Z => Y(14));
   Y_tri_15_inst : TBUF_X1 port map( A => n486, EN => n297, Z => Y(15));
   Y_tri_16_inst : TBUF_X1 port map( A => n485, EN => n297, Z => Y(16));
   Y_tri_17_inst : TBUF_X1 port map( A => n484, EN => n297, Z => Y(17));
   Y_tri_18_inst : TBUF_X1 port map( A => n483, EN => n297, Z => Y(18));
   Y_tri_19_inst : TBUF_X1 port map( A => n482, EN => n297, Z => Y(19));
   Y_tri_20_inst : TBUF_X1 port map( A => n481, EN => n297, Z => Y(20));
   Y_tri_21_inst : TBUF_X1 port map( A => n480, EN => n297, Z => Y(21));
   Y_tri_22_inst : TBUF_X1 port map( A => n479, EN => n297, Z => Y(22));
   Y_tri_23_inst : TBUF_X1 port map( A => n478, EN => n297, Z => Y(23));
   Y_tri_24_inst : TBUF_X1 port map( A => n477, EN => n298, Z => Y(24));
   Y_tri_25_inst : TBUF_X1 port map( A => n476, EN => n298, Z => Y(25));
   Y_tri_26_inst : TBUF_X1 port map( A => n475, EN => n298, Z => Y(26));
   Y_tri_27_inst : TBUF_X1 port map( A => n474, EN => n298, Z => Y(27));
   Y_tri_28_inst : TBUF_X1 port map( A => n473, EN => n298, Z => Y(28));
   Y_tri_29_inst : TBUF_X1 port map( A => n472, EN => n298, Z => Y(29));
   Y_tri_30_inst : TBUF_X1 port map( A => n471, EN => n298, Z => Y(30));
   Y_tri_31_inst : TBUF_X1 port map( A => n470, EN => n298, Z => Y(31));
   Y_tri_32_inst : TBUF_X1 port map( A => n469, EN => n298, Z => Y(32));
   Y_tri_33_inst : TBUF_X1 port map( A => n468, EN => n298, Z => Y(33));
   Y_tri_3_inst : TBUF_X1 port map( A => n499, EN => n296, Z => Y(3));
   Y_tri_5_inst : TBUF_X1 port map( A => n497, EN => n296, Z => Y(5));
   Y_tri_6_inst : TBUF_X1 port map( A => n496, EN => n296, Z => Y(6));
   Y_tri_7_inst : TBUF_X1 port map( A => n495, EN => n296, Z => Y(7));
   Y_tri_8_inst : TBUF_X1 port map( A => n494, EN => n296, Z => Y(8));
   Y_tri_9_inst : TBUF_X1 port map( A => n492, EN => n296, Z => Y(9));
   Y_tri_10_inst : TBUF_X1 port map( A => n491, EN => n296, Z => Y(10));
   Y_tri_11_inst : TBUF_X1 port map( A => n490, EN => n296, Z => Y(11));
   Y_tri_2_inst : TBUF_X1 port map( A => n500, EN => n296, Z => Y(2));
   Y_tri_1_inst : TBUF_X1 port map( A => n501, EN => n296, Z => Y(1));
   Y_tri_0_inst : TBUF_X1 port map( A => n502, EN => n296, Z => Y(0));
   Y_tri_4_inst : TBUF_X1 port map( A => n498, EN => n296, Z => Y(4));
   U2 : NOR3_X1 port map( A1 => SEL(0), A2 => SEL(2), A3 => n302, ZN => n434);
   U3 : NOR3_X1 port map( A1 => n302, A2 => SEL(2), A3 => n303, ZN => n432);
   U4 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n303, ZN => n433);
   U5 : NAND2_X1 port map( A1 => n371, A2 => n370, ZN => n469);
   U6 : AOI22_X1 port map( A1 => plusA(32), A2 => n280, B1 => plus2A(32), B2 =>
                           n274, ZN => n371);
   U7 : AOI22_X1 port map( A1 => minus2A(32), A2 => n292, B1 => minusA(32), B2 
                           => n286, ZN => n370);
   U8 : NAND2_X1 port map( A1 => n363, A2 => n362, ZN => n473);
   U9 : AOI22_X1 port map( A1 => plusA(28), A2 => n280, B1 => plus2A(28), B2 =>
                           n274, ZN => n363);
   U10 : AOI22_X1 port map( A1 => minus2A(28), A2 => n292, B1 => minusA(28), B2
                           => n286, ZN => n362);
   U11 : NAND2_X1 port map( A1 => n367, A2 => n366, ZN => n471);
   U12 : AOI22_X1 port map( A1 => plusA(30), A2 => n280, B1 => plus2A(30), B2 
                           => n274, ZN => n367);
   U13 : AOI22_X1 port map( A1 => minus2A(30), A2 => n292, B1 => minusA(30), B2
                           => n286, ZN => n366);
   U14 : NAND2_X1 port map( A1 => n359, A2 => n358, ZN => n475);
   U15 : AOI22_X1 port map( A1 => plusA(26), A2 => n280, B1 => plus2A(26), B2 
                           => n274, ZN => n359);
   U16 : AOI22_X1 port map( A1 => minus2A(26), A2 => n292, B1 => minusA(26), B2
                           => n286, ZN => n358);
   U17 : NAND2_X1 port map( A1 => n373, A2 => n372, ZN => n468);
   U18 : AOI22_X1 port map( A1 => plusA(33), A2 => n280, B1 => plus2A(33), B2 
                           => n274, ZN => n373);
   U19 : AOI22_X1 port map( A1 => minus2A(33), A2 => n292, B1 => minusA(33), B2
                           => n286, ZN => n372);
   U20 : NAND2_X1 port map( A1 => n365, A2 => n364, ZN => n472);
   U21 : AOI22_X1 port map( A1 => plusA(29), A2 => n280, B1 => plus2A(29), B2 
                           => n274, ZN => n365);
   U22 : AOI22_X1 port map( A1 => minus2A(29), A2 => n292, B1 => minusA(29), B2
                           => n286, ZN => n364);
   U23 : NAND2_X1 port map( A1 => n369, A2 => n368, ZN => n470);
   U24 : AOI22_X1 port map( A1 => plusA(31), A2 => n280, B1 => plus2A(31), B2 
                           => n274, ZN => n369);
   U25 : AOI22_X1 port map( A1 => minus2A(31), A2 => n292, B1 => minusA(31), B2
                           => n286, ZN => n368);
   U26 : NAND2_X1 port map( A1 => n361, A2 => n360, ZN => n474);
   U27 : AOI22_X1 port map( A1 => plusA(27), A2 => n280, B1 => plus2A(27), B2 
                           => n274, ZN => n361);
   U28 : AOI22_X1 port map( A1 => minus2A(27), A2 => n292, B1 => minusA(27), B2
                           => n286, ZN => n360);
   U29 : NAND2_X1 port map( A1 => n425, A2 => n424, ZN => n442);
   U30 : AOI22_X1 port map( A1 => plusA(59), A2 => n282, B1 => plus2A(59), B2 
                           => n276, ZN => n425);
   U31 : AOI22_X1 port map( A1 => minus2A(59), A2 => n294, B1 => minusA(59), B2
                           => n288, ZN => n424);
   U32 : NAND2_X1 port map( A1 => n423, A2 => n422, ZN => n443);
   U33 : AOI22_X1 port map( A1 => plusA(58), A2 => n282, B1 => plus2A(58), B2 
                           => n276, ZN => n423);
   U34 : AOI22_X1 port map( A1 => minus2A(58), A2 => n294, B1 => minusA(58), B2
                           => n288, ZN => n422);
   U35 : NAND2_X1 port map( A1 => n421, A2 => n420, ZN => n444);
   U36 : AOI22_X1 port map( A1 => plusA(57), A2 => n282, B1 => plus2A(57), B2 
                           => n276, ZN => n421);
   U37 : AOI22_X1 port map( A1 => minus2A(57), A2 => n294, B1 => minusA(57), B2
                           => n288, ZN => n420);
   U38 : NAND2_X1 port map( A1 => n419, A2 => n418, ZN => n445);
   U39 : AOI22_X1 port map( A1 => plusA(56), A2 => n282, B1 => plus2A(56), B2 
                           => n276, ZN => n419);
   U40 : AOI22_X1 port map( A1 => minus2A(56), A2 => n294, B1 => minusA(56), B2
                           => n288, ZN => n418);
   U41 : NAND2_X1 port map( A1 => n417, A2 => n416, ZN => n446);
   U42 : AOI22_X1 port map( A1 => plusA(55), A2 => n282, B1 => plus2A(55), B2 
                           => n276, ZN => n417);
   U43 : AOI22_X1 port map( A1 => minus2A(55), A2 => n294, B1 => minusA(55), B2
                           => n288, ZN => n416);
   U44 : NAND2_X1 port map( A1 => n415, A2 => n414, ZN => n447);
   U45 : AOI22_X1 port map( A1 => plusA(54), A2 => n282, B1 => plus2A(54), B2 
                           => n276, ZN => n415);
   U46 : AOI22_X1 port map( A1 => minus2A(54), A2 => n294, B1 => minusA(54), B2
                           => n288, ZN => n414);
   U47 : NAND2_X1 port map( A1 => n413, A2 => n412, ZN => n448);
   U48 : AOI22_X1 port map( A1 => plusA(53), A2 => n282, B1 => plus2A(53), B2 
                           => n276, ZN => n413);
   U49 : AOI22_X1 port map( A1 => minus2A(53), A2 => n294, B1 => minusA(53), B2
                           => n288, ZN => n412);
   U50 : NAND2_X1 port map( A1 => n411, A2 => n410, ZN => n449);
   U51 : AOI22_X1 port map( A1 => plusA(52), A2 => n282, B1 => plus2A(52), B2 
                           => n276, ZN => n411);
   U52 : AOI22_X1 port map( A1 => minus2A(52), A2 => n294, B1 => minusA(52), B2
                           => n288, ZN => n410);
   U53 : NAND2_X1 port map( A1 => n409, A2 => n408, ZN => n450);
   U54 : AOI22_X1 port map( A1 => plusA(51), A2 => n282, B1 => plus2A(51), B2 
                           => n276, ZN => n409);
   U55 : AOI22_X1 port map( A1 => minus2A(51), A2 => n294, B1 => minusA(51), B2
                           => n288, ZN => n408);
   U56 : NAND2_X1 port map( A1 => n407, A2 => n406, ZN => n451);
   U57 : AOI22_X1 port map( A1 => plusA(50), A2 => n282, B1 => plus2A(50), B2 
                           => n276, ZN => n407);
   U58 : AOI22_X1 port map( A1 => minus2A(50), A2 => n294, B1 => minusA(50), B2
                           => n288, ZN => n406);
   U59 : NAND2_X1 port map( A1 => n405, A2 => n404, ZN => n452);
   U60 : AOI22_X1 port map( A1 => plusA(49), A2 => n282, B1 => plus2A(49), B2 
                           => n276, ZN => n405);
   U61 : AOI22_X1 port map( A1 => minus2A(49), A2 => n294, B1 => minusA(49), B2
                           => n288, ZN => n404);
   U62 : NAND2_X1 port map( A1 => n403, A2 => n402, ZN => n453);
   U63 : AOI22_X1 port map( A1 => plusA(48), A2 => n282, B1 => plus2A(48), B2 
                           => n276, ZN => n403);
   U64 : AOI22_X1 port map( A1 => minus2A(48), A2 => n294, B1 => minusA(48), B2
                           => n288, ZN => n402);
   U65 : NAND2_X1 port map( A1 => n401, A2 => n400, ZN => n454);
   U66 : AOI22_X1 port map( A1 => plusA(47), A2 => n281, B1 => plus2A(47), B2 
                           => n275, ZN => n401);
   U67 : AOI22_X1 port map( A1 => minus2A(47), A2 => n293, B1 => minusA(47), B2
                           => n287, ZN => n400);
   U68 : NAND2_X1 port map( A1 => n399, A2 => n398, ZN => n455);
   U69 : AOI22_X1 port map( A1 => plusA(46), A2 => n281, B1 => plus2A(46), B2 
                           => n275, ZN => n399);
   U70 : AOI22_X1 port map( A1 => minus2A(46), A2 => n293, B1 => minusA(46), B2
                           => n287, ZN => n398);
   U71 : NAND2_X1 port map( A1 => n397, A2 => n396, ZN => n456);
   U72 : AOI22_X1 port map( A1 => plusA(45), A2 => n281, B1 => plus2A(45), B2 
                           => n275, ZN => n397);
   U73 : AOI22_X1 port map( A1 => minus2A(45), A2 => n293, B1 => minusA(45), B2
                           => n287, ZN => n396);
   U74 : NAND2_X1 port map( A1 => n395, A2 => n394, ZN => n457);
   U75 : AOI22_X1 port map( A1 => plusA(44), A2 => n281, B1 => plus2A(44), B2 
                           => n275, ZN => n395);
   U76 : AOI22_X1 port map( A1 => minus2A(44), A2 => n293, B1 => minusA(44), B2
                           => n287, ZN => n394);
   U77 : NAND2_X1 port map( A1 => n387, A2 => n386, ZN => n461);
   U78 : AOI22_X1 port map( A1 => plusA(40), A2 => n281, B1 => plus2A(40), B2 
                           => n275, ZN => n387);
   U79 : AOI22_X1 port map( A1 => minus2A(40), A2 => n293, B1 => minusA(40), B2
                           => n287, ZN => n386);
   U80 : NAND2_X1 port map( A1 => n379, A2 => n378, ZN => n465);
   U81 : AOI22_X1 port map( A1 => plusA(36), A2 => n281, B1 => plus2A(36), B2 
                           => n275, ZN => n379);
   U82 : AOI22_X1 port map( A1 => minus2A(36), A2 => n293, B1 => minusA(36), B2
                           => n287, ZN => n378);
   U83 : NAND2_X1 port map( A1 => n391, A2 => n390, ZN => n459);
   U84 : AOI22_X1 port map( A1 => plusA(42), A2 => n281, B1 => plus2A(42), B2 
                           => n275, ZN => n391);
   U85 : AOI22_X1 port map( A1 => minus2A(42), A2 => n293, B1 => minusA(42), B2
                           => n287, ZN => n390);
   U86 : NAND2_X1 port map( A1 => n383, A2 => n382, ZN => n463);
   U87 : AOI22_X1 port map( A1 => plusA(38), A2 => n281, B1 => plus2A(38), B2 
                           => n275, ZN => n383);
   U88 : AOI22_X1 port map( A1 => minus2A(38), A2 => n293, B1 => minusA(38), B2
                           => n287, ZN => n382);
   U89 : NAND2_X1 port map( A1 => n375, A2 => n374, ZN => n467);
   U90 : AOI22_X1 port map( A1 => plusA(34), A2 => n280, B1 => plus2A(34), B2 
                           => n274, ZN => n375);
   U91 : AOI22_X1 port map( A1 => minus2A(34), A2 => n292, B1 => minusA(34), B2
                           => n286, ZN => n374);
   U92 : NAND2_X1 port map( A1 => n389, A2 => n388, ZN => n460);
   U93 : AOI22_X1 port map( A1 => plusA(41), A2 => n281, B1 => plus2A(41), B2 
                           => n275, ZN => n389);
   U94 : AOI22_X1 port map( A1 => minus2A(41), A2 => n293, B1 => minusA(41), B2
                           => n287, ZN => n388);
   U95 : NAND2_X1 port map( A1 => n381, A2 => n380, ZN => n464);
   U96 : AOI22_X1 port map( A1 => plusA(37), A2 => n281, B1 => plus2A(37), B2 
                           => n275, ZN => n381);
   U97 : AOI22_X1 port map( A1 => minus2A(37), A2 => n293, B1 => minusA(37), B2
                           => n287, ZN => n380);
   U98 : NAND2_X1 port map( A1 => n393, A2 => n392, ZN => n458);
   U99 : AOI22_X1 port map( A1 => plusA(43), A2 => n281, B1 => plus2A(43), B2 
                           => n275, ZN => n393);
   U100 : AOI22_X1 port map( A1 => minus2A(43), A2 => n293, B1 => minusA(43), 
                           B2 => n287, ZN => n392);
   U101 : NAND2_X1 port map( A1 => n385, A2 => n384, ZN => n462);
   U102 : AOI22_X1 port map( A1 => plusA(39), A2 => n281, B1 => plus2A(39), B2 
                           => n275, ZN => n385);
   U103 : AOI22_X1 port map( A1 => minus2A(39), A2 => n293, B1 => minusA(39), 
                           B2 => n287, ZN => n384);
   U104 : NAND2_X1 port map( A1 => n377, A2 => n376, ZN => n466);
   U105 : AOI22_X1 port map( A1 => plusA(35), A2 => n280, B1 => plus2A(35), B2 
                           => n274, ZN => n377);
   U106 : AOI22_X1 port map( A1 => minus2A(35), A2 => n292, B1 => minusA(35), 
                           B2 => n286, ZN => n376);
   U107 : NAND2_X1 port map( A1 => n437, A2 => n436, ZN => n438);
   U108 : AOI22_X1 port map( A1 => plusA(63), A2 => n283, B1 => plus2A(63), B2 
                           => n277, ZN => n437);
   U109 : AOI22_X1 port map( A1 => minus2A(63), A2 => n295, B1 => minusA(63), 
                           B2 => n289, ZN => n436);
   U110 : NAND2_X1 port map( A1 => n431, A2 => n430, ZN => n439);
   U111 : AOI22_X1 port map( A1 => plusA(62), A2 => n283, B1 => plus2A(62), B2 
                           => n277, ZN => n431);
   U112 : AOI22_X1 port map( A1 => minus2A(62), A2 => n295, B1 => minusA(62), 
                           B2 => n289, ZN => n430);
   U113 : NAND2_X1 port map( A1 => n429, A2 => n428, ZN => n440);
   U114 : AOI22_X1 port map( A1 => plusA(61), A2 => n283, B1 => plus2A(61), B2 
                           => n277, ZN => n429);
   U115 : AOI22_X1 port map( A1 => minus2A(61), A2 => n295, B1 => minusA(61), 
                           B2 => n289, ZN => n428);
   U116 : NAND2_X1 port map( A1 => n427, A2 => n426, ZN => n441);
   U117 : AOI22_X1 port map( A1 => plusA(60), A2 => n283, B1 => plus2A(60), B2 
                           => n277, ZN => n427);
   U118 : AOI22_X1 port map( A1 => minus2A(60), A2 => n295, B1 => minusA(60), 
                           B2 => n289, ZN => n426);
   U119 : BUF_X1 port map( A => n493, Z => n296);
   U120 : BUF_X1 port map( A => n493, Z => n297);
   U121 : BUF_X1 port map( A => n433, Z => n279);
   U122 : BUF_X1 port map( A => n434, Z => n285);
   U123 : NAND2_X1 port map( A1 => n355, A2 => n354, ZN => n477);
   U124 : AOI22_X1 port map( A1 => plusA(24), A2 => n280, B1 => plus2A(24), B2 
                           => n274, ZN => n355);
   U125 : AOI22_X1 port map( A1 => minus2A(24), A2 => n292, B1 => minusA(24), 
                           B2 => n286, ZN => n354);
   U126 : NAND2_X1 port map( A1 => n357, A2 => n356, ZN => n476);
   U127 : AOI22_X1 port map( A1 => plusA(25), A2 => n280, B1 => plus2A(25), B2 
                           => n274, ZN => n357);
   U128 : AOI22_X1 port map( A1 => minus2A(25), A2 => n292, B1 => minusA(25), 
                           B2 => n286, ZN => n356);
   U129 : BUF_X1 port map( A => n493, Z => n298);
   U130 : BUF_X1 port map( A => n433, Z => n280);
   U131 : BUF_X1 port map( A => n434, Z => n286);
   U132 : BUF_X1 port map( A => n432, Z => n274);
   U133 : BUF_X1 port map( A => n432, Z => n273);
   U134 : BUF_X1 port map( A => n435, Z => n292);
   U135 : BUF_X1 port map( A => n435, Z => n291);
   U136 : BUF_X1 port map( A => n493, Z => n299);
   U137 : BUF_X1 port map( A => n433, Z => n281);
   U138 : BUF_X1 port map( A => n434, Z => n287);
   U139 : BUF_X1 port map( A => n432, Z => n275);
   U140 : BUF_X1 port map( A => n435, Z => n293);
   U141 : BUF_X1 port map( A => n493, Z => n300);
   U142 : BUF_X1 port map( A => n433, Z => n282);
   U143 : BUF_X1 port map( A => n434, Z => n288);
   U144 : BUF_X1 port map( A => n432, Z => n276);
   U145 : BUF_X1 port map( A => n435, Z => n294);
   U146 : BUF_X1 port map( A => n433, Z => n278);
   U147 : BUF_X1 port map( A => n434, Z => n284);
   U148 : BUF_X1 port map( A => n432, Z => n272);
   U149 : BUF_X1 port map( A => n435, Z => n290);
   U150 : NOR2_X1 port map( A1 => n323, A2 => n304, ZN => n493);
   U151 : INV_X1 port map( A => SEL(2), ZN => n304);
   U152 : NOR2_X1 port map( A1 => SEL(1), A2 => SEL(0), ZN => n323);
   U153 : INV_X1 port map( A => SEL(1), ZN => n302);
   U154 : INV_X1 port map( A => SEL(0), ZN => n303);
   U155 : NAND2_X1 port map( A1 => n353, A2 => n352, ZN => n478);
   U156 : AOI22_X1 port map( A1 => plusA(23), A2 => n279, B1 => plus2A(23), B2 
                           => n273, ZN => n353);
   U157 : AOI22_X1 port map( A1 => minus2A(23), A2 => n291, B1 => minusA(23), 
                           B2 => n285, ZN => n352);
   U158 : AND2_X1 port map( A1 => SEL(2), A2 => n323, ZN => n435);
   U159 : NAND2_X1 port map( A1 => n351, A2 => n350, ZN => n479);
   U160 : AOI22_X1 port map( A1 => plusA(22), A2 => n279, B1 => plus2A(22), B2 
                           => n273, ZN => n351);
   U161 : AOI22_X1 port map( A1 => minus2A(22), A2 => n291, B1 => minusA(22), 
                           B2 => n285, ZN => n350);
   U162 : NAND2_X1 port map( A1 => n349, A2 => n348, ZN => n480);
   U163 : AOI22_X1 port map( A1 => plusA(21), A2 => n279, B1 => plus2A(21), B2 
                           => n273, ZN => n349);
   U164 : AOI22_X1 port map( A1 => minus2A(21), A2 => n291, B1 => minusA(21), 
                           B2 => n285, ZN => n348);
   U165 : NAND2_X1 port map( A1 => n345, A2 => n344, ZN => n482);
   U166 : AOI22_X1 port map( A1 => plusA(19), A2 => n279, B1 => plus2A(19), B2 
                           => n273, ZN => n345);
   U167 : AOI22_X1 port map( A1 => minus2A(19), A2 => n291, B1 => minusA(19), 
                           B2 => n285, ZN => n344);
   U168 : NAND2_X1 port map( A1 => n343, A2 => n342, ZN => n483);
   U169 : AOI22_X1 port map( A1 => plusA(18), A2 => n279, B1 => plus2A(18), B2 
                           => n273, ZN => n343);
   U170 : AOI22_X1 port map( A1 => minus2A(18), A2 => n291, B1 => minusA(18), 
                           B2 => n285, ZN => n342);
   U171 : NAND2_X1 port map( A1 => n341, A2 => n340, ZN => n484);
   U172 : AOI22_X1 port map( A1 => plusA(17), A2 => n279, B1 => plus2A(17), B2 
                           => n273, ZN => n341);
   U173 : AOI22_X1 port map( A1 => minus2A(17), A2 => n291, B1 => minusA(17), 
                           B2 => n285, ZN => n340);
   U174 : NAND2_X1 port map( A1 => n337, A2 => n336, ZN => n486);
   U175 : AOI22_X1 port map( A1 => plusA(15), A2 => n279, B1 => plus2A(15), B2 
                           => n273, ZN => n337);
   U176 : AOI22_X1 port map( A1 => minus2A(15), A2 => n291, B1 => minusA(15), 
                           B2 => n285, ZN => n336);
   U177 : NAND2_X1 port map( A1 => n335, A2 => n334, ZN => n487);
   U178 : AOI22_X1 port map( A1 => plusA(14), A2 => n279, B1 => plus2A(14), B2 
                           => n273, ZN => n335);
   U179 : AOI22_X1 port map( A1 => minus2A(14), A2 => n291, B1 => minusA(14), 
                           B2 => n285, ZN => n334);
   U180 : NAND2_X1 port map( A1 => n333, A2 => n332, ZN => n488);
   U181 : AOI22_X1 port map( A1 => plusA(13), A2 => n279, B1 => plus2A(13), B2 
                           => n273, ZN => n333);
   U182 : AOI22_X1 port map( A1 => minus2A(13), A2 => n291, B1 => minusA(13), 
                           B2 => n285, ZN => n332);
   U183 : NAND2_X1 port map( A1 => n329, A2 => n328, ZN => n490);
   U184 : AOI22_X1 port map( A1 => plusA(11), A2 => n278, B1 => plus2A(11), B2 
                           => n272, ZN => n329);
   U185 : AOI22_X1 port map( A1 => minus2A(11), A2 => n290, B1 => minusA(11), 
                           B2 => n284, ZN => n328);
   U186 : NAND2_X1 port map( A1 => n327, A2 => n326, ZN => n491);
   U187 : AOI22_X1 port map( A1 => plusA(10), A2 => n278, B1 => plus2A(10), B2 
                           => n272, ZN => n327);
   U188 : AOI22_X1 port map( A1 => minus2A(10), A2 => n290, B1 => minusA(10), 
                           B2 => n284, ZN => n326);
   U189 : NAND2_X1 port map( A1 => n325, A2 => n324, ZN => n492);
   U190 : AOI22_X1 port map( A1 => plusA(9), A2 => n278, B1 => plus2A(9), B2 =>
                           n272, ZN => n325);
   U191 : AOI22_X1 port map( A1 => minus2A(9), A2 => n290, B1 => minusA(9), B2 
                           => n284, ZN => n324);
   U192 : NAND2_X1 port map( A1 => n320, A2 => n319, ZN => n495);
   U193 : AOI22_X1 port map( A1 => plusA(7), A2 => n278, B1 => plus2A(7), B2 =>
                           n272, ZN => n320);
   U194 : AOI22_X1 port map( A1 => minus2A(7), A2 => n290, B1 => minusA(7), B2 
                           => n284, ZN => n319);
   U195 : NAND2_X1 port map( A1 => n318, A2 => n317, ZN => n496);
   U196 : AOI22_X1 port map( A1 => plusA(6), A2 => n278, B1 => plus2A(6), B2 =>
                           n272, ZN => n318);
   U197 : AOI22_X1 port map( A1 => minus2A(6), A2 => n290, B1 => minusA(6), B2 
                           => n284, ZN => n317);
   U198 : NAND2_X1 port map( A1 => n316, A2 => n315, ZN => n497);
   U199 : AOI22_X1 port map( A1 => plusA(5), A2 => n278, B1 => plus2A(5), B2 =>
                           n272, ZN => n316);
   U200 : AOI22_X1 port map( A1 => minus2A(5), A2 => n290, B1 => minusA(5), B2 
                           => n284, ZN => n315);
   U201 : NAND2_X1 port map( A1 => n312, A2 => n311, ZN => n499);
   U202 : AOI22_X1 port map( A1 => plusA(3), A2 => n278, B1 => plus2A(3), B2 =>
                           n272, ZN => n312);
   U203 : AOI22_X1 port map( A1 => minus2A(3), A2 => n290, B1 => minusA(3), B2 
                           => n284, ZN => n311);
   U204 : NAND2_X1 port map( A1 => n347, A2 => n346, ZN => n481);
   U205 : AOI22_X1 port map( A1 => plusA(20), A2 => n279, B1 => plus2A(20), B2 
                           => n273, ZN => n347);
   U206 : AOI22_X1 port map( A1 => minus2A(20), A2 => n291, B1 => minusA(20), 
                           B2 => n285, ZN => n346);
   U207 : NAND2_X1 port map( A1 => n339, A2 => n338, ZN => n485);
   U208 : AOI22_X1 port map( A1 => plusA(16), A2 => n279, B1 => plus2A(16), B2 
                           => n273, ZN => n339);
   U209 : AOI22_X1 port map( A1 => minus2A(16), A2 => n291, B1 => minusA(16), 
                           B2 => n285, ZN => n338);
   U210 : NAND2_X1 port map( A1 => n331, A2 => n330, ZN => n489);
   U211 : AOI22_X1 port map( A1 => plusA(12), A2 => n279, B1 => plus2A(12), B2 
                           => n273, ZN => n331);
   U212 : AOI22_X1 port map( A1 => minus2A(12), A2 => n291, B1 => minusA(12), 
                           B2 => n285, ZN => n330);
   U213 : NAND2_X1 port map( A1 => n322, A2 => n321, ZN => n494);
   U214 : AOI22_X1 port map( A1 => plusA(8), A2 => n278, B1 => plus2A(8), B2 =>
                           n272, ZN => n322);
   U215 : AOI22_X1 port map( A1 => minus2A(8), A2 => n290, B1 => minusA(8), B2 
                           => n284, ZN => n321);
   U216 : NAND2_X1 port map( A1 => n314, A2 => n313, ZN => n498);
   U217 : AOI22_X1 port map( A1 => plusA(4), A2 => n278, B1 => plus2A(4), B2 =>
                           n272, ZN => n314);
   U218 : AOI22_X1 port map( A1 => minus2A(4), A2 => n290, B1 => minusA(4), B2 
                           => n284, ZN => n313);
   U219 : NAND2_X1 port map( A1 => n310, A2 => n309, ZN => n500);
   U220 : AOI22_X1 port map( A1 => plusA(2), A2 => n278, B1 => plus2A(2), B2 =>
                           n272, ZN => n310);
   U221 : AOI22_X1 port map( A1 => minus2A(2), A2 => n290, B1 => minusA(2), B2 
                           => n284, ZN => n309);
   U222 : NAND2_X1 port map( A1 => n308, A2 => n307, ZN => n501);
   U223 : AOI22_X1 port map( A1 => plusA(1), A2 => n278, B1 => plus2A(1), B2 =>
                           n272, ZN => n308);
   U224 : AOI22_X1 port map( A1 => minus2A(1), A2 => n290, B1 => minusA(1), B2 
                           => n284, ZN => n307);
   U225 : NAND2_X1 port map( A1 => n306, A2 => n305, ZN => n502);
   U226 : AOI22_X1 port map( A1 => plusA(0), A2 => n278, B1 => plus2A(0), B2 =>
                           n272, ZN => n306);
   U227 : AOI22_X1 port map( A1 => minus2A(0), A2 => n290, B1 => minusA(0), B2 
                           => n284, ZN => n305);
   U228 : CLKBUF_X1 port map( A => n432, Z => n277);
   U229 : CLKBUF_X1 port map( A => n433, Z => n283);
   U230 : CLKBUF_X1 port map( A => n434, Z => n289);
   U231 : CLKBUF_X1 port map( A => n435, Z => n295);
   U232 : CLKBUF_X1 port map( A => n493, Z => n301);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity MUX_GENERIC_N64_RADIX3_4 is

   port( plusA, minusA, plus2A, minus2A : in std_logic_vector (63 downto 0);  
         SEL : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (63 
         downto 0));

end MUX_GENERIC_N64_RADIX3_4;

architecture SYN_beh of MUX_GENERIC_N64_RADIX3_4 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component TBUF_X1
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   signal n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, 
      n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, 
      n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, 
      n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, 
      n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, 
      n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, 
      n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, 
      n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, 
      n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, 
      n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, 
      n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, 
      n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, 
      n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, 
      n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, 
      n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, 
      n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, 
      n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, 
      n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, 
      n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, 
      n499, n500, n501, n502 : std_logic;

begin
   
   Y_tri_60_inst : TBUF_X1 port map( A => n441, EN => n301, Z => Y(60));
   Y_tri_61_inst : TBUF_X1 port map( A => n440, EN => n301, Z => Y(61));
   Y_tri_62_inst : TBUF_X1 port map( A => n439, EN => n301, Z => Y(62));
   Y_tri_63_inst : TBUF_X1 port map( A => n438, EN => n301, Z => Y(63));
   Y_tri_53_inst : TBUF_X1 port map( A => n448, EN => n300, Z => Y(53));
   Y_tri_54_inst : TBUF_X1 port map( A => n447, EN => n300, Z => Y(54));
   Y_tri_55_inst : TBUF_X1 port map( A => n446, EN => n300, Z => Y(55));
   Y_tri_56_inst : TBUF_X1 port map( A => n445, EN => n300, Z => Y(56));
   Y_tri_57_inst : TBUF_X1 port map( A => n444, EN => n300, Z => Y(57));
   Y_tri_58_inst : TBUF_X1 port map( A => n443, EN => n300, Z => Y(58));
   Y_tri_59_inst : TBUF_X1 port map( A => n442, EN => n300, Z => Y(59));
   Y_tri_21_inst : TBUF_X1 port map( A => n480, EN => n297, Z => Y(21));
   Y_tri_22_inst : TBUF_X1 port map( A => n479, EN => n297, Z => Y(22));
   Y_tri_23_inst : TBUF_X1 port map( A => n478, EN => n297, Z => Y(23));
   Y_tri_26_inst : TBUF_X1 port map( A => n475, EN => n298, Z => Y(26));
   Y_tri_27_inst : TBUF_X1 port map( A => n474, EN => n298, Z => Y(27));
   Y_tri_28_inst : TBUF_X1 port map( A => n473, EN => n298, Z => Y(28));
   Y_tri_29_inst : TBUF_X1 port map( A => n472, EN => n298, Z => Y(29));
   Y_tri_30_inst : TBUF_X1 port map( A => n471, EN => n298, Z => Y(30));
   Y_tri_31_inst : TBUF_X1 port map( A => n470, EN => n298, Z => Y(31));
   Y_tri_32_inst : TBUF_X1 port map( A => n469, EN => n298, Z => Y(32));
   Y_tri_33_inst : TBUF_X1 port map( A => n468, EN => n298, Z => Y(33));
   Y_tri_34_inst : TBUF_X1 port map( A => n467, EN => n298, Z => Y(34));
   Y_tri_35_inst : TBUF_X1 port map( A => n466, EN => n298, Z => Y(35));
   Y_tri_36_inst : TBUF_X1 port map( A => n465, EN => n299, Z => Y(36));
   Y_tri_37_inst : TBUF_X1 port map( A => n464, EN => n299, Z => Y(37));
   Y_tri_38_inst : TBUF_X1 port map( A => n463, EN => n299, Z => Y(38));
   Y_tri_39_inst : TBUF_X1 port map( A => n462, EN => n299, Z => Y(39));
   Y_tri_40_inst : TBUF_X1 port map( A => n461, EN => n299, Z => Y(40));
   Y_tri_41_inst : TBUF_X1 port map( A => n460, EN => n299, Z => Y(41));
   Y_tri_42_inst : TBUF_X1 port map( A => n459, EN => n299, Z => Y(42));
   Y_tri_43_inst : TBUF_X1 port map( A => n458, EN => n299, Z => Y(43));
   Y_tri_44_inst : TBUF_X1 port map( A => n457, EN => n299, Z => Y(44));
   Y_tri_45_inst : TBUF_X1 port map( A => n456, EN => n299, Z => Y(45));
   Y_tri_46_inst : TBUF_X1 port map( A => n455, EN => n299, Z => Y(46));
   Y_tri_47_inst : TBUF_X1 port map( A => n454, EN => n299, Z => Y(47));
   Y_tri_48_inst : TBUF_X1 port map( A => n453, EN => n300, Z => Y(48));
   Y_tri_49_inst : TBUF_X1 port map( A => n452, EN => n300, Z => Y(49));
   Y_tri_50_inst : TBUF_X1 port map( A => n451, EN => n300, Z => Y(50));
   Y_tri_51_inst : TBUF_X1 port map( A => n450, EN => n300, Z => Y(51));
   Y_tri_52_inst : TBUF_X1 port map( A => n449, EN => n300, Z => Y(52));
   Y_tri_10_inst : TBUF_X1 port map( A => n491, EN => n296, Z => Y(10));
   Y_tri_11_inst : TBUF_X1 port map( A => n490, EN => n296, Z => Y(11));
   Y_tri_12_inst : TBUF_X1 port map( A => n489, EN => n297, Z => Y(12));
   Y_tri_13_inst : TBUF_X1 port map( A => n488, EN => n297, Z => Y(13));
   Y_tri_14_inst : TBUF_X1 port map( A => n487, EN => n297, Z => Y(14));
   Y_tri_15_inst : TBUF_X1 port map( A => n486, EN => n297, Z => Y(15));
   Y_tri_16_inst : TBUF_X1 port map( A => n485, EN => n297, Z => Y(16));
   Y_tri_17_inst : TBUF_X1 port map( A => n484, EN => n297, Z => Y(17));
   Y_tri_18_inst : TBUF_X1 port map( A => n483, EN => n297, Z => Y(18));
   Y_tri_19_inst : TBUF_X1 port map( A => n482, EN => n297, Z => Y(19));
   Y_tri_20_inst : TBUF_X1 port map( A => n481, EN => n297, Z => Y(20));
   Y_tri_24_inst : TBUF_X1 port map( A => n477, EN => n298, Z => Y(24));
   Y_tri_25_inst : TBUF_X1 port map( A => n476, EN => n298, Z => Y(25));
   Y_tri_0_inst : TBUF_X1 port map( A => n502, EN => n296, Z => Y(0));
   Y_tri_1_inst : TBUF_X1 port map( A => n501, EN => n296, Z => Y(1));
   Y_tri_2_inst : TBUF_X1 port map( A => n500, EN => n296, Z => Y(2));
   Y_tri_3_inst : TBUF_X1 port map( A => n499, EN => n296, Z => Y(3));
   Y_tri_4_inst : TBUF_X1 port map( A => n498, EN => n296, Z => Y(4));
   Y_tri_5_inst : TBUF_X1 port map( A => n497, EN => n296, Z => Y(5));
   Y_tri_6_inst : TBUF_X1 port map( A => n496, EN => n296, Z => Y(6));
   Y_tri_7_inst : TBUF_X1 port map( A => n495, EN => n296, Z => Y(7));
   Y_tri_8_inst : TBUF_X1 port map( A => n494, EN => n296, Z => Y(8));
   Y_tri_9_inst : TBUF_X1 port map( A => n492, EN => n296, Z => Y(9));
   U2 : NOR3_X1 port map( A1 => SEL(0), A2 => SEL(2), A3 => n302, ZN => n434);
   U3 : NOR3_X1 port map( A1 => n302, A2 => SEL(2), A3 => n303, ZN => n432);
   U4 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n303, ZN => n433);
   U5 : NAND2_X1 port map( A1 => n411, A2 => n410, ZN => n449);
   U6 : AOI22_X1 port map( A1 => plusA(52), A2 => n282, B1 => plus2A(52), B2 =>
                           n276, ZN => n411);
   U7 : AOI22_X1 port map( A1 => minus2A(52), A2 => n294, B1 => minusA(52), B2 
                           => n288, ZN => n410);
   U8 : NAND2_X1 port map( A1 => n409, A2 => n408, ZN => n450);
   U9 : AOI22_X1 port map( A1 => plusA(51), A2 => n282, B1 => plus2A(51), B2 =>
                           n276, ZN => n409);
   U10 : AOI22_X1 port map( A1 => minus2A(51), A2 => n294, B1 => minusA(51), B2
                           => n288, ZN => n408);
   U11 : NAND2_X1 port map( A1 => n407, A2 => n406, ZN => n451);
   U12 : AOI22_X1 port map( A1 => plusA(50), A2 => n282, B1 => plus2A(50), B2 
                           => n276, ZN => n407);
   U13 : AOI22_X1 port map( A1 => minus2A(50), A2 => n294, B1 => minusA(50), B2
                           => n288, ZN => n406);
   U14 : NAND2_X1 port map( A1 => n405, A2 => n404, ZN => n452);
   U15 : AOI22_X1 port map( A1 => plusA(49), A2 => n282, B1 => plus2A(49), B2 
                           => n276, ZN => n405);
   U16 : AOI22_X1 port map( A1 => minus2A(49), A2 => n294, B1 => minusA(49), B2
                           => n288, ZN => n404);
   U17 : NAND2_X1 port map( A1 => n403, A2 => n402, ZN => n453);
   U18 : AOI22_X1 port map( A1 => plusA(48), A2 => n282, B1 => plus2A(48), B2 
                           => n276, ZN => n403);
   U19 : AOI22_X1 port map( A1 => minus2A(48), A2 => n294, B1 => minusA(48), B2
                           => n288, ZN => n402);
   U20 : NAND2_X1 port map( A1 => n401, A2 => n400, ZN => n454);
   U21 : AOI22_X1 port map( A1 => plusA(47), A2 => n281, B1 => plus2A(47), B2 
                           => n275, ZN => n401);
   U22 : AOI22_X1 port map( A1 => minus2A(47), A2 => n293, B1 => minusA(47), B2
                           => n287, ZN => n400);
   U23 : NAND2_X1 port map( A1 => n399, A2 => n398, ZN => n455);
   U24 : AOI22_X1 port map( A1 => plusA(46), A2 => n281, B1 => plus2A(46), B2 
                           => n275, ZN => n399);
   U25 : AOI22_X1 port map( A1 => minus2A(46), A2 => n293, B1 => minusA(46), B2
                           => n287, ZN => n398);
   U26 : NAND2_X1 port map( A1 => n393, A2 => n392, ZN => n458);
   U27 : AOI22_X1 port map( A1 => plusA(43), A2 => n281, B1 => plus2A(43), B2 
                           => n275, ZN => n393);
   U28 : AOI22_X1 port map( A1 => minus2A(43), A2 => n293, B1 => minusA(43), B2
                           => n287, ZN => n392);
   U29 : NAND2_X1 port map( A1 => n387, A2 => n386, ZN => n461);
   U30 : AOI22_X1 port map( A1 => plusA(40), A2 => n281, B1 => plus2A(40), B2 
                           => n275, ZN => n387);
   U31 : AOI22_X1 port map( A1 => minus2A(40), A2 => n293, B1 => minusA(40), B2
                           => n287, ZN => n386);
   U32 : NAND2_X1 port map( A1 => n385, A2 => n384, ZN => n462);
   U33 : AOI22_X1 port map( A1 => plusA(39), A2 => n281, B1 => plus2A(39), B2 
                           => n275, ZN => n385);
   U34 : AOI22_X1 port map( A1 => minus2A(39), A2 => n293, B1 => minusA(39), B2
                           => n287, ZN => n384);
   U35 : NAND2_X1 port map( A1 => n383, A2 => n382, ZN => n463);
   U36 : AOI22_X1 port map( A1 => plusA(38), A2 => n281, B1 => plus2A(38), B2 
                           => n275, ZN => n383);
   U37 : AOI22_X1 port map( A1 => minus2A(38), A2 => n293, B1 => minusA(38), B2
                           => n287, ZN => n382);
   U38 : NAND2_X1 port map( A1 => n391, A2 => n390, ZN => n459);
   U39 : AOI22_X1 port map( A1 => plusA(42), A2 => n281, B1 => plus2A(42), B2 
                           => n275, ZN => n391);
   U40 : AOI22_X1 port map( A1 => minus2A(42), A2 => n293, B1 => minusA(42), B2
                           => n287, ZN => n390);
   U41 : NAND2_X1 port map( A1 => n375, A2 => n374, ZN => n467);
   U42 : AOI22_X1 port map( A1 => plusA(34), A2 => n280, B1 => plus2A(34), B2 
                           => n274, ZN => n375);
   U43 : AOI22_X1 port map( A1 => minus2A(34), A2 => n292, B1 => minusA(34), B2
                           => n286, ZN => n374);
   U44 : NAND2_X1 port map( A1 => n367, A2 => n366, ZN => n471);
   U45 : AOI22_X1 port map( A1 => plusA(30), A2 => n280, B1 => plus2A(30), B2 
                           => n274, ZN => n367);
   U46 : AOI22_X1 port map( A1 => minus2A(30), A2 => n292, B1 => minusA(30), B2
                           => n286, ZN => n366);
   U47 : NAND2_X1 port map( A1 => n395, A2 => n394, ZN => n457);
   U48 : AOI22_X1 port map( A1 => plusA(44), A2 => n281, B1 => plus2A(44), B2 
                           => n275, ZN => n395);
   U49 : AOI22_X1 port map( A1 => minus2A(44), A2 => n293, B1 => minusA(44), B2
                           => n287, ZN => n394);
   U50 : NAND2_X1 port map( A1 => n379, A2 => n378, ZN => n465);
   U51 : AOI22_X1 port map( A1 => plusA(36), A2 => n281, B1 => plus2A(36), B2 
                           => n275, ZN => n379);
   U52 : AOI22_X1 port map( A1 => minus2A(36), A2 => n293, B1 => minusA(36), B2
                           => n287, ZN => n378);
   U53 : NAND2_X1 port map( A1 => n371, A2 => n370, ZN => n469);
   U54 : AOI22_X1 port map( A1 => plusA(32), A2 => n280, B1 => plus2A(32), B2 
                           => n274, ZN => n371);
   U55 : AOI22_X1 port map( A1 => minus2A(32), A2 => n292, B1 => minusA(32), B2
                           => n286, ZN => n370);
   U56 : NAND2_X1 port map( A1 => n363, A2 => n362, ZN => n473);
   U57 : AOI22_X1 port map( A1 => plusA(28), A2 => n280, B1 => plus2A(28), B2 
                           => n274, ZN => n363);
   U58 : AOI22_X1 port map( A1 => minus2A(28), A2 => n292, B1 => minusA(28), B2
                           => n286, ZN => n362);
   U59 : NAND2_X1 port map( A1 => n377, A2 => n376, ZN => n466);
   U60 : AOI22_X1 port map( A1 => plusA(35), A2 => n280, B1 => plus2A(35), B2 
                           => n274, ZN => n377);
   U61 : AOI22_X1 port map( A1 => minus2A(35), A2 => n292, B1 => minusA(35), B2
                           => n286, ZN => n376);
   U62 : NAND2_X1 port map( A1 => n369, A2 => n368, ZN => n470);
   U63 : AOI22_X1 port map( A1 => plusA(31), A2 => n280, B1 => plus2A(31), B2 
                           => n274, ZN => n369);
   U64 : AOI22_X1 port map( A1 => minus2A(31), A2 => n292, B1 => minusA(31), B2
                           => n286, ZN => n368);
   U65 : NAND2_X1 port map( A1 => n397, A2 => n396, ZN => n456);
   U66 : AOI22_X1 port map( A1 => plusA(45), A2 => n281, B1 => plus2A(45), B2 
                           => n275, ZN => n397);
   U67 : AOI22_X1 port map( A1 => minus2A(45), A2 => n293, B1 => minusA(45), B2
                           => n287, ZN => n396);
   U68 : NAND2_X1 port map( A1 => n389, A2 => n388, ZN => n460);
   U69 : AOI22_X1 port map( A1 => plusA(41), A2 => n281, B1 => plus2A(41), B2 
                           => n275, ZN => n389);
   U70 : AOI22_X1 port map( A1 => minus2A(41), A2 => n293, B1 => minusA(41), B2
                           => n287, ZN => n388);
   U71 : NAND2_X1 port map( A1 => n381, A2 => n380, ZN => n464);
   U72 : AOI22_X1 port map( A1 => plusA(37), A2 => n281, B1 => plus2A(37), B2 
                           => n275, ZN => n381);
   U73 : AOI22_X1 port map( A1 => minus2A(37), A2 => n293, B1 => minusA(37), B2
                           => n287, ZN => n380);
   U74 : NAND2_X1 port map( A1 => n373, A2 => n372, ZN => n468);
   U75 : AOI22_X1 port map( A1 => plusA(33), A2 => n280, B1 => plus2A(33), B2 
                           => n274, ZN => n373);
   U76 : AOI22_X1 port map( A1 => minus2A(33), A2 => n292, B1 => minusA(33), B2
                           => n286, ZN => n372);
   U77 : NAND2_X1 port map( A1 => n365, A2 => n364, ZN => n472);
   U78 : AOI22_X1 port map( A1 => plusA(29), A2 => n280, B1 => plus2A(29), B2 
                           => n274, ZN => n365);
   U79 : AOI22_X1 port map( A1 => minus2A(29), A2 => n292, B1 => minusA(29), B2
                           => n286, ZN => n364);
   U80 : NAND2_X1 port map( A1 => n437, A2 => n436, ZN => n438);
   U81 : AOI22_X1 port map( A1 => plusA(63), A2 => n283, B1 => plus2A(63), B2 
                           => n277, ZN => n437);
   U82 : AOI22_X1 port map( A1 => minus2A(63), A2 => n295, B1 => minusA(63), B2
                           => n289, ZN => n436);
   U83 : NAND2_X1 port map( A1 => n431, A2 => n430, ZN => n439);
   U84 : AOI22_X1 port map( A1 => plusA(62), A2 => n283, B1 => plus2A(62), B2 
                           => n277, ZN => n431);
   U85 : AOI22_X1 port map( A1 => minus2A(62), A2 => n295, B1 => minusA(62), B2
                           => n289, ZN => n430);
   U86 : NAND2_X1 port map( A1 => n429, A2 => n428, ZN => n440);
   U87 : AOI22_X1 port map( A1 => plusA(61), A2 => n283, B1 => plus2A(61), B2 
                           => n277, ZN => n429);
   U88 : AOI22_X1 port map( A1 => minus2A(61), A2 => n295, B1 => minusA(61), B2
                           => n289, ZN => n428);
   U89 : NAND2_X1 port map( A1 => n427, A2 => n426, ZN => n441);
   U90 : AOI22_X1 port map( A1 => plusA(60), A2 => n283, B1 => plus2A(60), B2 
                           => n277, ZN => n427);
   U91 : AOI22_X1 port map( A1 => minus2A(60), A2 => n295, B1 => minusA(60), B2
                           => n289, ZN => n426);
   U92 : NAND2_X1 port map( A1 => n425, A2 => n424, ZN => n442);
   U93 : AOI22_X1 port map( A1 => plusA(59), A2 => n282, B1 => plus2A(59), B2 
                           => n276, ZN => n425);
   U94 : AOI22_X1 port map( A1 => minus2A(59), A2 => n294, B1 => minusA(59), B2
                           => n288, ZN => n424);
   U95 : NAND2_X1 port map( A1 => n423, A2 => n422, ZN => n443);
   U96 : AOI22_X1 port map( A1 => plusA(58), A2 => n282, B1 => plus2A(58), B2 
                           => n276, ZN => n423);
   U97 : AOI22_X1 port map( A1 => minus2A(58), A2 => n294, B1 => minusA(58), B2
                           => n288, ZN => n422);
   U98 : NAND2_X1 port map( A1 => n421, A2 => n420, ZN => n444);
   U99 : AOI22_X1 port map( A1 => plusA(57), A2 => n282, B1 => plus2A(57), B2 
                           => n276, ZN => n421);
   U100 : AOI22_X1 port map( A1 => minus2A(57), A2 => n294, B1 => minusA(57), 
                           B2 => n288, ZN => n420);
   U101 : NAND2_X1 port map( A1 => n419, A2 => n418, ZN => n445);
   U102 : AOI22_X1 port map( A1 => plusA(56), A2 => n282, B1 => plus2A(56), B2 
                           => n276, ZN => n419);
   U103 : AOI22_X1 port map( A1 => minus2A(56), A2 => n294, B1 => minusA(56), 
                           B2 => n288, ZN => n418);
   U104 : NAND2_X1 port map( A1 => n417, A2 => n416, ZN => n446);
   U105 : AOI22_X1 port map( A1 => plusA(55), A2 => n282, B1 => plus2A(55), B2 
                           => n276, ZN => n417);
   U106 : AOI22_X1 port map( A1 => minus2A(55), A2 => n294, B1 => minusA(55), 
                           B2 => n288, ZN => n416);
   U107 : NAND2_X1 port map( A1 => n415, A2 => n414, ZN => n447);
   U108 : AOI22_X1 port map( A1 => plusA(54), A2 => n282, B1 => plus2A(54), B2 
                           => n276, ZN => n415);
   U109 : AOI22_X1 port map( A1 => minus2A(54), A2 => n294, B1 => minusA(54), 
                           B2 => n288, ZN => n414);
   U110 : NAND2_X1 port map( A1 => n413, A2 => n412, ZN => n448);
   U111 : AOI22_X1 port map( A1 => plusA(53), A2 => n282, B1 => plus2A(53), B2 
                           => n276, ZN => n413);
   U112 : AOI22_X1 port map( A1 => minus2A(53), A2 => n294, B1 => minusA(53), 
                           B2 => n288, ZN => n412);
   U113 : BUF_X1 port map( A => n493, Z => n296);
   U114 : BUF_X1 port map( A => n493, Z => n297);
   U115 : BUF_X1 port map( A => n493, Z => n298);
   U116 : BUF_X1 port map( A => n433, Z => n280);
   U117 : BUF_X1 port map( A => n434, Z => n286);
   U118 : BUF_X1 port map( A => n432, Z => n274);
   U119 : BUF_X1 port map( A => n435, Z => n292);
   U120 : NAND2_X1 port map( A1 => n359, A2 => n358, ZN => n475);
   U121 : AOI22_X1 port map( A1 => plusA(26), A2 => n280, B1 => plus2A(26), B2 
                           => n274, ZN => n359);
   U122 : AOI22_X1 port map( A1 => minus2A(26), A2 => n292, B1 => minusA(26), 
                           B2 => n286, ZN => n358);
   U123 : NAND2_X1 port map( A1 => n361, A2 => n360, ZN => n474);
   U124 : AOI22_X1 port map( A1 => plusA(27), A2 => n280, B1 => plus2A(27), B2 
                           => n274, ZN => n361);
   U125 : AOI22_X1 port map( A1 => minus2A(27), A2 => n292, B1 => minusA(27), 
                           B2 => n286, ZN => n360);
   U126 : BUF_X1 port map( A => n493, Z => n299);
   U127 : BUF_X1 port map( A => n433, Z => n281);
   U128 : BUF_X1 port map( A => n434, Z => n287);
   U129 : BUF_X1 port map( A => n432, Z => n275);
   U130 : BUF_X1 port map( A => n435, Z => n293);
   U131 : BUF_X1 port map( A => n493, Z => n300);
   U132 : BUF_X1 port map( A => n433, Z => n282);
   U133 : BUF_X1 port map( A => n434, Z => n288);
   U134 : BUF_X1 port map( A => n432, Z => n276);
   U135 : BUF_X1 port map( A => n435, Z => n294);
   U136 : BUF_X1 port map( A => n433, Z => n279);
   U137 : BUF_X1 port map( A => n433, Z => n278);
   U138 : BUF_X1 port map( A => n434, Z => n285);
   U139 : BUF_X1 port map( A => n432, Z => n273);
   U140 : BUF_X1 port map( A => n434, Z => n284);
   U141 : BUF_X1 port map( A => n432, Z => n272);
   U142 : BUF_X1 port map( A => n435, Z => n291);
   U143 : BUF_X1 port map( A => n435, Z => n290);
   U144 : NOR2_X1 port map( A1 => n323, A2 => n304, ZN => n493);
   U145 : INV_X1 port map( A => SEL(2), ZN => n304);
   U146 : NOR2_X1 port map( A1 => SEL(1), A2 => SEL(0), ZN => n323);
   U147 : NAND2_X1 port map( A1 => n357, A2 => n356, ZN => n476);
   U148 : AOI22_X1 port map( A1 => plusA(25), A2 => n280, B1 => plus2A(25), B2 
                           => n274, ZN => n357);
   U149 : AOI22_X1 port map( A1 => minus2A(25), A2 => n292, B1 => minusA(25), 
                           B2 => n286, ZN => n356);
   U150 : AND2_X1 port map( A1 => SEL(2), A2 => n323, ZN => n435);
   U151 : INV_X1 port map( A => SEL(1), ZN => n302);
   U152 : INV_X1 port map( A => SEL(0), ZN => n303);
   U153 : NAND2_X1 port map( A1 => n355, A2 => n354, ZN => n477);
   U154 : AOI22_X1 port map( A1 => plusA(24), A2 => n280, B1 => plus2A(24), B2 
                           => n274, ZN => n355);
   U155 : AOI22_X1 port map( A1 => minus2A(24), A2 => n292, B1 => minusA(24), 
                           B2 => n286, ZN => n354);
   U156 : NAND2_X1 port map( A1 => n353, A2 => n352, ZN => n478);
   U157 : AOI22_X1 port map( A1 => plusA(23), A2 => n279, B1 => plus2A(23), B2 
                           => n273, ZN => n353);
   U158 : AOI22_X1 port map( A1 => minus2A(23), A2 => n291, B1 => minusA(23), 
                           B2 => n285, ZN => n352);
   U159 : NAND2_X1 port map( A1 => n351, A2 => n350, ZN => n479);
   U160 : AOI22_X1 port map( A1 => plusA(22), A2 => n279, B1 => plus2A(22), B2 
                           => n273, ZN => n351);
   U161 : AOI22_X1 port map( A1 => minus2A(22), A2 => n291, B1 => minusA(22), 
                           B2 => n285, ZN => n350);
   U162 : NAND2_X1 port map( A1 => n349, A2 => n348, ZN => n480);
   U163 : AOI22_X1 port map( A1 => plusA(21), A2 => n279, B1 => plus2A(21), B2 
                           => n273, ZN => n349);
   U164 : AOI22_X1 port map( A1 => minus2A(21), A2 => n291, B1 => minusA(21), 
                           B2 => n285, ZN => n348);
   U165 : NAND2_X1 port map( A1 => n345, A2 => n344, ZN => n482);
   U166 : AOI22_X1 port map( A1 => plusA(19), A2 => n279, B1 => plus2A(19), B2 
                           => n273, ZN => n345);
   U167 : AOI22_X1 port map( A1 => minus2A(19), A2 => n291, B1 => minusA(19), 
                           B2 => n285, ZN => n344);
   U168 : NAND2_X1 port map( A1 => n343, A2 => n342, ZN => n483);
   U169 : AOI22_X1 port map( A1 => plusA(18), A2 => n279, B1 => plus2A(18), B2 
                           => n273, ZN => n343);
   U170 : AOI22_X1 port map( A1 => minus2A(18), A2 => n291, B1 => minusA(18), 
                           B2 => n285, ZN => n342);
   U171 : NAND2_X1 port map( A1 => n341, A2 => n340, ZN => n484);
   U172 : AOI22_X1 port map( A1 => plusA(17), A2 => n279, B1 => plus2A(17), B2 
                           => n273, ZN => n341);
   U173 : AOI22_X1 port map( A1 => minus2A(17), A2 => n291, B1 => minusA(17), 
                           B2 => n285, ZN => n340);
   U174 : NAND2_X1 port map( A1 => n337, A2 => n336, ZN => n486);
   U175 : AOI22_X1 port map( A1 => plusA(15), A2 => n279, B1 => plus2A(15), B2 
                           => n273, ZN => n337);
   U176 : AOI22_X1 port map( A1 => minus2A(15), A2 => n291, B1 => minusA(15), 
                           B2 => n285, ZN => n336);
   U177 : NAND2_X1 port map( A1 => n335, A2 => n334, ZN => n487);
   U178 : AOI22_X1 port map( A1 => plusA(14), A2 => n279, B1 => plus2A(14), B2 
                           => n273, ZN => n335);
   U179 : AOI22_X1 port map( A1 => minus2A(14), A2 => n291, B1 => minusA(14), 
                           B2 => n285, ZN => n334);
   U180 : NAND2_X1 port map( A1 => n333, A2 => n332, ZN => n488);
   U181 : AOI22_X1 port map( A1 => plusA(13), A2 => n279, B1 => plus2A(13), B2 
                           => n273, ZN => n333);
   U182 : AOI22_X1 port map( A1 => minus2A(13), A2 => n291, B1 => minusA(13), 
                           B2 => n285, ZN => n332);
   U183 : NAND2_X1 port map( A1 => n329, A2 => n328, ZN => n490);
   U184 : AOI22_X1 port map( A1 => plusA(11), A2 => n278, B1 => plus2A(11), B2 
                           => n272, ZN => n329);
   U185 : AOI22_X1 port map( A1 => minus2A(11), A2 => n290, B1 => minusA(11), 
                           B2 => n284, ZN => n328);
   U186 : NAND2_X1 port map( A1 => n327, A2 => n326, ZN => n491);
   U187 : AOI22_X1 port map( A1 => plusA(10), A2 => n278, B1 => plus2A(10), B2 
                           => n272, ZN => n327);
   U188 : AOI22_X1 port map( A1 => minus2A(10), A2 => n290, B1 => minusA(10), 
                           B2 => n284, ZN => n326);
   U189 : NAND2_X1 port map( A1 => n325, A2 => n324, ZN => n492);
   U190 : AOI22_X1 port map( A1 => plusA(9), A2 => n278, B1 => plus2A(9), B2 =>
                           n272, ZN => n325);
   U191 : AOI22_X1 port map( A1 => minus2A(9), A2 => n290, B1 => minusA(9), B2 
                           => n284, ZN => n324);
   U192 : NAND2_X1 port map( A1 => n320, A2 => n319, ZN => n495);
   U193 : AOI22_X1 port map( A1 => plusA(7), A2 => n278, B1 => plus2A(7), B2 =>
                           n272, ZN => n320);
   U194 : AOI22_X1 port map( A1 => minus2A(7), A2 => n290, B1 => minusA(7), B2 
                           => n284, ZN => n319);
   U195 : NAND2_X1 port map( A1 => n318, A2 => n317, ZN => n496);
   U196 : AOI22_X1 port map( A1 => plusA(6), A2 => n278, B1 => plus2A(6), B2 =>
                           n272, ZN => n318);
   U197 : AOI22_X1 port map( A1 => minus2A(6), A2 => n290, B1 => minusA(6), B2 
                           => n284, ZN => n317);
   U198 : NAND2_X1 port map( A1 => n316, A2 => n315, ZN => n497);
   U199 : AOI22_X1 port map( A1 => plusA(5), A2 => n278, B1 => plus2A(5), B2 =>
                           n272, ZN => n316);
   U200 : AOI22_X1 port map( A1 => minus2A(5), A2 => n290, B1 => minusA(5), B2 
                           => n284, ZN => n315);
   U201 : NAND2_X1 port map( A1 => n312, A2 => n311, ZN => n499);
   U202 : AOI22_X1 port map( A1 => plusA(3), A2 => n278, B1 => plus2A(3), B2 =>
                           n272, ZN => n312);
   U203 : AOI22_X1 port map( A1 => minus2A(3), A2 => n290, B1 => minusA(3), B2 
                           => n284, ZN => n311);
   U204 : NAND2_X1 port map( A1 => n347, A2 => n346, ZN => n481);
   U205 : AOI22_X1 port map( A1 => plusA(20), A2 => n279, B1 => plus2A(20), B2 
                           => n273, ZN => n347);
   U206 : AOI22_X1 port map( A1 => minus2A(20), A2 => n291, B1 => minusA(20), 
                           B2 => n285, ZN => n346);
   U207 : NAND2_X1 port map( A1 => n339, A2 => n338, ZN => n485);
   U208 : AOI22_X1 port map( A1 => plusA(16), A2 => n279, B1 => plus2A(16), B2 
                           => n273, ZN => n339);
   U209 : AOI22_X1 port map( A1 => minus2A(16), A2 => n291, B1 => minusA(16), 
                           B2 => n285, ZN => n338);
   U210 : NAND2_X1 port map( A1 => n331, A2 => n330, ZN => n489);
   U211 : AOI22_X1 port map( A1 => plusA(12), A2 => n279, B1 => plus2A(12), B2 
                           => n273, ZN => n331);
   U212 : AOI22_X1 port map( A1 => minus2A(12), A2 => n291, B1 => minusA(12), 
                           B2 => n285, ZN => n330);
   U213 : NAND2_X1 port map( A1 => n322, A2 => n321, ZN => n494);
   U214 : AOI22_X1 port map( A1 => plusA(8), A2 => n278, B1 => plus2A(8), B2 =>
                           n272, ZN => n322);
   U215 : AOI22_X1 port map( A1 => minus2A(8), A2 => n290, B1 => minusA(8), B2 
                           => n284, ZN => n321);
   U216 : NAND2_X1 port map( A1 => n314, A2 => n313, ZN => n498);
   U217 : AOI22_X1 port map( A1 => plusA(4), A2 => n278, B1 => plus2A(4), B2 =>
                           n272, ZN => n314);
   U218 : AOI22_X1 port map( A1 => minus2A(4), A2 => n290, B1 => minusA(4), B2 
                           => n284, ZN => n313);
   U219 : NAND2_X1 port map( A1 => n310, A2 => n309, ZN => n500);
   U220 : AOI22_X1 port map( A1 => plusA(2), A2 => n278, B1 => plus2A(2), B2 =>
                           n272, ZN => n310);
   U221 : AOI22_X1 port map( A1 => minus2A(2), A2 => n290, B1 => minusA(2), B2 
                           => n284, ZN => n309);
   U222 : NAND2_X1 port map( A1 => n308, A2 => n307, ZN => n501);
   U223 : AOI22_X1 port map( A1 => plusA(1), A2 => n278, B1 => plus2A(1), B2 =>
                           n272, ZN => n308);
   U224 : AOI22_X1 port map( A1 => minus2A(1), A2 => n290, B1 => minusA(1), B2 
                           => n284, ZN => n307);
   U225 : NAND2_X1 port map( A1 => n306, A2 => n305, ZN => n502);
   U226 : AOI22_X1 port map( A1 => plusA(0), A2 => n278, B1 => plus2A(0), B2 =>
                           n272, ZN => n306);
   U227 : AOI22_X1 port map( A1 => minus2A(0), A2 => n290, B1 => minusA(0), B2 
                           => n284, ZN => n305);
   U228 : CLKBUF_X1 port map( A => n432, Z => n277);
   U229 : CLKBUF_X1 port map( A => n433, Z => n283);
   U230 : CLKBUF_X1 port map( A => n434, Z => n289);
   U231 : CLKBUF_X1 port map( A => n435, Z => n295);
   U232 : CLKBUF_X1 port map( A => n493, Z => n301);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity MUX_GENERIC_N64_RADIX3_3 is

   port( plusA, minusA, plus2A, minus2A : in std_logic_vector (63 downto 0);  
         SEL : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (63 
         downto 0));

end MUX_GENERIC_N64_RADIX3_3;

architecture SYN_beh of MUX_GENERIC_N64_RADIX3_3 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component TBUF_X1
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   signal n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, 
      n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, 
      n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, 
      n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, 
      n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, 
      n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, 
      n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, 
      n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, 
      n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, 
      n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, 
      n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, 
      n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, 
      n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, 
      n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, 
      n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, 
      n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, 
      n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, 
      n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, 
      n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, 
      n499, n500, n501, n502 : std_logic;

begin
   
   Y_tri_60_inst : TBUF_X1 port map( A => n441, EN => n301, Z => Y(60));
   Y_tri_61_inst : TBUF_X1 port map( A => n440, EN => n301, Z => Y(61));
   Y_tri_62_inst : TBUF_X1 port map( A => n439, EN => n301, Z => Y(62));
   Y_tri_63_inst : TBUF_X1 port map( A => n438, EN => n301, Z => Y(63));
   Y_tri_46_inst : TBUF_X1 port map( A => n455, EN => n299, Z => Y(46));
   Y_tri_47_inst : TBUF_X1 port map( A => n454, EN => n299, Z => Y(47));
   Y_tri_48_inst : TBUF_X1 port map( A => n453, EN => n300, Z => Y(48));
   Y_tri_49_inst : TBUF_X1 port map( A => n452, EN => n300, Z => Y(49));
   Y_tri_50_inst : TBUF_X1 port map( A => n451, EN => n300, Z => Y(50));
   Y_tri_51_inst : TBUF_X1 port map( A => n450, EN => n300, Z => Y(51));
   Y_tri_52_inst : TBUF_X1 port map( A => n449, EN => n300, Z => Y(52));
   Y_tri_53_inst : TBUF_X1 port map( A => n448, EN => n300, Z => Y(53));
   Y_tri_54_inst : TBUF_X1 port map( A => n447, EN => n300, Z => Y(54));
   Y_tri_55_inst : TBUF_X1 port map( A => n446, EN => n300, Z => Y(55));
   Y_tri_56_inst : TBUF_X1 port map( A => n445, EN => n300, Z => Y(56));
   Y_tri_57_inst : TBUF_X1 port map( A => n444, EN => n300, Z => Y(57));
   Y_tri_58_inst : TBUF_X1 port map( A => n443, EN => n300, Z => Y(58));
   Y_tri_59_inst : TBUF_X1 port map( A => n442, EN => n300, Z => Y(59));
   Y_tri_19_inst : TBUF_X1 port map( A => n482, EN => n297, Z => Y(19));
   Y_tri_20_inst : TBUF_X1 port map( A => n481, EN => n297, Z => Y(20));
   Y_tri_21_inst : TBUF_X1 port map( A => n480, EN => n297, Z => Y(21));
   Y_tri_22_inst : TBUF_X1 port map( A => n479, EN => n297, Z => Y(22));
   Y_tri_23_inst : TBUF_X1 port map( A => n478, EN => n297, Z => Y(23));
   Y_tri_24_inst : TBUF_X1 port map( A => n477, EN => n298, Z => Y(24));
   Y_tri_25_inst : TBUF_X1 port map( A => n476, EN => n298, Z => Y(25));
   Y_tri_26_inst : TBUF_X1 port map( A => n475, EN => n298, Z => Y(26));
   Y_tri_27_inst : TBUF_X1 port map( A => n474, EN => n298, Z => Y(27));
   Y_tri_28_inst : TBUF_X1 port map( A => n473, EN => n298, Z => Y(28));
   Y_tri_29_inst : TBUF_X1 port map( A => n472, EN => n298, Z => Y(29));
   Y_tri_30_inst : TBUF_X1 port map( A => n471, EN => n298, Z => Y(30));
   Y_tri_31_inst : TBUF_X1 port map( A => n470, EN => n298, Z => Y(31));
   Y_tri_32_inst : TBUF_X1 port map( A => n469, EN => n298, Z => Y(32));
   Y_tri_33_inst : TBUF_X1 port map( A => n468, EN => n298, Z => Y(33));
   Y_tri_34_inst : TBUF_X1 port map( A => n467, EN => n298, Z => Y(34));
   Y_tri_35_inst : TBUF_X1 port map( A => n466, EN => n298, Z => Y(35));
   Y_tri_36_inst : TBUF_X1 port map( A => n465, EN => n299, Z => Y(36));
   Y_tri_37_inst : TBUF_X1 port map( A => n464, EN => n299, Z => Y(37));
   Y_tri_38_inst : TBUF_X1 port map( A => n463, EN => n299, Z => Y(38));
   Y_tri_39_inst : TBUF_X1 port map( A => n462, EN => n299, Z => Y(39));
   Y_tri_40_inst : TBUF_X1 port map( A => n461, EN => n299, Z => Y(40));
   Y_tri_41_inst : TBUF_X1 port map( A => n460, EN => n299, Z => Y(41));
   Y_tri_42_inst : TBUF_X1 port map( A => n459, EN => n299, Z => Y(42));
   Y_tri_43_inst : TBUF_X1 port map( A => n458, EN => n299, Z => Y(43));
   Y_tri_44_inst : TBUF_X1 port map( A => n457, EN => n299, Z => Y(44));
   Y_tri_45_inst : TBUF_X1 port map( A => n456, EN => n299, Z => Y(45));
   Y_tri_8_inst : TBUF_X1 port map( A => n494, EN => n296, Z => Y(8));
   Y_tri_9_inst : TBUF_X1 port map( A => n492, EN => n296, Z => Y(9));
   Y_tri_10_inst : TBUF_X1 port map( A => n491, EN => n296, Z => Y(10));
   Y_tri_11_inst : TBUF_X1 port map( A => n490, EN => n296, Z => Y(11));
   Y_tri_12_inst : TBUF_X1 port map( A => n489, EN => n297, Z => Y(12));
   Y_tri_13_inst : TBUF_X1 port map( A => n488, EN => n297, Z => Y(13));
   Y_tri_14_inst : TBUF_X1 port map( A => n487, EN => n297, Z => Y(14));
   Y_tri_15_inst : TBUF_X1 port map( A => n486, EN => n297, Z => Y(15));
   Y_tri_16_inst : TBUF_X1 port map( A => n485, EN => n297, Z => Y(16));
   Y_tri_17_inst : TBUF_X1 port map( A => n484, EN => n297, Z => Y(17));
   Y_tri_18_inst : TBUF_X1 port map( A => n483, EN => n297, Z => Y(18));
   Y_tri_0_inst : TBUF_X1 port map( A => n502, EN => n296, Z => Y(0));
   Y_tri_1_inst : TBUF_X1 port map( A => n501, EN => n296, Z => Y(1));
   Y_tri_2_inst : TBUF_X1 port map( A => n500, EN => n296, Z => Y(2));
   Y_tri_3_inst : TBUF_X1 port map( A => n499, EN => n296, Z => Y(3));
   Y_tri_4_inst : TBUF_X1 port map( A => n498, EN => n296, Z => Y(4));
   Y_tri_5_inst : TBUF_X1 port map( A => n497, EN => n296, Z => Y(5));
   Y_tri_6_inst : TBUF_X1 port map( A => n496, EN => n296, Z => Y(6));
   Y_tri_7_inst : TBUF_X1 port map( A => n495, EN => n296, Z => Y(7));
   U2 : NOR3_X1 port map( A1 => SEL(0), A2 => SEL(2), A3 => n302, ZN => n434);
   U3 : NOR3_X1 port map( A1 => n302, A2 => SEL(2), A3 => n303, ZN => n432);
   U4 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n303, ZN => n433);
   U5 : NAND2_X1 port map( A1 => n395, A2 => n394, ZN => n457);
   U6 : AOI22_X1 port map( A1 => plusA(44), A2 => n281, B1 => plus2A(44), B2 =>
                           n275, ZN => n395);
   U7 : AOI22_X1 port map( A1 => minus2A(44), A2 => n293, B1 => minusA(44), B2 
                           => n287, ZN => n394);
   U8 : NAND2_X1 port map( A1 => n393, A2 => n392, ZN => n458);
   U9 : AOI22_X1 port map( A1 => plusA(43), A2 => n281, B1 => plus2A(43), B2 =>
                           n275, ZN => n393);
   U10 : AOI22_X1 port map( A1 => minus2A(43), A2 => n293, B1 => minusA(43), B2
                           => n287, ZN => n392);
   U11 : NAND2_X1 port map( A1 => n387, A2 => n386, ZN => n461);
   U12 : AOI22_X1 port map( A1 => plusA(40), A2 => n281, B1 => plus2A(40), B2 
                           => n275, ZN => n387);
   U13 : AOI22_X1 port map( A1 => minus2A(40), A2 => n293, B1 => minusA(40), B2
                           => n287, ZN => n386);
   U14 : NAND2_X1 port map( A1 => n385, A2 => n384, ZN => n462);
   U15 : AOI22_X1 port map( A1 => plusA(39), A2 => n281, B1 => plus2A(39), B2 
                           => n275, ZN => n385);
   U16 : AOI22_X1 port map( A1 => minus2A(39), A2 => n293, B1 => minusA(39), B2
                           => n287, ZN => n384);
   U17 : NAND2_X1 port map( A1 => n379, A2 => n378, ZN => n465);
   U18 : AOI22_X1 port map( A1 => plusA(36), A2 => n281, B1 => plus2A(36), B2 
                           => n275, ZN => n379);
   U19 : AOI22_X1 port map( A1 => minus2A(36), A2 => n293, B1 => minusA(36), B2
                           => n287, ZN => n378);
   U20 : NAND2_X1 port map( A1 => n377, A2 => n376, ZN => n466);
   U21 : AOI22_X1 port map( A1 => plusA(35), A2 => n280, B1 => plus2A(35), B2 
                           => n274, ZN => n377);
   U22 : AOI22_X1 port map( A1 => minus2A(35), A2 => n292, B1 => minusA(35), B2
                           => n286, ZN => n376);
   U23 : NAND2_X1 port map( A1 => n369, A2 => n368, ZN => n470);
   U24 : AOI22_X1 port map( A1 => plusA(31), A2 => n280, B1 => plus2A(31), B2 
                           => n274, ZN => n369);
   U25 : AOI22_X1 port map( A1 => minus2A(31), A2 => n292, B1 => minusA(31), B2
                           => n286, ZN => n368);
   U26 : NAND2_X1 port map( A1 => n397, A2 => n396, ZN => n456);
   U27 : AOI22_X1 port map( A1 => plusA(45), A2 => n281, B1 => plus2A(45), B2 
                           => n275, ZN => n397);
   U28 : AOI22_X1 port map( A1 => minus2A(45), A2 => n293, B1 => minusA(45), B2
                           => n287, ZN => n396);
   U29 : NAND2_X1 port map( A1 => n389, A2 => n388, ZN => n460);
   U30 : AOI22_X1 port map( A1 => plusA(41), A2 => n281, B1 => plus2A(41), B2 
                           => n275, ZN => n389);
   U31 : AOI22_X1 port map( A1 => minus2A(41), A2 => n293, B1 => minusA(41), B2
                           => n287, ZN => n388);
   U32 : NAND2_X1 port map( A1 => n381, A2 => n380, ZN => n464);
   U33 : AOI22_X1 port map( A1 => plusA(37), A2 => n281, B1 => plus2A(37), B2 
                           => n275, ZN => n381);
   U34 : AOI22_X1 port map( A1 => minus2A(37), A2 => n293, B1 => minusA(37), B2
                           => n287, ZN => n380);
   U35 : NAND2_X1 port map( A1 => n373, A2 => n372, ZN => n468);
   U36 : AOI22_X1 port map( A1 => plusA(33), A2 => n280, B1 => plus2A(33), B2 
                           => n274, ZN => n373);
   U37 : AOI22_X1 port map( A1 => minus2A(33), A2 => n292, B1 => minusA(33), B2
                           => n286, ZN => n372);
   U38 : NAND2_X1 port map( A1 => n371, A2 => n370, ZN => n469);
   U39 : AOI22_X1 port map( A1 => plusA(32), A2 => n280, B1 => plus2A(32), B2 
                           => n274, ZN => n371);
   U40 : AOI22_X1 port map( A1 => minus2A(32), A2 => n292, B1 => minusA(32), B2
                           => n286, ZN => n370);
   U41 : NAND2_X1 port map( A1 => n391, A2 => n390, ZN => n459);
   U42 : AOI22_X1 port map( A1 => plusA(42), A2 => n281, B1 => plus2A(42), B2 
                           => n275, ZN => n391);
   U43 : AOI22_X1 port map( A1 => minus2A(42), A2 => n293, B1 => minusA(42), B2
                           => n287, ZN => n390);
   U44 : NAND2_X1 port map( A1 => n383, A2 => n382, ZN => n463);
   U45 : AOI22_X1 port map( A1 => plusA(38), A2 => n281, B1 => plus2A(38), B2 
                           => n275, ZN => n383);
   U46 : AOI22_X1 port map( A1 => minus2A(38), A2 => n293, B1 => minusA(38), B2
                           => n287, ZN => n382);
   U47 : NAND2_X1 port map( A1 => n375, A2 => n374, ZN => n467);
   U48 : AOI22_X1 port map( A1 => plusA(34), A2 => n280, B1 => plus2A(34), B2 
                           => n274, ZN => n375);
   U49 : AOI22_X1 port map( A1 => minus2A(34), A2 => n292, B1 => minusA(34), B2
                           => n286, ZN => n374);
   U50 : NAND2_X1 port map( A1 => n367, A2 => n366, ZN => n471);
   U51 : AOI22_X1 port map( A1 => plusA(30), A2 => n280, B1 => plus2A(30), B2 
                           => n274, ZN => n367);
   U52 : AOI22_X1 port map( A1 => minus2A(30), A2 => n292, B1 => minusA(30), B2
                           => n286, ZN => n366);
   U53 : NAND2_X1 port map( A1 => n437, A2 => n436, ZN => n438);
   U54 : AOI22_X1 port map( A1 => plusA(63), A2 => n283, B1 => plus2A(63), B2 
                           => n277, ZN => n437);
   U55 : AOI22_X1 port map( A1 => minus2A(63), A2 => n295, B1 => minusA(63), B2
                           => n289, ZN => n436);
   U56 : NAND2_X1 port map( A1 => n431, A2 => n430, ZN => n439);
   U57 : AOI22_X1 port map( A1 => plusA(62), A2 => n283, B1 => plus2A(62), B2 
                           => n277, ZN => n431);
   U58 : AOI22_X1 port map( A1 => minus2A(62), A2 => n295, B1 => minusA(62), B2
                           => n289, ZN => n430);
   U59 : NAND2_X1 port map( A1 => n429, A2 => n428, ZN => n440);
   U60 : AOI22_X1 port map( A1 => plusA(61), A2 => n283, B1 => plus2A(61), B2 
                           => n277, ZN => n429);
   U61 : AOI22_X1 port map( A1 => minus2A(61), A2 => n295, B1 => minusA(61), B2
                           => n289, ZN => n428);
   U62 : NAND2_X1 port map( A1 => n427, A2 => n426, ZN => n441);
   U63 : AOI22_X1 port map( A1 => plusA(60), A2 => n283, B1 => plus2A(60), B2 
                           => n277, ZN => n427);
   U64 : AOI22_X1 port map( A1 => minus2A(60), A2 => n295, B1 => minusA(60), B2
                           => n289, ZN => n426);
   U65 : NAND2_X1 port map( A1 => n425, A2 => n424, ZN => n442);
   U66 : AOI22_X1 port map( A1 => plusA(59), A2 => n282, B1 => plus2A(59), B2 
                           => n276, ZN => n425);
   U67 : AOI22_X1 port map( A1 => minus2A(59), A2 => n294, B1 => minusA(59), B2
                           => n288, ZN => n424);
   U68 : NAND2_X1 port map( A1 => n423, A2 => n422, ZN => n443);
   U69 : AOI22_X1 port map( A1 => plusA(58), A2 => n282, B1 => plus2A(58), B2 
                           => n276, ZN => n423);
   U70 : AOI22_X1 port map( A1 => minus2A(58), A2 => n294, B1 => minusA(58), B2
                           => n288, ZN => n422);
   U71 : NAND2_X1 port map( A1 => n421, A2 => n420, ZN => n444);
   U72 : AOI22_X1 port map( A1 => plusA(57), A2 => n282, B1 => plus2A(57), B2 
                           => n276, ZN => n421);
   U73 : AOI22_X1 port map( A1 => minus2A(57), A2 => n294, B1 => minusA(57), B2
                           => n288, ZN => n420);
   U74 : NAND2_X1 port map( A1 => n419, A2 => n418, ZN => n445);
   U75 : AOI22_X1 port map( A1 => plusA(56), A2 => n282, B1 => plus2A(56), B2 
                           => n276, ZN => n419);
   U76 : AOI22_X1 port map( A1 => minus2A(56), A2 => n294, B1 => minusA(56), B2
                           => n288, ZN => n418);
   U77 : NAND2_X1 port map( A1 => n417, A2 => n416, ZN => n446);
   U78 : AOI22_X1 port map( A1 => plusA(55), A2 => n282, B1 => plus2A(55), B2 
                           => n276, ZN => n417);
   U79 : AOI22_X1 port map( A1 => minus2A(55), A2 => n294, B1 => minusA(55), B2
                           => n288, ZN => n416);
   U80 : NAND2_X1 port map( A1 => n415, A2 => n414, ZN => n447);
   U81 : AOI22_X1 port map( A1 => plusA(54), A2 => n282, B1 => plus2A(54), B2 
                           => n276, ZN => n415);
   U82 : AOI22_X1 port map( A1 => minus2A(54), A2 => n294, B1 => minusA(54), B2
                           => n288, ZN => n414);
   U83 : NAND2_X1 port map( A1 => n413, A2 => n412, ZN => n448);
   U84 : AOI22_X1 port map( A1 => plusA(53), A2 => n282, B1 => plus2A(53), B2 
                           => n276, ZN => n413);
   U85 : AOI22_X1 port map( A1 => minus2A(53), A2 => n294, B1 => minusA(53), B2
                           => n288, ZN => n412);
   U86 : NAND2_X1 port map( A1 => n411, A2 => n410, ZN => n449);
   U87 : AOI22_X1 port map( A1 => plusA(52), A2 => n282, B1 => plus2A(52), B2 
                           => n276, ZN => n411);
   U88 : AOI22_X1 port map( A1 => minus2A(52), A2 => n294, B1 => minusA(52), B2
                           => n288, ZN => n410);
   U89 : NAND2_X1 port map( A1 => n409, A2 => n408, ZN => n450);
   U90 : AOI22_X1 port map( A1 => plusA(51), A2 => n282, B1 => plus2A(51), B2 
                           => n276, ZN => n409);
   U91 : AOI22_X1 port map( A1 => minus2A(51), A2 => n294, B1 => minusA(51), B2
                           => n288, ZN => n408);
   U92 : NAND2_X1 port map( A1 => n407, A2 => n406, ZN => n451);
   U93 : AOI22_X1 port map( A1 => plusA(50), A2 => n282, B1 => plus2A(50), B2 
                           => n276, ZN => n407);
   U94 : AOI22_X1 port map( A1 => minus2A(50), A2 => n294, B1 => minusA(50), B2
                           => n288, ZN => n406);
   U95 : NAND2_X1 port map( A1 => n405, A2 => n404, ZN => n452);
   U96 : AOI22_X1 port map( A1 => plusA(49), A2 => n282, B1 => plus2A(49), B2 
                           => n276, ZN => n405);
   U97 : AOI22_X1 port map( A1 => minus2A(49), A2 => n294, B1 => minusA(49), B2
                           => n288, ZN => n404);
   U98 : NAND2_X1 port map( A1 => n403, A2 => n402, ZN => n453);
   U99 : AOI22_X1 port map( A1 => plusA(48), A2 => n282, B1 => plus2A(48), B2 
                           => n276, ZN => n403);
   U100 : AOI22_X1 port map( A1 => minus2A(48), A2 => n294, B1 => minusA(48), 
                           B2 => n288, ZN => n402);
   U101 : NAND2_X1 port map( A1 => n401, A2 => n400, ZN => n454);
   U102 : AOI22_X1 port map( A1 => plusA(47), A2 => n281, B1 => plus2A(47), B2 
                           => n275, ZN => n401);
   U103 : AOI22_X1 port map( A1 => minus2A(47), A2 => n293, B1 => minusA(47), 
                           B2 => n287, ZN => n400);
   U104 : NAND2_X1 port map( A1 => n399, A2 => n398, ZN => n455);
   U105 : AOI22_X1 port map( A1 => plusA(46), A2 => n281, B1 => plus2A(46), B2 
                           => n275, ZN => n399);
   U106 : AOI22_X1 port map( A1 => minus2A(46), A2 => n293, B1 => minusA(46), 
                           B2 => n287, ZN => n398);
   U107 : BUF_X1 port map( A => n493, Z => n296);
   U108 : BUF_X1 port map( A => n493, Z => n297);
   U109 : BUF_X1 port map( A => n493, Z => n298);
   U110 : BUF_X1 port map( A => n433, Z => n280);
   U111 : BUF_X1 port map( A => n434, Z => n286);
   U112 : BUF_X1 port map( A => n432, Z => n274);
   U113 : BUF_X1 port map( A => n435, Z => n292);
   U114 : NAND2_X1 port map( A1 => n365, A2 => n364, ZN => n472);
   U115 : AOI22_X1 port map( A1 => plusA(29), A2 => n280, B1 => plus2A(29), B2 
                           => n274, ZN => n365);
   U116 : AOI22_X1 port map( A1 => minus2A(29), A2 => n292, B1 => minusA(29), 
                           B2 => n286, ZN => n364);
   U117 : NAND2_X1 port map( A1 => n363, A2 => n362, ZN => n473);
   U118 : AOI22_X1 port map( A1 => plusA(28), A2 => n280, B1 => plus2A(28), B2 
                           => n274, ZN => n363);
   U119 : AOI22_X1 port map( A1 => minus2A(28), A2 => n292, B1 => minusA(28), 
                           B2 => n286, ZN => n362);
   U120 : BUF_X1 port map( A => n493, Z => n299);
   U121 : BUF_X1 port map( A => n433, Z => n281);
   U122 : BUF_X1 port map( A => n434, Z => n287);
   U123 : BUF_X1 port map( A => n432, Z => n275);
   U124 : BUF_X1 port map( A => n435, Z => n293);
   U125 : BUF_X1 port map( A => n493, Z => n300);
   U126 : BUF_X1 port map( A => n433, Z => n282);
   U127 : BUF_X1 port map( A => n434, Z => n288);
   U128 : BUF_X1 port map( A => n432, Z => n276);
   U129 : BUF_X1 port map( A => n435, Z => n294);
   U130 : BUF_X1 port map( A => n433, Z => n279);
   U131 : BUF_X1 port map( A => n433, Z => n278);
   U132 : BUF_X1 port map( A => n434, Z => n285);
   U133 : BUF_X1 port map( A => n432, Z => n273);
   U134 : BUF_X1 port map( A => n434, Z => n284);
   U135 : BUF_X1 port map( A => n432, Z => n272);
   U136 : BUF_X1 port map( A => n435, Z => n291);
   U137 : BUF_X1 port map( A => n435, Z => n290);
   U138 : NOR2_X1 port map( A1 => n323, A2 => n304, ZN => n493);
   U139 : INV_X1 port map( A => SEL(2), ZN => n304);
   U140 : NOR2_X1 port map( A1 => SEL(1), A2 => SEL(0), ZN => n323);
   U141 : AND2_X1 port map( A1 => SEL(2), A2 => n323, ZN => n435);
   U142 : INV_X1 port map( A => SEL(1), ZN => n302);
   U143 : INV_X1 port map( A => SEL(0), ZN => n303);
   U144 : NAND2_X1 port map( A1 => n361, A2 => n360, ZN => n474);
   U145 : AOI22_X1 port map( A1 => plusA(27), A2 => n280, B1 => plus2A(27), B2 
                           => n274, ZN => n361);
   U146 : AOI22_X1 port map( A1 => minus2A(27), A2 => n292, B1 => minusA(27), 
                           B2 => n286, ZN => n360);
   U147 : NAND2_X1 port map( A1 => n359, A2 => n358, ZN => n475);
   U148 : AOI22_X1 port map( A1 => plusA(26), A2 => n280, B1 => plus2A(26), B2 
                           => n274, ZN => n359);
   U149 : AOI22_X1 port map( A1 => minus2A(26), A2 => n292, B1 => minusA(26), 
                           B2 => n286, ZN => n358);
   U150 : NAND2_X1 port map( A1 => n357, A2 => n356, ZN => n476);
   U151 : AOI22_X1 port map( A1 => plusA(25), A2 => n280, B1 => plus2A(25), B2 
                           => n274, ZN => n357);
   U152 : AOI22_X1 port map( A1 => minus2A(25), A2 => n292, B1 => minusA(25), 
                           B2 => n286, ZN => n356);
   U153 : NAND2_X1 port map( A1 => n353, A2 => n352, ZN => n478);
   U154 : AOI22_X1 port map( A1 => plusA(23), A2 => n279, B1 => plus2A(23), B2 
                           => n273, ZN => n353);
   U155 : AOI22_X1 port map( A1 => minus2A(23), A2 => n291, B1 => minusA(23), 
                           B2 => n285, ZN => n352);
   U156 : NAND2_X1 port map( A1 => n351, A2 => n350, ZN => n479);
   U157 : AOI22_X1 port map( A1 => plusA(22), A2 => n279, B1 => plus2A(22), B2 
                           => n273, ZN => n351);
   U158 : AOI22_X1 port map( A1 => minus2A(22), A2 => n291, B1 => minusA(22), 
                           B2 => n285, ZN => n350);
   U159 : NAND2_X1 port map( A1 => n349, A2 => n348, ZN => n480);
   U160 : AOI22_X1 port map( A1 => plusA(21), A2 => n279, B1 => plus2A(21), B2 
                           => n273, ZN => n349);
   U161 : AOI22_X1 port map( A1 => minus2A(21), A2 => n291, B1 => minusA(21), 
                           B2 => n285, ZN => n348);
   U162 : NAND2_X1 port map( A1 => n345, A2 => n344, ZN => n482);
   U163 : AOI22_X1 port map( A1 => plusA(19), A2 => n279, B1 => plus2A(19), B2 
                           => n273, ZN => n345);
   U164 : AOI22_X1 port map( A1 => minus2A(19), A2 => n291, B1 => minusA(19), 
                           B2 => n285, ZN => n344);
   U165 : NAND2_X1 port map( A1 => n343, A2 => n342, ZN => n483);
   U166 : AOI22_X1 port map( A1 => plusA(18), A2 => n279, B1 => plus2A(18), B2 
                           => n273, ZN => n343);
   U167 : AOI22_X1 port map( A1 => minus2A(18), A2 => n291, B1 => minusA(18), 
                           B2 => n285, ZN => n342);
   U168 : NAND2_X1 port map( A1 => n341, A2 => n340, ZN => n484);
   U169 : AOI22_X1 port map( A1 => plusA(17), A2 => n279, B1 => plus2A(17), B2 
                           => n273, ZN => n341);
   U170 : AOI22_X1 port map( A1 => minus2A(17), A2 => n291, B1 => minusA(17), 
                           B2 => n285, ZN => n340);
   U171 : NAND2_X1 port map( A1 => n337, A2 => n336, ZN => n486);
   U172 : AOI22_X1 port map( A1 => plusA(15), A2 => n279, B1 => plus2A(15), B2 
                           => n273, ZN => n337);
   U173 : AOI22_X1 port map( A1 => minus2A(15), A2 => n291, B1 => minusA(15), 
                           B2 => n285, ZN => n336);
   U174 : NAND2_X1 port map( A1 => n335, A2 => n334, ZN => n487);
   U175 : AOI22_X1 port map( A1 => plusA(14), A2 => n279, B1 => plus2A(14), B2 
                           => n273, ZN => n335);
   U176 : AOI22_X1 port map( A1 => minus2A(14), A2 => n291, B1 => minusA(14), 
                           B2 => n285, ZN => n334);
   U177 : NAND2_X1 port map( A1 => n333, A2 => n332, ZN => n488);
   U178 : AOI22_X1 port map( A1 => plusA(13), A2 => n279, B1 => plus2A(13), B2 
                           => n273, ZN => n333);
   U179 : AOI22_X1 port map( A1 => minus2A(13), A2 => n291, B1 => minusA(13), 
                           B2 => n285, ZN => n332);
   U180 : NAND2_X1 port map( A1 => n329, A2 => n328, ZN => n490);
   U181 : AOI22_X1 port map( A1 => plusA(11), A2 => n278, B1 => plus2A(11), B2 
                           => n272, ZN => n329);
   U182 : AOI22_X1 port map( A1 => minus2A(11), A2 => n290, B1 => minusA(11), 
                           B2 => n284, ZN => n328);
   U183 : NAND2_X1 port map( A1 => n327, A2 => n326, ZN => n491);
   U184 : AOI22_X1 port map( A1 => plusA(10), A2 => n278, B1 => plus2A(10), B2 
                           => n272, ZN => n327);
   U185 : AOI22_X1 port map( A1 => minus2A(10), A2 => n290, B1 => minusA(10), 
                           B2 => n284, ZN => n326);
   U186 : NAND2_X1 port map( A1 => n325, A2 => n324, ZN => n492);
   U187 : AOI22_X1 port map( A1 => plusA(9), A2 => n278, B1 => plus2A(9), B2 =>
                           n272, ZN => n325);
   U188 : AOI22_X1 port map( A1 => minus2A(9), A2 => n290, B1 => minusA(9), B2 
                           => n284, ZN => n324);
   U189 : NAND2_X1 port map( A1 => n320, A2 => n319, ZN => n495);
   U190 : AOI22_X1 port map( A1 => plusA(7), A2 => n278, B1 => plus2A(7), B2 =>
                           n272, ZN => n320);
   U191 : AOI22_X1 port map( A1 => minus2A(7), A2 => n290, B1 => minusA(7), B2 
                           => n284, ZN => n319);
   U192 : NAND2_X1 port map( A1 => n318, A2 => n317, ZN => n496);
   U193 : AOI22_X1 port map( A1 => plusA(6), A2 => n278, B1 => plus2A(6), B2 =>
                           n272, ZN => n318);
   U194 : AOI22_X1 port map( A1 => minus2A(6), A2 => n290, B1 => minusA(6), B2 
                           => n284, ZN => n317);
   U195 : NAND2_X1 port map( A1 => n316, A2 => n315, ZN => n497);
   U196 : AOI22_X1 port map( A1 => plusA(5), A2 => n278, B1 => plus2A(5), B2 =>
                           n272, ZN => n316);
   U197 : AOI22_X1 port map( A1 => minus2A(5), A2 => n290, B1 => minusA(5), B2 
                           => n284, ZN => n315);
   U198 : NAND2_X1 port map( A1 => n312, A2 => n311, ZN => n499);
   U199 : AOI22_X1 port map( A1 => plusA(3), A2 => n278, B1 => plus2A(3), B2 =>
                           n272, ZN => n312);
   U200 : AOI22_X1 port map( A1 => minus2A(3), A2 => n290, B1 => minusA(3), B2 
                           => n284, ZN => n311);
   U201 : NAND2_X1 port map( A1 => n355, A2 => n354, ZN => n477);
   U202 : AOI22_X1 port map( A1 => plusA(24), A2 => n280, B1 => plus2A(24), B2 
                           => n274, ZN => n355);
   U203 : AOI22_X1 port map( A1 => minus2A(24), A2 => n292, B1 => minusA(24), 
                           B2 => n286, ZN => n354);
   U204 : NAND2_X1 port map( A1 => n347, A2 => n346, ZN => n481);
   U205 : AOI22_X1 port map( A1 => plusA(20), A2 => n279, B1 => plus2A(20), B2 
                           => n273, ZN => n347);
   U206 : AOI22_X1 port map( A1 => minus2A(20), A2 => n291, B1 => minusA(20), 
                           B2 => n285, ZN => n346);
   U207 : NAND2_X1 port map( A1 => n339, A2 => n338, ZN => n485);
   U208 : AOI22_X1 port map( A1 => plusA(16), A2 => n279, B1 => plus2A(16), B2 
                           => n273, ZN => n339);
   U209 : AOI22_X1 port map( A1 => minus2A(16), A2 => n291, B1 => minusA(16), 
                           B2 => n285, ZN => n338);
   U210 : NAND2_X1 port map( A1 => n331, A2 => n330, ZN => n489);
   U211 : AOI22_X1 port map( A1 => plusA(12), A2 => n279, B1 => plus2A(12), B2 
                           => n273, ZN => n331);
   U212 : AOI22_X1 port map( A1 => minus2A(12), A2 => n291, B1 => minusA(12), 
                           B2 => n285, ZN => n330);
   U213 : NAND2_X1 port map( A1 => n322, A2 => n321, ZN => n494);
   U214 : AOI22_X1 port map( A1 => plusA(8), A2 => n278, B1 => plus2A(8), B2 =>
                           n272, ZN => n322);
   U215 : AOI22_X1 port map( A1 => minus2A(8), A2 => n290, B1 => minusA(8), B2 
                           => n284, ZN => n321);
   U216 : NAND2_X1 port map( A1 => n314, A2 => n313, ZN => n498);
   U217 : AOI22_X1 port map( A1 => plusA(4), A2 => n278, B1 => plus2A(4), B2 =>
                           n272, ZN => n314);
   U218 : AOI22_X1 port map( A1 => minus2A(4), A2 => n290, B1 => minusA(4), B2 
                           => n284, ZN => n313);
   U219 : NAND2_X1 port map( A1 => n310, A2 => n309, ZN => n500);
   U220 : AOI22_X1 port map( A1 => plusA(2), A2 => n278, B1 => plus2A(2), B2 =>
                           n272, ZN => n310);
   U221 : AOI22_X1 port map( A1 => minus2A(2), A2 => n290, B1 => minusA(2), B2 
                           => n284, ZN => n309);
   U222 : NAND2_X1 port map( A1 => n308, A2 => n307, ZN => n501);
   U223 : AOI22_X1 port map( A1 => plusA(1), A2 => n278, B1 => plus2A(1), B2 =>
                           n272, ZN => n308);
   U224 : AOI22_X1 port map( A1 => minus2A(1), A2 => n290, B1 => minusA(1), B2 
                           => n284, ZN => n307);
   U225 : NAND2_X1 port map( A1 => n306, A2 => n305, ZN => n502);
   U226 : AOI22_X1 port map( A1 => plusA(0), A2 => n278, B1 => plus2A(0), B2 =>
                           n272, ZN => n306);
   U227 : AOI22_X1 port map( A1 => minus2A(0), A2 => n290, B1 => minusA(0), B2 
                           => n284, ZN => n305);
   U228 : CLKBUF_X1 port map( A => n432, Z => n277);
   U229 : CLKBUF_X1 port map( A => n433, Z => n283);
   U230 : CLKBUF_X1 port map( A => n434, Z => n289);
   U231 : CLKBUF_X1 port map( A => n435, Z => n295);
   U232 : CLKBUF_X1 port map( A => n493, Z => n301);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity MUX_GENERIC_N64_RADIX3_2 is

   port( plusA, minusA, plus2A, minus2A : in std_logic_vector (63 downto 0);  
         SEL : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (63 
         downto 0));

end MUX_GENERIC_N64_RADIX3_2;

architecture SYN_beh of MUX_GENERIC_N64_RADIX3_2 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component TBUF_X1
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   signal n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, 
      n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, 
      n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, 
      n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, 
      n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, 
      n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, 
      n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, 
      n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, 
      n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, 
      n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, 
      n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, 
      n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, 
      n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, 
      n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, 
      n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, 
      n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, 
      n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, 
      n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, 
      n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, 
      n499, n500, n501, n502 : std_logic;

begin
   
   Y_tri_60_inst : TBUF_X1 port map( A => n441, EN => n301, Z => Y(60));
   Y_tri_61_inst : TBUF_X1 port map( A => n440, EN => n301, Z => Y(61));
   Y_tri_62_inst : TBUF_X1 port map( A => n439, EN => n301, Z => Y(62));
   Y_tri_63_inst : TBUF_X1 port map( A => n438, EN => n301, Z => Y(63));
   Y_tri_42_inst : TBUF_X1 port map( A => n459, EN => n299, Z => Y(42));
   Y_tri_43_inst : TBUF_X1 port map( A => n458, EN => n299, Z => Y(43));
   Y_tri_44_inst : TBUF_X1 port map( A => n457, EN => n299, Z => Y(44));
   Y_tri_45_inst : TBUF_X1 port map( A => n456, EN => n299, Z => Y(45));
   Y_tri_46_inst : TBUF_X1 port map( A => n455, EN => n299, Z => Y(46));
   Y_tri_47_inst : TBUF_X1 port map( A => n454, EN => n299, Z => Y(47));
   Y_tri_48_inst : TBUF_X1 port map( A => n453, EN => n300, Z => Y(48));
   Y_tri_49_inst : TBUF_X1 port map( A => n452, EN => n300, Z => Y(49));
   Y_tri_50_inst : TBUF_X1 port map( A => n451, EN => n300, Z => Y(50));
   Y_tri_51_inst : TBUF_X1 port map( A => n450, EN => n300, Z => Y(51));
   Y_tri_52_inst : TBUF_X1 port map( A => n449, EN => n300, Z => Y(52));
   Y_tri_53_inst : TBUF_X1 port map( A => n448, EN => n300, Z => Y(53));
   Y_tri_54_inst : TBUF_X1 port map( A => n447, EN => n300, Z => Y(54));
   Y_tri_55_inst : TBUF_X1 port map( A => n446, EN => n300, Z => Y(55));
   Y_tri_56_inst : TBUF_X1 port map( A => n445, EN => n300, Z => Y(56));
   Y_tri_57_inst : TBUF_X1 port map( A => n444, EN => n300, Z => Y(57));
   Y_tri_58_inst : TBUF_X1 port map( A => n443, EN => n300, Z => Y(58));
   Y_tri_59_inst : TBUF_X1 port map( A => n442, EN => n300, Z => Y(59));
   Y_tri_17_inst : TBUF_X1 port map( A => n484, EN => n297, Z => Y(17));
   Y_tri_18_inst : TBUF_X1 port map( A => n483, EN => n297, Z => Y(18));
   Y_tri_19_inst : TBUF_X1 port map( A => n482, EN => n297, Z => Y(19));
   Y_tri_20_inst : TBUF_X1 port map( A => n481, EN => n297, Z => Y(20));
   Y_tri_21_inst : TBUF_X1 port map( A => n480, EN => n297, Z => Y(21));
   Y_tri_22_inst : TBUF_X1 port map( A => n479, EN => n297, Z => Y(22));
   Y_tri_23_inst : TBUF_X1 port map( A => n478, EN => n297, Z => Y(23));
   Y_tri_24_inst : TBUF_X1 port map( A => n477, EN => n298, Z => Y(24));
   Y_tri_25_inst : TBUF_X1 port map( A => n476, EN => n298, Z => Y(25));
   Y_tri_26_inst : TBUF_X1 port map( A => n475, EN => n298, Z => Y(26));
   Y_tri_27_inst : TBUF_X1 port map( A => n474, EN => n298, Z => Y(27));
   Y_tri_28_inst : TBUF_X1 port map( A => n473, EN => n298, Z => Y(28));
   Y_tri_29_inst : TBUF_X1 port map( A => n472, EN => n298, Z => Y(29));
   Y_tri_30_inst : TBUF_X1 port map( A => n471, EN => n298, Z => Y(30));
   Y_tri_31_inst : TBUF_X1 port map( A => n470, EN => n298, Z => Y(31));
   Y_tri_32_inst : TBUF_X1 port map( A => n469, EN => n298, Z => Y(32));
   Y_tri_33_inst : TBUF_X1 port map( A => n468, EN => n298, Z => Y(33));
   Y_tri_34_inst : TBUF_X1 port map( A => n467, EN => n298, Z => Y(34));
   Y_tri_35_inst : TBUF_X1 port map( A => n466, EN => n298, Z => Y(35));
   Y_tri_36_inst : TBUF_X1 port map( A => n465, EN => n299, Z => Y(36));
   Y_tri_37_inst : TBUF_X1 port map( A => n464, EN => n299, Z => Y(37));
   Y_tri_38_inst : TBUF_X1 port map( A => n463, EN => n299, Z => Y(38));
   Y_tri_39_inst : TBUF_X1 port map( A => n462, EN => n299, Z => Y(39));
   Y_tri_40_inst : TBUF_X1 port map( A => n461, EN => n299, Z => Y(40));
   Y_tri_41_inst : TBUF_X1 port map( A => n460, EN => n299, Z => Y(41));
   Y_tri_6_inst : TBUF_X1 port map( A => n496, EN => n296, Z => Y(6));
   Y_tri_7_inst : TBUF_X1 port map( A => n495, EN => n296, Z => Y(7));
   Y_tri_8_inst : TBUF_X1 port map( A => n494, EN => n296, Z => Y(8));
   Y_tri_9_inst : TBUF_X1 port map( A => n492, EN => n296, Z => Y(9));
   Y_tri_10_inst : TBUF_X1 port map( A => n491, EN => n296, Z => Y(10));
   Y_tri_11_inst : TBUF_X1 port map( A => n490, EN => n296, Z => Y(11));
   Y_tri_12_inst : TBUF_X1 port map( A => n489, EN => n297, Z => Y(12));
   Y_tri_13_inst : TBUF_X1 port map( A => n488, EN => n297, Z => Y(13));
   Y_tri_14_inst : TBUF_X1 port map( A => n487, EN => n297, Z => Y(14));
   Y_tri_15_inst : TBUF_X1 port map( A => n486, EN => n297, Z => Y(15));
   Y_tri_16_inst : TBUF_X1 port map( A => n485, EN => n297, Z => Y(16));
   Y_tri_0_inst : TBUF_X1 port map( A => n502, EN => n296, Z => Y(0));
   Y_tri_1_inst : TBUF_X1 port map( A => n501, EN => n296, Z => Y(1));
   Y_tri_2_inst : TBUF_X1 port map( A => n500, EN => n296, Z => Y(2));
   Y_tri_3_inst : TBUF_X1 port map( A => n499, EN => n296, Z => Y(3));
   Y_tri_4_inst : TBUF_X1 port map( A => n498, EN => n296, Z => Y(4));
   Y_tri_5_inst : TBUF_X1 port map( A => n497, EN => n296, Z => Y(5));
   U2 : NOR3_X1 port map( A1 => SEL(0), A2 => SEL(2), A3 => n302, ZN => n434);
   U3 : NOR3_X1 port map( A1 => n302, A2 => SEL(2), A3 => n303, ZN => n432);
   U4 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n303, ZN => n433);
   U5 : NAND2_X1 port map( A1 => n389, A2 => n388, ZN => n460);
   U6 : AOI22_X1 port map( A1 => plusA(41), A2 => n281, B1 => plus2A(41), B2 =>
                           n275, ZN => n389);
   U7 : AOI22_X1 port map( A1 => minus2A(41), A2 => n293, B1 => minusA(41), B2 
                           => n287, ZN => n388);
   U8 : NAND2_X1 port map( A1 => n387, A2 => n386, ZN => n461);
   U9 : AOI22_X1 port map( A1 => plusA(40), A2 => n281, B1 => plus2A(40), B2 =>
                           n275, ZN => n387);
   U10 : AOI22_X1 port map( A1 => minus2A(40), A2 => n293, B1 => minusA(40), B2
                           => n287, ZN => n386);
   U11 : NAND2_X1 port map( A1 => n385, A2 => n384, ZN => n462);
   U12 : AOI22_X1 port map( A1 => plusA(39), A2 => n281, B1 => plus2A(39), B2 
                           => n275, ZN => n385);
   U13 : AOI22_X1 port map( A1 => minus2A(39), A2 => n293, B1 => minusA(39), B2
                           => n287, ZN => n384);
   U14 : NAND2_X1 port map( A1 => n379, A2 => n378, ZN => n465);
   U15 : AOI22_X1 port map( A1 => plusA(36), A2 => n281, B1 => plus2A(36), B2 
                           => n275, ZN => n379);
   U16 : AOI22_X1 port map( A1 => minus2A(36), A2 => n293, B1 => minusA(36), B2
                           => n287, ZN => n378);
   U17 : NAND2_X1 port map( A1 => n377, A2 => n376, ZN => n466);
   U18 : AOI22_X1 port map( A1 => plusA(35), A2 => n280, B1 => plus2A(35), B2 
                           => n274, ZN => n377);
   U19 : AOI22_X1 port map( A1 => minus2A(35), A2 => n292, B1 => minusA(35), B2
                           => n286, ZN => n376);
   U20 : NAND2_X1 port map( A1 => n381, A2 => n380, ZN => n464);
   U21 : AOI22_X1 port map( A1 => plusA(37), A2 => n281, B1 => plus2A(37), B2 
                           => n275, ZN => n381);
   U22 : AOI22_X1 port map( A1 => minus2A(37), A2 => n293, B1 => minusA(37), B2
                           => n287, ZN => n380);
   U23 : NAND2_X1 port map( A1 => n373, A2 => n372, ZN => n468);
   U24 : AOI22_X1 port map( A1 => plusA(33), A2 => n280, B1 => plus2A(33), B2 
                           => n274, ZN => n373);
   U25 : AOI22_X1 port map( A1 => minus2A(33), A2 => n292, B1 => minusA(33), B2
                           => n286, ZN => n372);
   U26 : NAND2_X1 port map( A1 => n383, A2 => n382, ZN => n463);
   U27 : AOI22_X1 port map( A1 => plusA(38), A2 => n281, B1 => plus2A(38), B2 
                           => n275, ZN => n383);
   U28 : AOI22_X1 port map( A1 => minus2A(38), A2 => n293, B1 => minusA(38), B2
                           => n287, ZN => n382);
   U29 : NAND2_X1 port map( A1 => n375, A2 => n374, ZN => n467);
   U30 : AOI22_X1 port map( A1 => plusA(34), A2 => n280, B1 => plus2A(34), B2 
                           => n274, ZN => n375);
   U31 : AOI22_X1 port map( A1 => minus2A(34), A2 => n292, B1 => minusA(34), B2
                           => n286, ZN => n374);
   U32 : NAND2_X1 port map( A1 => n371, A2 => n370, ZN => n469);
   U33 : AOI22_X1 port map( A1 => plusA(32), A2 => n280, B1 => plus2A(32), B2 
                           => n274, ZN => n371);
   U34 : AOI22_X1 port map( A1 => minus2A(32), A2 => n292, B1 => minusA(32), B2
                           => n286, ZN => n370);
   U35 : NAND2_X1 port map( A1 => n437, A2 => n436, ZN => n438);
   U36 : AOI22_X1 port map( A1 => plusA(63), A2 => n283, B1 => plus2A(63), B2 
                           => n277, ZN => n437);
   U37 : AOI22_X1 port map( A1 => minus2A(63), A2 => n295, B1 => minusA(63), B2
                           => n289, ZN => n436);
   U38 : NAND2_X1 port map( A1 => n431, A2 => n430, ZN => n439);
   U39 : AOI22_X1 port map( A1 => plusA(62), A2 => n283, B1 => plus2A(62), B2 
                           => n277, ZN => n431);
   U40 : AOI22_X1 port map( A1 => minus2A(62), A2 => n295, B1 => minusA(62), B2
                           => n289, ZN => n430);
   U41 : NAND2_X1 port map( A1 => n429, A2 => n428, ZN => n440);
   U42 : AOI22_X1 port map( A1 => plusA(61), A2 => n283, B1 => plus2A(61), B2 
                           => n277, ZN => n429);
   U43 : AOI22_X1 port map( A1 => minus2A(61), A2 => n295, B1 => minusA(61), B2
                           => n289, ZN => n428);
   U44 : NAND2_X1 port map( A1 => n427, A2 => n426, ZN => n441);
   U45 : AOI22_X1 port map( A1 => plusA(60), A2 => n283, B1 => plus2A(60), B2 
                           => n277, ZN => n427);
   U46 : AOI22_X1 port map( A1 => minus2A(60), A2 => n295, B1 => minusA(60), B2
                           => n289, ZN => n426);
   U47 : NAND2_X1 port map( A1 => n425, A2 => n424, ZN => n442);
   U48 : AOI22_X1 port map( A1 => plusA(59), A2 => n282, B1 => plus2A(59), B2 
                           => n276, ZN => n425);
   U49 : AOI22_X1 port map( A1 => minus2A(59), A2 => n294, B1 => minusA(59), B2
                           => n288, ZN => n424);
   U50 : NAND2_X1 port map( A1 => n423, A2 => n422, ZN => n443);
   U51 : AOI22_X1 port map( A1 => plusA(58), A2 => n282, B1 => plus2A(58), B2 
                           => n276, ZN => n423);
   U52 : AOI22_X1 port map( A1 => minus2A(58), A2 => n294, B1 => minusA(58), B2
                           => n288, ZN => n422);
   U53 : NAND2_X1 port map( A1 => n421, A2 => n420, ZN => n444);
   U54 : AOI22_X1 port map( A1 => plusA(57), A2 => n282, B1 => plus2A(57), B2 
                           => n276, ZN => n421);
   U55 : AOI22_X1 port map( A1 => minus2A(57), A2 => n294, B1 => minusA(57), B2
                           => n288, ZN => n420);
   U56 : NAND2_X1 port map( A1 => n419, A2 => n418, ZN => n445);
   U57 : AOI22_X1 port map( A1 => plusA(56), A2 => n282, B1 => plus2A(56), B2 
                           => n276, ZN => n419);
   U58 : AOI22_X1 port map( A1 => minus2A(56), A2 => n294, B1 => minusA(56), B2
                           => n288, ZN => n418);
   U59 : NAND2_X1 port map( A1 => n417, A2 => n416, ZN => n446);
   U60 : AOI22_X1 port map( A1 => plusA(55), A2 => n282, B1 => plus2A(55), B2 
                           => n276, ZN => n417);
   U61 : AOI22_X1 port map( A1 => minus2A(55), A2 => n294, B1 => minusA(55), B2
                           => n288, ZN => n416);
   U62 : NAND2_X1 port map( A1 => n415, A2 => n414, ZN => n447);
   U63 : AOI22_X1 port map( A1 => plusA(54), A2 => n282, B1 => plus2A(54), B2 
                           => n276, ZN => n415);
   U64 : AOI22_X1 port map( A1 => minus2A(54), A2 => n294, B1 => minusA(54), B2
                           => n288, ZN => n414);
   U65 : NAND2_X1 port map( A1 => n413, A2 => n412, ZN => n448);
   U66 : AOI22_X1 port map( A1 => plusA(53), A2 => n282, B1 => plus2A(53), B2 
                           => n276, ZN => n413);
   U67 : AOI22_X1 port map( A1 => minus2A(53), A2 => n294, B1 => minusA(53), B2
                           => n288, ZN => n412);
   U68 : NAND2_X1 port map( A1 => n411, A2 => n410, ZN => n449);
   U69 : AOI22_X1 port map( A1 => plusA(52), A2 => n282, B1 => plus2A(52), B2 
                           => n276, ZN => n411);
   U70 : AOI22_X1 port map( A1 => minus2A(52), A2 => n294, B1 => minusA(52), B2
                           => n288, ZN => n410);
   U71 : NAND2_X1 port map( A1 => n409, A2 => n408, ZN => n450);
   U72 : AOI22_X1 port map( A1 => plusA(51), A2 => n282, B1 => plus2A(51), B2 
                           => n276, ZN => n409);
   U73 : AOI22_X1 port map( A1 => minus2A(51), A2 => n294, B1 => minusA(51), B2
                           => n288, ZN => n408);
   U74 : NAND2_X1 port map( A1 => n407, A2 => n406, ZN => n451);
   U75 : AOI22_X1 port map( A1 => plusA(50), A2 => n282, B1 => plus2A(50), B2 
                           => n276, ZN => n407);
   U76 : AOI22_X1 port map( A1 => minus2A(50), A2 => n294, B1 => minusA(50), B2
                           => n288, ZN => n406);
   U77 : NAND2_X1 port map( A1 => n405, A2 => n404, ZN => n452);
   U78 : AOI22_X1 port map( A1 => plusA(49), A2 => n282, B1 => plus2A(49), B2 
                           => n276, ZN => n405);
   U79 : AOI22_X1 port map( A1 => minus2A(49), A2 => n294, B1 => minusA(49), B2
                           => n288, ZN => n404);
   U80 : NAND2_X1 port map( A1 => n403, A2 => n402, ZN => n453);
   U81 : AOI22_X1 port map( A1 => plusA(48), A2 => n282, B1 => plus2A(48), B2 
                           => n276, ZN => n403);
   U82 : AOI22_X1 port map( A1 => minus2A(48), A2 => n294, B1 => minusA(48), B2
                           => n288, ZN => n402);
   U83 : NAND2_X1 port map( A1 => n401, A2 => n400, ZN => n454);
   U84 : AOI22_X1 port map( A1 => plusA(47), A2 => n281, B1 => plus2A(47), B2 
                           => n275, ZN => n401);
   U85 : AOI22_X1 port map( A1 => minus2A(47), A2 => n293, B1 => minusA(47), B2
                           => n287, ZN => n400);
   U86 : NAND2_X1 port map( A1 => n399, A2 => n398, ZN => n455);
   U87 : AOI22_X1 port map( A1 => plusA(46), A2 => n281, B1 => plus2A(46), B2 
                           => n275, ZN => n399);
   U88 : AOI22_X1 port map( A1 => minus2A(46), A2 => n293, B1 => minusA(46), B2
                           => n287, ZN => n398);
   U89 : NAND2_X1 port map( A1 => n397, A2 => n396, ZN => n456);
   U90 : AOI22_X1 port map( A1 => plusA(45), A2 => n281, B1 => plus2A(45), B2 
                           => n275, ZN => n397);
   U91 : AOI22_X1 port map( A1 => minus2A(45), A2 => n293, B1 => minusA(45), B2
                           => n287, ZN => n396);
   U92 : NAND2_X1 port map( A1 => n391, A2 => n390, ZN => n459);
   U93 : AOI22_X1 port map( A1 => plusA(42), A2 => n281, B1 => plus2A(42), B2 
                           => n275, ZN => n391);
   U94 : AOI22_X1 port map( A1 => minus2A(42), A2 => n293, B1 => minusA(42), B2
                           => n287, ZN => n390);
   U95 : NAND2_X1 port map( A1 => n393, A2 => n392, ZN => n458);
   U96 : AOI22_X1 port map( A1 => plusA(43), A2 => n281, B1 => plus2A(43), B2 
                           => n275, ZN => n393);
   U97 : AOI22_X1 port map( A1 => minus2A(43), A2 => n293, B1 => minusA(43), B2
                           => n287, ZN => n392);
   U98 : NAND2_X1 port map( A1 => n395, A2 => n394, ZN => n457);
   U99 : AOI22_X1 port map( A1 => plusA(44), A2 => n281, B1 => plus2A(44), B2 
                           => n275, ZN => n395);
   U100 : AOI22_X1 port map( A1 => minus2A(44), A2 => n293, B1 => minusA(44), 
                           B2 => n287, ZN => n394);
   U101 : BUF_X1 port map( A => n493, Z => n296);
   U102 : BUF_X1 port map( A => n493, Z => n297);
   U103 : BUF_X1 port map( A => n493, Z => n298);
   U104 : BUF_X1 port map( A => n433, Z => n280);
   U105 : BUF_X1 port map( A => n434, Z => n286);
   U106 : NAND2_X1 port map( A1 => n369, A2 => n368, ZN => n470);
   U107 : AOI22_X1 port map( A1 => plusA(31), A2 => n280, B1 => plus2A(31), B2 
                           => n274, ZN => n369);
   U108 : AOI22_X1 port map( A1 => minus2A(31), A2 => n292, B1 => minusA(31), 
                           B2 => n286, ZN => n368);
   U109 : NAND2_X1 port map( A1 => n367, A2 => n366, ZN => n471);
   U110 : AOI22_X1 port map( A1 => plusA(30), A2 => n280, B1 => plus2A(30), B2 
                           => n274, ZN => n367);
   U111 : AOI22_X1 port map( A1 => minus2A(30), A2 => n292, B1 => minusA(30), 
                           B2 => n286, ZN => n366);
   U112 : BUF_X1 port map( A => n493, Z => n299);
   U113 : BUF_X1 port map( A => n433, Z => n281);
   U114 : BUF_X1 port map( A => n434, Z => n287);
   U115 : BUF_X1 port map( A => n432, Z => n275);
   U116 : BUF_X1 port map( A => n432, Z => n274);
   U117 : BUF_X1 port map( A => n435, Z => n293);
   U118 : BUF_X1 port map( A => n435, Z => n292);
   U119 : BUF_X1 port map( A => n493, Z => n300);
   U120 : BUF_X1 port map( A => n433, Z => n282);
   U121 : BUF_X1 port map( A => n434, Z => n288);
   U122 : BUF_X1 port map( A => n432, Z => n276);
   U123 : BUF_X1 port map( A => n435, Z => n294);
   U124 : BUF_X1 port map( A => n433, Z => n279);
   U125 : BUF_X1 port map( A => n433, Z => n278);
   U126 : BUF_X1 port map( A => n434, Z => n285);
   U127 : BUF_X1 port map( A => n432, Z => n273);
   U128 : BUF_X1 port map( A => n434, Z => n284);
   U129 : BUF_X1 port map( A => n432, Z => n272);
   U130 : BUF_X1 port map( A => n435, Z => n291);
   U131 : BUF_X1 port map( A => n435, Z => n290);
   U132 : NOR2_X1 port map( A1 => n323, A2 => n304, ZN => n493);
   U133 : INV_X1 port map( A => SEL(2), ZN => n304);
   U134 : NOR2_X1 port map( A1 => SEL(1), A2 => SEL(0), ZN => n323);
   U135 : INV_X1 port map( A => SEL(1), ZN => n302);
   U136 : INV_X1 port map( A => SEL(0), ZN => n303);
   U137 : NAND2_X1 port map( A1 => n365, A2 => n364, ZN => n472);
   U138 : AOI22_X1 port map( A1 => plusA(29), A2 => n280, B1 => plus2A(29), B2 
                           => n274, ZN => n365);
   U139 : AOI22_X1 port map( A1 => minus2A(29), A2 => n292, B1 => minusA(29), 
                           B2 => n286, ZN => n364);
   U140 : AND2_X1 port map( A1 => SEL(2), A2 => n323, ZN => n435);
   U141 : NAND2_X1 port map( A1 => n363, A2 => n362, ZN => n473);
   U142 : AOI22_X1 port map( A1 => plusA(28), A2 => n280, B1 => plus2A(28), B2 
                           => n274, ZN => n363);
   U143 : AOI22_X1 port map( A1 => minus2A(28), A2 => n292, B1 => minusA(28), 
                           B2 => n286, ZN => n362);
   U144 : NAND2_X1 port map( A1 => n361, A2 => n360, ZN => n474);
   U145 : AOI22_X1 port map( A1 => plusA(27), A2 => n280, B1 => plus2A(27), B2 
                           => n274, ZN => n361);
   U146 : AOI22_X1 port map( A1 => minus2A(27), A2 => n292, B1 => minusA(27), 
                           B2 => n286, ZN => n360);
   U147 : NAND2_X1 port map( A1 => n359, A2 => n358, ZN => n475);
   U148 : AOI22_X1 port map( A1 => plusA(26), A2 => n280, B1 => plus2A(26), B2 
                           => n274, ZN => n359);
   U149 : AOI22_X1 port map( A1 => minus2A(26), A2 => n292, B1 => minusA(26), 
                           B2 => n286, ZN => n358);
   U150 : NAND2_X1 port map( A1 => n357, A2 => n356, ZN => n476);
   U151 : AOI22_X1 port map( A1 => plusA(25), A2 => n280, B1 => plus2A(25), B2 
                           => n274, ZN => n357);
   U152 : AOI22_X1 port map( A1 => minus2A(25), A2 => n292, B1 => minusA(25), 
                           B2 => n286, ZN => n356);
   U153 : NAND2_X1 port map( A1 => n353, A2 => n352, ZN => n478);
   U154 : AOI22_X1 port map( A1 => plusA(23), A2 => n279, B1 => plus2A(23), B2 
                           => n273, ZN => n353);
   U155 : AOI22_X1 port map( A1 => minus2A(23), A2 => n291, B1 => minusA(23), 
                           B2 => n285, ZN => n352);
   U156 : NAND2_X1 port map( A1 => n351, A2 => n350, ZN => n479);
   U157 : AOI22_X1 port map( A1 => plusA(22), A2 => n279, B1 => plus2A(22), B2 
                           => n273, ZN => n351);
   U158 : AOI22_X1 port map( A1 => minus2A(22), A2 => n291, B1 => minusA(22), 
                           B2 => n285, ZN => n350);
   U159 : NAND2_X1 port map( A1 => n349, A2 => n348, ZN => n480);
   U160 : AOI22_X1 port map( A1 => plusA(21), A2 => n279, B1 => plus2A(21), B2 
                           => n273, ZN => n349);
   U161 : AOI22_X1 port map( A1 => minus2A(21), A2 => n291, B1 => minusA(21), 
                           B2 => n285, ZN => n348);
   U162 : NAND2_X1 port map( A1 => n345, A2 => n344, ZN => n482);
   U163 : AOI22_X1 port map( A1 => plusA(19), A2 => n279, B1 => plus2A(19), B2 
                           => n273, ZN => n345);
   U164 : AOI22_X1 port map( A1 => minus2A(19), A2 => n291, B1 => minusA(19), 
                           B2 => n285, ZN => n344);
   U165 : NAND2_X1 port map( A1 => n343, A2 => n342, ZN => n483);
   U166 : AOI22_X1 port map( A1 => plusA(18), A2 => n279, B1 => plus2A(18), B2 
                           => n273, ZN => n343);
   U167 : AOI22_X1 port map( A1 => minus2A(18), A2 => n291, B1 => minusA(18), 
                           B2 => n285, ZN => n342);
   U168 : NAND2_X1 port map( A1 => n341, A2 => n340, ZN => n484);
   U169 : AOI22_X1 port map( A1 => plusA(17), A2 => n279, B1 => plus2A(17), B2 
                           => n273, ZN => n341);
   U170 : AOI22_X1 port map( A1 => minus2A(17), A2 => n291, B1 => minusA(17), 
                           B2 => n285, ZN => n340);
   U171 : NAND2_X1 port map( A1 => n337, A2 => n336, ZN => n486);
   U172 : AOI22_X1 port map( A1 => plusA(15), A2 => n279, B1 => plus2A(15), B2 
                           => n273, ZN => n337);
   U173 : AOI22_X1 port map( A1 => minus2A(15), A2 => n291, B1 => minusA(15), 
                           B2 => n285, ZN => n336);
   U174 : NAND2_X1 port map( A1 => n335, A2 => n334, ZN => n487);
   U175 : AOI22_X1 port map( A1 => plusA(14), A2 => n279, B1 => plus2A(14), B2 
                           => n273, ZN => n335);
   U176 : AOI22_X1 port map( A1 => minus2A(14), A2 => n291, B1 => minusA(14), 
                           B2 => n285, ZN => n334);
   U177 : NAND2_X1 port map( A1 => n333, A2 => n332, ZN => n488);
   U178 : AOI22_X1 port map( A1 => plusA(13), A2 => n279, B1 => plus2A(13), B2 
                           => n273, ZN => n333);
   U179 : AOI22_X1 port map( A1 => minus2A(13), A2 => n291, B1 => minusA(13), 
                           B2 => n285, ZN => n332);
   U180 : NAND2_X1 port map( A1 => n329, A2 => n328, ZN => n490);
   U181 : AOI22_X1 port map( A1 => plusA(11), A2 => n278, B1 => plus2A(11), B2 
                           => n272, ZN => n329);
   U182 : AOI22_X1 port map( A1 => minus2A(11), A2 => n290, B1 => minusA(11), 
                           B2 => n284, ZN => n328);
   U183 : NAND2_X1 port map( A1 => n327, A2 => n326, ZN => n491);
   U184 : AOI22_X1 port map( A1 => plusA(10), A2 => n278, B1 => plus2A(10), B2 
                           => n272, ZN => n327);
   U185 : AOI22_X1 port map( A1 => minus2A(10), A2 => n290, B1 => minusA(10), 
                           B2 => n284, ZN => n326);
   U186 : NAND2_X1 port map( A1 => n325, A2 => n324, ZN => n492);
   U187 : AOI22_X1 port map( A1 => plusA(9), A2 => n278, B1 => plus2A(9), B2 =>
                           n272, ZN => n325);
   U188 : AOI22_X1 port map( A1 => minus2A(9), A2 => n290, B1 => minusA(9), B2 
                           => n284, ZN => n324);
   U189 : NAND2_X1 port map( A1 => n320, A2 => n319, ZN => n495);
   U190 : AOI22_X1 port map( A1 => plusA(7), A2 => n278, B1 => plus2A(7), B2 =>
                           n272, ZN => n320);
   U191 : AOI22_X1 port map( A1 => minus2A(7), A2 => n290, B1 => minusA(7), B2 
                           => n284, ZN => n319);
   U192 : NAND2_X1 port map( A1 => n318, A2 => n317, ZN => n496);
   U193 : AOI22_X1 port map( A1 => plusA(6), A2 => n278, B1 => plus2A(6), B2 =>
                           n272, ZN => n318);
   U194 : AOI22_X1 port map( A1 => minus2A(6), A2 => n290, B1 => minusA(6), B2 
                           => n284, ZN => n317);
   U195 : NAND2_X1 port map( A1 => n316, A2 => n315, ZN => n497);
   U196 : AOI22_X1 port map( A1 => plusA(5), A2 => n278, B1 => plus2A(5), B2 =>
                           n272, ZN => n316);
   U197 : AOI22_X1 port map( A1 => minus2A(5), A2 => n290, B1 => minusA(5), B2 
                           => n284, ZN => n315);
   U198 : NAND2_X1 port map( A1 => n312, A2 => n311, ZN => n499);
   U199 : AOI22_X1 port map( A1 => plusA(3), A2 => n278, B1 => plus2A(3), B2 =>
                           n272, ZN => n312);
   U200 : AOI22_X1 port map( A1 => minus2A(3), A2 => n290, B1 => minusA(3), B2 
                           => n284, ZN => n311);
   U201 : NAND2_X1 port map( A1 => n355, A2 => n354, ZN => n477);
   U202 : AOI22_X1 port map( A1 => plusA(24), A2 => n280, B1 => plus2A(24), B2 
                           => n274, ZN => n355);
   U203 : AOI22_X1 port map( A1 => minus2A(24), A2 => n292, B1 => minusA(24), 
                           B2 => n286, ZN => n354);
   U204 : NAND2_X1 port map( A1 => n347, A2 => n346, ZN => n481);
   U205 : AOI22_X1 port map( A1 => plusA(20), A2 => n279, B1 => plus2A(20), B2 
                           => n273, ZN => n347);
   U206 : AOI22_X1 port map( A1 => minus2A(20), A2 => n291, B1 => minusA(20), 
                           B2 => n285, ZN => n346);
   U207 : NAND2_X1 port map( A1 => n339, A2 => n338, ZN => n485);
   U208 : AOI22_X1 port map( A1 => plusA(16), A2 => n279, B1 => plus2A(16), B2 
                           => n273, ZN => n339);
   U209 : AOI22_X1 port map( A1 => minus2A(16), A2 => n291, B1 => minusA(16), 
                           B2 => n285, ZN => n338);
   U210 : NAND2_X1 port map( A1 => n331, A2 => n330, ZN => n489);
   U211 : AOI22_X1 port map( A1 => plusA(12), A2 => n279, B1 => plus2A(12), B2 
                           => n273, ZN => n331);
   U212 : AOI22_X1 port map( A1 => minus2A(12), A2 => n291, B1 => minusA(12), 
                           B2 => n285, ZN => n330);
   U213 : NAND2_X1 port map( A1 => n322, A2 => n321, ZN => n494);
   U214 : AOI22_X1 port map( A1 => plusA(8), A2 => n278, B1 => plus2A(8), B2 =>
                           n272, ZN => n322);
   U215 : AOI22_X1 port map( A1 => minus2A(8), A2 => n290, B1 => minusA(8), B2 
                           => n284, ZN => n321);
   U216 : NAND2_X1 port map( A1 => n314, A2 => n313, ZN => n498);
   U217 : AOI22_X1 port map( A1 => plusA(4), A2 => n278, B1 => plus2A(4), B2 =>
                           n272, ZN => n314);
   U218 : AOI22_X1 port map( A1 => minus2A(4), A2 => n290, B1 => minusA(4), B2 
                           => n284, ZN => n313);
   U219 : NAND2_X1 port map( A1 => n310, A2 => n309, ZN => n500);
   U220 : AOI22_X1 port map( A1 => plusA(2), A2 => n278, B1 => plus2A(2), B2 =>
                           n272, ZN => n310);
   U221 : AOI22_X1 port map( A1 => minus2A(2), A2 => n290, B1 => minusA(2), B2 
                           => n284, ZN => n309);
   U222 : NAND2_X1 port map( A1 => n308, A2 => n307, ZN => n501);
   U223 : AOI22_X1 port map( A1 => plusA(1), A2 => n278, B1 => plus2A(1), B2 =>
                           n272, ZN => n308);
   U224 : AOI22_X1 port map( A1 => minus2A(1), A2 => n290, B1 => minusA(1), B2 
                           => n284, ZN => n307);
   U225 : NAND2_X1 port map( A1 => n306, A2 => n305, ZN => n502);
   U226 : AOI22_X1 port map( A1 => plusA(0), A2 => n278, B1 => plus2A(0), B2 =>
                           n272, ZN => n306);
   U227 : AOI22_X1 port map( A1 => minus2A(0), A2 => n290, B1 => minusA(0), B2 
                           => n284, ZN => n305);
   U228 : CLKBUF_X1 port map( A => n432, Z => n277);
   U229 : CLKBUF_X1 port map( A => n433, Z => n283);
   U230 : CLKBUF_X1 port map( A => n434, Z => n289);
   U231 : CLKBUF_X1 port map( A => n435, Z => n295);
   U232 : CLKBUF_X1 port map( A => n493, Z => n301);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity MUX_GENERIC_N64_RADIX3_1 is

   port( plusA, minusA, plus2A, minus2A : in std_logic_vector (63 downto 0);  
         SEL : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (63 
         downto 0));

end MUX_GENERIC_N64_RADIX3_1;

architecture SYN_beh of MUX_GENERIC_N64_RADIX3_1 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component TBUF_X1
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   signal n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, 
      n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, 
      n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, 
      n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, 
      n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, 
      n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, 
      n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, 
      n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, 
      n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, 
      n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, 
      n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, 
      n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, 
      n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, 
      n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, 
      n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, 
      n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, 
      n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, 
      n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, 
      n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, 
      n499, n500, n501, n502 : std_logic;

begin
   
   Y_tri_61_inst : TBUF_X1 port map( A => n440, EN => n301, Z => Y(61));
   Y_tri_62_inst : TBUF_X1 port map( A => n439, EN => n301, Z => Y(62));
   Y_tri_63_inst : TBUF_X1 port map( A => n438, EN => n301, Z => Y(63));
   Y_tri_60_inst : TBUF_X1 port map( A => n441, EN => n301, Z => Y(60));
   Y_tri_26_inst : TBUF_X1 port map( A => n475, EN => n298, Z => Y(26));
   Y_tri_27_inst : TBUF_X1 port map( A => n474, EN => n298, Z => Y(27));
   Y_tri_28_inst : TBUF_X1 port map( A => n473, EN => n298, Z => Y(28));
   Y_tri_29_inst : TBUF_X1 port map( A => n472, EN => n298, Z => Y(29));
   Y_tri_35_inst : TBUF_X1 port map( A => n466, EN => n298, Z => Y(35));
   Y_tri_36_inst : TBUF_X1 port map( A => n465, EN => n299, Z => Y(36));
   Y_tri_37_inst : TBUF_X1 port map( A => n464, EN => n299, Z => Y(37));
   Y_tri_38_inst : TBUF_X1 port map( A => n463, EN => n299, Z => Y(38));
   Y_tri_39_inst : TBUF_X1 port map( A => n462, EN => n299, Z => Y(39));
   Y_tri_40_inst : TBUF_X1 port map( A => n461, EN => n299, Z => Y(40));
   Y_tri_41_inst : TBUF_X1 port map( A => n460, EN => n299, Z => Y(41));
   Y_tri_42_inst : TBUF_X1 port map( A => n459, EN => n299, Z => Y(42));
   Y_tri_43_inst : TBUF_X1 port map( A => n458, EN => n299, Z => Y(43));
   Y_tri_44_inst : TBUF_X1 port map( A => n457, EN => n299, Z => Y(44));
   Y_tri_45_inst : TBUF_X1 port map( A => n456, EN => n299, Z => Y(45));
   Y_tri_46_inst : TBUF_X1 port map( A => n455, EN => n299, Z => Y(46));
   Y_tri_47_inst : TBUF_X1 port map( A => n454, EN => n299, Z => Y(47));
   Y_tri_48_inst : TBUF_X1 port map( A => n453, EN => n300, Z => Y(48));
   Y_tri_49_inst : TBUF_X1 port map( A => n452, EN => n300, Z => Y(49));
   Y_tri_50_inst : TBUF_X1 port map( A => n451, EN => n300, Z => Y(50));
   Y_tri_51_inst : TBUF_X1 port map( A => n450, EN => n300, Z => Y(51));
   Y_tri_52_inst : TBUF_X1 port map( A => n449, EN => n300, Z => Y(52));
   Y_tri_53_inst : TBUF_X1 port map( A => n448, EN => n300, Z => Y(53));
   Y_tri_54_inst : TBUF_X1 port map( A => n447, EN => n300, Z => Y(54));
   Y_tri_55_inst : TBUF_X1 port map( A => n446, EN => n300, Z => Y(55));
   Y_tri_56_inst : TBUF_X1 port map( A => n445, EN => n300, Z => Y(56));
   Y_tri_57_inst : TBUF_X1 port map( A => n444, EN => n300, Z => Y(57));
   Y_tri_58_inst : TBUF_X1 port map( A => n443, EN => n300, Z => Y(58));
   Y_tri_59_inst : TBUF_X1 port map( A => n442, EN => n300, Z => Y(59));
   Y_tri_15_inst : TBUF_X1 port map( A => n486, EN => n297, Z => Y(15));
   Y_tri_16_inst : TBUF_X1 port map( A => n485, EN => n297, Z => Y(16));
   Y_tri_17_inst : TBUF_X1 port map( A => n484, EN => n297, Z => Y(17));
   Y_tri_18_inst : TBUF_X1 port map( A => n483, EN => n297, Z => Y(18));
   Y_tri_19_inst : TBUF_X1 port map( A => n482, EN => n297, Z => Y(19));
   Y_tri_20_inst : TBUF_X1 port map( A => n481, EN => n297, Z => Y(20));
   Y_tri_21_inst : TBUF_X1 port map( A => n480, EN => n297, Z => Y(21));
   Y_tri_22_inst : TBUF_X1 port map( A => n479, EN => n297, Z => Y(22));
   Y_tri_23_inst : TBUF_X1 port map( A => n478, EN => n297, Z => Y(23));
   Y_tri_24_inst : TBUF_X1 port map( A => n477, EN => n298, Z => Y(24));
   Y_tri_25_inst : TBUF_X1 port map( A => n476, EN => n298, Z => Y(25));
   Y_tri_30_inst : TBUF_X1 port map( A => n471, EN => n298, Z => Y(30));
   Y_tri_31_inst : TBUF_X1 port map( A => n470, EN => n298, Z => Y(31));
   Y_tri_32_inst : TBUF_X1 port map( A => n469, EN => n298, Z => Y(32));
   Y_tri_33_inst : TBUF_X1 port map( A => n468, EN => n298, Z => Y(33));
   Y_tri_34_inst : TBUF_X1 port map( A => n467, EN => n298, Z => Y(34));
   Y_tri_4_inst : TBUF_X1 port map( A => n498, EN => n296, Z => Y(4));
   Y_tri_5_inst : TBUF_X1 port map( A => n497, EN => n296, Z => Y(5));
   Y_tri_6_inst : TBUF_X1 port map( A => n496, EN => n296, Z => Y(6));
   Y_tri_7_inst : TBUF_X1 port map( A => n495, EN => n296, Z => Y(7));
   Y_tri_8_inst : TBUF_X1 port map( A => n494, EN => n296, Z => Y(8));
   Y_tri_9_inst : TBUF_X1 port map( A => n492, EN => n296, Z => Y(9));
   Y_tri_10_inst : TBUF_X1 port map( A => n491, EN => n296, Z => Y(10));
   Y_tri_11_inst : TBUF_X1 port map( A => n490, EN => n296, Z => Y(11));
   Y_tri_12_inst : TBUF_X1 port map( A => n489, EN => n297, Z => Y(12));
   Y_tri_13_inst : TBUF_X1 port map( A => n488, EN => n297, Z => Y(13));
   Y_tri_14_inst : TBUF_X1 port map( A => n487, EN => n297, Z => Y(14));
   Y_tri_1_inst : TBUF_X1 port map( A => n501, EN => n296, Z => Y(1));
   Y_tri_2_inst : TBUF_X1 port map( A => n500, EN => n296, Z => Y(2));
   Y_tri_3_inst : TBUF_X1 port map( A => n499, EN => n296, Z => Y(3));
   Y_tri_0_inst : TBUF_X1 port map( A => n502, EN => n296, Z => Y(0));
   U2 : NOR3_X1 port map( A1 => SEL(0), A2 => SEL(2), A3 => n302, ZN => n434);
   U3 : NOR3_X1 port map( A1 => n302, A2 => SEL(2), A3 => n303, ZN => n432);
   U4 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n303, ZN => n433);
   U5 : NAND2_X1 port map( A1 => n375, A2 => n374, ZN => n467);
   U6 : AOI22_X1 port map( A1 => plusA(34), A2 => n280, B1 => plus2A(34), B2 =>
                           n274, ZN => n375);
   U7 : AOI22_X1 port map( A1 => minus2A(34), A2 => n292, B1 => minusA(34), B2 
                           => n286, ZN => n374);
   U8 : NAND2_X1 port map( A1 => n427, A2 => n426, ZN => n441);
   U9 : AOI22_X1 port map( A1 => plusA(60), A2 => n283, B1 => plus2A(60), B2 =>
                           n277, ZN => n427);
   U10 : AOI22_X1 port map( A1 => minus2A(60), A2 => n295, B1 => minusA(60), B2
                           => n289, ZN => n426);
   U11 : NAND2_X1 port map( A1 => n425, A2 => n424, ZN => n442);
   U12 : AOI22_X1 port map( A1 => plusA(59), A2 => n282, B1 => plus2A(59), B2 
                           => n276, ZN => n425);
   U13 : AOI22_X1 port map( A1 => minus2A(59), A2 => n294, B1 => minusA(59), B2
                           => n288, ZN => n424);
   U14 : NAND2_X1 port map( A1 => n423, A2 => n422, ZN => n443);
   U15 : AOI22_X1 port map( A1 => plusA(58), A2 => n282, B1 => plus2A(58), B2 
                           => n276, ZN => n423);
   U16 : AOI22_X1 port map( A1 => minus2A(58), A2 => n294, B1 => minusA(58), B2
                           => n288, ZN => n422);
   U17 : NAND2_X1 port map( A1 => n421, A2 => n420, ZN => n444);
   U18 : AOI22_X1 port map( A1 => plusA(57), A2 => n282, B1 => plus2A(57), B2 
                           => n276, ZN => n421);
   U19 : AOI22_X1 port map( A1 => minus2A(57), A2 => n294, B1 => minusA(57), B2
                           => n288, ZN => n420);
   U20 : NAND2_X1 port map( A1 => n419, A2 => n418, ZN => n445);
   U21 : AOI22_X1 port map( A1 => plusA(56), A2 => n282, B1 => plus2A(56), B2 
                           => n276, ZN => n419);
   U22 : AOI22_X1 port map( A1 => minus2A(56), A2 => n294, B1 => minusA(56), B2
                           => n288, ZN => n418);
   U23 : NAND2_X1 port map( A1 => n417, A2 => n416, ZN => n446);
   U24 : AOI22_X1 port map( A1 => plusA(55), A2 => n282, B1 => plus2A(55), B2 
                           => n276, ZN => n417);
   U25 : AOI22_X1 port map( A1 => minus2A(55), A2 => n294, B1 => minusA(55), B2
                           => n288, ZN => n416);
   U26 : NAND2_X1 port map( A1 => n415, A2 => n414, ZN => n447);
   U27 : AOI22_X1 port map( A1 => plusA(54), A2 => n282, B1 => plus2A(54), B2 
                           => n276, ZN => n415);
   U28 : AOI22_X1 port map( A1 => minus2A(54), A2 => n294, B1 => minusA(54), B2
                           => n288, ZN => n414);
   U29 : NAND2_X1 port map( A1 => n413, A2 => n412, ZN => n448);
   U30 : AOI22_X1 port map( A1 => plusA(53), A2 => n282, B1 => plus2A(53), B2 
                           => n276, ZN => n413);
   U31 : AOI22_X1 port map( A1 => minus2A(53), A2 => n294, B1 => minusA(53), B2
                           => n288, ZN => n412);
   U32 : NAND2_X1 port map( A1 => n411, A2 => n410, ZN => n449);
   U33 : AOI22_X1 port map( A1 => plusA(52), A2 => n282, B1 => plus2A(52), B2 
                           => n276, ZN => n411);
   U34 : AOI22_X1 port map( A1 => minus2A(52), A2 => n294, B1 => minusA(52), B2
                           => n288, ZN => n410);
   U35 : NAND2_X1 port map( A1 => n409, A2 => n408, ZN => n450);
   U36 : AOI22_X1 port map( A1 => plusA(51), A2 => n282, B1 => plus2A(51), B2 
                           => n276, ZN => n409);
   U37 : AOI22_X1 port map( A1 => minus2A(51), A2 => n294, B1 => minusA(51), B2
                           => n288, ZN => n408);
   U38 : NAND2_X1 port map( A1 => n407, A2 => n406, ZN => n451);
   U39 : AOI22_X1 port map( A1 => plusA(50), A2 => n282, B1 => plus2A(50), B2 
                           => n276, ZN => n407);
   U40 : AOI22_X1 port map( A1 => minus2A(50), A2 => n294, B1 => minusA(50), B2
                           => n288, ZN => n406);
   U41 : NAND2_X1 port map( A1 => n405, A2 => n404, ZN => n452);
   U42 : AOI22_X1 port map( A1 => plusA(49), A2 => n282, B1 => plus2A(49), B2 
                           => n276, ZN => n405);
   U43 : AOI22_X1 port map( A1 => minus2A(49), A2 => n294, B1 => minusA(49), B2
                           => n288, ZN => n404);
   U44 : NAND2_X1 port map( A1 => n401, A2 => n400, ZN => n454);
   U45 : AOI22_X1 port map( A1 => plusA(47), A2 => n281, B1 => plus2A(47), B2 
                           => n275, ZN => n401);
   U46 : AOI22_X1 port map( A1 => minus2A(47), A2 => n293, B1 => minusA(47), B2
                           => n287, ZN => n400);
   U47 : NAND2_X1 port map( A1 => n393, A2 => n392, ZN => n458);
   U48 : AOI22_X1 port map( A1 => plusA(43), A2 => n281, B1 => plus2A(43), B2 
                           => n275, ZN => n393);
   U49 : AOI22_X1 port map( A1 => minus2A(43), A2 => n293, B1 => minusA(43), B2
                           => n287, ZN => n392);
   U50 : NAND2_X1 port map( A1 => n385, A2 => n384, ZN => n462);
   U51 : AOI22_X1 port map( A1 => plusA(39), A2 => n281, B1 => plus2A(39), B2 
                           => n275, ZN => n385);
   U52 : AOI22_X1 port map( A1 => minus2A(39), A2 => n293, B1 => minusA(39), B2
                           => n287, ZN => n384);
   U53 : NAND2_X1 port map( A1 => n377, A2 => n376, ZN => n466);
   U54 : AOI22_X1 port map( A1 => plusA(35), A2 => n280, B1 => plus2A(35), B2 
                           => n274, ZN => n377);
   U55 : AOI22_X1 port map( A1 => minus2A(35), A2 => n292, B1 => minusA(35), B2
                           => n286, ZN => n376);
   U56 : NAND2_X1 port map( A1 => n397, A2 => n396, ZN => n456);
   U57 : AOI22_X1 port map( A1 => plusA(45), A2 => n281, B1 => plus2A(45), B2 
                           => n275, ZN => n397);
   U58 : AOI22_X1 port map( A1 => minus2A(45), A2 => n293, B1 => minusA(45), B2
                           => n287, ZN => n396);
   U59 : NAND2_X1 port map( A1 => n389, A2 => n388, ZN => n460);
   U60 : AOI22_X1 port map( A1 => plusA(41), A2 => n281, B1 => plus2A(41), B2 
                           => n275, ZN => n389);
   U61 : AOI22_X1 port map( A1 => minus2A(41), A2 => n293, B1 => minusA(41), B2
                           => n287, ZN => n388);
   U62 : NAND2_X1 port map( A1 => n381, A2 => n380, ZN => n464);
   U63 : AOI22_X1 port map( A1 => plusA(37), A2 => n281, B1 => plus2A(37), B2 
                           => n275, ZN => n381);
   U64 : AOI22_X1 port map( A1 => minus2A(37), A2 => n293, B1 => minusA(37), B2
                           => n287, ZN => n380);
   U65 : NAND2_X1 port map( A1 => n403, A2 => n402, ZN => n453);
   U66 : AOI22_X1 port map( A1 => plusA(48), A2 => n282, B1 => plus2A(48), B2 
                           => n276, ZN => n403);
   U67 : AOI22_X1 port map( A1 => minus2A(48), A2 => n294, B1 => minusA(48), B2
                           => n288, ZN => n402);
   U68 : NAND2_X1 port map( A1 => n395, A2 => n394, ZN => n457);
   U69 : AOI22_X1 port map( A1 => plusA(44), A2 => n281, B1 => plus2A(44), B2 
                           => n275, ZN => n395);
   U70 : AOI22_X1 port map( A1 => minus2A(44), A2 => n293, B1 => minusA(44), B2
                           => n287, ZN => n394);
   U71 : NAND2_X1 port map( A1 => n387, A2 => n386, ZN => n461);
   U72 : AOI22_X1 port map( A1 => plusA(40), A2 => n281, B1 => plus2A(40), B2 
                           => n275, ZN => n387);
   U73 : AOI22_X1 port map( A1 => minus2A(40), A2 => n293, B1 => minusA(40), B2
                           => n287, ZN => n386);
   U74 : NAND2_X1 port map( A1 => n379, A2 => n378, ZN => n465);
   U75 : AOI22_X1 port map( A1 => plusA(36), A2 => n281, B1 => plus2A(36), B2 
                           => n275, ZN => n379);
   U76 : AOI22_X1 port map( A1 => minus2A(36), A2 => n293, B1 => minusA(36), B2
                           => n287, ZN => n378);
   U77 : NAND2_X1 port map( A1 => n399, A2 => n398, ZN => n455);
   U78 : AOI22_X1 port map( A1 => plusA(46), A2 => n281, B1 => plus2A(46), B2 
                           => n275, ZN => n399);
   U79 : AOI22_X1 port map( A1 => minus2A(46), A2 => n293, B1 => minusA(46), B2
                           => n287, ZN => n398);
   U80 : NAND2_X1 port map( A1 => n391, A2 => n390, ZN => n459);
   U81 : AOI22_X1 port map( A1 => plusA(42), A2 => n281, B1 => plus2A(42), B2 
                           => n275, ZN => n391);
   U82 : AOI22_X1 port map( A1 => minus2A(42), A2 => n293, B1 => minusA(42), B2
                           => n287, ZN => n390);
   U83 : NAND2_X1 port map( A1 => n383, A2 => n382, ZN => n463);
   U84 : AOI22_X1 port map( A1 => plusA(38), A2 => n281, B1 => plus2A(38), B2 
                           => n275, ZN => n383);
   U85 : AOI22_X1 port map( A1 => minus2A(38), A2 => n293, B1 => minusA(38), B2
                           => n287, ZN => n382);
   U86 : NAND2_X1 port map( A1 => n437, A2 => n436, ZN => n438);
   U87 : AOI22_X1 port map( A1 => plusA(63), A2 => n283, B1 => plus2A(63), B2 
                           => n277, ZN => n437);
   U88 : AOI22_X1 port map( A1 => minus2A(63), A2 => n295, B1 => minusA(63), B2
                           => n289, ZN => n436);
   U89 : NAND2_X1 port map( A1 => n429, A2 => n428, ZN => n440);
   U90 : AOI22_X1 port map( A1 => plusA(61), A2 => n283, B1 => plus2A(61), B2 
                           => n277, ZN => n429);
   U91 : AOI22_X1 port map( A1 => minus2A(61), A2 => n295, B1 => minusA(61), B2
                           => n289, ZN => n428);
   U92 : NAND2_X1 port map( A1 => n431, A2 => n430, ZN => n439);
   U93 : AOI22_X1 port map( A1 => plusA(62), A2 => n283, B1 => plus2A(62), B2 
                           => n277, ZN => n431);
   U94 : AOI22_X1 port map( A1 => minus2A(62), A2 => n295, B1 => minusA(62), B2
                           => n289, ZN => n430);
   U95 : BUF_X1 port map( A => n493, Z => n296);
   U96 : BUF_X1 port map( A => n493, Z => n297);
   U97 : BUF_X1 port map( A => n493, Z => n298);
   U98 : NAND2_X1 port map( A1 => n373, A2 => n372, ZN => n468);
   U99 : AOI22_X1 port map( A1 => plusA(33), A2 => n280, B1 => plus2A(33), B2 
                           => n274, ZN => n373);
   U100 : AOI22_X1 port map( A1 => minus2A(33), A2 => n292, B1 => minusA(33), 
                           B2 => n286, ZN => n372);
   U101 : NAND2_X1 port map( A1 => n371, A2 => n370, ZN => n469);
   U102 : AOI22_X1 port map( A1 => plusA(32), A2 => n280, B1 => plus2A(32), B2 
                           => n274, ZN => n371);
   U103 : AOI22_X1 port map( A1 => minus2A(32), A2 => n292, B1 => minusA(32), 
                           B2 => n286, ZN => n370);
   U104 : BUF_X1 port map( A => n493, Z => n299);
   U105 : BUF_X1 port map( A => n433, Z => n281);
   U106 : BUF_X1 port map( A => n433, Z => n280);
   U107 : BUF_X1 port map( A => n434, Z => n287);
   U108 : BUF_X1 port map( A => n432, Z => n275);
   U109 : BUF_X1 port map( A => n434, Z => n286);
   U110 : BUF_X1 port map( A => n432, Z => n274);
   U111 : BUF_X1 port map( A => n435, Z => n293);
   U112 : BUF_X1 port map( A => n435, Z => n292);
   U113 : BUF_X1 port map( A => n493, Z => n300);
   U114 : BUF_X1 port map( A => n433, Z => n282);
   U115 : BUF_X1 port map( A => n434, Z => n288);
   U116 : BUF_X1 port map( A => n432, Z => n276);
   U117 : BUF_X1 port map( A => n435, Z => n294);
   U118 : BUF_X1 port map( A => n433, Z => n279);
   U119 : BUF_X1 port map( A => n433, Z => n278);
   U120 : BUF_X1 port map( A => n434, Z => n285);
   U121 : BUF_X1 port map( A => n432, Z => n273);
   U122 : BUF_X1 port map( A => n434, Z => n284);
   U123 : BUF_X1 port map( A => n432, Z => n272);
   U124 : BUF_X1 port map( A => n435, Z => n291);
   U125 : BUF_X1 port map( A => n435, Z => n290);
   U126 : NOR2_X1 port map( A1 => n323, A2 => n304, ZN => n493);
   U127 : INV_X1 port map( A => SEL(2), ZN => n304);
   U128 : NOR2_X1 port map( A1 => SEL(1), A2 => SEL(0), ZN => n323);
   U129 : NAND2_X1 port map( A1 => n369, A2 => n368, ZN => n470);
   U130 : AOI22_X1 port map( A1 => plusA(31), A2 => n280, B1 => plus2A(31), B2 
                           => n274, ZN => n369);
   U131 : AOI22_X1 port map( A1 => minus2A(31), A2 => n292, B1 => minusA(31), 
                           B2 => n286, ZN => n368);
   U132 : AND2_X1 port map( A1 => SEL(2), A2 => n323, ZN => n435);
   U133 : INV_X1 port map( A => SEL(1), ZN => n302);
   U134 : INV_X1 port map( A => SEL(0), ZN => n303);
   U135 : NAND2_X1 port map( A1 => n367, A2 => n366, ZN => n471);
   U136 : AOI22_X1 port map( A1 => plusA(30), A2 => n280, B1 => plus2A(30), B2 
                           => n274, ZN => n367);
   U137 : AOI22_X1 port map( A1 => minus2A(30), A2 => n292, B1 => minusA(30), 
                           B2 => n286, ZN => n366);
   U138 : NAND2_X1 port map( A1 => n365, A2 => n364, ZN => n472);
   U139 : AOI22_X1 port map( A1 => plusA(29), A2 => n280, B1 => plus2A(29), B2 
                           => n274, ZN => n365);
   U140 : AOI22_X1 port map( A1 => minus2A(29), A2 => n292, B1 => minusA(29), 
                           B2 => n286, ZN => n364);
   U141 : NAND2_X1 port map( A1 => n361, A2 => n360, ZN => n474);
   U142 : AOI22_X1 port map( A1 => plusA(27), A2 => n280, B1 => plus2A(27), B2 
                           => n274, ZN => n361);
   U143 : AOI22_X1 port map( A1 => minus2A(27), A2 => n292, B1 => minusA(27), 
                           B2 => n286, ZN => n360);
   U144 : NAND2_X1 port map( A1 => n359, A2 => n358, ZN => n475);
   U145 : AOI22_X1 port map( A1 => plusA(26), A2 => n280, B1 => plus2A(26), B2 
                           => n274, ZN => n359);
   U146 : AOI22_X1 port map( A1 => minus2A(26), A2 => n292, B1 => minusA(26), 
                           B2 => n286, ZN => n358);
   U147 : NAND2_X1 port map( A1 => n357, A2 => n356, ZN => n476);
   U148 : AOI22_X1 port map( A1 => plusA(25), A2 => n280, B1 => plus2A(25), B2 
                           => n274, ZN => n357);
   U149 : AOI22_X1 port map( A1 => minus2A(25), A2 => n292, B1 => minusA(25), 
                           B2 => n286, ZN => n356);
   U150 : NAND2_X1 port map( A1 => n353, A2 => n352, ZN => n478);
   U151 : AOI22_X1 port map( A1 => plusA(23), A2 => n279, B1 => plus2A(23), B2 
                           => n273, ZN => n353);
   U152 : AOI22_X1 port map( A1 => minus2A(23), A2 => n291, B1 => minusA(23), 
                           B2 => n285, ZN => n352);
   U153 : NAND2_X1 port map( A1 => n351, A2 => n350, ZN => n479);
   U154 : AOI22_X1 port map( A1 => plusA(22), A2 => n279, B1 => plus2A(22), B2 
                           => n273, ZN => n351);
   U155 : AOI22_X1 port map( A1 => minus2A(22), A2 => n291, B1 => minusA(22), 
                           B2 => n285, ZN => n350);
   U156 : NAND2_X1 port map( A1 => n349, A2 => n348, ZN => n480);
   U157 : AOI22_X1 port map( A1 => plusA(21), A2 => n279, B1 => plus2A(21), B2 
                           => n273, ZN => n349);
   U158 : AOI22_X1 port map( A1 => minus2A(21), A2 => n291, B1 => minusA(21), 
                           B2 => n285, ZN => n348);
   U159 : NAND2_X1 port map( A1 => n345, A2 => n344, ZN => n482);
   U160 : AOI22_X1 port map( A1 => plusA(19), A2 => n279, B1 => plus2A(19), B2 
                           => n273, ZN => n345);
   U161 : AOI22_X1 port map( A1 => minus2A(19), A2 => n291, B1 => minusA(19), 
                           B2 => n285, ZN => n344);
   U162 : NAND2_X1 port map( A1 => n343, A2 => n342, ZN => n483);
   U163 : AOI22_X1 port map( A1 => plusA(18), A2 => n279, B1 => plus2A(18), B2 
                           => n273, ZN => n343);
   U164 : AOI22_X1 port map( A1 => minus2A(18), A2 => n291, B1 => minusA(18), 
                           B2 => n285, ZN => n342);
   U165 : NAND2_X1 port map( A1 => n341, A2 => n340, ZN => n484);
   U166 : AOI22_X1 port map( A1 => plusA(17), A2 => n279, B1 => plus2A(17), B2 
                           => n273, ZN => n341);
   U167 : AOI22_X1 port map( A1 => minus2A(17), A2 => n291, B1 => minusA(17), 
                           B2 => n285, ZN => n340);
   U168 : NAND2_X1 port map( A1 => n337, A2 => n336, ZN => n486);
   U169 : AOI22_X1 port map( A1 => plusA(15), A2 => n279, B1 => plus2A(15), B2 
                           => n273, ZN => n337);
   U170 : AOI22_X1 port map( A1 => minus2A(15), A2 => n291, B1 => minusA(15), 
                           B2 => n285, ZN => n336);
   U171 : NAND2_X1 port map( A1 => n335, A2 => n334, ZN => n487);
   U172 : AOI22_X1 port map( A1 => plusA(14), A2 => n279, B1 => plus2A(14), B2 
                           => n273, ZN => n335);
   U173 : AOI22_X1 port map( A1 => minus2A(14), A2 => n291, B1 => minusA(14), 
                           B2 => n285, ZN => n334);
   U174 : NAND2_X1 port map( A1 => n333, A2 => n332, ZN => n488);
   U175 : AOI22_X1 port map( A1 => plusA(13), A2 => n279, B1 => plus2A(13), B2 
                           => n273, ZN => n333);
   U176 : AOI22_X1 port map( A1 => minus2A(13), A2 => n291, B1 => minusA(13), 
                           B2 => n285, ZN => n332);
   U177 : NAND2_X1 port map( A1 => n329, A2 => n328, ZN => n490);
   U178 : AOI22_X1 port map( A1 => plusA(11), A2 => n278, B1 => plus2A(11), B2 
                           => n272, ZN => n329);
   U179 : AOI22_X1 port map( A1 => minus2A(11), A2 => n290, B1 => minusA(11), 
                           B2 => n284, ZN => n328);
   U180 : NAND2_X1 port map( A1 => n327, A2 => n326, ZN => n491);
   U181 : AOI22_X1 port map( A1 => plusA(10), A2 => n278, B1 => plus2A(10), B2 
                           => n272, ZN => n327);
   U182 : AOI22_X1 port map( A1 => minus2A(10), A2 => n290, B1 => minusA(10), 
                           B2 => n284, ZN => n326);
   U183 : NAND2_X1 port map( A1 => n325, A2 => n324, ZN => n492);
   U184 : AOI22_X1 port map( A1 => plusA(9), A2 => n278, B1 => plus2A(9), B2 =>
                           n272, ZN => n325);
   U185 : AOI22_X1 port map( A1 => minus2A(9), A2 => n290, B1 => minusA(9), B2 
                           => n284, ZN => n324);
   U186 : NAND2_X1 port map( A1 => n320, A2 => n319, ZN => n495);
   U187 : AOI22_X1 port map( A1 => plusA(7), A2 => n278, B1 => plus2A(7), B2 =>
                           n272, ZN => n320);
   U188 : AOI22_X1 port map( A1 => minus2A(7), A2 => n290, B1 => minusA(7), B2 
                           => n284, ZN => n319);
   U189 : NAND2_X1 port map( A1 => n318, A2 => n317, ZN => n496);
   U190 : AOI22_X1 port map( A1 => plusA(6), A2 => n278, B1 => plus2A(6), B2 =>
                           n272, ZN => n318);
   U191 : AOI22_X1 port map( A1 => minus2A(6), A2 => n290, B1 => minusA(6), B2 
                           => n284, ZN => n317);
   U192 : NAND2_X1 port map( A1 => n316, A2 => n315, ZN => n497);
   U193 : AOI22_X1 port map( A1 => plusA(5), A2 => n278, B1 => plus2A(5), B2 =>
                           n272, ZN => n316);
   U194 : AOI22_X1 port map( A1 => minus2A(5), A2 => n290, B1 => minusA(5), B2 
                           => n284, ZN => n315);
   U195 : NAND2_X1 port map( A1 => n312, A2 => n311, ZN => n499);
   U196 : AOI22_X1 port map( A1 => plusA(3), A2 => n278, B1 => plus2A(3), B2 =>
                           n272, ZN => n312);
   U197 : AOI22_X1 port map( A1 => minus2A(3), A2 => n290, B1 => minusA(3), B2 
                           => n284, ZN => n311);
   U198 : NAND2_X1 port map( A1 => n363, A2 => n362, ZN => n473);
   U199 : AOI22_X1 port map( A1 => plusA(28), A2 => n280, B1 => plus2A(28), B2 
                           => n274, ZN => n363);
   U200 : AOI22_X1 port map( A1 => minus2A(28), A2 => n292, B1 => minusA(28), 
                           B2 => n286, ZN => n362);
   U201 : NAND2_X1 port map( A1 => n355, A2 => n354, ZN => n477);
   U202 : AOI22_X1 port map( A1 => plusA(24), A2 => n280, B1 => plus2A(24), B2 
                           => n274, ZN => n355);
   U203 : AOI22_X1 port map( A1 => minus2A(24), A2 => n292, B1 => minusA(24), 
                           B2 => n286, ZN => n354);
   U204 : NAND2_X1 port map( A1 => n347, A2 => n346, ZN => n481);
   U205 : AOI22_X1 port map( A1 => plusA(20), A2 => n279, B1 => plus2A(20), B2 
                           => n273, ZN => n347);
   U206 : AOI22_X1 port map( A1 => minus2A(20), A2 => n291, B1 => minusA(20), 
                           B2 => n285, ZN => n346);
   U207 : NAND2_X1 port map( A1 => n339, A2 => n338, ZN => n485);
   U208 : AOI22_X1 port map( A1 => plusA(16), A2 => n279, B1 => plus2A(16), B2 
                           => n273, ZN => n339);
   U209 : AOI22_X1 port map( A1 => minus2A(16), A2 => n291, B1 => minusA(16), 
                           B2 => n285, ZN => n338);
   U210 : NAND2_X1 port map( A1 => n331, A2 => n330, ZN => n489);
   U211 : AOI22_X1 port map( A1 => plusA(12), A2 => n279, B1 => plus2A(12), B2 
                           => n273, ZN => n331);
   U212 : AOI22_X1 port map( A1 => minus2A(12), A2 => n291, B1 => minusA(12), 
                           B2 => n285, ZN => n330);
   U213 : NAND2_X1 port map( A1 => n322, A2 => n321, ZN => n494);
   U214 : AOI22_X1 port map( A1 => plusA(8), A2 => n278, B1 => plus2A(8), B2 =>
                           n272, ZN => n322);
   U215 : AOI22_X1 port map( A1 => minus2A(8), A2 => n290, B1 => minusA(8), B2 
                           => n284, ZN => n321);
   U216 : NAND2_X1 port map( A1 => n314, A2 => n313, ZN => n498);
   U217 : AOI22_X1 port map( A1 => plusA(4), A2 => n278, B1 => plus2A(4), B2 =>
                           n272, ZN => n314);
   U218 : AOI22_X1 port map( A1 => minus2A(4), A2 => n290, B1 => minusA(4), B2 
                           => n284, ZN => n313);
   U219 : NAND2_X1 port map( A1 => n310, A2 => n309, ZN => n500);
   U220 : AOI22_X1 port map( A1 => plusA(2), A2 => n278, B1 => plus2A(2), B2 =>
                           n272, ZN => n310);
   U221 : AOI22_X1 port map( A1 => minus2A(2), A2 => n290, B1 => minusA(2), B2 
                           => n284, ZN => n309);
   U222 : NAND2_X1 port map( A1 => n308, A2 => n307, ZN => n501);
   U223 : AOI22_X1 port map( A1 => plusA(1), A2 => n278, B1 => plus2A(1), B2 =>
                           n272, ZN => n308);
   U224 : AOI22_X1 port map( A1 => minus2A(1), A2 => n290, B1 => minusA(1), B2 
                           => n284, ZN => n307);
   U225 : NAND2_X1 port map( A1 => n306, A2 => n305, ZN => n502);
   U226 : AOI22_X1 port map( A1 => plusA(0), A2 => n278, B1 => plus2A(0), B2 =>
                           n272, ZN => n306);
   U227 : AOI22_X1 port map( A1 => minus2A(0), A2 => n290, B1 => minusA(0), B2 
                           => n284, ZN => n305);
   U228 : CLKBUF_X1 port map( A => n432, Z => n277);
   U229 : CLKBUF_X1 port map( A => n433, Z => n283);
   U230 : CLKBUF_X1 port map( A => n434, Z => n289);
   U231 : CLKBUF_X1 port map( A => n435, Z => n295);
   U232 : CLKBUF_X1 port map( A => n493, Z => n301);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity encoder_N64_RADIX3_15 is

   port( X : in std_logic_vector (2 downto 0);  Z : out std_logic_vector (2 
         downto 0));

end encoder_N64_RADIX3_15;

architecture SYN_beh of encoder_N64_RADIX3_15 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7, n8, n9, n10, n11, n12, n13, n15, n16 : std_logic;

begin
   
   U1 : AND2_X2 port map( A1 => n6, A2 => n12, ZN => Z(2));
   U2 : OR2_X1 port map( A1 => X(0), A2 => X(1), ZN => n8);
   U3 : OR2_X1 port map( A1 => X(0), A2 => X(1), ZN => n5);
   U4 : OR2_X1 port map( A1 => X(0), A2 => X(1), ZN => n11);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n10, ZN => n6);
   U6 : NAND2_X1 port map( A1 => X(0), A2 => X(1), ZN => n7);
   U7 : AOI21_X1 port map( B1 => n16, B2 => n10, A => X(2), ZN => Z(0));
   U8 : NAND2_X1 port map( A1 => n11, A2 => n7, ZN => n9);
   U9 : NAND2_X1 port map( A1 => X(0), A2 => X(1), ZN => n10);
   U10 : NAND2_X1 port map( A1 => n8, A2 => n15, ZN => n16);
   U11 : AND2_X1 port map( A1 => n15, A2 => X(2), ZN => n12);
   U12 : INV_X1 port map( A => X(2), ZN => n13);
   U13 : NAND2_X1 port map( A1 => X(0), A2 => X(1), ZN => n15);
   U14 : OAI22_X1 port map( A1 => n9, A2 => n13, B1 => n10, B2 => X(2), ZN => 
                           Z(1));

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity encoder_N64_RADIX3_14 is

   port( X : in std_logic_vector (2 downto 0);  Z : out std_logic_vector (2 
         downto 0));

end encoder_N64_RADIX3_14;

architecture SYN_beh of encoder_N64_RADIX3_14 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7, n8, n9, n11, n12 : std_logic;

begin
   
   U2 : AND3_X2 port map( A1 => X(2), A2 => n7, A3 => n12, ZN => Z(2));
   U1 : NAND2_X1 port map( A1 => X(1), A2 => X(0), ZN => n5);
   U3 : NAND2_X1 port map( A1 => X(1), A2 => X(0), ZN => n6);
   U4 : NAND2_X1 port map( A1 => X(1), A2 => X(0), ZN => n7);
   U5 : OAI21_X1 port map( B1 => X(1), B2 => X(0), A => n11, ZN => n8);
   U6 : OAI22_X1 port map( A1 => n8, A2 => n9, B1 => X(2), B2 => n7, ZN => Z(1)
                           );
   U7 : INV_X1 port map( A => X(2), ZN => n9);
   U8 : AOI21_X1 port map( B1 => n8, B2 => n5, A => X(2), ZN => Z(0));
   U9 : OAI21_X1 port map( B1 => X(1), B2 => X(0), A => n6, ZN => n12);
   U10 : NAND2_X1 port map( A1 => X(1), A2 => X(0), ZN => n11);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity encoder_N64_RADIX3_13 is

   port( X : in std_logic_vector (2 downto 0);  Z : out std_logic_vector (2 
         downto 0));

end encoder_N64_RADIX3_13;

architecture SYN_beh of encoder_N64_RADIX3_13 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n7, n8 : std_logic;

begin
   
   U2 : AND3_X2 port map( A1 => X(2), A2 => n7, A3 => n8, ZN => Z(2));
   U1 : OAI22_X1 port map( A1 => n8, A2 => n5, B1 => X(2), B2 => n7, ZN => Z(1)
                           );
   U3 : INV_X1 port map( A => X(2), ZN => n5);
   U4 : AOI21_X1 port map( B1 => n8, B2 => n7, A => X(2), ZN => Z(0));
   U5 : OAI21_X1 port map( B1 => X(1), B2 => X(0), A => n7, ZN => n8);
   U6 : NAND2_X1 port map( A1 => X(1), A2 => X(0), ZN => n7);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity encoder_N64_RADIX3_12 is

   port( X : in std_logic_vector (2 downto 0);  Z : out std_logic_vector (2 
         downto 0));

end encoder_N64_RADIX3_12;

architecture SYN_beh of encoder_N64_RADIX3_12 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n7, n8 : std_logic;

begin
   
   U1 : AND3_X1 port map( A1 => X(2), A2 => n7, A3 => n8, ZN => Z(2));
   U2 : OAI22_X1 port map( A1 => n8, A2 => n5, B1 => X(2), B2 => n7, ZN => Z(1)
                           );
   U3 : INV_X1 port map( A => X(2), ZN => n5);
   U4 : AOI21_X1 port map( B1 => n8, B2 => n7, A => X(2), ZN => Z(0));
   U5 : OAI21_X1 port map( B1 => X(1), B2 => X(0), A => n7, ZN => n8);
   U6 : NAND2_X1 port map( A1 => X(1), A2 => X(0), ZN => n7);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity encoder_N64_RADIX3_11 is

   port( X : in std_logic_vector (2 downto 0);  Z : out std_logic_vector (2 
         downto 0));

end encoder_N64_RADIX3_11;

architecture SYN_beh of encoder_N64_RADIX3_11 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n7, n8 : std_logic;

begin
   
   U1 : OAI22_X1 port map( A1 => n8, A2 => n5, B1 => X(2), B2 => n7, ZN => Z(1)
                           );
   U2 : INV_X1 port map( A => X(2), ZN => n5);
   U3 : AOI21_X1 port map( B1 => n8, B2 => n7, A => X(2), ZN => Z(0));
   U4 : OAI21_X1 port map( B1 => X(1), B2 => X(0), A => n7, ZN => n8);
   U5 : AND3_X1 port map( A1 => X(2), A2 => n7, A3 => n8, ZN => Z(2));
   U6 : NAND2_X1 port map( A1 => X(1), A2 => X(0), ZN => n7);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity encoder_N64_RADIX3_10 is

   port( X : in std_logic_vector (2 downto 0);  Z : out std_logic_vector (2 
         downto 0));

end encoder_N64_RADIX3_10;

architecture SYN_beh of encoder_N64_RADIX3_10 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n7, n8 : std_logic;

begin
   
   U1 : OAI22_X1 port map( A1 => n8, A2 => n5, B1 => X(2), B2 => n7, ZN => Z(1)
                           );
   U2 : INV_X1 port map( A => X(2), ZN => n5);
   U3 : AOI21_X1 port map( B1 => n8, B2 => n7, A => X(2), ZN => Z(0));
   U4 : OAI21_X1 port map( B1 => X(1), B2 => X(0), A => n7, ZN => n8);
   U5 : AND3_X1 port map( A1 => X(2), A2 => n7, A3 => n8, ZN => Z(2));
   U6 : NAND2_X1 port map( A1 => X(1), A2 => X(0), ZN => n7);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity encoder_N64_RADIX3_9 is

   port( X : in std_logic_vector (2 downto 0);  Z : out std_logic_vector (2 
         downto 0));

end encoder_N64_RADIX3_9;

architecture SYN_beh of encoder_N64_RADIX3_9 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n7, n8 : std_logic;

begin
   
   U1 : OAI22_X1 port map( A1 => n8, A2 => n5, B1 => X(2), B2 => n7, ZN => Z(1)
                           );
   U2 : INV_X1 port map( A => X(2), ZN => n5);
   U3 : AOI21_X1 port map( B1 => n8, B2 => n7, A => X(2), ZN => Z(0));
   U4 : OAI21_X1 port map( B1 => X(1), B2 => X(0), A => n7, ZN => n8);
   U5 : AND3_X1 port map( A1 => X(2), A2 => n7, A3 => n8, ZN => Z(2));
   U6 : NAND2_X1 port map( A1 => X(1), A2 => X(0), ZN => n7);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity encoder_N64_RADIX3_8 is

   port( X : in std_logic_vector (2 downto 0);  Z : out std_logic_vector (2 
         downto 0));

end encoder_N64_RADIX3_8;

architecture SYN_beh of encoder_N64_RADIX3_8 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n7, n8 : std_logic;

begin
   
   U1 : OAI22_X1 port map( A1 => n8, A2 => n5, B1 => X(2), B2 => n7, ZN => Z(1)
                           );
   U2 : INV_X1 port map( A => X(2), ZN => n5);
   U3 : AOI21_X1 port map( B1 => n8, B2 => n7, A => X(2), ZN => Z(0));
   U4 : OAI21_X1 port map( B1 => X(1), B2 => X(0), A => n7, ZN => n8);
   U5 : AND3_X1 port map( A1 => X(2), A2 => n7, A3 => n8, ZN => Z(2));
   U6 : NAND2_X1 port map( A1 => X(1), A2 => X(0), ZN => n7);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity encoder_N64_RADIX3_7 is

   port( X : in std_logic_vector (2 downto 0);  Z : out std_logic_vector (2 
         downto 0));

end encoder_N64_RADIX3_7;

architecture SYN_beh of encoder_N64_RADIX3_7 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n7, n8 : std_logic;

begin
   
   U1 : OAI22_X1 port map( A1 => n8, A2 => n5, B1 => X(2), B2 => n7, ZN => Z(1)
                           );
   U2 : INV_X1 port map( A => X(2), ZN => n5);
   U3 : AOI21_X1 port map( B1 => n8, B2 => n7, A => X(2), ZN => Z(0));
   U4 : OAI21_X1 port map( B1 => X(1), B2 => X(0), A => n7, ZN => n8);
   U5 : AND3_X1 port map( A1 => X(2), A2 => n7, A3 => n8, ZN => Z(2));
   U6 : NAND2_X1 port map( A1 => X(1), A2 => X(0), ZN => n7);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity encoder_N64_RADIX3_6 is

   port( X : in std_logic_vector (2 downto 0);  Z : out std_logic_vector (2 
         downto 0));

end encoder_N64_RADIX3_6;

architecture SYN_beh of encoder_N64_RADIX3_6 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n7, n8 : std_logic;

begin
   
   U1 : OAI22_X1 port map( A1 => n8, A2 => n5, B1 => X(2), B2 => n7, ZN => Z(1)
                           );
   U2 : INV_X1 port map( A => X(2), ZN => n5);
   U3 : AOI21_X1 port map( B1 => n8, B2 => n7, A => X(2), ZN => Z(0));
   U4 : OAI21_X1 port map( B1 => X(1), B2 => X(0), A => n7, ZN => n8);
   U5 : AND3_X1 port map( A1 => X(2), A2 => n7, A3 => n8, ZN => Z(2));
   U6 : NAND2_X1 port map( A1 => X(1), A2 => X(0), ZN => n7);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity encoder_N64_RADIX3_5 is

   port( X : in std_logic_vector (2 downto 0);  Z : out std_logic_vector (2 
         downto 0));

end encoder_N64_RADIX3_5;

architecture SYN_beh of encoder_N64_RADIX3_5 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n7, n8 : std_logic;

begin
   
   U1 : OAI22_X1 port map( A1 => n8, A2 => n5, B1 => X(2), B2 => n7, ZN => Z(1)
                           );
   U2 : INV_X1 port map( A => X(2), ZN => n5);
   U3 : AOI21_X1 port map( B1 => n8, B2 => n7, A => X(2), ZN => Z(0));
   U4 : OAI21_X1 port map( B1 => X(1), B2 => X(0), A => n7, ZN => n8);
   U5 : AND3_X1 port map( A1 => X(2), A2 => n7, A3 => n8, ZN => Z(2));
   U6 : NAND2_X1 port map( A1 => X(1), A2 => X(0), ZN => n7);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity encoder_N64_RADIX3_4 is

   port( X : in std_logic_vector (2 downto 0);  Z : out std_logic_vector (2 
         downto 0));

end encoder_N64_RADIX3_4;

architecture SYN_beh of encoder_N64_RADIX3_4 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n7, n8 : std_logic;

begin
   
   U1 : OAI22_X1 port map( A1 => n8, A2 => n5, B1 => X(2), B2 => n7, ZN => Z(1)
                           );
   U2 : INV_X1 port map( A => X(2), ZN => n5);
   U3 : AOI21_X1 port map( B1 => n8, B2 => n7, A => X(2), ZN => Z(0));
   U4 : OAI21_X1 port map( B1 => X(1), B2 => X(0), A => n7, ZN => n8);
   U5 : AND3_X1 port map( A1 => X(2), A2 => n7, A3 => n8, ZN => Z(2));
   U6 : NAND2_X1 port map( A1 => X(1), A2 => X(0), ZN => n7);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity encoder_N64_RADIX3_3 is

   port( X : in std_logic_vector (2 downto 0);  Z : out std_logic_vector (2 
         downto 0));

end encoder_N64_RADIX3_3;

architecture SYN_beh of encoder_N64_RADIX3_3 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n7, n8 : std_logic;

begin
   
   U1 : OAI22_X1 port map( A1 => n8, A2 => n5, B1 => X(2), B2 => n7, ZN => Z(1)
                           );
   U2 : INV_X1 port map( A => X(2), ZN => n5);
   U3 : AOI21_X1 port map( B1 => n8, B2 => n7, A => X(2), ZN => Z(0));
   U4 : OAI21_X1 port map( B1 => X(1), B2 => X(0), A => n7, ZN => n8);
   U5 : AND3_X1 port map( A1 => X(2), A2 => n7, A3 => n8, ZN => Z(2));
   U6 : NAND2_X1 port map( A1 => X(1), A2 => X(0), ZN => n7);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity encoder_N64_RADIX3_2 is

   port( X : in std_logic_vector (2 downto 0);  Z : out std_logic_vector (2 
         downto 0));

end encoder_N64_RADIX3_2;

architecture SYN_beh of encoder_N64_RADIX3_2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n7, n8 : std_logic;

begin
   
   U1 : OAI22_X1 port map( A1 => n8, A2 => n5, B1 => X(2), B2 => n7, ZN => Z(1)
                           );
   U2 : INV_X1 port map( A => X(2), ZN => n5);
   U3 : AOI21_X1 port map( B1 => n8, B2 => n7, A => X(2), ZN => Z(0));
   U4 : OAI21_X1 port map( B1 => X(1), B2 => X(0), A => n7, ZN => n8);
   U5 : AND3_X1 port map( A1 => X(2), A2 => n7, A3 => n8, ZN => Z(2));
   U6 : NAND2_X1 port map( A1 => X(1), A2 => X(0), ZN => n7);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity encoder_N64_RADIX3_1 is

   port( X : in std_logic_vector (2 downto 0);  Z : out std_logic_vector (2 
         downto 0));

end encoder_N64_RADIX3_1;

architecture SYN_beh of encoder_N64_RADIX3_1 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n7, n8 : std_logic;

begin
   
   U1 : OAI22_X1 port map( A1 => n8, A2 => n5, B1 => X(2), B2 => n7, ZN => Z(1)
                           );
   U2 : INV_X1 port map( A => X(2), ZN => n5);
   U3 : AOI21_X1 port map( B1 => n8, B2 => n7, A => X(2), ZN => Z(0));
   U4 : OAI21_X1 port map( B1 => X(1), B2 => X(0), A => n7, ZN => n8);
   U5 : AND3_X1 port map( A1 => X(2), A2 => n7, A3 => n8, ZN => Z(2));
   U6 : NAND2_X1 port map( A1 => X(1), A2 => X(0), ZN => n7);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_1_DW01_sub_0 is

   port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (63 downto 0);  CO : out std_logic);

end complementer_N64_1_DW01_sub_0;

architecture SYN_rpl of complementer_N64_1_DW01_sub_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal DIFF_62_port, DIFF_63_port, DIFF_31_port, DIFF_32_port, DIFF_33_port,
      DIFF_34_port, DIFF_35_port, DIFF_36_port, DIFF_37_port, DIFF_38_port, 
      DIFF_39_port, DIFF_40_port, DIFF_41_port, DIFF_42_port, DIFF_43_port, 
      DIFF_44_port, DIFF_45_port, DIFF_46_port, DIFF_47_port, DIFF_48_port, 
      DIFF_49_port, DIFF_50_port, DIFF_51_port, DIFF_52_port, DIFF_53_port, 
      DIFF_54_port, DIFF_55_port, DIFF_56_port, DIFF_57_port, DIFF_58_port, 
      DIFF_59_port, DIFF_60_port, DIFF_61_port, DIFF_3_port, DIFF_4_port, 
      DIFF_5_port, DIFF_6_port, DIFF_7_port, DIFF_8_port, DIFF_9_port, 
      DIFF_10_port, DIFF_11_port, DIFF_12_port, DIFF_13_port, DIFF_14_port, 
      DIFF_15_port, DIFF_16_port, DIFF_17_port, DIFF_18_port, DIFF_19_port, 
      DIFF_20_port, DIFF_21_port, DIFF_22_port, DIFF_23_port, DIFF_24_port, 
      DIFF_25_port, DIFF_26_port, DIFF_27_port, DIFF_28_port, DIFF_29_port, 
      DIFF_30_port, DIFF_2_port, DIFF_1_port, n190, n191, n192, n194, n195, 
      n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, 
      n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, 
      n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, 
      n232, n233, n234, n235, n237, n238, n239, n241, n242, n243, n245, n246, 
      n247, n249, n250, n189, n193, n236, n240, n244, n248, n251 : std_logic;

begin
   DIFF <= ( DIFF_63_port, DIFF_62_port, DIFF_61_port, DIFF_60_port, 
      DIFF_59_port, DIFF_58_port, DIFF_57_port, DIFF_56_port, DIFF_55_port, 
      DIFF_54_port, DIFF_53_port, DIFF_52_port, DIFF_51_port, DIFF_50_port, 
      DIFF_49_port, DIFF_48_port, DIFF_47_port, DIFF_46_port, DIFF_45_port, 
      DIFF_44_port, DIFF_43_port, DIFF_42_port, DIFF_41_port, DIFF_40_port, 
      DIFF_39_port, DIFF_38_port, DIFF_37_port, DIFF_36_port, DIFF_35_port, 
      DIFF_34_port, DIFF_33_port, DIFF_32_port, DIFF_31_port, DIFF_30_port, 
      DIFF_29_port, DIFF_28_port, DIFF_27_port, DIFF_26_port, DIFF_25_port, 
      DIFF_24_port, DIFF_23_port, DIFF_22_port, DIFF_21_port, DIFF_20_port, 
      DIFF_19_port, DIFF_18_port, DIFF_17_port, DIFF_16_port, DIFF_15_port, 
      DIFF_14_port, DIFF_13_port, DIFF_12_port, DIFF_11_port, DIFF_10_port, 
      DIFF_9_port, DIFF_8_port, DIFF_7_port, DIFF_6_port, DIFF_5_port, 
      DIFF_4_port, DIFF_3_port, DIFF_2_port, DIFF_1_port, B(0) );
   
   U81 : XOR2_X1 port map( A => n190, B => B(9), Z => DIFF_9_port);
   U82 : XOR2_X1 port map( A => n192, B => B(7), Z => DIFF_7_port);
   U84 : XOR2_X1 port map( A => n195, B => B(63), Z => DIFF_63_port);
   U85 : XOR2_X1 port map( A => n196, B => B(62), Z => DIFF_62_port);
   U86 : XOR2_X1 port map( A => n194, B => B(5), Z => DIFF_5_port);
   U87 : XOR2_X1 port map( A => n198, B => B(59), Z => DIFF_59_port);
   U88 : XOR2_X1 port map( A => n201, B => B(58), Z => DIFF_58_port);
   U89 : XOR2_X1 port map( A => n200, B => B(57), Z => DIFF_57_port);
   U90 : XOR2_X1 port map( A => n202, B => B(55), Z => DIFF_55_port);
   U91 : XOR2_X1 port map( A => n205, B => B(54), Z => DIFF_54_port);
   U92 : XOR2_X1 port map( A => n204, B => B(53), Z => DIFF_53_port);
   U93 : XOR2_X1 port map( A => n206, B => B(51), Z => DIFF_51_port);
   U94 : XOR2_X1 port map( A => n209, B => B(50), Z => DIFF_50_port);
   U95 : XOR2_X1 port map( A => n208, B => B(49), Z => DIFF_49_port);
   U96 : XOR2_X1 port map( A => n212, B => B(47), Z => DIFF_47_port);
   U97 : XOR2_X1 port map( A => n215, B => B(46), Z => DIFF_46_port);
   U98 : XOR2_X1 port map( A => n214, B => B(45), Z => DIFF_45_port);
   U99 : XOR2_X1 port map( A => n216, B => B(43), Z => DIFF_43_port);
   U100 : XOR2_X1 port map( A => n219, B => B(42), Z => DIFF_42_port);
   U101 : XOR2_X1 port map( A => n218, B => B(41), Z => DIFF_41_port);
   U102 : XOR2_X1 port map( A => n211, B => B(3), Z => DIFF_3_port);
   U103 : XOR2_X1 port map( A => n220, B => B(39), Z => DIFF_39_port);
   U104 : XOR2_X1 port map( A => n223, B => B(38), Z => DIFF_38_port);
   U105 : XOR2_X1 port map( A => n222, B => B(37), Z => DIFF_37_port);
   U106 : XOR2_X1 port map( A => n224, B => B(35), Z => DIFF_35_port);
   U107 : XOR2_X1 port map( A => n227, B => B(34), Z => DIFF_34_port);
   U108 : XOR2_X1 port map( A => n226, B => B(33), Z => DIFF_33_port);
   U109 : XOR2_X1 port map( A => n228, B => B(31), Z => DIFF_31_port);
   U110 : XOR2_X1 port map( A => n231, B => B(30), Z => DIFF_30_port);
   U111 : XOR2_X1 port map( A => n230, B => B(29), Z => DIFF_29_port);
   U112 : XOR2_X1 port map( A => n233, B => B(27), Z => DIFF_27_port);
   U114 : XOR2_X1 port map( A => n235, B => B(25), Z => DIFF_25_port);
   U115 : XOR2_X1 port map( A => n237, B => B(23), Z => DIFF_23_port);
   U117 : XOR2_X1 port map( A => n239, B => B(21), Z => DIFF_21_port);
   U118 : XOR2_X1 port map( A => B(1), B => B(0), Z => DIFF_1_port);
   U119 : XOR2_X1 port map( A => n241, B => B(19), Z => DIFF_19_port);
   U121 : XOR2_X1 port map( A => n243, B => B(17), Z => DIFF_17_port);
   U122 : XOR2_X1 port map( A => n245, B => B(15), Z => DIFF_15_port);
   U124 : XOR2_X1 port map( A => n247, B => B(13), Z => DIFF_13_port);
   U125 : XOR2_X1 port map( A => n249, B => B(11), Z => DIFF_11_port);
   U1 : NAND2_X1 port map( A1 => n197, A2 => n251, ZN => n196);
   U2 : NOR2_X1 port map( A1 => B(55), A2 => n202, ZN => n203);
   U3 : NOR2_X1 port map( A1 => B(51), A2 => n206, ZN => n207);
   U4 : NOR2_X1 port map( A1 => B(47), A2 => n212, ZN => n213);
   U5 : NOR2_X1 port map( A1 => B(43), A2 => n216, ZN => n217);
   U6 : OR3_X1 port map( A1 => B(53), A2 => B(54), A3 => n204, ZN => n202);
   U7 : OR3_X1 port map( A1 => B(49), A2 => B(50), A3 => n208, ZN => n206);
   U8 : OR3_X1 port map( A1 => B(45), A2 => B(46), A3 => n214, ZN => n212);
   U9 : OR3_X1 port map( A1 => B(41), A2 => B(42), A3 => n218, ZN => n216);
   U10 : OR3_X1 port map( A1 => B(55), A2 => B(56), A3 => n202, ZN => n200);
   U11 : OR3_X1 port map( A1 => B(51), A2 => B(52), A3 => n206, ZN => n204);
   U12 : OR3_X1 port map( A1 => B(47), A2 => B(48), A3 => n212, ZN => n208);
   U13 : OR3_X1 port map( A1 => B(43), A2 => B(44), A3 => n216, ZN => n214);
   U14 : OR2_X1 port map( A1 => n204, A2 => B(53), ZN => n205);
   U15 : OR2_X1 port map( A1 => n208, A2 => B(49), ZN => n209);
   U16 : OR2_X1 port map( A1 => n214, A2 => B(45), ZN => n215);
   U17 : OR2_X1 port map( A1 => n218, A2 => B(41), ZN => n219);
   U18 : NOR3_X1 port map( A1 => B(59), A2 => B(60), A3 => n198, ZN => n197);
   U19 : NOR2_X1 port map( A1 => B(59), A2 => n198, ZN => n199);
   U20 : OR3_X1 port map( A1 => B(57), A2 => B(58), A3 => n200, ZN => n198);
   U21 : OR2_X1 port map( A1 => n196, A2 => B(62), ZN => n195);
   U22 : OR2_X1 port map( A1 => n200, A2 => B(57), ZN => n201);
   U23 : NOR2_X1 port map( A1 => B(39), A2 => n220, ZN => n221);
   U24 : OR3_X1 port map( A1 => B(39), A2 => B(40), A3 => n220, ZN => n218);
   U25 : OR3_X1 port map( A1 => B(37), A2 => B(38), A3 => n222, ZN => n220);
   U26 : OR2_X1 port map( A1 => n222, A2 => B(37), ZN => n223);
   U27 : XNOR2_X1 port map( A => B(60), B => n199, ZN => DIFF_60_port);
   U28 : NOR2_X1 port map( A1 => B(35), A2 => n224, ZN => n225);
   U29 : XNOR2_X1 port map( A => B(56), B => n203, ZN => DIFF_56_port);
   U30 : XNOR2_X1 port map( A => B(52), B => n207, ZN => DIFF_52_port);
   U31 : OR3_X1 port map( A1 => B(35), A2 => B(36), A3 => n224, ZN => n222);
   U32 : XNOR2_X1 port map( A => B(48), B => n213, ZN => DIFF_48_port);
   U33 : XNOR2_X1 port map( A => B(44), B => n217, ZN => DIFF_44_port);
   U34 : XNOR2_X1 port map( A => B(40), B => n221, ZN => DIFF_40_port);
   U35 : XNOR2_X1 port map( A => B(36), B => n225, ZN => DIFF_36_port);
   U36 : XNOR2_X1 port map( A => n197, B => B(61), ZN => DIFF_61_port);
   U37 : XNOR2_X1 port map( A => B(32), B => n229, ZN => DIFF_32_port);
   U38 : OR3_X1 port map( A1 => B(33), A2 => B(34), A3 => n226, ZN => n224);
   U39 : OR2_X1 port map( A1 => n226, A2 => B(33), ZN => n227);
   U40 : NOR2_X1 port map( A1 => B(31), A2 => n228, ZN => n229);
   U41 : OR3_X1 port map( A1 => B(31), A2 => B(32), A3 => n228, ZN => n226);
   U42 : XNOR2_X1 port map( A => n189, B => B(26), ZN => DIFF_26_port);
   U43 : NOR2_X1 port map( A1 => n235, A2 => B(25), ZN => n189);
   U44 : XNOR2_X1 port map( A => n193, B => B(22), ZN => DIFF_22_port);
   U45 : NOR2_X1 port map( A1 => n239, A2 => B(21), ZN => n193);
   U46 : XNOR2_X1 port map( A => n236, B => B(18), ZN => DIFF_18_port);
   U47 : NOR2_X1 port map( A1 => n243, A2 => B(17), ZN => n236);
   U48 : XNOR2_X1 port map( A => n240, B => B(14), ZN => DIFF_14_port);
   U49 : NOR2_X1 port map( A1 => n247, A2 => B(13), ZN => n240);
   U50 : XNOR2_X1 port map( A => n244, B => B(10), ZN => DIFF_10_port);
   U51 : NOR2_X1 port map( A1 => n190, A2 => B(9), ZN => n244);
   U52 : XNOR2_X1 port map( A => n248, B => B(6), ZN => DIFF_6_port);
   U53 : NOR2_X1 port map( A1 => n194, A2 => B(5), ZN => n248);
   U54 : XNOR2_X1 port map( A => B(28), B => n234, ZN => DIFF_28_port);
   U55 : NOR2_X1 port map( A1 => B(27), A2 => n233, ZN => n234);
   U56 : XNOR2_X1 port map( A => B(24), B => n238, ZN => DIFF_24_port);
   U57 : NOR2_X1 port map( A1 => B(23), A2 => n237, ZN => n238);
   U58 : XNOR2_X1 port map( A => B(20), B => n242, ZN => DIFF_20_port);
   U59 : NOR2_X1 port map( A1 => B(19), A2 => n241, ZN => n242);
   U60 : XNOR2_X1 port map( A => B(16), B => n246, ZN => DIFF_16_port);
   U61 : NOR2_X1 port map( A1 => B(15), A2 => n245, ZN => n246);
   U62 : XNOR2_X1 port map( A => B(12), B => n250, ZN => DIFF_12_port);
   U63 : NOR2_X1 port map( A1 => B(11), A2 => n249, ZN => n250);
   U64 : XNOR2_X1 port map( A => B(8), B => n191, ZN => DIFF_8_port);
   U65 : NOR2_X1 port map( A1 => B(7), A2 => n192, ZN => n191);
   U66 : XNOR2_X1 port map( A => B(2), B => n232, ZN => DIFF_2_port);
   U67 : NOR2_X1 port map( A1 => B(0), A2 => B(1), ZN => n232);
   U68 : XNOR2_X1 port map( A => B(4), B => n210, ZN => DIFF_4_port);
   U69 : NOR2_X1 port map( A1 => B(3), A2 => n211, ZN => n210);
   U70 : OR3_X1 port map( A1 => B(5), A2 => B(6), A3 => n194, ZN => n192);
   U71 : OR3_X1 port map( A1 => B(10), A2 => B(9), A3 => n190, ZN => n249);
   U72 : OR3_X1 port map( A1 => B(13), A2 => B(14), A3 => n247, ZN => n245);
   U73 : OR3_X1 port map( A1 => B(17), A2 => B(18), A3 => n243, ZN => n241);
   U74 : OR3_X1 port map( A1 => B(21), A2 => B(22), A3 => n239, ZN => n237);
   U75 : OR3_X1 port map( A1 => B(25), A2 => B(26), A3 => n235, ZN => n233);
   U76 : OR3_X1 port map( A1 => B(29), A2 => B(30), A3 => n230, ZN => n228);
   U77 : OR3_X1 port map( A1 => B(7), A2 => B(8), A3 => n192, ZN => n190);
   U78 : OR3_X1 port map( A1 => B(11), A2 => B(12), A3 => n249, ZN => n247);
   U79 : OR3_X1 port map( A1 => B(15), A2 => B(16), A3 => n245, ZN => n243);
   U80 : OR3_X1 port map( A1 => B(19), A2 => B(20), A3 => n241, ZN => n239);
   U83 : OR3_X1 port map( A1 => B(23), A2 => B(24), A3 => n237, ZN => n235);
   U113 : OR3_X1 port map( A1 => B(27), A2 => B(28), A3 => n233, ZN => n230);
   U116 : OR3_X1 port map( A1 => B(3), A2 => B(4), A3 => n211, ZN => n194);
   U120 : OR2_X1 port map( A1 => n230, A2 => B(29), ZN => n231);
   U123 : OR3_X1 port map( A1 => B(1), A2 => B(2), A3 => B(0), ZN => n211);
   U126 : INV_X1 port map( A => B(61), ZN => n251);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_2_DW01_sub_0 is

   port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (63 downto 0);  CO : out std_logic);

end complementer_N64_2_DW01_sub_0;

architecture SYN_rpl of complementer_N64_2_DW01_sub_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal DIFF_62_port, DIFF_61_port, DIFF_60_port, DIFF_59_port, DIFF_58_port,
      DIFF_57_port, DIFF_56_port, DIFF_55_port, DIFF_54_port, DIFF_53_port, 
      DIFF_52_port, DIFF_51_port, DIFF_50_port, DIFF_49_port, DIFF_48_port, 
      DIFF_47_port, DIFF_46_port, DIFF_45_port, DIFF_44_port, DIFF_43_port, 
      DIFF_42_port, DIFF_41_port, DIFF_40_port, DIFF_39_port, DIFF_38_port, 
      DIFF_37_port, DIFF_36_port, DIFF_35_port, DIFF_34_port, DIFF_33_port, 
      DIFF_32_port, DIFF_31_port, DIFF_30_port, DIFF_29_port, DIFF_28_port, 
      DIFF_27_port, DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, 
      DIFF_22_port, DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, 
      DIFF_17_port, DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, 
      DIFF_12_port, DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, 
      DIFF_7_port, DIFF_6_port, DIFF_5_port, DIFF_4_port, DIFF_3_port, 
      DIFF_2_port, DIFF_1_port, DIFF_63_port, n190, n191, n192, n193, n194, 
      n196, n197, n198, n199, n200, n202, n203, n204, n206, n207, n208, n210, 
      n211, n212, n213, n214, n216, n217, n218, n220, n221, n222, n224, n225, 
      n226, n228, n229, n230, n232, n233, n234, n235, n236, n237, n238, n239, 
      n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, 
      n189, n195, n201, n205, n209, n215, n219, n223, n227, n231 : std_logic;

begin
   DIFF <= ( DIFF_63_port, DIFF_62_port, DIFF_61_port, DIFF_60_port, 
      DIFF_59_port, DIFF_58_port, DIFF_57_port, DIFF_56_port, DIFF_55_port, 
      DIFF_54_port, DIFF_53_port, DIFF_52_port, DIFF_51_port, DIFF_50_port, 
      DIFF_49_port, DIFF_48_port, DIFF_47_port, DIFF_46_port, DIFF_45_port, 
      DIFF_44_port, DIFF_43_port, DIFF_42_port, DIFF_41_port, DIFF_40_port, 
      DIFF_39_port, DIFF_38_port, DIFF_37_port, DIFF_36_port, DIFF_35_port, 
      DIFF_34_port, DIFF_33_port, DIFF_32_port, DIFF_31_port, DIFF_30_port, 
      DIFF_29_port, DIFF_28_port, DIFF_27_port, DIFF_26_port, DIFF_25_port, 
      DIFF_24_port, DIFF_23_port, DIFF_22_port, DIFF_21_port, DIFF_20_port, 
      DIFF_19_port, DIFF_18_port, DIFF_17_port, DIFF_16_port, DIFF_15_port, 
      DIFF_14_port, DIFF_13_port, DIFF_12_port, DIFF_11_port, DIFF_10_port, 
      DIFF_9_port, DIFF_8_port, DIFF_7_port, DIFF_6_port, DIFF_5_port, 
      DIFF_4_port, DIFF_3_port, DIFF_2_port, DIFF_1_port, B(0) );
   
   U81 : XOR2_X1 port map( A => n190, B => B(9), Z => DIFF_9_port);
   U82 : XOR2_X1 port map( A => n192, B => B(7), Z => DIFF_7_port);
   U83 : XOR2_X1 port map( A => n193, B => B(6), Z => DIFF_6_port);
   U85 : XOR2_X1 port map( A => n196, B => B(62), Z => DIFF_62_port);
   U86 : XOR2_X1 port map( A => n194, B => B(5), Z => DIFF_5_port);
   U87 : XOR2_X1 port map( A => n198, B => B(59), Z => DIFF_59_port);
   U89 : XOR2_X1 port map( A => n200, B => B(57), Z => DIFF_57_port);
   U90 : XOR2_X1 port map( A => n202, B => B(55), Z => DIFF_55_port);
   U92 : XOR2_X1 port map( A => n204, B => B(53), Z => DIFF_53_port);
   U93 : XOR2_X1 port map( A => n206, B => B(51), Z => DIFF_51_port);
   U95 : XOR2_X1 port map( A => n208, B => B(49), Z => DIFF_49_port);
   U96 : XOR2_X1 port map( A => n212, B => B(47), Z => DIFF_47_port);
   U98 : XOR2_X1 port map( A => n214, B => B(45), Z => DIFF_45_port);
   U99 : XOR2_X1 port map( A => n216, B => B(43), Z => DIFF_43_port);
   U101 : XOR2_X1 port map( A => n218, B => B(41), Z => DIFF_41_port);
   U102 : XOR2_X1 port map( A => n211, B => B(3), Z => DIFF_3_port);
   U103 : XOR2_X1 port map( A => n220, B => B(39), Z => DIFF_39_port);
   U105 : XOR2_X1 port map( A => n222, B => B(37), Z => DIFF_37_port);
   U106 : XOR2_X1 port map( A => n224, B => B(35), Z => DIFF_35_port);
   U108 : XOR2_X1 port map( A => n226, B => B(33), Z => DIFF_33_port);
   U109 : XOR2_X1 port map( A => n228, B => B(31), Z => DIFF_31_port);
   U111 : XOR2_X1 port map( A => n230, B => B(29), Z => DIFF_29_port);
   U112 : XOR2_X1 port map( A => n233, B => B(27), Z => DIFF_27_port);
   U113 : XOR2_X1 port map( A => n236, B => B(26), Z => DIFF_26_port);
   U114 : XOR2_X1 port map( A => n235, B => B(25), Z => DIFF_25_port);
   U115 : XOR2_X1 port map( A => n237, B => B(23), Z => DIFF_23_port);
   U116 : XOR2_X1 port map( A => n240, B => B(22), Z => DIFF_22_port);
   U117 : XOR2_X1 port map( A => n239, B => B(21), Z => DIFF_21_port);
   U118 : XOR2_X1 port map( A => B(1), B => B(0), Z => DIFF_1_port);
   U119 : XOR2_X1 port map( A => n241, B => B(19), Z => DIFF_19_port);
   U120 : XOR2_X1 port map( A => n244, B => B(18), Z => DIFF_18_port);
   U121 : XOR2_X1 port map( A => n243, B => B(17), Z => DIFF_17_port);
   U122 : XOR2_X1 port map( A => n245, B => B(15), Z => DIFF_15_port);
   U123 : XOR2_X1 port map( A => n248, B => B(14), Z => DIFF_14_port);
   U124 : XOR2_X1 port map( A => n247, B => B(13), Z => DIFF_13_port);
   U125 : XOR2_X1 port map( A => n249, B => B(11), Z => DIFF_11_port);
   U126 : XOR2_X1 port map( A => n251, B => B(10), Z => DIFF_10_port);
   U1 : XOR2_X1 port map( A => n197, B => n231, Z => DIFF_61_port);
   U2 : NAND2_X1 port map( A1 => n197, A2 => n231, ZN => n196);
   U3 : XNOR2_X1 port map( A => n189, B => B(54), ZN => DIFF_54_port);
   U4 : NOR2_X1 port map( A1 => n204, A2 => B(53), ZN => n189);
   U5 : XNOR2_X1 port map( A => n195, B => B(58), ZN => DIFF_58_port);
   U6 : NOR2_X1 port map( A1 => n200, A2 => B(57), ZN => n195);
   U7 : XNOR2_X1 port map( A => B(60), B => n199, ZN => DIFF_60_port);
   U8 : NOR2_X1 port map( A1 => B(59), A2 => n198, ZN => n199);
   U9 : XNOR2_X1 port map( A => B(56), B => n203, ZN => DIFF_56_port);
   U10 : NOR2_X1 port map( A1 => B(55), A2 => n202, ZN => n203);
   U11 : XNOR2_X1 port map( A => B(52), B => n207, ZN => DIFF_52_port);
   U12 : NOR2_X1 port map( A1 => B(51), A2 => n206, ZN => n207);
   U13 : XNOR2_X1 port map( A => B(48), B => n213, ZN => DIFF_48_port);
   U14 : NOR2_X1 port map( A1 => B(47), A2 => n212, ZN => n213);
   U15 : XNOR2_X1 port map( A => B(44), B => n217, ZN => DIFF_44_port);
   U16 : NOR2_X1 port map( A1 => B(43), A2 => n216, ZN => n217);
   U17 : OR3_X1 port map( A1 => B(57), A2 => B(58), A3 => n200, ZN => n198);
   U18 : OR3_X1 port map( A1 => B(41), A2 => B(42), A3 => n218, ZN => n216);
   U19 : OR3_X1 port map( A1 => B(45), A2 => B(46), A3 => n214, ZN => n212);
   U20 : OR3_X1 port map( A1 => B(49), A2 => B(50), A3 => n208, ZN => n206);
   U21 : OR3_X1 port map( A1 => B(53), A2 => B(54), A3 => n204, ZN => n202);
   U22 : OR3_X1 port map( A1 => B(43), A2 => B(44), A3 => n216, ZN => n214);
   U23 : OR3_X1 port map( A1 => B(47), A2 => B(48), A3 => n212, ZN => n208);
   U24 : OR3_X1 port map( A1 => B(51), A2 => B(52), A3 => n206, ZN => n204);
   U25 : OR3_X1 port map( A1 => B(55), A2 => B(56), A3 => n202, ZN => n200);
   U26 : XNOR2_X1 port map( A => n201, B => B(50), ZN => DIFF_50_port);
   U27 : NOR2_X1 port map( A1 => n208, A2 => B(49), ZN => n201);
   U28 : XNOR2_X1 port map( A => n205, B => B(46), ZN => DIFF_46_port);
   U29 : NOR2_X1 port map( A1 => n214, A2 => B(45), ZN => n205);
   U30 : XNOR2_X1 port map( A => n209, B => B(42), ZN => DIFF_42_port);
   U31 : NOR2_X1 port map( A1 => n218, A2 => B(41), ZN => n209);
   U32 : NOR3_X1 port map( A1 => B(59), A2 => B(60), A3 => n198, ZN => n197);
   U33 : XNOR2_X1 port map( A => B(40), B => n221, ZN => DIFF_40_port);
   U34 : NOR2_X1 port map( A1 => B(39), A2 => n220, ZN => n221);
   U35 : OR3_X1 port map( A1 => B(39), A2 => B(40), A3 => n220, ZN => n218);
   U36 : XNOR2_X1 port map( A => n215, B => B(63), ZN => DIFF_63_port);
   U37 : NOR2_X1 port map( A1 => n196, A2 => B(62), ZN => n215);
   U38 : OR3_X1 port map( A1 => B(37), A2 => B(38), A3 => n222, ZN => n220);
   U39 : XNOR2_X1 port map( A => n219, B => B(38), ZN => DIFF_38_port);
   U40 : NOR2_X1 port map( A1 => n222, A2 => B(37), ZN => n219);
   U41 : XNOR2_X1 port map( A => B(36), B => n225, ZN => DIFF_36_port);
   U42 : NOR2_X1 port map( A1 => B(35), A2 => n224, ZN => n225);
   U43 : OR3_X1 port map( A1 => B(35), A2 => B(36), A3 => n224, ZN => n222);
   U44 : XNOR2_X1 port map( A => n223, B => B(34), ZN => DIFF_34_port);
   U45 : NOR2_X1 port map( A1 => n226, A2 => B(33), ZN => n223);
   U46 : OR3_X1 port map( A1 => B(33), A2 => B(34), A3 => n226, ZN => n224);
   U47 : XNOR2_X1 port map( A => B(32), B => n229, ZN => DIFF_32_port);
   U48 : NOR2_X1 port map( A1 => B(31), A2 => n228, ZN => n229);
   U49 : OR3_X1 port map( A1 => B(31), A2 => B(32), A3 => n228, ZN => n226);
   U50 : XNOR2_X1 port map( A => n227, B => B(30), ZN => DIFF_30_port);
   U51 : NOR2_X1 port map( A1 => n230, A2 => B(29), ZN => n227);
   U52 : OR3_X1 port map( A1 => B(29), A2 => B(30), A3 => n230, ZN => n228);
   U53 : NOR2_X1 port map( A1 => B(27), A2 => n233, ZN => n234);
   U54 : NOR2_X1 port map( A1 => B(23), A2 => n237, ZN => n238);
   U55 : NOR2_X1 port map( A1 => B(19), A2 => n241, ZN => n242);
   U56 : NOR2_X1 port map( A1 => B(15), A2 => n245, ZN => n246);
   U57 : NOR2_X1 port map( A1 => B(11), A2 => n249, ZN => n250);
   U58 : NOR2_X1 port map( A1 => B(7), A2 => n192, ZN => n191);
   U59 : NOR2_X1 port map( A1 => B(3), A2 => n211, ZN => n210);
   U60 : OR3_X1 port map( A1 => B(25), A2 => B(26), A3 => n235, ZN => n233);
   U61 : OR3_X1 port map( A1 => B(21), A2 => B(22), A3 => n239, ZN => n237);
   U62 : OR3_X1 port map( A1 => B(17), A2 => B(18), A3 => n243, ZN => n241);
   U63 : OR3_X1 port map( A1 => B(13), A2 => B(14), A3 => n247, ZN => n245);
   U64 : OR3_X1 port map( A1 => B(10), A2 => B(9), A3 => n190, ZN => n249);
   U65 : OR3_X1 port map( A1 => B(5), A2 => B(6), A3 => n194, ZN => n192);
   U66 : OR3_X1 port map( A1 => B(27), A2 => B(28), A3 => n233, ZN => n230);
   U67 : OR3_X1 port map( A1 => B(23), A2 => B(24), A3 => n237, ZN => n235);
   U68 : OR3_X1 port map( A1 => B(19), A2 => B(20), A3 => n241, ZN => n239);
   U69 : OR3_X1 port map( A1 => B(15), A2 => B(16), A3 => n245, ZN => n243);
   U70 : OR3_X1 port map( A1 => B(11), A2 => B(12), A3 => n249, ZN => n247);
   U71 : OR3_X1 port map( A1 => B(7), A2 => B(8), A3 => n192, ZN => n190);
   U72 : OR3_X1 port map( A1 => B(3), A2 => B(4), A3 => n211, ZN => n194);
   U73 : XNOR2_X1 port map( A => B(28), B => n234, ZN => DIFF_28_port);
   U74 : XNOR2_X1 port map( A => B(24), B => n238, ZN => DIFF_24_port);
   U75 : XNOR2_X1 port map( A => B(20), B => n242, ZN => DIFF_20_port);
   U76 : XNOR2_X1 port map( A => B(16), B => n246, ZN => DIFF_16_port);
   U77 : XNOR2_X1 port map( A => B(12), B => n250, ZN => DIFF_12_port);
   U78 : XNOR2_X1 port map( A => B(8), B => n191, ZN => DIFF_8_port);
   U79 : XNOR2_X1 port map( A => B(4), B => n210, ZN => DIFF_4_port);
   U80 : XNOR2_X1 port map( A => B(2), B => n232, ZN => DIFF_2_port);
   U84 : OR2_X1 port map( A1 => n235, A2 => B(25), ZN => n236);
   U88 : OR2_X1 port map( A1 => n239, A2 => B(21), ZN => n240);
   U91 : OR2_X1 port map( A1 => n243, A2 => B(17), ZN => n244);
   U94 : OR2_X1 port map( A1 => n247, A2 => B(13), ZN => n248);
   U97 : OR2_X1 port map( A1 => n190, A2 => B(9), ZN => n251);
   U100 : OR2_X1 port map( A1 => n194, A2 => B(5), ZN => n193);
   U104 : OR3_X1 port map( A1 => B(1), A2 => B(2), A3 => B(0), ZN => n211);
   U107 : NOR2_X1 port map( A1 => B(0), A2 => B(1), ZN => n232);
   U110 : INV_X1 port map( A => B(61), ZN => n231);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_3_DW01_sub_0 is

   port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (63 downto 0);  CO : out std_logic);

end complementer_N64_3_DW01_sub_0;

architecture SYN_rpl of complementer_N64_3_DW01_sub_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal DIFF_62_port, DIFF_63_port, DIFF_29_port, DIFF_30_port, DIFF_31_port,
      DIFF_32_port, DIFF_33_port, DIFF_34_port, DIFF_35_port, DIFF_36_port, 
      DIFF_37_port, DIFF_38_port, DIFF_39_port, DIFF_40_port, DIFF_41_port, 
      DIFF_42_port, DIFF_43_port, DIFF_44_port, DIFF_45_port, DIFF_46_port, 
      DIFF_47_port, DIFF_48_port, DIFF_49_port, DIFF_50_port, DIFF_51_port, 
      DIFF_52_port, DIFF_53_port, DIFF_54_port, DIFF_55_port, DIFF_56_port, 
      DIFF_57_port, DIFF_58_port, DIFF_59_port, DIFF_60_port, DIFF_61_port, 
      DIFF_3_port, DIFF_4_port, DIFF_5_port, DIFF_6_port, DIFF_7_port, 
      DIFF_8_port, DIFF_9_port, DIFF_10_port, DIFF_11_port, DIFF_12_port, 
      DIFF_13_port, DIFF_14_port, DIFF_15_port, DIFF_16_port, DIFF_17_port, 
      DIFF_18_port, DIFF_19_port, DIFF_20_port, DIFF_21_port, DIFF_22_port, 
      DIFF_23_port, DIFF_24_port, DIFF_25_port, DIFF_26_port, DIFF_27_port, 
      DIFF_28_port, DIFF_2_port, DIFF_1_port, n190, n191, n192, n194, n195, 
      n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, 
      n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, 
      n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, 
      n232, n233, n234, n235, n237, n238, n239, n241, n242, n243, n245, n246, 
      n247, n249, n250, n189, n193, n236, n240, n244, n248, n251 : std_logic;

begin
   DIFF <= ( DIFF_63_port, DIFF_62_port, DIFF_61_port, DIFF_60_port, 
      DIFF_59_port, DIFF_58_port, DIFF_57_port, DIFF_56_port, DIFF_55_port, 
      DIFF_54_port, DIFF_53_port, DIFF_52_port, DIFF_51_port, DIFF_50_port, 
      DIFF_49_port, DIFF_48_port, DIFF_47_port, DIFF_46_port, DIFF_45_port, 
      DIFF_44_port, DIFF_43_port, DIFF_42_port, DIFF_41_port, DIFF_40_port, 
      DIFF_39_port, DIFF_38_port, DIFF_37_port, DIFF_36_port, DIFF_35_port, 
      DIFF_34_port, DIFF_33_port, DIFF_32_port, DIFF_31_port, DIFF_30_port, 
      DIFF_29_port, DIFF_28_port, DIFF_27_port, DIFF_26_port, DIFF_25_port, 
      DIFF_24_port, DIFF_23_port, DIFF_22_port, DIFF_21_port, DIFF_20_port, 
      DIFF_19_port, DIFF_18_port, DIFF_17_port, DIFF_16_port, DIFF_15_port, 
      DIFF_14_port, DIFF_13_port, DIFF_12_port, DIFF_11_port, DIFF_10_port, 
      DIFF_9_port, DIFF_8_port, DIFF_7_port, DIFF_6_port, DIFF_5_port, 
      DIFF_4_port, DIFF_3_port, DIFF_2_port, DIFF_1_port, B(0) );
   
   U81 : XOR2_X1 port map( A => n190, B => B(9), Z => DIFF_9_port);
   U82 : XOR2_X1 port map( A => n192, B => B(7), Z => DIFF_7_port);
   U84 : XOR2_X1 port map( A => n195, B => B(63), Z => DIFF_63_port);
   U85 : XOR2_X1 port map( A => n196, B => B(62), Z => DIFF_62_port);
   U86 : XOR2_X1 port map( A => n194, B => B(5), Z => DIFF_5_port);
   U87 : XOR2_X1 port map( A => n198, B => B(59), Z => DIFF_59_port);
   U88 : XOR2_X1 port map( A => n201, B => B(58), Z => DIFF_58_port);
   U89 : XOR2_X1 port map( A => n200, B => B(57), Z => DIFF_57_port);
   U90 : XOR2_X1 port map( A => n202, B => B(55), Z => DIFF_55_port);
   U91 : XOR2_X1 port map( A => n205, B => B(54), Z => DIFF_54_port);
   U92 : XOR2_X1 port map( A => n204, B => B(53), Z => DIFF_53_port);
   U93 : XOR2_X1 port map( A => n206, B => B(51), Z => DIFF_51_port);
   U94 : XOR2_X1 port map( A => n209, B => B(50), Z => DIFF_50_port);
   U95 : XOR2_X1 port map( A => n208, B => B(49), Z => DIFF_49_port);
   U96 : XOR2_X1 port map( A => n212, B => B(47), Z => DIFF_47_port);
   U97 : XOR2_X1 port map( A => n215, B => B(46), Z => DIFF_46_port);
   U98 : XOR2_X1 port map( A => n214, B => B(45), Z => DIFF_45_port);
   U99 : XOR2_X1 port map( A => n216, B => B(43), Z => DIFF_43_port);
   U100 : XOR2_X1 port map( A => n219, B => B(42), Z => DIFF_42_port);
   U101 : XOR2_X1 port map( A => n218, B => B(41), Z => DIFF_41_port);
   U102 : XOR2_X1 port map( A => n211, B => B(3), Z => DIFF_3_port);
   U103 : XOR2_X1 port map( A => n220, B => B(39), Z => DIFF_39_port);
   U104 : XOR2_X1 port map( A => n223, B => B(38), Z => DIFF_38_port);
   U105 : XOR2_X1 port map( A => n222, B => B(37), Z => DIFF_37_port);
   U106 : XOR2_X1 port map( A => n224, B => B(35), Z => DIFF_35_port);
   U107 : XOR2_X1 port map( A => n227, B => B(34), Z => DIFF_34_port);
   U108 : XOR2_X1 port map( A => n226, B => B(33), Z => DIFF_33_port);
   U109 : XOR2_X1 port map( A => n228, B => B(31), Z => DIFF_31_port);
   U110 : XOR2_X1 port map( A => n231, B => B(30), Z => DIFF_30_port);
   U111 : XOR2_X1 port map( A => n230, B => B(29), Z => DIFF_29_port);
   U112 : XOR2_X1 port map( A => n233, B => B(27), Z => DIFF_27_port);
   U114 : XOR2_X1 port map( A => n235, B => B(25), Z => DIFF_25_port);
   U115 : XOR2_X1 port map( A => n237, B => B(23), Z => DIFF_23_port);
   U117 : XOR2_X1 port map( A => n239, B => B(21), Z => DIFF_21_port);
   U118 : XOR2_X1 port map( A => B(1), B => B(0), Z => DIFF_1_port);
   U119 : XOR2_X1 port map( A => n241, B => B(19), Z => DIFF_19_port);
   U121 : XOR2_X1 port map( A => n243, B => B(17), Z => DIFF_17_port);
   U122 : XOR2_X1 port map( A => n245, B => B(15), Z => DIFF_15_port);
   U124 : XOR2_X1 port map( A => n247, B => B(13), Z => DIFF_13_port);
   U125 : XOR2_X1 port map( A => n249, B => B(11), Z => DIFF_11_port);
   U1 : NAND2_X1 port map( A1 => n197, A2 => n251, ZN => n196);
   U2 : NOR3_X1 port map( A1 => B(59), A2 => B(60), A3 => n198, ZN => n197);
   U3 : NOR2_X1 port map( A1 => B(59), A2 => n198, ZN => n199);
   U4 : NOR2_X1 port map( A1 => B(55), A2 => n202, ZN => n203);
   U5 : NOR2_X1 port map( A1 => B(51), A2 => n206, ZN => n207);
   U6 : NOR2_X1 port map( A1 => B(47), A2 => n212, ZN => n213);
   U7 : NOR2_X1 port map( A1 => B(43), A2 => n216, ZN => n217);
   U8 : NOR2_X1 port map( A1 => B(39), A2 => n220, ZN => n221);
   U9 : OR3_X1 port map( A1 => B(57), A2 => B(58), A3 => n200, ZN => n198);
   U10 : OR3_X1 port map( A1 => B(53), A2 => B(54), A3 => n204, ZN => n202);
   U11 : OR3_X1 port map( A1 => B(49), A2 => B(50), A3 => n208, ZN => n206);
   U12 : OR3_X1 port map( A1 => B(45), A2 => B(46), A3 => n214, ZN => n212);
   U13 : OR3_X1 port map( A1 => B(41), A2 => B(42), A3 => n218, ZN => n216);
   U14 : OR3_X1 port map( A1 => B(55), A2 => B(56), A3 => n202, ZN => n200);
   U15 : OR3_X1 port map( A1 => B(51), A2 => B(52), A3 => n206, ZN => n204);
   U16 : OR3_X1 port map( A1 => B(47), A2 => B(48), A3 => n212, ZN => n208);
   U17 : OR3_X1 port map( A1 => B(43), A2 => B(44), A3 => n216, ZN => n214);
   U18 : OR3_X1 port map( A1 => B(39), A2 => B(40), A3 => n220, ZN => n218);
   U19 : OR2_X1 port map( A1 => n204, A2 => B(53), ZN => n205);
   U20 : OR2_X1 port map( A1 => n208, A2 => B(49), ZN => n209);
   U21 : OR2_X1 port map( A1 => n214, A2 => B(45), ZN => n215);
   U22 : OR2_X1 port map( A1 => n218, A2 => B(41), ZN => n219);
   U23 : OR2_X1 port map( A1 => n200, A2 => B(57), ZN => n201);
   U24 : OR2_X1 port map( A1 => n222, A2 => B(37), ZN => n223);
   U25 : OR3_X1 port map( A1 => B(37), A2 => B(38), A3 => n222, ZN => n220);
   U26 : OR2_X1 port map( A1 => n196, A2 => B(62), ZN => n195);
   U27 : NOR2_X1 port map( A1 => B(35), A2 => n224, ZN => n225);
   U28 : OR3_X1 port map( A1 => B(35), A2 => B(36), A3 => n224, ZN => n222);
   U29 : XNOR2_X1 port map( A => B(40), B => n221, ZN => DIFF_40_port);
   U30 : XNOR2_X1 port map( A => B(36), B => n225, ZN => DIFF_36_port);
   U31 : OR3_X1 port map( A1 => B(33), A2 => B(34), A3 => n226, ZN => n224);
   U32 : XNOR2_X1 port map( A => B(32), B => n229, ZN => DIFF_32_port);
   U33 : OR2_X1 port map( A1 => n226, A2 => B(33), ZN => n227);
   U34 : XNOR2_X1 port map( A => n197, B => B(61), ZN => DIFF_61_port);
   U35 : XNOR2_X1 port map( A => B(60), B => n199, ZN => DIFF_60_port);
   U36 : XNOR2_X1 port map( A => B(56), B => n203, ZN => DIFF_56_port);
   U37 : XNOR2_X1 port map( A => B(52), B => n207, ZN => DIFF_52_port);
   U38 : XNOR2_X1 port map( A => B(48), B => n213, ZN => DIFF_48_port);
   U39 : XNOR2_X1 port map( A => B(44), B => n217, ZN => DIFF_44_port);
   U40 : NOR2_X1 port map( A1 => B(31), A2 => n228, ZN => n229);
   U41 : OR3_X1 port map( A1 => B(31), A2 => B(32), A3 => n228, ZN => n226);
   U42 : OR3_X1 port map( A1 => B(29), A2 => B(30), A3 => n230, ZN => n228);
   U43 : OR2_X1 port map( A1 => n230, A2 => B(29), ZN => n231);
   U44 : XNOR2_X1 port map( A => B(28), B => n234, ZN => DIFF_28_port);
   U45 : XNOR2_X1 port map( A => n189, B => B(26), ZN => DIFF_26_port);
   U46 : NOR2_X1 port map( A1 => n235, A2 => B(25), ZN => n189);
   U47 : XNOR2_X1 port map( A => n193, B => B(22), ZN => DIFF_22_port);
   U48 : NOR2_X1 port map( A1 => n239, A2 => B(21), ZN => n193);
   U49 : XNOR2_X1 port map( A => n236, B => B(18), ZN => DIFF_18_port);
   U50 : NOR2_X1 port map( A1 => n243, A2 => B(17), ZN => n236);
   U51 : XNOR2_X1 port map( A => n240, B => B(14), ZN => DIFF_14_port);
   U52 : NOR2_X1 port map( A1 => n247, A2 => B(13), ZN => n240);
   U53 : XNOR2_X1 port map( A => n244, B => B(10), ZN => DIFF_10_port);
   U54 : NOR2_X1 port map( A1 => n190, A2 => B(9), ZN => n244);
   U55 : XNOR2_X1 port map( A => n248, B => B(6), ZN => DIFF_6_port);
   U56 : NOR2_X1 port map( A1 => n194, A2 => B(5), ZN => n248);
   U57 : NOR2_X1 port map( A1 => B(27), A2 => n233, ZN => n234);
   U58 : XNOR2_X1 port map( A => B(24), B => n238, ZN => DIFF_24_port);
   U59 : NOR2_X1 port map( A1 => B(23), A2 => n237, ZN => n238);
   U60 : XNOR2_X1 port map( A => B(20), B => n242, ZN => DIFF_20_port);
   U61 : NOR2_X1 port map( A1 => B(19), A2 => n241, ZN => n242);
   U62 : XNOR2_X1 port map( A => B(16), B => n246, ZN => DIFF_16_port);
   U63 : NOR2_X1 port map( A1 => B(15), A2 => n245, ZN => n246);
   U64 : XNOR2_X1 port map( A => B(12), B => n250, ZN => DIFF_12_port);
   U65 : NOR2_X1 port map( A1 => B(11), A2 => n249, ZN => n250);
   U66 : XNOR2_X1 port map( A => B(8), B => n191, ZN => DIFF_8_port);
   U67 : NOR2_X1 port map( A1 => B(7), A2 => n192, ZN => n191);
   U68 : XNOR2_X1 port map( A => B(2), B => n232, ZN => DIFF_2_port);
   U69 : NOR2_X1 port map( A1 => B(0), A2 => B(1), ZN => n232);
   U70 : XNOR2_X1 port map( A => B(4), B => n210, ZN => DIFF_4_port);
   U71 : NOR2_X1 port map( A1 => B(3), A2 => n211, ZN => n210);
   U72 : OR3_X1 port map( A1 => B(5), A2 => B(6), A3 => n194, ZN => n192);
   U73 : OR3_X1 port map( A1 => B(10), A2 => B(9), A3 => n190, ZN => n249);
   U74 : OR3_X1 port map( A1 => B(13), A2 => B(14), A3 => n247, ZN => n245);
   U75 : OR3_X1 port map( A1 => B(17), A2 => B(18), A3 => n243, ZN => n241);
   U76 : OR3_X1 port map( A1 => B(21), A2 => B(22), A3 => n239, ZN => n237);
   U77 : OR3_X1 port map( A1 => B(25), A2 => B(26), A3 => n235, ZN => n233);
   U78 : OR3_X1 port map( A1 => B(7), A2 => B(8), A3 => n192, ZN => n190);
   U79 : OR3_X1 port map( A1 => B(11), A2 => B(12), A3 => n249, ZN => n247);
   U80 : OR3_X1 port map( A1 => B(15), A2 => B(16), A3 => n245, ZN => n243);
   U83 : OR3_X1 port map( A1 => B(19), A2 => B(20), A3 => n241, ZN => n239);
   U113 : OR3_X1 port map( A1 => B(23), A2 => B(24), A3 => n237, ZN => n235);
   U116 : OR3_X1 port map( A1 => B(27), A2 => B(28), A3 => n233, ZN => n230);
   U120 : OR3_X1 port map( A1 => B(3), A2 => B(4), A3 => n211, ZN => n194);
   U123 : OR3_X1 port map( A1 => B(1), A2 => B(2), A3 => B(0), ZN => n211);
   U126 : INV_X1 port map( A => B(61), ZN => n251);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_4_DW01_sub_0 is

   port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (63 downto 0);  CO : out std_logic);

end complementer_N64_4_DW01_sub_0;

architecture SYN_rpl of complementer_N64_4_DW01_sub_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal DIFF_62_port, DIFF_61_port, DIFF_60_port, DIFF_59_port, DIFF_58_port,
      DIFF_57_port, DIFF_56_port, DIFF_55_port, DIFF_54_port, DIFF_53_port, 
      DIFF_52_port, DIFF_51_port, DIFF_50_port, DIFF_49_port, DIFF_48_port, 
      DIFF_47_port, DIFF_46_port, DIFF_45_port, DIFF_44_port, DIFF_43_port, 
      DIFF_42_port, DIFF_41_port, DIFF_40_port, DIFF_39_port, DIFF_38_port, 
      DIFF_37_port, DIFF_36_port, DIFF_35_port, DIFF_34_port, DIFF_33_port, 
      DIFF_32_port, DIFF_31_port, DIFF_30_port, DIFF_29_port, DIFF_28_port, 
      DIFF_27_port, DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, 
      DIFF_22_port, DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, 
      DIFF_17_port, DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, 
      DIFF_12_port, DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, 
      DIFF_7_port, DIFF_6_port, DIFF_5_port, DIFF_4_port, DIFF_3_port, 
      DIFF_2_port, DIFF_1_port, DIFF_63_port, n190, n191, n192, n193, n194, 
      n196, n197, n198, n199, n200, n202, n203, n204, n206, n207, n208, n210, 
      n211, n212, n213, n214, n216, n217, n218, n220, n221, n222, n224, n225, 
      n226, n228, n229, n230, n232, n233, n234, n235, n236, n237, n238, n239, 
      n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, 
      n189, n195, n201, n205, n209, n215, n219, n223, n227, n231 : std_logic;

begin
   DIFF <= ( DIFF_63_port, DIFF_62_port, DIFF_61_port, DIFF_60_port, 
      DIFF_59_port, DIFF_58_port, DIFF_57_port, DIFF_56_port, DIFF_55_port, 
      DIFF_54_port, DIFF_53_port, DIFF_52_port, DIFF_51_port, DIFF_50_port, 
      DIFF_49_port, DIFF_48_port, DIFF_47_port, DIFF_46_port, DIFF_45_port, 
      DIFF_44_port, DIFF_43_port, DIFF_42_port, DIFF_41_port, DIFF_40_port, 
      DIFF_39_port, DIFF_38_port, DIFF_37_port, DIFF_36_port, DIFF_35_port, 
      DIFF_34_port, DIFF_33_port, DIFF_32_port, DIFF_31_port, DIFF_30_port, 
      DIFF_29_port, DIFF_28_port, DIFF_27_port, DIFF_26_port, DIFF_25_port, 
      DIFF_24_port, DIFF_23_port, DIFF_22_port, DIFF_21_port, DIFF_20_port, 
      DIFF_19_port, DIFF_18_port, DIFF_17_port, DIFF_16_port, DIFF_15_port, 
      DIFF_14_port, DIFF_13_port, DIFF_12_port, DIFF_11_port, DIFF_10_port, 
      DIFF_9_port, DIFF_8_port, DIFF_7_port, DIFF_6_port, DIFF_5_port, 
      DIFF_4_port, DIFF_3_port, DIFF_2_port, DIFF_1_port, B(0) );
   
   U81 : XOR2_X1 port map( A => n190, B => B(9), Z => DIFF_9_port);
   U82 : XOR2_X1 port map( A => n192, B => B(7), Z => DIFF_7_port);
   U83 : XOR2_X1 port map( A => n193, B => B(6), Z => DIFF_6_port);
   U85 : XOR2_X1 port map( A => n196, B => B(62), Z => DIFF_62_port);
   U86 : XOR2_X1 port map( A => n194, B => B(5), Z => DIFF_5_port);
   U87 : XOR2_X1 port map( A => n198, B => B(59), Z => DIFF_59_port);
   U89 : XOR2_X1 port map( A => n200, B => B(57), Z => DIFF_57_port);
   U90 : XOR2_X1 port map( A => n202, B => B(55), Z => DIFF_55_port);
   U92 : XOR2_X1 port map( A => n204, B => B(53), Z => DIFF_53_port);
   U93 : XOR2_X1 port map( A => n206, B => B(51), Z => DIFF_51_port);
   U95 : XOR2_X1 port map( A => n208, B => B(49), Z => DIFF_49_port);
   U96 : XOR2_X1 port map( A => n212, B => B(47), Z => DIFF_47_port);
   U98 : XOR2_X1 port map( A => n214, B => B(45), Z => DIFF_45_port);
   U99 : XOR2_X1 port map( A => n216, B => B(43), Z => DIFF_43_port);
   U101 : XOR2_X1 port map( A => n218, B => B(41), Z => DIFF_41_port);
   U102 : XOR2_X1 port map( A => n211, B => B(3), Z => DIFF_3_port);
   U103 : XOR2_X1 port map( A => n220, B => B(39), Z => DIFF_39_port);
   U105 : XOR2_X1 port map( A => n222, B => B(37), Z => DIFF_37_port);
   U106 : XOR2_X1 port map( A => n224, B => B(35), Z => DIFF_35_port);
   U108 : XOR2_X1 port map( A => n226, B => B(33), Z => DIFF_33_port);
   U109 : XOR2_X1 port map( A => n228, B => B(31), Z => DIFF_31_port);
   U111 : XOR2_X1 port map( A => n230, B => B(29), Z => DIFF_29_port);
   U112 : XOR2_X1 port map( A => n233, B => B(27), Z => DIFF_27_port);
   U113 : XOR2_X1 port map( A => n236, B => B(26), Z => DIFF_26_port);
   U114 : XOR2_X1 port map( A => n235, B => B(25), Z => DIFF_25_port);
   U115 : XOR2_X1 port map( A => n237, B => B(23), Z => DIFF_23_port);
   U116 : XOR2_X1 port map( A => n240, B => B(22), Z => DIFF_22_port);
   U117 : XOR2_X1 port map( A => n239, B => B(21), Z => DIFF_21_port);
   U118 : XOR2_X1 port map( A => B(1), B => B(0), Z => DIFF_1_port);
   U119 : XOR2_X1 port map( A => n241, B => B(19), Z => DIFF_19_port);
   U120 : XOR2_X1 port map( A => n244, B => B(18), Z => DIFF_18_port);
   U121 : XOR2_X1 port map( A => n243, B => B(17), Z => DIFF_17_port);
   U122 : XOR2_X1 port map( A => n245, B => B(15), Z => DIFF_15_port);
   U123 : XOR2_X1 port map( A => n248, B => B(14), Z => DIFF_14_port);
   U124 : XOR2_X1 port map( A => n247, B => B(13), Z => DIFF_13_port);
   U125 : XOR2_X1 port map( A => n249, B => B(11), Z => DIFF_11_port);
   U126 : XOR2_X1 port map( A => n251, B => B(10), Z => DIFF_10_port);
   U1 : XNOR2_X1 port map( A => B(40), B => n221, ZN => DIFF_40_port);
   U2 : NOR2_X1 port map( A1 => B(39), A2 => n220, ZN => n221);
   U3 : OR3_X1 port map( A1 => B(39), A2 => B(40), A3 => n220, ZN => n218);
   U4 : NOR3_X1 port map( A1 => B(59), A2 => B(60), A3 => n198, ZN => n197);
   U5 : XNOR2_X1 port map( A => n189, B => B(58), ZN => DIFF_58_port);
   U6 : NOR2_X1 port map( A1 => n200, A2 => B(57), ZN => n189);
   U7 : XNOR2_X1 port map( A => n195, B => B(54), ZN => DIFF_54_port);
   U8 : NOR2_X1 port map( A1 => n204, A2 => B(53), ZN => n195);
   U9 : XNOR2_X1 port map( A => n201, B => B(50), ZN => DIFF_50_port);
   U10 : NOR2_X1 port map( A1 => n208, A2 => B(49), ZN => n201);
   U11 : XNOR2_X1 port map( A => n205, B => B(46), ZN => DIFF_46_port);
   U12 : NOR2_X1 port map( A1 => n214, A2 => B(45), ZN => n205);
   U13 : XNOR2_X1 port map( A => n209, B => B(42), ZN => DIFF_42_port);
   U14 : NOR2_X1 port map( A1 => n218, A2 => B(41), ZN => n209);
   U15 : XNOR2_X1 port map( A => B(52), B => n207, ZN => DIFF_52_port);
   U16 : NOR2_X1 port map( A1 => B(51), A2 => n206, ZN => n207);
   U17 : XNOR2_X1 port map( A => B(48), B => n213, ZN => DIFF_48_port);
   U18 : NOR2_X1 port map( A1 => B(47), A2 => n212, ZN => n213);
   U19 : XNOR2_X1 port map( A => B(44), B => n217, ZN => DIFF_44_port);
   U20 : NOR2_X1 port map( A1 => B(43), A2 => n216, ZN => n217);
   U21 : XNOR2_X1 port map( A => B(56), B => n203, ZN => DIFF_56_port);
   U22 : NOR2_X1 port map( A1 => B(55), A2 => n202, ZN => n203);
   U23 : XNOR2_X1 port map( A => B(60), B => n199, ZN => DIFF_60_port);
   U24 : NOR2_X1 port map( A1 => B(59), A2 => n198, ZN => n199);
   U25 : XOR2_X1 port map( A => n197, B => n231, Z => DIFF_61_port);
   U26 : NAND2_X1 port map( A1 => n197, A2 => n231, ZN => n196);
   U27 : OR3_X1 port map( A1 => B(57), A2 => B(58), A3 => n200, ZN => n198);
   U28 : OR3_X1 port map( A1 => B(41), A2 => B(42), A3 => n218, ZN => n216);
   U29 : OR3_X1 port map( A1 => B(45), A2 => B(46), A3 => n214, ZN => n212);
   U30 : OR3_X1 port map( A1 => B(49), A2 => B(50), A3 => n208, ZN => n206);
   U31 : OR3_X1 port map( A1 => B(53), A2 => B(54), A3 => n204, ZN => n202);
   U32 : OR3_X1 port map( A1 => B(43), A2 => B(44), A3 => n216, ZN => n214);
   U33 : OR3_X1 port map( A1 => B(47), A2 => B(48), A3 => n212, ZN => n208);
   U34 : OR3_X1 port map( A1 => B(51), A2 => B(52), A3 => n206, ZN => n204);
   U35 : OR3_X1 port map( A1 => B(55), A2 => B(56), A3 => n202, ZN => n200);
   U36 : XNOR2_X1 port map( A => n215, B => B(38), ZN => DIFF_38_port);
   U37 : NOR2_X1 port map( A1 => n222, A2 => B(37), ZN => n215);
   U38 : OR3_X1 port map( A1 => B(37), A2 => B(38), A3 => n222, ZN => n220);
   U39 : XNOR2_X1 port map( A => n219, B => B(63), ZN => DIFF_63_port);
   U40 : NOR2_X1 port map( A1 => n196, A2 => B(62), ZN => n219);
   U41 : XNOR2_X1 port map( A => B(36), B => n225, ZN => DIFF_36_port);
   U42 : NOR2_X1 port map( A1 => B(35), A2 => n224, ZN => n225);
   U43 : OR3_X1 port map( A1 => B(35), A2 => B(36), A3 => n224, ZN => n222);
   U44 : OR3_X1 port map( A1 => B(33), A2 => B(34), A3 => n226, ZN => n224);
   U45 : XNOR2_X1 port map( A => n223, B => B(34), ZN => DIFF_34_port);
   U46 : NOR2_X1 port map( A1 => n226, A2 => B(33), ZN => n223);
   U47 : XNOR2_X1 port map( A => B(32), B => n229, ZN => DIFF_32_port);
   U48 : NOR2_X1 port map( A1 => B(31), A2 => n228, ZN => n229);
   U49 : OR3_X1 port map( A1 => B(31), A2 => B(32), A3 => n228, ZN => n226);
   U50 : OR3_X1 port map( A1 => B(29), A2 => B(30), A3 => n230, ZN => n228);
   U51 : XNOR2_X1 port map( A => n227, B => B(30), ZN => DIFF_30_port);
   U52 : NOR2_X1 port map( A1 => n230, A2 => B(29), ZN => n227);
   U53 : OR3_X1 port map( A1 => B(27), A2 => B(28), A3 => n233, ZN => n230);
   U54 : XNOR2_X1 port map( A => B(28), B => n234, ZN => DIFF_28_port);
   U55 : NOR2_X1 port map( A1 => B(27), A2 => n233, ZN => n234);
   U56 : NOR2_X1 port map( A1 => B(23), A2 => n237, ZN => n238);
   U57 : NOR2_X1 port map( A1 => B(19), A2 => n241, ZN => n242);
   U58 : NOR2_X1 port map( A1 => B(15), A2 => n245, ZN => n246);
   U59 : NOR2_X1 port map( A1 => B(11), A2 => n249, ZN => n250);
   U60 : NOR2_X1 port map( A1 => B(7), A2 => n192, ZN => n191);
   U61 : NOR2_X1 port map( A1 => B(3), A2 => n211, ZN => n210);
   U62 : OR3_X1 port map( A1 => B(25), A2 => B(26), A3 => n235, ZN => n233);
   U63 : OR3_X1 port map( A1 => B(21), A2 => B(22), A3 => n239, ZN => n237);
   U64 : OR3_X1 port map( A1 => B(17), A2 => B(18), A3 => n243, ZN => n241);
   U65 : OR3_X1 port map( A1 => B(13), A2 => B(14), A3 => n247, ZN => n245);
   U66 : OR3_X1 port map( A1 => B(10), A2 => B(9), A3 => n190, ZN => n249);
   U67 : OR3_X1 port map( A1 => B(5), A2 => B(6), A3 => n194, ZN => n192);
   U68 : OR3_X1 port map( A1 => B(23), A2 => B(24), A3 => n237, ZN => n235);
   U69 : OR3_X1 port map( A1 => B(19), A2 => B(20), A3 => n241, ZN => n239);
   U70 : OR3_X1 port map( A1 => B(15), A2 => B(16), A3 => n245, ZN => n243);
   U71 : OR3_X1 port map( A1 => B(11), A2 => B(12), A3 => n249, ZN => n247);
   U72 : OR3_X1 port map( A1 => B(7), A2 => B(8), A3 => n192, ZN => n190);
   U73 : OR3_X1 port map( A1 => B(3), A2 => B(4), A3 => n211, ZN => n194);
   U74 : XNOR2_X1 port map( A => B(24), B => n238, ZN => DIFF_24_port);
   U75 : XNOR2_X1 port map( A => B(20), B => n242, ZN => DIFF_20_port);
   U76 : XNOR2_X1 port map( A => B(16), B => n246, ZN => DIFF_16_port);
   U77 : XNOR2_X1 port map( A => B(12), B => n250, ZN => DIFF_12_port);
   U78 : XNOR2_X1 port map( A => B(8), B => n191, ZN => DIFF_8_port);
   U79 : XNOR2_X1 port map( A => B(4), B => n210, ZN => DIFF_4_port);
   U80 : XNOR2_X1 port map( A => B(2), B => n232, ZN => DIFF_2_port);
   U84 : OR2_X1 port map( A1 => n235, A2 => B(25), ZN => n236);
   U88 : OR2_X1 port map( A1 => n239, A2 => B(21), ZN => n240);
   U91 : OR2_X1 port map( A1 => n243, A2 => B(17), ZN => n244);
   U94 : OR2_X1 port map( A1 => n247, A2 => B(13), ZN => n248);
   U97 : OR2_X1 port map( A1 => n190, A2 => B(9), ZN => n251);
   U100 : OR2_X1 port map( A1 => n194, A2 => B(5), ZN => n193);
   U104 : OR3_X1 port map( A1 => B(1), A2 => B(2), A3 => B(0), ZN => n211);
   U107 : NOR2_X1 port map( A1 => B(0), A2 => B(1), ZN => n232);
   U110 : INV_X1 port map( A => B(61), ZN => n231);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_5_DW01_sub_0 is

   port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (63 downto 0);  CO : out std_logic);

end complementer_N64_5_DW01_sub_0;

architecture SYN_rpl of complementer_N64_5_DW01_sub_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal DIFF_62_port, DIFF_63_port, DIFF_27_port, DIFF_28_port, DIFF_29_port,
      DIFF_30_port, DIFF_31_port, DIFF_32_port, DIFF_33_port, DIFF_34_port, 
      DIFF_35_port, DIFF_36_port, DIFF_37_port, DIFF_38_port, DIFF_39_port, 
      DIFF_40_port, DIFF_41_port, DIFF_42_port, DIFF_43_port, DIFF_44_port, 
      DIFF_45_port, DIFF_46_port, DIFF_47_port, DIFF_48_port, DIFF_49_port, 
      DIFF_50_port, DIFF_51_port, DIFF_52_port, DIFF_53_port, DIFF_54_port, 
      DIFF_55_port, DIFF_56_port, DIFF_57_port, DIFF_58_port, DIFF_59_port, 
      DIFF_60_port, DIFF_61_port, DIFF_3_port, DIFF_4_port, DIFF_5_port, 
      DIFF_6_port, DIFF_7_port, DIFF_8_port, DIFF_9_port, DIFF_10_port, 
      DIFF_11_port, DIFF_12_port, DIFF_13_port, DIFF_14_port, DIFF_15_port, 
      DIFF_16_port, DIFF_17_port, DIFF_18_port, DIFF_19_port, DIFF_20_port, 
      DIFF_21_port, DIFF_22_port, DIFF_23_port, DIFF_24_port, DIFF_25_port, 
      DIFF_26_port, DIFF_2_port, DIFF_1_port, n190, n191, n192, n194, n196, 
      n197, n198, n199, n200, n202, n203, n204, n206, n207, n208, n210, n211, 
      n212, n213, n214, n216, n217, n218, n220, n221, n222, n224, n225, n226, 
      n228, n229, n230, n232, n233, n234, n235, n236, n237, n238, n239, n241, 
      n242, n243, n245, n246, n247, n249, n250, n189, n193, n195, n201, n205, 
      n209, n215, n219, n223, n227, n231, n240, n244, n248, n251 : std_logic;

begin
   DIFF <= ( DIFF_63_port, DIFF_62_port, DIFF_61_port, DIFF_60_port, 
      DIFF_59_port, DIFF_58_port, DIFF_57_port, DIFF_56_port, DIFF_55_port, 
      DIFF_54_port, DIFF_53_port, DIFF_52_port, DIFF_51_port, DIFF_50_port, 
      DIFF_49_port, DIFF_48_port, DIFF_47_port, DIFF_46_port, DIFF_45_port, 
      DIFF_44_port, DIFF_43_port, DIFF_42_port, DIFF_41_port, DIFF_40_port, 
      DIFF_39_port, DIFF_38_port, DIFF_37_port, DIFF_36_port, DIFF_35_port, 
      DIFF_34_port, DIFF_33_port, DIFF_32_port, DIFF_31_port, DIFF_30_port, 
      DIFF_29_port, DIFF_28_port, DIFF_27_port, DIFF_26_port, DIFF_25_port, 
      DIFF_24_port, DIFF_23_port, DIFF_22_port, DIFF_21_port, DIFF_20_port, 
      DIFF_19_port, DIFF_18_port, DIFF_17_port, DIFF_16_port, DIFF_15_port, 
      DIFF_14_port, DIFF_13_port, DIFF_12_port, DIFF_11_port, DIFF_10_port, 
      DIFF_9_port, DIFF_8_port, DIFF_7_port, DIFF_6_port, DIFF_5_port, 
      DIFF_4_port, DIFF_3_port, DIFF_2_port, DIFF_1_port, B(0) );
   
   U81 : XOR2_X1 port map( A => n190, B => B(9), Z => DIFF_9_port);
   U82 : XOR2_X1 port map( A => n192, B => B(7), Z => DIFF_7_port);
   U85 : XOR2_X1 port map( A => n196, B => B(62), Z => DIFF_62_port);
   U86 : XOR2_X1 port map( A => n194, B => B(5), Z => DIFF_5_port);
   U87 : XOR2_X1 port map( A => n198, B => B(59), Z => DIFF_59_port);
   U89 : XOR2_X1 port map( A => n200, B => B(57), Z => DIFF_57_port);
   U90 : XOR2_X1 port map( A => n202, B => B(55), Z => DIFF_55_port);
   U92 : XOR2_X1 port map( A => n204, B => B(53), Z => DIFF_53_port);
   U93 : XOR2_X1 port map( A => n206, B => B(51), Z => DIFF_51_port);
   U95 : XOR2_X1 port map( A => n208, B => B(49), Z => DIFF_49_port);
   U96 : XOR2_X1 port map( A => n212, B => B(47), Z => DIFF_47_port);
   U98 : XOR2_X1 port map( A => n214, B => B(45), Z => DIFF_45_port);
   U99 : XOR2_X1 port map( A => n216, B => B(43), Z => DIFF_43_port);
   U101 : XOR2_X1 port map( A => n218, B => B(41), Z => DIFF_41_port);
   U102 : XOR2_X1 port map( A => n211, B => B(3), Z => DIFF_3_port);
   U103 : XOR2_X1 port map( A => n220, B => B(39), Z => DIFF_39_port);
   U105 : XOR2_X1 port map( A => n222, B => B(37), Z => DIFF_37_port);
   U106 : XOR2_X1 port map( A => n224, B => B(35), Z => DIFF_35_port);
   U108 : XOR2_X1 port map( A => n226, B => B(33), Z => DIFF_33_port);
   U109 : XOR2_X1 port map( A => n228, B => B(31), Z => DIFF_31_port);
   U111 : XOR2_X1 port map( A => n230, B => B(29), Z => DIFF_29_port);
   U112 : XOR2_X1 port map( A => n233, B => B(27), Z => DIFF_27_port);
   U113 : XOR2_X1 port map( A => n236, B => B(26), Z => DIFF_26_port);
   U114 : XOR2_X1 port map( A => n235, B => B(25), Z => DIFF_25_port);
   U115 : XOR2_X1 port map( A => n237, B => B(23), Z => DIFF_23_port);
   U117 : XOR2_X1 port map( A => n239, B => B(21), Z => DIFF_21_port);
   U118 : XOR2_X1 port map( A => B(1), B => B(0), Z => DIFF_1_port);
   U119 : XOR2_X1 port map( A => n241, B => B(19), Z => DIFF_19_port);
   U121 : XOR2_X1 port map( A => n243, B => B(17), Z => DIFF_17_port);
   U122 : XOR2_X1 port map( A => n245, B => B(15), Z => DIFF_15_port);
   U124 : XOR2_X1 port map( A => n247, B => B(13), Z => DIFF_13_port);
   U125 : XOR2_X1 port map( A => n249, B => B(11), Z => DIFF_11_port);
   U1 : XNOR2_X1 port map( A => n189, B => B(42), ZN => DIFF_42_port);
   U2 : NOR2_X1 port map( A1 => n218, A2 => B(41), ZN => n189);
   U3 : XNOR2_X1 port map( A => n193, B => B(38), ZN => DIFF_38_port);
   U4 : NOR2_X1 port map( A1 => n222, A2 => B(37), ZN => n193);
   U5 : XNOR2_X1 port map( A => B(44), B => n217, ZN => DIFF_44_port);
   U6 : NOR2_X1 port map( A1 => B(43), A2 => n216, ZN => n217);
   U7 : XNOR2_X1 port map( A => B(40), B => n221, ZN => DIFF_40_port);
   U8 : NOR2_X1 port map( A1 => B(39), A2 => n220, ZN => n221);
   U9 : OR3_X1 port map( A1 => B(37), A2 => B(38), A3 => n222, ZN => n220);
   U10 : OR3_X1 port map( A1 => B(41), A2 => B(42), A3 => n218, ZN => n216);
   U11 : OR3_X1 port map( A1 => B(39), A2 => B(40), A3 => n220, ZN => n218);
   U12 : OR3_X1 port map( A1 => B(43), A2 => B(44), A3 => n216, ZN => n214);
   U13 : XNOR2_X1 port map( A => n195, B => B(58), ZN => DIFF_58_port);
   U14 : NOR2_X1 port map( A1 => n200, A2 => B(57), ZN => n195);
   U15 : XNOR2_X1 port map( A => n201, B => B(54), ZN => DIFF_54_port);
   U16 : NOR2_X1 port map( A1 => n204, A2 => B(53), ZN => n201);
   U17 : XNOR2_X1 port map( A => n205, B => B(50), ZN => DIFF_50_port);
   U18 : NOR2_X1 port map( A1 => n208, A2 => B(49), ZN => n205);
   U19 : XNOR2_X1 port map( A => n209, B => B(46), ZN => DIFF_46_port);
   U20 : NOR2_X1 port map( A1 => n214, A2 => B(45), ZN => n209);
   U21 : XNOR2_X1 port map( A => B(56), B => n203, ZN => DIFF_56_port);
   U22 : NOR2_X1 port map( A1 => B(55), A2 => n202, ZN => n203);
   U23 : XNOR2_X1 port map( A => B(52), B => n207, ZN => DIFF_52_port);
   U24 : NOR2_X1 port map( A1 => B(51), A2 => n206, ZN => n207);
   U25 : XNOR2_X1 port map( A => B(48), B => n213, ZN => DIFF_48_port);
   U26 : NOR2_X1 port map( A1 => B(47), A2 => n212, ZN => n213);
   U27 : XOR2_X1 port map( A => n197, B => n251, Z => DIFF_61_port);
   U28 : NAND2_X1 port map( A1 => n197, A2 => n251, ZN => n196);
   U29 : OR3_X1 port map( A1 => B(57), A2 => B(58), A3 => n200, ZN => n198);
   U30 : OR3_X1 port map( A1 => B(45), A2 => B(46), A3 => n214, ZN => n212);
   U31 : OR3_X1 port map( A1 => B(49), A2 => B(50), A3 => n208, ZN => n206);
   U32 : OR3_X1 port map( A1 => B(53), A2 => B(54), A3 => n204, ZN => n202);
   U33 : OR3_X1 port map( A1 => B(47), A2 => B(48), A3 => n212, ZN => n208);
   U34 : OR3_X1 port map( A1 => B(51), A2 => B(52), A3 => n206, ZN => n204);
   U35 : OR3_X1 port map( A1 => B(55), A2 => B(56), A3 => n202, ZN => n200);
   U36 : XNOR2_X1 port map( A => B(36), B => n225, ZN => DIFF_36_port);
   U37 : NOR2_X1 port map( A1 => B(35), A2 => n224, ZN => n225);
   U38 : OR3_X1 port map( A1 => B(35), A2 => B(36), A3 => n224, ZN => n222);
   U39 : NOR3_X1 port map( A1 => B(59), A2 => B(60), A3 => n198, ZN => n197);
   U40 : XNOR2_X1 port map( A => n215, B => B(63), ZN => DIFF_63_port);
   U41 : NOR2_X1 port map( A1 => n196, A2 => B(62), ZN => n215);
   U42 : XNOR2_X1 port map( A => B(60), B => n199, ZN => DIFF_60_port);
   U43 : NOR2_X1 port map( A1 => B(59), A2 => n198, ZN => n199);
   U44 : OR3_X1 port map( A1 => B(33), A2 => B(34), A3 => n226, ZN => n224);
   U45 : XNOR2_X1 port map( A => n219, B => B(34), ZN => DIFF_34_port);
   U46 : NOR2_X1 port map( A1 => n226, A2 => B(33), ZN => n219);
   U47 : XNOR2_X1 port map( A => B(32), B => n229, ZN => DIFF_32_port);
   U48 : NOR2_X1 port map( A1 => B(31), A2 => n228, ZN => n229);
   U49 : OR3_X1 port map( A1 => B(31), A2 => B(32), A3 => n228, ZN => n226);
   U50 : OR3_X1 port map( A1 => B(29), A2 => B(30), A3 => n230, ZN => n228);
   U51 : XNOR2_X1 port map( A => n223, B => B(30), ZN => DIFF_30_port);
   U52 : NOR2_X1 port map( A1 => n230, A2 => B(29), ZN => n223);
   U53 : XNOR2_X1 port map( A => B(28), B => n234, ZN => DIFF_28_port);
   U54 : NOR2_X1 port map( A1 => B(27), A2 => n233, ZN => n234);
   U55 : OR3_X1 port map( A1 => B(27), A2 => B(28), A3 => n233, ZN => n230);
   U56 : XNOR2_X1 port map( A => n227, B => B(22), ZN => DIFF_22_port);
   U57 : NOR2_X1 port map( A1 => n239, A2 => B(21), ZN => n227);
   U58 : XNOR2_X1 port map( A => n231, B => B(18), ZN => DIFF_18_port);
   U59 : NOR2_X1 port map( A1 => n243, A2 => B(17), ZN => n231);
   U60 : XNOR2_X1 port map( A => n240, B => B(14), ZN => DIFF_14_port);
   U61 : NOR2_X1 port map( A1 => n247, A2 => B(13), ZN => n240);
   U62 : XNOR2_X1 port map( A => n244, B => B(10), ZN => DIFF_10_port);
   U63 : NOR2_X1 port map( A1 => n190, A2 => B(9), ZN => n244);
   U64 : XNOR2_X1 port map( A => n248, B => B(6), ZN => DIFF_6_port);
   U65 : NOR2_X1 port map( A1 => n194, A2 => B(5), ZN => n248);
   U66 : XNOR2_X1 port map( A => B(24), B => n238, ZN => DIFF_24_port);
   U67 : NOR2_X1 port map( A1 => B(23), A2 => n237, ZN => n238);
   U68 : XNOR2_X1 port map( A => B(20), B => n242, ZN => DIFF_20_port);
   U69 : NOR2_X1 port map( A1 => B(19), A2 => n241, ZN => n242);
   U70 : XNOR2_X1 port map( A => B(16), B => n246, ZN => DIFF_16_port);
   U71 : NOR2_X1 port map( A1 => B(15), A2 => n245, ZN => n246);
   U72 : XNOR2_X1 port map( A => B(12), B => n250, ZN => DIFF_12_port);
   U73 : NOR2_X1 port map( A1 => B(11), A2 => n249, ZN => n250);
   U74 : XNOR2_X1 port map( A => B(8), B => n191, ZN => DIFF_8_port);
   U75 : NOR2_X1 port map( A1 => B(7), A2 => n192, ZN => n191);
   U76 : XNOR2_X1 port map( A => B(2), B => n232, ZN => DIFF_2_port);
   U77 : NOR2_X1 port map( A1 => B(0), A2 => B(1), ZN => n232);
   U78 : XNOR2_X1 port map( A => B(4), B => n210, ZN => DIFF_4_port);
   U79 : NOR2_X1 port map( A1 => B(3), A2 => n211, ZN => n210);
   U80 : OR3_X1 port map( A1 => B(5), A2 => B(6), A3 => n194, ZN => n192);
   U83 : OR3_X1 port map( A1 => B(10), A2 => B(9), A3 => n190, ZN => n249);
   U84 : OR3_X1 port map( A1 => B(13), A2 => B(14), A3 => n247, ZN => n245);
   U88 : OR3_X1 port map( A1 => B(17), A2 => B(18), A3 => n243, ZN => n241);
   U91 : OR3_X1 port map( A1 => B(21), A2 => B(22), A3 => n239, ZN => n237);
   U94 : OR3_X1 port map( A1 => B(25), A2 => B(26), A3 => n235, ZN => n233);
   U97 : OR3_X1 port map( A1 => B(7), A2 => B(8), A3 => n192, ZN => n190);
   U100 : OR3_X1 port map( A1 => B(11), A2 => B(12), A3 => n249, ZN => n247);
   U104 : OR3_X1 port map( A1 => B(15), A2 => B(16), A3 => n245, ZN => n243);
   U107 : OR3_X1 port map( A1 => B(19), A2 => B(20), A3 => n241, ZN => n239);
   U110 : OR3_X1 port map( A1 => B(23), A2 => B(24), A3 => n237, ZN => n235);
   U116 : OR3_X1 port map( A1 => B(3), A2 => B(4), A3 => n211, ZN => n194);
   U120 : OR2_X1 port map( A1 => n235, A2 => B(25), ZN => n236);
   U123 : OR3_X1 port map( A1 => B(1), A2 => B(2), A3 => B(0), ZN => n211);
   U126 : INV_X1 port map( A => B(61), ZN => n251);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_6_DW01_sub_0 is

   port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (63 downto 0);  CO : out std_logic);

end complementer_N64_6_DW01_sub_0;

architecture SYN_rpl of complementer_N64_6_DW01_sub_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal DIFF_62_port, DIFF_61_port, DIFF_60_port, DIFF_59_port, DIFF_58_port,
      DIFF_57_port, DIFF_56_port, DIFF_55_port, DIFF_54_port, DIFF_53_port, 
      DIFF_52_port, DIFF_51_port, DIFF_50_port, DIFF_49_port, DIFF_48_port, 
      DIFF_47_port, DIFF_46_port, DIFF_45_port, DIFF_44_port, DIFF_43_port, 
      DIFF_42_port, DIFF_41_port, DIFF_40_port, DIFF_39_port, DIFF_38_port, 
      DIFF_37_port, DIFF_36_port, DIFF_35_port, DIFF_34_port, DIFF_33_port, 
      DIFF_32_port, DIFF_31_port, DIFF_30_port, DIFF_29_port, DIFF_28_port, 
      DIFF_27_port, DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, 
      DIFF_22_port, DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, 
      DIFF_17_port, DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, 
      DIFF_12_port, DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, 
      DIFF_7_port, DIFF_6_port, DIFF_5_port, DIFF_4_port, DIFF_3_port, 
      DIFF_2_port, DIFF_1_port, DIFF_63_port, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, 
      n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, 
      n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, 
      n231, n232, n233, n234, n235, n237, n238, n239, n240, n241, n242, n243, 
      n244, n245, n246, n247, n248, n249, n250, n251, n189, n236 : std_logic;

begin
   DIFF <= ( DIFF_63_port, DIFF_62_port, DIFF_61_port, DIFF_60_port, 
      DIFF_59_port, DIFF_58_port, DIFF_57_port, DIFF_56_port, DIFF_55_port, 
      DIFF_54_port, DIFF_53_port, DIFF_52_port, DIFF_51_port, DIFF_50_port, 
      DIFF_49_port, DIFF_48_port, DIFF_47_port, DIFF_46_port, DIFF_45_port, 
      DIFF_44_port, DIFF_43_port, DIFF_42_port, DIFF_41_port, DIFF_40_port, 
      DIFF_39_port, DIFF_38_port, DIFF_37_port, DIFF_36_port, DIFF_35_port, 
      DIFF_34_port, DIFF_33_port, DIFF_32_port, DIFF_31_port, DIFF_30_port, 
      DIFF_29_port, DIFF_28_port, DIFF_27_port, DIFF_26_port, DIFF_25_port, 
      DIFF_24_port, DIFF_23_port, DIFF_22_port, DIFF_21_port, DIFF_20_port, 
      DIFF_19_port, DIFF_18_port, DIFF_17_port, DIFF_16_port, DIFF_15_port, 
      DIFF_14_port, DIFF_13_port, DIFF_12_port, DIFF_11_port, DIFF_10_port, 
      DIFF_9_port, DIFF_8_port, DIFF_7_port, DIFF_6_port, DIFF_5_port, 
      DIFF_4_port, DIFF_3_port, DIFF_2_port, DIFF_1_port, B(0) );
   
   U81 : XOR2_X1 port map( A => n190, B => B(9), Z => DIFF_9_port);
   U82 : XOR2_X1 port map( A => n192, B => B(7), Z => DIFF_7_port);
   U83 : XOR2_X1 port map( A => n193, B => B(6), Z => DIFF_6_port);
   U84 : XOR2_X1 port map( A => n195, B => B(63), Z => DIFF_63_port);
   U85 : XOR2_X1 port map( A => n196, B => B(62), Z => DIFF_62_port);
   U86 : XOR2_X1 port map( A => n194, B => B(5), Z => DIFF_5_port);
   U87 : XOR2_X1 port map( A => n198, B => B(59), Z => DIFF_59_port);
   U88 : XOR2_X1 port map( A => n201, B => B(58), Z => DIFF_58_port);
   U89 : XOR2_X1 port map( A => n200, B => B(57), Z => DIFF_57_port);
   U90 : XOR2_X1 port map( A => n202, B => B(55), Z => DIFF_55_port);
   U91 : XOR2_X1 port map( A => n205, B => B(54), Z => DIFF_54_port);
   U92 : XOR2_X1 port map( A => n204, B => B(53), Z => DIFF_53_port);
   U93 : XOR2_X1 port map( A => n206, B => B(51), Z => DIFF_51_port);
   U94 : XOR2_X1 port map( A => n209, B => B(50), Z => DIFF_50_port);
   U95 : XOR2_X1 port map( A => n208, B => B(49), Z => DIFF_49_port);
   U96 : XOR2_X1 port map( A => n212, B => B(47), Z => DIFF_47_port);
   U97 : XOR2_X1 port map( A => n215, B => B(46), Z => DIFF_46_port);
   U98 : XOR2_X1 port map( A => n214, B => B(45), Z => DIFF_45_port);
   U99 : XOR2_X1 port map( A => n216, B => B(43), Z => DIFF_43_port);
   U100 : XOR2_X1 port map( A => n219, B => B(42), Z => DIFF_42_port);
   U101 : XOR2_X1 port map( A => n218, B => B(41), Z => DIFF_41_port);
   U102 : XOR2_X1 port map( A => n211, B => B(3), Z => DIFF_3_port);
   U103 : XOR2_X1 port map( A => n220, B => B(39), Z => DIFF_39_port);
   U104 : XOR2_X1 port map( A => n223, B => B(38), Z => DIFF_38_port);
   U105 : XOR2_X1 port map( A => n222, B => B(37), Z => DIFF_37_port);
   U106 : XOR2_X1 port map( A => n224, B => B(35), Z => DIFF_35_port);
   U107 : XOR2_X1 port map( A => n227, B => B(34), Z => DIFF_34_port);
   U108 : XOR2_X1 port map( A => n226, B => B(33), Z => DIFF_33_port);
   U109 : XOR2_X1 port map( A => n228, B => B(31), Z => DIFF_31_port);
   U110 : XOR2_X1 port map( A => n231, B => B(30), Z => DIFF_30_port);
   U111 : XOR2_X1 port map( A => n230, B => B(29), Z => DIFF_29_port);
   U112 : XOR2_X1 port map( A => n233, B => B(27), Z => DIFF_27_port);
   U114 : XOR2_X1 port map( A => n235, B => B(25), Z => DIFF_25_port);
   U115 : XOR2_X1 port map( A => n237, B => B(23), Z => DIFF_23_port);
   U116 : XOR2_X1 port map( A => n240, B => B(22), Z => DIFF_22_port);
   U117 : XOR2_X1 port map( A => n239, B => B(21), Z => DIFF_21_port);
   U118 : XOR2_X1 port map( A => B(1), B => B(0), Z => DIFF_1_port);
   U119 : XOR2_X1 port map( A => n241, B => B(19), Z => DIFF_19_port);
   U120 : XOR2_X1 port map( A => n244, B => B(18), Z => DIFF_18_port);
   U121 : XOR2_X1 port map( A => n243, B => B(17), Z => DIFF_17_port);
   U122 : XOR2_X1 port map( A => n245, B => B(15), Z => DIFF_15_port);
   U123 : XOR2_X1 port map( A => n248, B => B(14), Z => DIFF_14_port);
   U124 : XOR2_X1 port map( A => n247, B => B(13), Z => DIFF_13_port);
   U125 : XOR2_X1 port map( A => n249, B => B(11), Z => DIFF_11_port);
   U126 : XOR2_X1 port map( A => n251, B => B(10), Z => DIFF_10_port);
   U1 : NAND2_X1 port map( A1 => n197, A2 => n236, ZN => n196);
   U2 : OR3_X1 port map( A1 => B(57), A2 => B(58), A3 => n200, ZN => n198);
   U3 : OR2_X1 port map( A1 => n200, A2 => B(57), ZN => n201);
   U4 : NOR2_X1 port map( A1 => B(43), A2 => n216, ZN => n217);
   U5 : NOR2_X1 port map( A1 => B(39), A2 => n220, ZN => n221);
   U6 : NOR2_X1 port map( A1 => B(35), A2 => n224, ZN => n225);
   U7 : OR3_X1 port map( A1 => B(41), A2 => B(42), A3 => n218, ZN => n216);
   U8 : OR3_X1 port map( A1 => B(37), A2 => B(38), A3 => n222, ZN => n220);
   U9 : OR3_X1 port map( A1 => B(43), A2 => B(44), A3 => n216, ZN => n214);
   U10 : OR3_X1 port map( A1 => B(39), A2 => B(40), A3 => n220, ZN => n218);
   U11 : OR3_X1 port map( A1 => B(35), A2 => B(36), A3 => n224, ZN => n222);
   U12 : OR2_X1 port map( A1 => n218, A2 => B(41), ZN => n219);
   U13 : OR2_X1 port map( A1 => n222, A2 => B(37), ZN => n223);
   U14 : NOR3_X1 port map( A1 => B(59), A2 => B(60), A3 => n198, ZN => n197);
   U15 : NOR2_X1 port map( A1 => B(59), A2 => n198, ZN => n199);
   U16 : NOR2_X1 port map( A1 => B(55), A2 => n202, ZN => n203);
   U17 : NOR2_X1 port map( A1 => B(51), A2 => n206, ZN => n207);
   U18 : NOR2_X1 port map( A1 => B(47), A2 => n212, ZN => n213);
   U19 : OR3_X1 port map( A1 => B(53), A2 => B(54), A3 => n204, ZN => n202);
   U20 : OR3_X1 port map( A1 => B(49), A2 => B(50), A3 => n208, ZN => n206);
   U21 : OR3_X1 port map( A1 => B(45), A2 => B(46), A3 => n214, ZN => n212);
   U22 : OR3_X1 port map( A1 => B(55), A2 => B(56), A3 => n202, ZN => n200);
   U23 : OR3_X1 port map( A1 => B(51), A2 => B(52), A3 => n206, ZN => n204);
   U24 : OR3_X1 port map( A1 => B(47), A2 => B(48), A3 => n212, ZN => n208);
   U25 : OR2_X1 port map( A1 => n204, A2 => B(53), ZN => n205);
   U26 : OR2_X1 port map( A1 => n208, A2 => B(49), ZN => n209);
   U27 : OR2_X1 port map( A1 => n214, A2 => B(45), ZN => n215);
   U28 : OR2_X1 port map( A1 => n196, A2 => B(62), ZN => n195);
   U29 : OR3_X1 port map( A1 => B(33), A2 => B(34), A3 => n226, ZN => n224);
   U30 : OR2_X1 port map( A1 => n226, A2 => B(33), ZN => n227);
   U31 : NOR2_X1 port map( A1 => B(31), A2 => n228, ZN => n229);
   U32 : XNOR2_X1 port map( A => B(44), B => n217, ZN => DIFF_44_port);
   U33 : XNOR2_X1 port map( A => B(40), B => n221, ZN => DIFF_40_port);
   U34 : XNOR2_X1 port map( A => B(36), B => n225, ZN => DIFF_36_port);
   U35 : OR3_X1 port map( A1 => B(31), A2 => B(32), A3 => n228, ZN => n226);
   U36 : XNOR2_X1 port map( A => B(32), B => n229, ZN => DIFF_32_port);
   U37 : XNOR2_X1 port map( A => n197, B => B(61), ZN => DIFF_61_port);
   U38 : XNOR2_X1 port map( A => B(60), B => n199, ZN => DIFF_60_port);
   U39 : XNOR2_X1 port map( A => B(56), B => n203, ZN => DIFF_56_port);
   U40 : XNOR2_X1 port map( A => B(52), B => n207, ZN => DIFF_52_port);
   U41 : XNOR2_X1 port map( A => B(48), B => n213, ZN => DIFF_48_port);
   U42 : OR3_X1 port map( A1 => B(29), A2 => B(30), A3 => n230, ZN => n228);
   U43 : XNOR2_X1 port map( A => B(28), B => n234, ZN => DIFF_28_port);
   U44 : OR2_X1 port map( A1 => n230, A2 => B(29), ZN => n231);
   U45 : NOR2_X1 port map( A1 => B(27), A2 => n233, ZN => n234);
   U46 : OR3_X1 port map( A1 => B(27), A2 => B(28), A3 => n233, ZN => n230);
   U47 : XNOR2_X1 port map( A => n189, B => B(26), ZN => DIFF_26_port);
   U48 : NOR2_X1 port map( A1 => n235, A2 => B(25), ZN => n189);
   U49 : OR3_X1 port map( A1 => B(25), A2 => B(26), A3 => n235, ZN => n233);
   U50 : NOR2_X1 port map( A1 => B(23), A2 => n237, ZN => n238);
   U51 : NOR2_X1 port map( A1 => B(19), A2 => n241, ZN => n242);
   U52 : NOR2_X1 port map( A1 => B(15), A2 => n245, ZN => n246);
   U53 : NOR2_X1 port map( A1 => B(11), A2 => n249, ZN => n250);
   U54 : NOR2_X1 port map( A1 => B(7), A2 => n192, ZN => n191);
   U55 : NOR2_X1 port map( A1 => B(3), A2 => n211, ZN => n210);
   U56 : OR3_X1 port map( A1 => B(21), A2 => B(22), A3 => n239, ZN => n237);
   U57 : OR3_X1 port map( A1 => B(17), A2 => B(18), A3 => n243, ZN => n241);
   U58 : OR3_X1 port map( A1 => B(13), A2 => B(14), A3 => n247, ZN => n245);
   U59 : OR3_X1 port map( A1 => B(10), A2 => B(9), A3 => n190, ZN => n249);
   U60 : OR3_X1 port map( A1 => B(5), A2 => B(6), A3 => n194, ZN => n192);
   U61 : OR3_X1 port map( A1 => B(23), A2 => B(24), A3 => n237, ZN => n235);
   U62 : OR3_X1 port map( A1 => B(19), A2 => B(20), A3 => n241, ZN => n239);
   U63 : OR3_X1 port map( A1 => B(15), A2 => B(16), A3 => n245, ZN => n243);
   U64 : OR3_X1 port map( A1 => B(11), A2 => B(12), A3 => n249, ZN => n247);
   U65 : OR3_X1 port map( A1 => B(7), A2 => B(8), A3 => n192, ZN => n190);
   U66 : OR3_X1 port map( A1 => B(3), A2 => B(4), A3 => n211, ZN => n194);
   U67 : XNOR2_X1 port map( A => B(24), B => n238, ZN => DIFF_24_port);
   U68 : XNOR2_X1 port map( A => B(20), B => n242, ZN => DIFF_20_port);
   U69 : XNOR2_X1 port map( A => B(16), B => n246, ZN => DIFF_16_port);
   U70 : XNOR2_X1 port map( A => B(12), B => n250, ZN => DIFF_12_port);
   U71 : XNOR2_X1 port map( A => B(8), B => n191, ZN => DIFF_8_port);
   U72 : XNOR2_X1 port map( A => B(4), B => n210, ZN => DIFF_4_port);
   U73 : XNOR2_X1 port map( A => B(2), B => n232, ZN => DIFF_2_port);
   U74 : OR2_X1 port map( A1 => n239, A2 => B(21), ZN => n240);
   U75 : OR2_X1 port map( A1 => n243, A2 => B(17), ZN => n244);
   U76 : OR2_X1 port map( A1 => n247, A2 => B(13), ZN => n248);
   U77 : OR2_X1 port map( A1 => n190, A2 => B(9), ZN => n251);
   U78 : OR2_X1 port map( A1 => n194, A2 => B(5), ZN => n193);
   U79 : OR3_X1 port map( A1 => B(1), A2 => B(2), A3 => B(0), ZN => n211);
   U80 : NOR2_X1 port map( A1 => B(0), A2 => B(1), ZN => n232);
   U113 : INV_X1 port map( A => B(61), ZN => n236);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_7_DW01_sub_0 is

   port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (63 downto 0);  CO : out std_logic);

end complementer_N64_7_DW01_sub_0;

architecture SYN_rpl of complementer_N64_7_DW01_sub_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal DIFF_62_port, DIFF_63_port, DIFF_25_port, DIFF_26_port, DIFF_27_port,
      DIFF_28_port, DIFF_29_port, DIFF_30_port, DIFF_31_port, DIFF_32_port, 
      DIFF_33_port, DIFF_34_port, DIFF_35_port, DIFF_36_port, DIFF_37_port, 
      DIFF_38_port, DIFF_39_port, DIFF_40_port, DIFF_41_port, DIFF_42_port, 
      DIFF_43_port, DIFF_44_port, DIFF_45_port, DIFF_46_port, DIFF_47_port, 
      DIFF_48_port, DIFF_49_port, DIFF_50_port, DIFF_51_port, DIFF_52_port, 
      DIFF_53_port, DIFF_54_port, DIFF_55_port, DIFF_56_port, DIFF_57_port, 
      DIFF_58_port, DIFF_59_port, DIFF_60_port, DIFF_61_port, DIFF_3_port, 
      DIFF_4_port, DIFF_5_port, DIFF_6_port, DIFF_7_port, DIFF_8_port, 
      DIFF_9_port, DIFF_10_port, DIFF_11_port, DIFF_12_port, DIFF_13_port, 
      DIFF_14_port, DIFF_15_port, DIFF_16_port, DIFF_17_port, DIFF_18_port, 
      DIFF_19_port, DIFF_20_port, DIFF_21_port, DIFF_22_port, DIFF_23_port, 
      DIFF_24_port, DIFF_2_port, DIFF_1_port, n190, n191, n192, n194, n195, 
      n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, 
      n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, 
      n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, 
      n232, n233, n234, n235, n236, n237, n238, n239, n241, n242, n243, n245, 
      n246, n247, n249, n250, n189, n193, n240, n244, n248, n251 : std_logic;

begin
   DIFF <= ( DIFF_63_port, DIFF_62_port, DIFF_61_port, DIFF_60_port, 
      DIFF_59_port, DIFF_58_port, DIFF_57_port, DIFF_56_port, DIFF_55_port, 
      DIFF_54_port, DIFF_53_port, DIFF_52_port, DIFF_51_port, DIFF_50_port, 
      DIFF_49_port, DIFF_48_port, DIFF_47_port, DIFF_46_port, DIFF_45_port, 
      DIFF_44_port, DIFF_43_port, DIFF_42_port, DIFF_41_port, DIFF_40_port, 
      DIFF_39_port, DIFF_38_port, DIFF_37_port, DIFF_36_port, DIFF_35_port, 
      DIFF_34_port, DIFF_33_port, DIFF_32_port, DIFF_31_port, DIFF_30_port, 
      DIFF_29_port, DIFF_28_port, DIFF_27_port, DIFF_26_port, DIFF_25_port, 
      DIFF_24_port, DIFF_23_port, DIFF_22_port, DIFF_21_port, DIFF_20_port, 
      DIFF_19_port, DIFF_18_port, DIFF_17_port, DIFF_16_port, DIFF_15_port, 
      DIFF_14_port, DIFF_13_port, DIFF_12_port, DIFF_11_port, DIFF_10_port, 
      DIFF_9_port, DIFF_8_port, DIFF_7_port, DIFF_6_port, DIFF_5_port, 
      DIFF_4_port, DIFF_3_port, DIFF_2_port, DIFF_1_port, B(0) );
   
   U81 : XOR2_X1 port map( A => n190, B => B(9), Z => DIFF_9_port);
   U82 : XOR2_X1 port map( A => n192, B => B(7), Z => DIFF_7_port);
   U84 : XOR2_X1 port map( A => n195, B => B(63), Z => DIFF_63_port);
   U85 : XOR2_X1 port map( A => n196, B => B(62), Z => DIFF_62_port);
   U86 : XOR2_X1 port map( A => n194, B => B(5), Z => DIFF_5_port);
   U87 : XOR2_X1 port map( A => n198, B => B(59), Z => DIFF_59_port);
   U88 : XOR2_X1 port map( A => n201, B => B(58), Z => DIFF_58_port);
   U89 : XOR2_X1 port map( A => n200, B => B(57), Z => DIFF_57_port);
   U90 : XOR2_X1 port map( A => n202, B => B(55), Z => DIFF_55_port);
   U91 : XOR2_X1 port map( A => n205, B => B(54), Z => DIFF_54_port);
   U92 : XOR2_X1 port map( A => n204, B => B(53), Z => DIFF_53_port);
   U93 : XOR2_X1 port map( A => n206, B => B(51), Z => DIFF_51_port);
   U94 : XOR2_X1 port map( A => n209, B => B(50), Z => DIFF_50_port);
   U95 : XOR2_X1 port map( A => n208, B => B(49), Z => DIFF_49_port);
   U96 : XOR2_X1 port map( A => n212, B => B(47), Z => DIFF_47_port);
   U97 : XOR2_X1 port map( A => n215, B => B(46), Z => DIFF_46_port);
   U98 : XOR2_X1 port map( A => n214, B => B(45), Z => DIFF_45_port);
   U99 : XOR2_X1 port map( A => n216, B => B(43), Z => DIFF_43_port);
   U100 : XOR2_X1 port map( A => n219, B => B(42), Z => DIFF_42_port);
   U101 : XOR2_X1 port map( A => n218, B => B(41), Z => DIFF_41_port);
   U102 : XOR2_X1 port map( A => n211, B => B(3), Z => DIFF_3_port);
   U103 : XOR2_X1 port map( A => n220, B => B(39), Z => DIFF_39_port);
   U104 : XOR2_X1 port map( A => n223, B => B(38), Z => DIFF_38_port);
   U105 : XOR2_X1 port map( A => n222, B => B(37), Z => DIFF_37_port);
   U106 : XOR2_X1 port map( A => n224, B => B(35), Z => DIFF_35_port);
   U107 : XOR2_X1 port map( A => n227, B => B(34), Z => DIFF_34_port);
   U108 : XOR2_X1 port map( A => n226, B => B(33), Z => DIFF_33_port);
   U109 : XOR2_X1 port map( A => n228, B => B(31), Z => DIFF_31_port);
   U110 : XOR2_X1 port map( A => n231, B => B(30), Z => DIFF_30_port);
   U111 : XOR2_X1 port map( A => n230, B => B(29), Z => DIFF_29_port);
   U112 : XOR2_X1 port map( A => n233, B => B(27), Z => DIFF_27_port);
   U113 : XOR2_X1 port map( A => n236, B => B(26), Z => DIFF_26_port);
   U114 : XOR2_X1 port map( A => n235, B => B(25), Z => DIFF_25_port);
   U115 : XOR2_X1 port map( A => n237, B => B(23), Z => DIFF_23_port);
   U117 : XOR2_X1 port map( A => n239, B => B(21), Z => DIFF_21_port);
   U118 : XOR2_X1 port map( A => B(1), B => B(0), Z => DIFF_1_port);
   U119 : XOR2_X1 port map( A => n241, B => B(19), Z => DIFF_19_port);
   U121 : XOR2_X1 port map( A => n243, B => B(17), Z => DIFF_17_port);
   U122 : XOR2_X1 port map( A => n245, B => B(15), Z => DIFF_15_port);
   U124 : XOR2_X1 port map( A => n247, B => B(13), Z => DIFF_13_port);
   U125 : XOR2_X1 port map( A => n249, B => B(11), Z => DIFF_11_port);
   U1 : NAND2_X1 port map( A1 => n197, A2 => n251, ZN => n196);
   U2 : NOR2_X1 port map( A1 => B(47), A2 => n212, ZN => n213);
   U3 : NOR2_X1 port map( A1 => B(43), A2 => n216, ZN => n217);
   U4 : NOR2_X1 port map( A1 => B(39), A2 => n220, ZN => n221);
   U5 : NOR2_X1 port map( A1 => B(35), A2 => n224, ZN => n225);
   U6 : OR3_X1 port map( A1 => B(45), A2 => B(46), A3 => n214, ZN => n212);
   U7 : OR3_X1 port map( A1 => B(41), A2 => B(42), A3 => n218, ZN => n216);
   U8 : OR3_X1 port map( A1 => B(37), A2 => B(38), A3 => n222, ZN => n220);
   U9 : OR3_X1 port map( A1 => B(33), A2 => B(34), A3 => n226, ZN => n224);
   U10 : OR3_X1 port map( A1 => B(47), A2 => B(48), A3 => n212, ZN => n208);
   U11 : OR3_X1 port map( A1 => B(43), A2 => B(44), A3 => n216, ZN => n214);
   U12 : OR3_X1 port map( A1 => B(39), A2 => B(40), A3 => n220, ZN => n218);
   U13 : OR3_X1 port map( A1 => B(35), A2 => B(36), A3 => n224, ZN => n222);
   U14 : OR2_X1 port map( A1 => n214, A2 => B(45), ZN => n215);
   U15 : OR2_X1 port map( A1 => n218, A2 => B(41), ZN => n219);
   U16 : OR2_X1 port map( A1 => n222, A2 => B(37), ZN => n223);
   U17 : OR2_X1 port map( A1 => n226, A2 => B(33), ZN => n227);
   U18 : NOR3_X1 port map( A1 => B(59), A2 => B(60), A3 => n198, ZN => n197);
   U19 : NOR2_X1 port map( A1 => B(55), A2 => n202, ZN => n203);
   U20 : NOR2_X1 port map( A1 => B(51), A2 => n206, ZN => n207);
   U21 : NOR2_X1 port map( A1 => B(59), A2 => n198, ZN => n199);
   U22 : OR3_X1 port map( A1 => B(57), A2 => B(58), A3 => n200, ZN => n198);
   U23 : OR3_X1 port map( A1 => B(53), A2 => B(54), A3 => n204, ZN => n202);
   U24 : OR3_X1 port map( A1 => B(49), A2 => B(50), A3 => n208, ZN => n206);
   U25 : OR3_X1 port map( A1 => B(55), A2 => B(56), A3 => n202, ZN => n200);
   U26 : OR3_X1 port map( A1 => B(51), A2 => B(52), A3 => n206, ZN => n204);
   U27 : OR2_X1 port map( A1 => n196, A2 => B(62), ZN => n195);
   U28 : OR2_X1 port map( A1 => n204, A2 => B(53), ZN => n205);
   U29 : OR2_X1 port map( A1 => n208, A2 => B(49), ZN => n209);
   U30 : OR2_X1 port map( A1 => n200, A2 => B(57), ZN => n201);
   U31 : NOR2_X1 port map( A1 => B(31), A2 => n228, ZN => n229);
   U32 : OR3_X1 port map( A1 => B(31), A2 => B(32), A3 => n228, ZN => n226);
   U33 : XNOR2_X1 port map( A => B(52), B => n207, ZN => DIFF_52_port);
   U34 : XNOR2_X1 port map( A => B(48), B => n213, ZN => DIFF_48_port);
   U35 : XNOR2_X1 port map( A => B(40), B => n221, ZN => DIFF_40_port);
   U36 : OR3_X1 port map( A1 => B(29), A2 => B(30), A3 => n230, ZN => n228);
   U37 : XNOR2_X1 port map( A => B(44), B => n217, ZN => DIFF_44_port);
   U38 : XNOR2_X1 port map( A => B(36), B => n225, ZN => DIFF_36_port);
   U39 : XNOR2_X1 port map( A => B(32), B => n229, ZN => DIFF_32_port);
   U40 : XNOR2_X1 port map( A => B(28), B => n234, ZN => DIFF_28_port);
   U41 : OR2_X1 port map( A1 => n230, A2 => B(29), ZN => n231);
   U42 : XNOR2_X1 port map( A => n197, B => B(61), ZN => DIFF_61_port);
   U43 : XNOR2_X1 port map( A => B(60), B => n199, ZN => DIFF_60_port);
   U44 : XNOR2_X1 port map( A => B(56), B => n203, ZN => DIFF_56_port);
   U45 : NOR2_X1 port map( A1 => B(27), A2 => n233, ZN => n234);
   U46 : OR3_X1 port map( A1 => B(27), A2 => B(28), A3 => n233, ZN => n230);
   U47 : OR3_X1 port map( A1 => B(25), A2 => B(26), A3 => n235, ZN => n233);
   U48 : OR2_X1 port map( A1 => n235, A2 => B(25), ZN => n236);
   U49 : XNOR2_X1 port map( A => B(24), B => n238, ZN => DIFF_24_port);
   U50 : XNOR2_X1 port map( A => n189, B => B(22), ZN => DIFF_22_port);
   U51 : NOR2_X1 port map( A1 => n239, A2 => B(21), ZN => n189);
   U52 : XNOR2_X1 port map( A => n193, B => B(18), ZN => DIFF_18_port);
   U53 : NOR2_X1 port map( A1 => n243, A2 => B(17), ZN => n193);
   U54 : XNOR2_X1 port map( A => n240, B => B(14), ZN => DIFF_14_port);
   U55 : NOR2_X1 port map( A1 => n247, A2 => B(13), ZN => n240);
   U56 : XNOR2_X1 port map( A => n244, B => B(10), ZN => DIFF_10_port);
   U57 : NOR2_X1 port map( A1 => n190, A2 => B(9), ZN => n244);
   U58 : XNOR2_X1 port map( A => n248, B => B(6), ZN => DIFF_6_port);
   U59 : NOR2_X1 port map( A1 => n194, A2 => B(5), ZN => n248);
   U60 : NOR2_X1 port map( A1 => B(23), A2 => n237, ZN => n238);
   U61 : XNOR2_X1 port map( A => B(20), B => n242, ZN => DIFF_20_port);
   U62 : NOR2_X1 port map( A1 => B(19), A2 => n241, ZN => n242);
   U63 : XNOR2_X1 port map( A => B(16), B => n246, ZN => DIFF_16_port);
   U64 : NOR2_X1 port map( A1 => B(15), A2 => n245, ZN => n246);
   U65 : XNOR2_X1 port map( A => B(12), B => n250, ZN => DIFF_12_port);
   U66 : NOR2_X1 port map( A1 => B(11), A2 => n249, ZN => n250);
   U67 : XNOR2_X1 port map( A => B(8), B => n191, ZN => DIFF_8_port);
   U68 : NOR2_X1 port map( A1 => B(7), A2 => n192, ZN => n191);
   U69 : XNOR2_X1 port map( A => B(2), B => n232, ZN => DIFF_2_port);
   U70 : NOR2_X1 port map( A1 => B(0), A2 => B(1), ZN => n232);
   U71 : XNOR2_X1 port map( A => B(4), B => n210, ZN => DIFF_4_port);
   U72 : NOR2_X1 port map( A1 => B(3), A2 => n211, ZN => n210);
   U73 : OR3_X1 port map( A1 => B(5), A2 => B(6), A3 => n194, ZN => n192);
   U74 : OR3_X1 port map( A1 => B(10), A2 => B(9), A3 => n190, ZN => n249);
   U75 : OR3_X1 port map( A1 => B(13), A2 => B(14), A3 => n247, ZN => n245);
   U76 : OR3_X1 port map( A1 => B(17), A2 => B(18), A3 => n243, ZN => n241);
   U77 : OR3_X1 port map( A1 => B(21), A2 => B(22), A3 => n239, ZN => n237);
   U78 : OR3_X1 port map( A1 => B(7), A2 => B(8), A3 => n192, ZN => n190);
   U79 : OR3_X1 port map( A1 => B(11), A2 => B(12), A3 => n249, ZN => n247);
   U80 : OR3_X1 port map( A1 => B(15), A2 => B(16), A3 => n245, ZN => n243);
   U83 : OR3_X1 port map( A1 => B(19), A2 => B(20), A3 => n241, ZN => n239);
   U116 : OR3_X1 port map( A1 => B(23), A2 => B(24), A3 => n237, ZN => n235);
   U120 : OR3_X1 port map( A1 => B(3), A2 => B(4), A3 => n211, ZN => n194);
   U123 : OR3_X1 port map( A1 => B(1), A2 => B(2), A3 => B(0), ZN => n211);
   U126 : INV_X1 port map( A => B(61), ZN => n251);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_8_DW01_sub_0 is

   port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (63 downto 0);  CO : out std_logic);

end complementer_N64_8_DW01_sub_0;

architecture SYN_rpl of complementer_N64_8_DW01_sub_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal DIFF_62_port, DIFF_61_port, DIFF_60_port, DIFF_59_port, DIFF_58_port,
      DIFF_57_port, DIFF_56_port, DIFF_55_port, DIFF_54_port, DIFF_53_port, 
      DIFF_52_port, DIFF_51_port, DIFF_50_port, DIFF_49_port, DIFF_48_port, 
      DIFF_47_port, DIFF_46_port, DIFF_45_port, DIFF_44_port, DIFF_43_port, 
      DIFF_42_port, DIFF_41_port, DIFF_40_port, DIFF_39_port, DIFF_38_port, 
      DIFF_37_port, DIFF_36_port, DIFF_35_port, DIFF_34_port, DIFF_33_port, 
      DIFF_32_port, DIFF_31_port, DIFF_30_port, DIFF_29_port, DIFF_28_port, 
      DIFF_27_port, DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, 
      DIFF_22_port, DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, 
      DIFF_17_port, DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, 
      DIFF_12_port, DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, 
      DIFF_7_port, DIFF_6_port, DIFF_5_port, DIFF_4_port, DIFF_3_port, 
      DIFF_2_port, DIFF_1_port, DIFF_63_port, n190, n191, n192, n193, n194, 
      n196, n197, n198, n199, n200, n202, n203, n204, n206, n207, n208, n210, 
      n211, n212, n213, n214, n216, n217, n218, n220, n221, n222, n224, n225, 
      n226, n228, n229, n230, n232, n233, n234, n235, n237, n238, n239, n240, 
      n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n189, 
      n195, n201, n205, n209, n215, n219, n223, n227, n231, n236 : std_logic;

begin
   DIFF <= ( DIFF_63_port, DIFF_62_port, DIFF_61_port, DIFF_60_port, 
      DIFF_59_port, DIFF_58_port, DIFF_57_port, DIFF_56_port, DIFF_55_port, 
      DIFF_54_port, DIFF_53_port, DIFF_52_port, DIFF_51_port, DIFF_50_port, 
      DIFF_49_port, DIFF_48_port, DIFF_47_port, DIFF_46_port, DIFF_45_port, 
      DIFF_44_port, DIFF_43_port, DIFF_42_port, DIFF_41_port, DIFF_40_port, 
      DIFF_39_port, DIFF_38_port, DIFF_37_port, DIFF_36_port, DIFF_35_port, 
      DIFF_34_port, DIFF_33_port, DIFF_32_port, DIFF_31_port, DIFF_30_port, 
      DIFF_29_port, DIFF_28_port, DIFF_27_port, DIFF_26_port, DIFF_25_port, 
      DIFF_24_port, DIFF_23_port, DIFF_22_port, DIFF_21_port, DIFF_20_port, 
      DIFF_19_port, DIFF_18_port, DIFF_17_port, DIFF_16_port, DIFF_15_port, 
      DIFF_14_port, DIFF_13_port, DIFF_12_port, DIFF_11_port, DIFF_10_port, 
      DIFF_9_port, DIFF_8_port, DIFF_7_port, DIFF_6_port, DIFF_5_port, 
      DIFF_4_port, DIFF_3_port, DIFF_2_port, DIFF_1_port, B(0) );
   
   U81 : XOR2_X1 port map( A => n190, B => B(9), Z => DIFF_9_port);
   U82 : XOR2_X1 port map( A => n192, B => B(7), Z => DIFF_7_port);
   U83 : XOR2_X1 port map( A => n193, B => B(6), Z => DIFF_6_port);
   U85 : XOR2_X1 port map( A => n196, B => B(62), Z => DIFF_62_port);
   U86 : XOR2_X1 port map( A => n194, B => B(5), Z => DIFF_5_port);
   U87 : XOR2_X1 port map( A => n198, B => B(59), Z => DIFF_59_port);
   U89 : XOR2_X1 port map( A => n200, B => B(57), Z => DIFF_57_port);
   U90 : XOR2_X1 port map( A => n202, B => B(55), Z => DIFF_55_port);
   U92 : XOR2_X1 port map( A => n204, B => B(53), Z => DIFF_53_port);
   U93 : XOR2_X1 port map( A => n206, B => B(51), Z => DIFF_51_port);
   U95 : XOR2_X1 port map( A => n208, B => B(49), Z => DIFF_49_port);
   U96 : XOR2_X1 port map( A => n212, B => B(47), Z => DIFF_47_port);
   U98 : XOR2_X1 port map( A => n214, B => B(45), Z => DIFF_45_port);
   U99 : XOR2_X1 port map( A => n216, B => B(43), Z => DIFF_43_port);
   U101 : XOR2_X1 port map( A => n218, B => B(41), Z => DIFF_41_port);
   U102 : XOR2_X1 port map( A => n211, B => B(3), Z => DIFF_3_port);
   U103 : XOR2_X1 port map( A => n220, B => B(39), Z => DIFF_39_port);
   U105 : XOR2_X1 port map( A => n222, B => B(37), Z => DIFF_37_port);
   U106 : XOR2_X1 port map( A => n224, B => B(35), Z => DIFF_35_port);
   U108 : XOR2_X1 port map( A => n226, B => B(33), Z => DIFF_33_port);
   U109 : XOR2_X1 port map( A => n228, B => B(31), Z => DIFF_31_port);
   U111 : XOR2_X1 port map( A => n230, B => B(29), Z => DIFF_29_port);
   U112 : XOR2_X1 port map( A => n233, B => B(27), Z => DIFF_27_port);
   U114 : XOR2_X1 port map( A => n235, B => B(25), Z => DIFF_25_port);
   U115 : XOR2_X1 port map( A => n237, B => B(23), Z => DIFF_23_port);
   U116 : XOR2_X1 port map( A => n240, B => B(22), Z => DIFF_22_port);
   U117 : XOR2_X1 port map( A => n239, B => B(21), Z => DIFF_21_port);
   U118 : XOR2_X1 port map( A => B(1), B => B(0), Z => DIFF_1_port);
   U119 : XOR2_X1 port map( A => n241, B => B(19), Z => DIFF_19_port);
   U120 : XOR2_X1 port map( A => n244, B => B(18), Z => DIFF_18_port);
   U121 : XOR2_X1 port map( A => n243, B => B(17), Z => DIFF_17_port);
   U122 : XOR2_X1 port map( A => n245, B => B(15), Z => DIFF_15_port);
   U123 : XOR2_X1 port map( A => n248, B => B(14), Z => DIFF_14_port);
   U124 : XOR2_X1 port map( A => n247, B => B(13), Z => DIFF_13_port);
   U125 : XOR2_X1 port map( A => n249, B => B(11), Z => DIFF_11_port);
   U126 : XOR2_X1 port map( A => n251, B => B(10), Z => DIFF_10_port);
   U1 : XOR2_X1 port map( A => n197, B => n236, Z => DIFF_61_port);
   U2 : NAND2_X1 port map( A1 => n197, A2 => n236, ZN => n196);
   U3 : XNOR2_X1 port map( A => n189, B => B(50), ZN => DIFF_50_port);
   U4 : NOR2_X1 port map( A1 => n208, A2 => B(49), ZN => n189);
   U5 : XNOR2_X1 port map( A => n195, B => B(46), ZN => DIFF_46_port);
   U6 : NOR2_X1 port map( A1 => n214, A2 => B(45), ZN => n195);
   U7 : XNOR2_X1 port map( A => n201, B => B(42), ZN => DIFF_42_port);
   U8 : NOR2_X1 port map( A1 => n218, A2 => B(41), ZN => n201);
   U9 : XNOR2_X1 port map( A => B(52), B => n207, ZN => DIFF_52_port);
   U10 : NOR2_X1 port map( A1 => B(51), A2 => n206, ZN => n207);
   U11 : XNOR2_X1 port map( A => B(48), B => n213, ZN => DIFF_48_port);
   U12 : NOR2_X1 port map( A1 => B(47), A2 => n212, ZN => n213);
   U13 : XNOR2_X1 port map( A => B(44), B => n217, ZN => DIFF_44_port);
   U14 : NOR2_X1 port map( A1 => B(43), A2 => n216, ZN => n217);
   U15 : XNOR2_X1 port map( A => B(40), B => n221, ZN => DIFF_40_port);
   U16 : NOR2_X1 port map( A1 => B(39), A2 => n220, ZN => n221);
   U17 : XNOR2_X1 port map( A => B(36), B => n225, ZN => DIFF_36_port);
   U18 : NOR2_X1 port map( A1 => B(35), A2 => n224, ZN => n225);
   U19 : OR3_X1 port map( A1 => B(33), A2 => B(34), A3 => n226, ZN => n224);
   U20 : OR3_X1 port map( A1 => B(37), A2 => B(38), A3 => n222, ZN => n220);
   U21 : OR3_X1 port map( A1 => B(41), A2 => B(42), A3 => n218, ZN => n216);
   U22 : OR3_X1 port map( A1 => B(45), A2 => B(46), A3 => n214, ZN => n212);
   U23 : OR3_X1 port map( A1 => B(49), A2 => B(50), A3 => n208, ZN => n206);
   U24 : OR3_X1 port map( A1 => B(35), A2 => B(36), A3 => n224, ZN => n222);
   U25 : OR3_X1 port map( A1 => B(39), A2 => B(40), A3 => n220, ZN => n218);
   U26 : OR3_X1 port map( A1 => B(43), A2 => B(44), A3 => n216, ZN => n214);
   U27 : OR3_X1 port map( A1 => B(47), A2 => B(48), A3 => n212, ZN => n208);
   U28 : XNOR2_X1 port map( A => n205, B => B(38), ZN => DIFF_38_port);
   U29 : NOR2_X1 port map( A1 => n222, A2 => B(37), ZN => n205);
   U30 : XNOR2_X1 port map( A => n209, B => B(34), ZN => DIFF_34_port);
   U31 : NOR2_X1 port map( A1 => n226, A2 => B(33), ZN => n209);
   U32 : NOR3_X1 port map( A1 => B(59), A2 => B(60), A3 => n198, ZN => n197);
   U33 : XNOR2_X1 port map( A => n215, B => B(54), ZN => DIFF_54_port);
   U34 : NOR2_X1 port map( A1 => n204, A2 => B(53), ZN => n215);
   U35 : XNOR2_X1 port map( A => B(60), B => n199, ZN => DIFF_60_port);
   U36 : NOR2_X1 port map( A1 => B(59), A2 => n198, ZN => n199);
   U37 : XNOR2_X1 port map( A => B(56), B => n203, ZN => DIFF_56_port);
   U38 : NOR2_X1 port map( A1 => B(55), A2 => n202, ZN => n203);
   U39 : OR3_X1 port map( A1 => B(57), A2 => B(58), A3 => n200, ZN => n198);
   U40 : OR3_X1 port map( A1 => B(53), A2 => B(54), A3 => n204, ZN => n202);
   U41 : OR3_X1 port map( A1 => B(51), A2 => B(52), A3 => n206, ZN => n204);
   U42 : OR3_X1 port map( A1 => B(55), A2 => B(56), A3 => n202, ZN => n200);
   U43 : XNOR2_X1 port map( A => n219, B => B(58), ZN => DIFF_58_port);
   U44 : NOR2_X1 port map( A1 => n200, A2 => B(57), ZN => n219);
   U45 : XNOR2_X1 port map( A => B(32), B => n229, ZN => DIFF_32_port);
   U46 : NOR2_X1 port map( A1 => B(31), A2 => n228, ZN => n229);
   U47 : OR3_X1 port map( A1 => B(31), A2 => B(32), A3 => n228, ZN => n226);
   U48 : XNOR2_X1 port map( A => n223, B => B(63), ZN => DIFF_63_port);
   U49 : NOR2_X1 port map( A1 => n196, A2 => B(62), ZN => n223);
   U50 : OR3_X1 port map( A1 => B(29), A2 => B(30), A3 => n230, ZN => n228);
   U51 : XNOR2_X1 port map( A => n227, B => B(30), ZN => DIFF_30_port);
   U52 : NOR2_X1 port map( A1 => n230, A2 => B(29), ZN => n227);
   U53 : XNOR2_X1 port map( A => B(28), B => n234, ZN => DIFF_28_port);
   U54 : NOR2_X1 port map( A1 => B(27), A2 => n233, ZN => n234);
   U55 : OR3_X1 port map( A1 => B(27), A2 => B(28), A3 => n233, ZN => n230);
   U56 : OR3_X1 port map( A1 => B(25), A2 => B(26), A3 => n235, ZN => n233);
   U57 : XNOR2_X1 port map( A => n231, B => B(26), ZN => DIFF_26_port);
   U58 : NOR2_X1 port map( A1 => n235, A2 => B(25), ZN => n231);
   U59 : OR3_X1 port map( A1 => B(23), A2 => B(24), A3 => n237, ZN => n235);
   U60 : XNOR2_X1 port map( A => B(24), B => n238, ZN => DIFF_24_port);
   U61 : NOR2_X1 port map( A1 => B(23), A2 => n237, ZN => n238);
   U62 : NOR2_X1 port map( A1 => B(19), A2 => n241, ZN => n242);
   U63 : NOR2_X1 port map( A1 => B(15), A2 => n245, ZN => n246);
   U64 : NOR2_X1 port map( A1 => B(11), A2 => n249, ZN => n250);
   U65 : NOR2_X1 port map( A1 => B(7), A2 => n192, ZN => n191);
   U66 : NOR2_X1 port map( A1 => B(3), A2 => n211, ZN => n210);
   U67 : OR3_X1 port map( A1 => B(21), A2 => B(22), A3 => n239, ZN => n237);
   U68 : OR3_X1 port map( A1 => B(17), A2 => B(18), A3 => n243, ZN => n241);
   U69 : OR3_X1 port map( A1 => B(13), A2 => B(14), A3 => n247, ZN => n245);
   U70 : OR3_X1 port map( A1 => B(10), A2 => B(9), A3 => n190, ZN => n249);
   U71 : OR3_X1 port map( A1 => B(5), A2 => B(6), A3 => n194, ZN => n192);
   U72 : OR3_X1 port map( A1 => B(19), A2 => B(20), A3 => n241, ZN => n239);
   U73 : OR3_X1 port map( A1 => B(15), A2 => B(16), A3 => n245, ZN => n243);
   U74 : OR3_X1 port map( A1 => B(11), A2 => B(12), A3 => n249, ZN => n247);
   U75 : OR3_X1 port map( A1 => B(7), A2 => B(8), A3 => n192, ZN => n190);
   U76 : OR3_X1 port map( A1 => B(3), A2 => B(4), A3 => n211, ZN => n194);
   U77 : XNOR2_X1 port map( A => B(20), B => n242, ZN => DIFF_20_port);
   U78 : XNOR2_X1 port map( A => B(16), B => n246, ZN => DIFF_16_port);
   U79 : XNOR2_X1 port map( A => B(12), B => n250, ZN => DIFF_12_port);
   U80 : XNOR2_X1 port map( A => B(8), B => n191, ZN => DIFF_8_port);
   U84 : XNOR2_X1 port map( A => B(4), B => n210, ZN => DIFF_4_port);
   U88 : XNOR2_X1 port map( A => B(2), B => n232, ZN => DIFF_2_port);
   U91 : OR2_X1 port map( A1 => n239, A2 => B(21), ZN => n240);
   U94 : OR2_X1 port map( A1 => n243, A2 => B(17), ZN => n244);
   U97 : OR2_X1 port map( A1 => n247, A2 => B(13), ZN => n248);
   U100 : OR2_X1 port map( A1 => n190, A2 => B(9), ZN => n251);
   U104 : OR2_X1 port map( A1 => n194, A2 => B(5), ZN => n193);
   U107 : OR3_X1 port map( A1 => B(1), A2 => B(2), A3 => B(0), ZN => n211);
   U110 : NOR2_X1 port map( A1 => B(0), A2 => B(1), ZN => n232);
   U113 : INV_X1 port map( A => B(61), ZN => n236);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_9_DW01_sub_0 is

   port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (63 downto 0);  CO : out std_logic);

end complementer_N64_9_DW01_sub_0;

architecture SYN_rpl of complementer_N64_9_DW01_sub_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal DIFF_62_port, DIFF_63_port, DIFF_23_port, DIFF_24_port, DIFF_25_port,
      DIFF_26_port, DIFF_27_port, DIFF_28_port, DIFF_29_port, DIFF_30_port, 
      DIFF_31_port, DIFF_32_port, DIFF_33_port, DIFF_34_port, DIFF_35_port, 
      DIFF_36_port, DIFF_37_port, DIFF_38_port, DIFF_39_port, DIFF_40_port, 
      DIFF_41_port, DIFF_42_port, DIFF_43_port, DIFF_44_port, DIFF_45_port, 
      DIFF_46_port, DIFF_47_port, DIFF_48_port, DIFF_49_port, DIFF_50_port, 
      DIFF_51_port, DIFF_52_port, DIFF_53_port, DIFF_54_port, DIFF_55_port, 
      DIFF_56_port, DIFF_57_port, DIFF_58_port, DIFF_59_port, DIFF_60_port, 
      DIFF_61_port, DIFF_3_port, DIFF_4_port, DIFF_5_port, DIFF_6_port, 
      DIFF_7_port, DIFF_8_port, DIFF_9_port, DIFF_10_port, DIFF_11_port, 
      DIFF_12_port, DIFF_13_port, DIFF_14_port, DIFF_15_port, DIFF_16_port, 
      DIFF_17_port, DIFF_18_port, DIFF_19_port, DIFF_20_port, DIFF_21_port, 
      DIFF_22_port, DIFF_2_port, DIFF_1_port, n190, n191, n192, n194, n195, 
      n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, 
      n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, 
      n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, 
      n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, 
      n245, n246, n247, n249, n250, n189, n193, n244, n248, n251 : std_logic;

begin
   DIFF <= ( DIFF_63_port, DIFF_62_port, DIFF_61_port, DIFF_60_port, 
      DIFF_59_port, DIFF_58_port, DIFF_57_port, DIFF_56_port, DIFF_55_port, 
      DIFF_54_port, DIFF_53_port, DIFF_52_port, DIFF_51_port, DIFF_50_port, 
      DIFF_49_port, DIFF_48_port, DIFF_47_port, DIFF_46_port, DIFF_45_port, 
      DIFF_44_port, DIFF_43_port, DIFF_42_port, DIFF_41_port, DIFF_40_port, 
      DIFF_39_port, DIFF_38_port, DIFF_37_port, DIFF_36_port, DIFF_35_port, 
      DIFF_34_port, DIFF_33_port, DIFF_32_port, DIFF_31_port, DIFF_30_port, 
      DIFF_29_port, DIFF_28_port, DIFF_27_port, DIFF_26_port, DIFF_25_port, 
      DIFF_24_port, DIFF_23_port, DIFF_22_port, DIFF_21_port, DIFF_20_port, 
      DIFF_19_port, DIFF_18_port, DIFF_17_port, DIFF_16_port, DIFF_15_port, 
      DIFF_14_port, DIFF_13_port, DIFF_12_port, DIFF_11_port, DIFF_10_port, 
      DIFF_9_port, DIFF_8_port, DIFF_7_port, DIFF_6_port, DIFF_5_port, 
      DIFF_4_port, DIFF_3_port, DIFF_2_port, DIFF_1_port, B(0) );
   
   U81 : XOR2_X1 port map( A => n190, B => B(9), Z => DIFF_9_port);
   U82 : XOR2_X1 port map( A => n192, B => B(7), Z => DIFF_7_port);
   U84 : XOR2_X1 port map( A => n195, B => B(63), Z => DIFF_63_port);
   U85 : XOR2_X1 port map( A => n196, B => B(62), Z => DIFF_62_port);
   U86 : XOR2_X1 port map( A => n194, B => B(5), Z => DIFF_5_port);
   U87 : XOR2_X1 port map( A => n198, B => B(59), Z => DIFF_59_port);
   U88 : XOR2_X1 port map( A => n201, B => B(58), Z => DIFF_58_port);
   U89 : XOR2_X1 port map( A => n200, B => B(57), Z => DIFF_57_port);
   U90 : XOR2_X1 port map( A => n202, B => B(55), Z => DIFF_55_port);
   U91 : XOR2_X1 port map( A => n205, B => B(54), Z => DIFF_54_port);
   U92 : XOR2_X1 port map( A => n204, B => B(53), Z => DIFF_53_port);
   U93 : XOR2_X1 port map( A => n206, B => B(51), Z => DIFF_51_port);
   U94 : XOR2_X1 port map( A => n209, B => B(50), Z => DIFF_50_port);
   U95 : XOR2_X1 port map( A => n208, B => B(49), Z => DIFF_49_port);
   U96 : XOR2_X1 port map( A => n212, B => B(47), Z => DIFF_47_port);
   U97 : XOR2_X1 port map( A => n215, B => B(46), Z => DIFF_46_port);
   U98 : XOR2_X1 port map( A => n214, B => B(45), Z => DIFF_45_port);
   U99 : XOR2_X1 port map( A => n216, B => B(43), Z => DIFF_43_port);
   U100 : XOR2_X1 port map( A => n219, B => B(42), Z => DIFF_42_port);
   U101 : XOR2_X1 port map( A => n218, B => B(41), Z => DIFF_41_port);
   U102 : XOR2_X1 port map( A => n211, B => B(3), Z => DIFF_3_port);
   U103 : XOR2_X1 port map( A => n220, B => B(39), Z => DIFF_39_port);
   U104 : XOR2_X1 port map( A => n223, B => B(38), Z => DIFF_38_port);
   U105 : XOR2_X1 port map( A => n222, B => B(37), Z => DIFF_37_port);
   U106 : XOR2_X1 port map( A => n224, B => B(35), Z => DIFF_35_port);
   U107 : XOR2_X1 port map( A => n227, B => B(34), Z => DIFF_34_port);
   U108 : XOR2_X1 port map( A => n226, B => B(33), Z => DIFF_33_port);
   U109 : XOR2_X1 port map( A => n228, B => B(31), Z => DIFF_31_port);
   U110 : XOR2_X1 port map( A => n231, B => B(30), Z => DIFF_30_port);
   U111 : XOR2_X1 port map( A => n230, B => B(29), Z => DIFF_29_port);
   U112 : XOR2_X1 port map( A => n233, B => B(27), Z => DIFF_27_port);
   U113 : XOR2_X1 port map( A => n236, B => B(26), Z => DIFF_26_port);
   U114 : XOR2_X1 port map( A => n235, B => B(25), Z => DIFF_25_port);
   U115 : XOR2_X1 port map( A => n237, B => B(23), Z => DIFF_23_port);
   U116 : XOR2_X1 port map( A => n240, B => B(22), Z => DIFF_22_port);
   U117 : XOR2_X1 port map( A => n239, B => B(21), Z => DIFF_21_port);
   U118 : XOR2_X1 port map( A => B(1), B => B(0), Z => DIFF_1_port);
   U119 : XOR2_X1 port map( A => n241, B => B(19), Z => DIFF_19_port);
   U121 : XOR2_X1 port map( A => n243, B => B(17), Z => DIFF_17_port);
   U122 : XOR2_X1 port map( A => n245, B => B(15), Z => DIFF_15_port);
   U124 : XOR2_X1 port map( A => n247, B => B(13), Z => DIFF_13_port);
   U125 : XOR2_X1 port map( A => n249, B => B(11), Z => DIFF_11_port);
   U1 : NAND2_X1 port map( A1 => n197, A2 => n251, ZN => n196);
   U2 : NOR2_X1 port map( A1 => B(51), A2 => n206, ZN => n207);
   U3 : NOR2_X1 port map( A1 => B(47), A2 => n212, ZN => n213);
   U4 : NOR2_X1 port map( A1 => B(43), A2 => n216, ZN => n217);
   U5 : NOR2_X1 port map( A1 => B(39), A2 => n220, ZN => n221);
   U6 : NOR2_X1 port map( A1 => B(35), A2 => n224, ZN => n225);
   U7 : NOR2_X1 port map( A1 => B(31), A2 => n228, ZN => n229);
   U8 : NOR2_X1 port map( A1 => B(55), A2 => n202, ZN => n203);
   U9 : OR3_X1 port map( A1 => B(53), A2 => B(54), A3 => n204, ZN => n202);
   U10 : OR3_X1 port map( A1 => B(49), A2 => B(50), A3 => n208, ZN => n206);
   U11 : OR3_X1 port map( A1 => B(45), A2 => B(46), A3 => n214, ZN => n212);
   U12 : OR3_X1 port map( A1 => B(41), A2 => B(42), A3 => n218, ZN => n216);
   U13 : OR3_X1 port map( A1 => B(37), A2 => B(38), A3 => n222, ZN => n220);
   U14 : OR3_X1 port map( A1 => B(33), A2 => B(34), A3 => n226, ZN => n224);
   U15 : OR3_X1 port map( A1 => B(51), A2 => B(52), A3 => n206, ZN => n204);
   U16 : OR3_X1 port map( A1 => B(47), A2 => B(48), A3 => n212, ZN => n208);
   U17 : OR3_X1 port map( A1 => B(43), A2 => B(44), A3 => n216, ZN => n214);
   U18 : OR3_X1 port map( A1 => B(39), A2 => B(40), A3 => n220, ZN => n218);
   U19 : OR3_X1 port map( A1 => B(35), A2 => B(36), A3 => n224, ZN => n222);
   U20 : OR3_X1 port map( A1 => B(31), A2 => B(32), A3 => n228, ZN => n226);
   U21 : OR2_X1 port map( A1 => n204, A2 => B(53), ZN => n205);
   U22 : OR2_X1 port map( A1 => n208, A2 => B(49), ZN => n209);
   U23 : OR2_X1 port map( A1 => n214, A2 => B(45), ZN => n215);
   U24 : OR2_X1 port map( A1 => n218, A2 => B(41), ZN => n219);
   U25 : OR2_X1 port map( A1 => n222, A2 => B(37), ZN => n223);
   U26 : OR2_X1 port map( A1 => n226, A2 => B(33), ZN => n227);
   U27 : NOR3_X1 port map( A1 => B(59), A2 => B(60), A3 => n198, ZN => n197);
   U28 : NOR2_X1 port map( A1 => B(59), A2 => n198, ZN => n199);
   U29 : OR2_X1 port map( A1 => n230, A2 => B(29), ZN => n231);
   U30 : OR3_X1 port map( A1 => B(29), A2 => B(30), A3 => n230, ZN => n228);
   U31 : OR3_X1 port map( A1 => B(55), A2 => B(56), A3 => n202, ZN => n200);
   U32 : OR3_X1 port map( A1 => B(57), A2 => B(58), A3 => n200, ZN => n198);
   U33 : OR2_X1 port map( A1 => n196, A2 => B(62), ZN => n195);
   U34 : OR2_X1 port map( A1 => n200, A2 => B(57), ZN => n201);
   U35 : NOR2_X1 port map( A1 => B(27), A2 => n233, ZN => n234);
   U36 : OR3_X1 port map( A1 => B(27), A2 => B(28), A3 => n233, ZN => n230);
   U37 : XNOR2_X1 port map( A => B(32), B => n229, ZN => DIFF_32_port);
   U38 : XNOR2_X1 port map( A => B(28), B => n234, ZN => DIFF_28_port);
   U39 : XNOR2_X1 port map( A => B(56), B => n203, ZN => DIFF_56_port);
   U40 : XNOR2_X1 port map( A => B(52), B => n207, ZN => DIFF_52_port);
   U41 : XNOR2_X1 port map( A => B(48), B => n213, ZN => DIFF_48_port);
   U42 : XNOR2_X1 port map( A => B(44), B => n217, ZN => DIFF_44_port);
   U43 : XNOR2_X1 port map( A => B(40), B => n221, ZN => DIFF_40_port);
   U44 : XNOR2_X1 port map( A => B(36), B => n225, ZN => DIFF_36_port);
   U45 : XNOR2_X1 port map( A => n197, B => B(61), ZN => DIFF_61_port);
   U46 : XNOR2_X1 port map( A => B(60), B => n199, ZN => DIFF_60_port);
   U47 : OR3_X1 port map( A1 => B(25), A2 => B(26), A3 => n235, ZN => n233);
   U48 : XNOR2_X1 port map( A => B(24), B => n238, ZN => DIFF_24_port);
   U49 : OR2_X1 port map( A1 => n235, A2 => B(25), ZN => n236);
   U50 : NOR2_X1 port map( A1 => B(23), A2 => n237, ZN => n238);
   U51 : OR3_X1 port map( A1 => B(23), A2 => B(24), A3 => n237, ZN => n235);
   U52 : XNOR2_X1 port map( A => n189, B => B(18), ZN => DIFF_18_port);
   U53 : NOR2_X1 port map( A1 => n243, A2 => B(17), ZN => n189);
   U54 : XNOR2_X1 port map( A => n193, B => B(14), ZN => DIFF_14_port);
   U55 : NOR2_X1 port map( A1 => n247, A2 => B(13), ZN => n193);
   U56 : XNOR2_X1 port map( A => n244, B => B(10), ZN => DIFF_10_port);
   U57 : NOR2_X1 port map( A1 => n190, A2 => B(9), ZN => n244);
   U58 : XNOR2_X1 port map( A => n248, B => B(6), ZN => DIFF_6_port);
   U59 : NOR2_X1 port map( A1 => n194, A2 => B(5), ZN => n248);
   U60 : XNOR2_X1 port map( A => B(20), B => n242, ZN => DIFF_20_port);
   U61 : NOR2_X1 port map( A1 => B(19), A2 => n241, ZN => n242);
   U62 : XNOR2_X1 port map( A => B(16), B => n246, ZN => DIFF_16_port);
   U63 : NOR2_X1 port map( A1 => B(15), A2 => n245, ZN => n246);
   U64 : XNOR2_X1 port map( A => B(12), B => n250, ZN => DIFF_12_port);
   U65 : NOR2_X1 port map( A1 => B(11), A2 => n249, ZN => n250);
   U66 : XNOR2_X1 port map( A => B(8), B => n191, ZN => DIFF_8_port);
   U67 : NOR2_X1 port map( A1 => B(7), A2 => n192, ZN => n191);
   U68 : XNOR2_X1 port map( A => B(2), B => n232, ZN => DIFF_2_port);
   U69 : NOR2_X1 port map( A1 => B(0), A2 => B(1), ZN => n232);
   U70 : XNOR2_X1 port map( A => B(4), B => n210, ZN => DIFF_4_port);
   U71 : NOR2_X1 port map( A1 => B(3), A2 => n211, ZN => n210);
   U72 : OR3_X1 port map( A1 => B(5), A2 => B(6), A3 => n194, ZN => n192);
   U73 : OR3_X1 port map( A1 => B(10), A2 => B(9), A3 => n190, ZN => n249);
   U74 : OR3_X1 port map( A1 => B(13), A2 => B(14), A3 => n247, ZN => n245);
   U75 : OR3_X1 port map( A1 => B(17), A2 => B(18), A3 => n243, ZN => n241);
   U76 : OR3_X1 port map( A1 => B(21), A2 => B(22), A3 => n239, ZN => n237);
   U77 : OR3_X1 port map( A1 => B(7), A2 => B(8), A3 => n192, ZN => n190);
   U78 : OR3_X1 port map( A1 => B(11), A2 => B(12), A3 => n249, ZN => n247);
   U79 : OR3_X1 port map( A1 => B(15), A2 => B(16), A3 => n245, ZN => n243);
   U80 : OR3_X1 port map( A1 => B(19), A2 => B(20), A3 => n241, ZN => n239);
   U83 : OR3_X1 port map( A1 => B(3), A2 => B(4), A3 => n211, ZN => n194);
   U120 : OR2_X1 port map( A1 => n239, A2 => B(21), ZN => n240);
   U123 : OR3_X1 port map( A1 => B(1), A2 => B(2), A3 => B(0), ZN => n211);
   U126 : INV_X1 port map( A => B(61), ZN => n251);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_10_DW01_sub_0 is

   port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (63 downto 0);  CO : out std_logic);

end complementer_N64_10_DW01_sub_0;

architecture SYN_rpl of complementer_N64_10_DW01_sub_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal DIFF_62_port, DIFF_61_port, DIFF_60_port, DIFF_59_port, DIFF_58_port,
      DIFF_57_port, DIFF_56_port, DIFF_55_port, DIFF_54_port, DIFF_53_port, 
      DIFF_52_port, DIFF_51_port, DIFF_50_port, DIFF_49_port, DIFF_48_port, 
      DIFF_47_port, DIFF_46_port, DIFF_45_port, DIFF_44_port, DIFF_43_port, 
      DIFF_42_port, DIFF_41_port, DIFF_40_port, DIFF_39_port, DIFF_38_port, 
      DIFF_37_port, DIFF_36_port, DIFF_35_port, DIFF_34_port, DIFF_33_port, 
      DIFF_32_port, DIFF_31_port, DIFF_30_port, DIFF_29_port, DIFF_28_port, 
      DIFF_27_port, DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, 
      DIFF_22_port, DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, 
      DIFF_17_port, DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, 
      DIFF_12_port, DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, 
      DIFF_7_port, DIFF_6_port, DIFF_5_port, DIFF_4_port, DIFF_3_port, 
      DIFF_2_port, DIFF_1_port, DIFF_63_port, n190, n191, n192, n193, n194, 
      n196, n197, n198, n199, n200, n202, n203, n204, n206, n207, n208, n210, 
      n211, n212, n213, n214, n216, n217, n218, n220, n221, n222, n224, n225, 
      n226, n228, n229, n230, n232, n233, n234, n235, n237, n238, n239, n241, 
      n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n189, n195, 
      n201, n205, n209, n215, n219, n223, n227, n231, n236, n240 : std_logic;

begin
   DIFF <= ( DIFF_63_port, DIFF_62_port, DIFF_61_port, DIFF_60_port, 
      DIFF_59_port, DIFF_58_port, DIFF_57_port, DIFF_56_port, DIFF_55_port, 
      DIFF_54_port, DIFF_53_port, DIFF_52_port, DIFF_51_port, DIFF_50_port, 
      DIFF_49_port, DIFF_48_port, DIFF_47_port, DIFF_46_port, DIFF_45_port, 
      DIFF_44_port, DIFF_43_port, DIFF_42_port, DIFF_41_port, DIFF_40_port, 
      DIFF_39_port, DIFF_38_port, DIFF_37_port, DIFF_36_port, DIFF_35_port, 
      DIFF_34_port, DIFF_33_port, DIFF_32_port, DIFF_31_port, DIFF_30_port, 
      DIFF_29_port, DIFF_28_port, DIFF_27_port, DIFF_26_port, DIFF_25_port, 
      DIFF_24_port, DIFF_23_port, DIFF_22_port, DIFF_21_port, DIFF_20_port, 
      DIFF_19_port, DIFF_18_port, DIFF_17_port, DIFF_16_port, DIFF_15_port, 
      DIFF_14_port, DIFF_13_port, DIFF_12_port, DIFF_11_port, DIFF_10_port, 
      DIFF_9_port, DIFF_8_port, DIFF_7_port, DIFF_6_port, DIFF_5_port, 
      DIFF_4_port, DIFF_3_port, DIFF_2_port, DIFF_1_port, B(0) );
   
   U81 : XOR2_X1 port map( A => n190, B => B(9), Z => DIFF_9_port);
   U82 : XOR2_X1 port map( A => n192, B => B(7), Z => DIFF_7_port);
   U83 : XOR2_X1 port map( A => n193, B => B(6), Z => DIFF_6_port);
   U85 : XOR2_X1 port map( A => n196, B => B(62), Z => DIFF_62_port);
   U86 : XOR2_X1 port map( A => n194, B => B(5), Z => DIFF_5_port);
   U87 : XOR2_X1 port map( A => n198, B => B(59), Z => DIFF_59_port);
   U89 : XOR2_X1 port map( A => n200, B => B(57), Z => DIFF_57_port);
   U90 : XOR2_X1 port map( A => n202, B => B(55), Z => DIFF_55_port);
   U92 : XOR2_X1 port map( A => n204, B => B(53), Z => DIFF_53_port);
   U93 : XOR2_X1 port map( A => n206, B => B(51), Z => DIFF_51_port);
   U95 : XOR2_X1 port map( A => n208, B => B(49), Z => DIFF_49_port);
   U96 : XOR2_X1 port map( A => n212, B => B(47), Z => DIFF_47_port);
   U98 : XOR2_X1 port map( A => n214, B => B(45), Z => DIFF_45_port);
   U99 : XOR2_X1 port map( A => n216, B => B(43), Z => DIFF_43_port);
   U101 : XOR2_X1 port map( A => n218, B => B(41), Z => DIFF_41_port);
   U102 : XOR2_X1 port map( A => n211, B => B(3), Z => DIFF_3_port);
   U103 : XOR2_X1 port map( A => n220, B => B(39), Z => DIFF_39_port);
   U105 : XOR2_X1 port map( A => n222, B => B(37), Z => DIFF_37_port);
   U106 : XOR2_X1 port map( A => n224, B => B(35), Z => DIFF_35_port);
   U108 : XOR2_X1 port map( A => n226, B => B(33), Z => DIFF_33_port);
   U109 : XOR2_X1 port map( A => n228, B => B(31), Z => DIFF_31_port);
   U111 : XOR2_X1 port map( A => n230, B => B(29), Z => DIFF_29_port);
   U112 : XOR2_X1 port map( A => n233, B => B(27), Z => DIFF_27_port);
   U114 : XOR2_X1 port map( A => n235, B => B(25), Z => DIFF_25_port);
   U115 : XOR2_X1 port map( A => n237, B => B(23), Z => DIFF_23_port);
   U117 : XOR2_X1 port map( A => n239, B => B(21), Z => DIFF_21_port);
   U118 : XOR2_X1 port map( A => B(1), B => B(0), Z => DIFF_1_port);
   U119 : XOR2_X1 port map( A => n241, B => B(19), Z => DIFF_19_port);
   U120 : XOR2_X1 port map( A => n244, B => B(18), Z => DIFF_18_port);
   U121 : XOR2_X1 port map( A => n243, B => B(17), Z => DIFF_17_port);
   U122 : XOR2_X1 port map( A => n245, B => B(15), Z => DIFF_15_port);
   U123 : XOR2_X1 port map( A => n248, B => B(14), Z => DIFF_14_port);
   U124 : XOR2_X1 port map( A => n247, B => B(13), Z => DIFF_13_port);
   U125 : XOR2_X1 port map( A => n249, B => B(11), Z => DIFF_11_port);
   U126 : XOR2_X1 port map( A => n251, B => B(10), Z => DIFF_10_port);
   U1 : XNOR2_X1 port map( A => B(32), B => n229, ZN => DIFF_32_port);
   U2 : NOR2_X1 port map( A1 => B(31), A2 => n228, ZN => n229);
   U3 : OR3_X1 port map( A1 => B(31), A2 => B(32), A3 => n228, ZN => n226);
   U4 : XNOR2_X1 port map( A => n189, B => B(50), ZN => DIFF_50_port);
   U5 : NOR2_X1 port map( A1 => n208, A2 => B(49), ZN => n189);
   U6 : XNOR2_X1 port map( A => n195, B => B(46), ZN => DIFF_46_port);
   U7 : NOR2_X1 port map( A1 => n214, A2 => B(45), ZN => n195);
   U8 : XNOR2_X1 port map( A => n201, B => B(42), ZN => DIFF_42_port);
   U9 : NOR2_X1 port map( A1 => n218, A2 => B(41), ZN => n201);
   U10 : XNOR2_X1 port map( A => n205, B => B(38), ZN => DIFF_38_port);
   U11 : NOR2_X1 port map( A1 => n222, A2 => B(37), ZN => n205);
   U12 : XNOR2_X1 port map( A => n209, B => B(34), ZN => DIFF_34_port);
   U13 : NOR2_X1 port map( A1 => n226, A2 => B(33), ZN => n209);
   U14 : XNOR2_X1 port map( A => n215, B => B(54), ZN => DIFF_54_port);
   U15 : NOR2_X1 port map( A1 => n204, A2 => B(53), ZN => n215);
   U16 : XNOR2_X1 port map( A => B(36), B => n225, ZN => DIFF_36_port);
   U17 : NOR2_X1 port map( A1 => B(35), A2 => n224, ZN => n225);
   U18 : XNOR2_X1 port map( A => B(52), B => n207, ZN => DIFF_52_port);
   U19 : NOR2_X1 port map( A1 => B(51), A2 => n206, ZN => n207);
   U20 : XNOR2_X1 port map( A => B(48), B => n213, ZN => DIFF_48_port);
   U21 : NOR2_X1 port map( A1 => B(47), A2 => n212, ZN => n213);
   U22 : XNOR2_X1 port map( A => B(44), B => n217, ZN => DIFF_44_port);
   U23 : NOR2_X1 port map( A1 => B(43), A2 => n216, ZN => n217);
   U24 : XNOR2_X1 port map( A => B(40), B => n221, ZN => DIFF_40_port);
   U25 : NOR2_X1 port map( A1 => B(39), A2 => n220, ZN => n221);
   U26 : OR3_X1 port map( A1 => B(57), A2 => B(58), A3 => n200, ZN => n198);
   U27 : OR3_X1 port map( A1 => B(33), A2 => B(34), A3 => n226, ZN => n224);
   U28 : OR3_X1 port map( A1 => B(37), A2 => B(38), A3 => n222, ZN => n220);
   U29 : OR3_X1 port map( A1 => B(41), A2 => B(42), A3 => n218, ZN => n216);
   U30 : OR3_X1 port map( A1 => B(45), A2 => B(46), A3 => n214, ZN => n212);
   U31 : OR3_X1 port map( A1 => B(49), A2 => B(50), A3 => n208, ZN => n206);
   U32 : OR3_X1 port map( A1 => B(53), A2 => B(54), A3 => n204, ZN => n202);
   U33 : OR3_X1 port map( A1 => B(35), A2 => B(36), A3 => n224, ZN => n222);
   U34 : OR3_X1 port map( A1 => B(39), A2 => B(40), A3 => n220, ZN => n218);
   U35 : OR3_X1 port map( A1 => B(43), A2 => B(44), A3 => n216, ZN => n214);
   U36 : OR3_X1 port map( A1 => B(47), A2 => B(48), A3 => n212, ZN => n208);
   U37 : OR3_X1 port map( A1 => B(51), A2 => B(52), A3 => n206, ZN => n204);
   U38 : XNOR2_X1 port map( A => n219, B => B(58), ZN => DIFF_58_port);
   U39 : NOR2_X1 port map( A1 => n200, A2 => B(57), ZN => n219);
   U40 : NOR3_X1 port map( A1 => B(59), A2 => B(60), A3 => n198, ZN => n197);
   U41 : XNOR2_X1 port map( A => B(60), B => n199, ZN => DIFF_60_port);
   U42 : NOR2_X1 port map( A1 => B(59), A2 => n198, ZN => n199);
   U43 : XOR2_X1 port map( A => n197, B => n240, Z => DIFF_61_port);
   U44 : NAND2_X1 port map( A1 => n197, A2 => n240, ZN => n196);
   U45 : XNOR2_X1 port map( A => n223, B => B(30), ZN => DIFF_30_port);
   U46 : NOR2_X1 port map( A1 => n230, A2 => B(29), ZN => n223);
   U47 : OR3_X1 port map( A1 => B(29), A2 => B(30), A3 => n230, ZN => n228);
   U48 : XNOR2_X1 port map( A => B(56), B => n203, ZN => DIFF_56_port);
   U49 : NOR2_X1 port map( A1 => B(55), A2 => n202, ZN => n203);
   U50 : OR3_X1 port map( A1 => B(55), A2 => B(56), A3 => n202, ZN => n200);
   U51 : XNOR2_X1 port map( A => n227, B => B(63), ZN => DIFF_63_port);
   U52 : NOR2_X1 port map( A1 => n196, A2 => B(62), ZN => n227);
   U53 : XNOR2_X1 port map( A => B(28), B => n234, ZN => DIFF_28_port);
   U54 : NOR2_X1 port map( A1 => B(27), A2 => n233, ZN => n234);
   U55 : OR3_X1 port map( A1 => B(27), A2 => B(28), A3 => n233, ZN => n230);
   U56 : XNOR2_X1 port map( A => n231, B => B(26), ZN => DIFF_26_port);
   U57 : NOR2_X1 port map( A1 => n235, A2 => B(25), ZN => n231);
   U58 : OR3_X1 port map( A1 => B(25), A2 => B(26), A3 => n235, ZN => n233);
   U59 : XNOR2_X1 port map( A => B(24), B => n238, ZN => DIFF_24_port);
   U60 : NOR2_X1 port map( A1 => B(23), A2 => n237, ZN => n238);
   U61 : OR3_X1 port map( A1 => B(23), A2 => B(24), A3 => n237, ZN => n235);
   U62 : XNOR2_X1 port map( A => n236, B => B(22), ZN => DIFF_22_port);
   U63 : NOR2_X1 port map( A1 => n239, A2 => B(21), ZN => n236);
   U64 : OR3_X1 port map( A1 => B(21), A2 => B(22), A3 => n239, ZN => n237);
   U65 : NOR2_X1 port map( A1 => B(19), A2 => n241, ZN => n242);
   U66 : NOR2_X1 port map( A1 => B(15), A2 => n245, ZN => n246);
   U67 : NOR2_X1 port map( A1 => B(11), A2 => n249, ZN => n250);
   U68 : NOR2_X1 port map( A1 => B(7), A2 => n192, ZN => n191);
   U69 : NOR2_X1 port map( A1 => B(3), A2 => n211, ZN => n210);
   U70 : OR3_X1 port map( A1 => B(17), A2 => B(18), A3 => n243, ZN => n241);
   U71 : OR3_X1 port map( A1 => B(13), A2 => B(14), A3 => n247, ZN => n245);
   U72 : OR3_X1 port map( A1 => B(10), A2 => B(9), A3 => n190, ZN => n249);
   U73 : OR3_X1 port map( A1 => B(5), A2 => B(6), A3 => n194, ZN => n192);
   U74 : OR3_X1 port map( A1 => B(19), A2 => B(20), A3 => n241, ZN => n239);
   U75 : OR3_X1 port map( A1 => B(15), A2 => B(16), A3 => n245, ZN => n243);
   U76 : OR3_X1 port map( A1 => B(11), A2 => B(12), A3 => n249, ZN => n247);
   U77 : OR3_X1 port map( A1 => B(7), A2 => B(8), A3 => n192, ZN => n190);
   U78 : OR3_X1 port map( A1 => B(3), A2 => B(4), A3 => n211, ZN => n194);
   U79 : XNOR2_X1 port map( A => B(20), B => n242, ZN => DIFF_20_port);
   U80 : XNOR2_X1 port map( A => B(16), B => n246, ZN => DIFF_16_port);
   U84 : XNOR2_X1 port map( A => B(12), B => n250, ZN => DIFF_12_port);
   U88 : XNOR2_X1 port map( A => B(8), B => n191, ZN => DIFF_8_port);
   U91 : XNOR2_X1 port map( A => B(4), B => n210, ZN => DIFF_4_port);
   U94 : XNOR2_X1 port map( A => B(2), B => n232, ZN => DIFF_2_port);
   U97 : OR2_X1 port map( A1 => n243, A2 => B(17), ZN => n244);
   U100 : OR2_X1 port map( A1 => n247, A2 => B(13), ZN => n248);
   U104 : OR2_X1 port map( A1 => n190, A2 => B(9), ZN => n251);
   U107 : OR2_X1 port map( A1 => n194, A2 => B(5), ZN => n193);
   U110 : OR3_X1 port map( A1 => B(1), A2 => B(2), A3 => B(0), ZN => n211);
   U113 : NOR2_X1 port map( A1 => B(0), A2 => B(1), ZN => n232);
   U116 : INV_X1 port map( A => B(61), ZN => n240);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_11_DW01_sub_0 is

   port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (63 downto 0);  CO : out std_logic);

end complementer_N64_11_DW01_sub_0;

architecture SYN_rpl of complementer_N64_11_DW01_sub_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal DIFF_62_port, DIFF_63_port, DIFF_21_port, DIFF_22_port, DIFF_23_port,
      DIFF_24_port, DIFF_25_port, DIFF_26_port, DIFF_27_port, DIFF_28_port, 
      DIFF_29_port, DIFF_30_port, DIFF_31_port, DIFF_32_port, DIFF_33_port, 
      DIFF_34_port, DIFF_35_port, DIFF_36_port, DIFF_37_port, DIFF_38_port, 
      DIFF_39_port, DIFF_40_port, DIFF_41_port, DIFF_42_port, DIFF_43_port, 
      DIFF_44_port, DIFF_45_port, DIFF_46_port, DIFF_47_port, DIFF_48_port, 
      DIFF_49_port, DIFF_50_port, DIFF_51_port, DIFF_52_port, DIFF_53_port, 
      DIFF_54_port, DIFF_55_port, DIFF_56_port, DIFF_57_port, DIFF_58_port, 
      DIFF_59_port, DIFF_60_port, DIFF_61_port, DIFF_3_port, DIFF_4_port, 
      DIFF_5_port, DIFF_6_port, DIFF_7_port, DIFF_8_port, DIFF_9_port, 
      DIFF_10_port, DIFF_11_port, DIFF_12_port, DIFF_13_port, DIFF_14_port, 
      DIFF_15_port, DIFF_16_port, DIFF_17_port, DIFF_18_port, DIFF_19_port, 
      DIFF_20_port, DIFF_2_port, DIFF_1_port, n190, n191, n192, n194, n195, 
      n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, 
      n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, 
      n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, 
      n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, 
      n245, n246, n247, n249, n250, n189, n193, n244, n248, n251 : std_logic;

begin
   DIFF <= ( DIFF_63_port, DIFF_62_port, DIFF_61_port, DIFF_60_port, 
      DIFF_59_port, DIFF_58_port, DIFF_57_port, DIFF_56_port, DIFF_55_port, 
      DIFF_54_port, DIFF_53_port, DIFF_52_port, DIFF_51_port, DIFF_50_port, 
      DIFF_49_port, DIFF_48_port, DIFF_47_port, DIFF_46_port, DIFF_45_port, 
      DIFF_44_port, DIFF_43_port, DIFF_42_port, DIFF_41_port, DIFF_40_port, 
      DIFF_39_port, DIFF_38_port, DIFF_37_port, DIFF_36_port, DIFF_35_port, 
      DIFF_34_port, DIFF_33_port, DIFF_32_port, DIFF_31_port, DIFF_30_port, 
      DIFF_29_port, DIFF_28_port, DIFF_27_port, DIFF_26_port, DIFF_25_port, 
      DIFF_24_port, DIFF_23_port, DIFF_22_port, DIFF_21_port, DIFF_20_port, 
      DIFF_19_port, DIFF_18_port, DIFF_17_port, DIFF_16_port, DIFF_15_port, 
      DIFF_14_port, DIFF_13_port, DIFF_12_port, DIFF_11_port, DIFF_10_port, 
      DIFF_9_port, DIFF_8_port, DIFF_7_port, DIFF_6_port, DIFF_5_port, 
      DIFF_4_port, DIFF_3_port, DIFF_2_port, DIFF_1_port, B(0) );
   
   U81 : XOR2_X1 port map( A => n190, B => B(9), Z => DIFF_9_port);
   U82 : XOR2_X1 port map( A => n192, B => B(7), Z => DIFF_7_port);
   U84 : XOR2_X1 port map( A => n195, B => B(63), Z => DIFF_63_port);
   U85 : XOR2_X1 port map( A => n196, B => B(62), Z => DIFF_62_port);
   U86 : XOR2_X1 port map( A => n194, B => B(5), Z => DIFF_5_port);
   U87 : XOR2_X1 port map( A => n198, B => B(59), Z => DIFF_59_port);
   U88 : XOR2_X1 port map( A => n201, B => B(58), Z => DIFF_58_port);
   U89 : XOR2_X1 port map( A => n200, B => B(57), Z => DIFF_57_port);
   U90 : XOR2_X1 port map( A => n202, B => B(55), Z => DIFF_55_port);
   U91 : XOR2_X1 port map( A => n205, B => B(54), Z => DIFF_54_port);
   U92 : XOR2_X1 port map( A => n204, B => B(53), Z => DIFF_53_port);
   U93 : XOR2_X1 port map( A => n206, B => B(51), Z => DIFF_51_port);
   U94 : XOR2_X1 port map( A => n209, B => B(50), Z => DIFF_50_port);
   U95 : XOR2_X1 port map( A => n208, B => B(49), Z => DIFF_49_port);
   U96 : XOR2_X1 port map( A => n212, B => B(47), Z => DIFF_47_port);
   U97 : XOR2_X1 port map( A => n215, B => B(46), Z => DIFF_46_port);
   U98 : XOR2_X1 port map( A => n214, B => B(45), Z => DIFF_45_port);
   U99 : XOR2_X1 port map( A => n216, B => B(43), Z => DIFF_43_port);
   U100 : XOR2_X1 port map( A => n219, B => B(42), Z => DIFF_42_port);
   U101 : XOR2_X1 port map( A => n218, B => B(41), Z => DIFF_41_port);
   U102 : XOR2_X1 port map( A => n211, B => B(3), Z => DIFF_3_port);
   U103 : XOR2_X1 port map( A => n220, B => B(39), Z => DIFF_39_port);
   U104 : XOR2_X1 port map( A => n223, B => B(38), Z => DIFF_38_port);
   U105 : XOR2_X1 port map( A => n222, B => B(37), Z => DIFF_37_port);
   U106 : XOR2_X1 port map( A => n224, B => B(35), Z => DIFF_35_port);
   U107 : XOR2_X1 port map( A => n227, B => B(34), Z => DIFF_34_port);
   U108 : XOR2_X1 port map( A => n226, B => B(33), Z => DIFF_33_port);
   U109 : XOR2_X1 port map( A => n228, B => B(31), Z => DIFF_31_port);
   U110 : XOR2_X1 port map( A => n231, B => B(30), Z => DIFF_30_port);
   U111 : XOR2_X1 port map( A => n230, B => B(29), Z => DIFF_29_port);
   U112 : XOR2_X1 port map( A => n233, B => B(27), Z => DIFF_27_port);
   U113 : XOR2_X1 port map( A => n236, B => B(26), Z => DIFF_26_port);
   U114 : XOR2_X1 port map( A => n235, B => B(25), Z => DIFF_25_port);
   U115 : XOR2_X1 port map( A => n237, B => B(23), Z => DIFF_23_port);
   U116 : XOR2_X1 port map( A => n240, B => B(22), Z => DIFF_22_port);
   U117 : XOR2_X1 port map( A => n239, B => B(21), Z => DIFF_21_port);
   U118 : XOR2_X1 port map( A => B(1), B => B(0), Z => DIFF_1_port);
   U119 : XOR2_X1 port map( A => n241, B => B(19), Z => DIFF_19_port);
   U121 : XOR2_X1 port map( A => n243, B => B(17), Z => DIFF_17_port);
   U122 : XOR2_X1 port map( A => n245, B => B(15), Z => DIFF_15_port);
   U124 : XOR2_X1 port map( A => n247, B => B(13), Z => DIFF_13_port);
   U125 : XOR2_X1 port map( A => n249, B => B(11), Z => DIFF_11_port);
   U1 : NOR2_X1 port map( A1 => B(51), A2 => n206, ZN => n207);
   U2 : NOR2_X1 port map( A1 => B(59), A2 => n198, ZN => n199);
   U3 : OR3_X1 port map( A1 => B(51), A2 => B(52), A3 => n206, ZN => n204);
   U4 : OR2_X1 port map( A1 => n204, A2 => B(53), ZN => n205);
   U5 : NAND2_X1 port map( A1 => n197, A2 => n251, ZN => n196);
   U6 : NOR2_X1 port map( A1 => B(31), A2 => n228, ZN => n229);
   U7 : NOR2_X1 port map( A1 => B(27), A2 => n233, ZN => n234);
   U8 : OR3_X1 port map( A1 => B(29), A2 => B(30), A3 => n230, ZN => n228);
   U9 : OR3_X1 port map( A1 => B(31), A2 => B(32), A3 => n228, ZN => n226);
   U10 : OR3_X1 port map( A1 => B(27), A2 => B(28), A3 => n233, ZN => n230);
   U11 : OR2_X1 port map( A1 => n230, A2 => B(29), ZN => n231);
   U12 : NOR2_X1 port map( A1 => B(47), A2 => n212, ZN => n213);
   U13 : NOR2_X1 port map( A1 => B(43), A2 => n216, ZN => n217);
   U14 : NOR2_X1 port map( A1 => B(39), A2 => n220, ZN => n221);
   U15 : NOR2_X1 port map( A1 => B(35), A2 => n224, ZN => n225);
   U16 : NOR2_X1 port map( A1 => B(55), A2 => n202, ZN => n203);
   U17 : OR3_X1 port map( A1 => B(57), A2 => B(58), A3 => n200, ZN => n198);
   U18 : OR3_X1 port map( A1 => B(49), A2 => B(50), A3 => n208, ZN => n206);
   U19 : OR3_X1 port map( A1 => B(45), A2 => B(46), A3 => n214, ZN => n212);
   U20 : OR3_X1 port map( A1 => B(41), A2 => B(42), A3 => n218, ZN => n216);
   U21 : OR3_X1 port map( A1 => B(37), A2 => B(38), A3 => n222, ZN => n220);
   U22 : OR3_X1 port map( A1 => B(33), A2 => B(34), A3 => n226, ZN => n224);
   U23 : OR3_X1 port map( A1 => B(53), A2 => B(54), A3 => n204, ZN => n202);
   U24 : OR3_X1 port map( A1 => B(47), A2 => B(48), A3 => n212, ZN => n208);
   U25 : OR3_X1 port map( A1 => B(43), A2 => B(44), A3 => n216, ZN => n214);
   U26 : OR3_X1 port map( A1 => B(39), A2 => B(40), A3 => n220, ZN => n218);
   U27 : OR3_X1 port map( A1 => B(35), A2 => B(36), A3 => n224, ZN => n222);
   U28 : OR3_X1 port map( A1 => B(55), A2 => B(56), A3 => n202, ZN => n200);
   U29 : OR2_X1 port map( A1 => n208, A2 => B(49), ZN => n209);
   U30 : OR2_X1 port map( A1 => n214, A2 => B(45), ZN => n215);
   U31 : OR2_X1 port map( A1 => n218, A2 => B(41), ZN => n219);
   U32 : OR2_X1 port map( A1 => n222, A2 => B(37), ZN => n223);
   U33 : OR2_X1 port map( A1 => n226, A2 => B(33), ZN => n227);
   U34 : OR2_X1 port map( A1 => n200, A2 => B(57), ZN => n201);
   U35 : NOR3_X1 port map( A1 => B(59), A2 => B(60), A3 => n198, ZN => n197);
   U36 : OR2_X1 port map( A1 => n196, A2 => B(62), ZN => n195);
   U37 : OR3_X1 port map( A1 => B(25), A2 => B(26), A3 => n235, ZN => n233);
   U38 : XNOR2_X1 port map( A => B(36), B => n225, ZN => DIFF_36_port);
   U39 : XNOR2_X1 port map( A => B(32), B => n229, ZN => DIFF_32_port);
   U40 : XNOR2_X1 port map( A => B(28), B => n234, ZN => DIFF_28_port);
   U41 : XNOR2_X1 port map( A => B(24), B => n238, ZN => DIFF_24_port);
   U42 : OR2_X1 port map( A1 => n235, A2 => B(25), ZN => n236);
   U43 : XNOR2_X1 port map( A => n197, B => B(61), ZN => DIFF_61_port);
   U44 : XNOR2_X1 port map( A => B(60), B => n199, ZN => DIFF_60_port);
   U45 : XNOR2_X1 port map( A => B(56), B => n203, ZN => DIFF_56_port);
   U46 : XNOR2_X1 port map( A => B(52), B => n207, ZN => DIFF_52_port);
   U47 : XNOR2_X1 port map( A => B(48), B => n213, ZN => DIFF_48_port);
   U48 : XNOR2_X1 port map( A => B(44), B => n217, ZN => DIFF_44_port);
   U49 : XNOR2_X1 port map( A => B(40), B => n221, ZN => DIFF_40_port);
   U50 : NOR2_X1 port map( A1 => B(23), A2 => n237, ZN => n238);
   U51 : OR3_X1 port map( A1 => B(23), A2 => B(24), A3 => n237, ZN => n235);
   U52 : OR3_X1 port map( A1 => B(21), A2 => B(22), A3 => n239, ZN => n237);
   U53 : OR2_X1 port map( A1 => n239, A2 => B(21), ZN => n240);
   U54 : XNOR2_X1 port map( A => B(20), B => n242, ZN => DIFF_20_port);
   U55 : XNOR2_X1 port map( A => n189, B => B(18), ZN => DIFF_18_port);
   U56 : NOR2_X1 port map( A1 => n243, A2 => B(17), ZN => n189);
   U57 : XNOR2_X1 port map( A => n193, B => B(14), ZN => DIFF_14_port);
   U58 : NOR2_X1 port map( A1 => n247, A2 => B(13), ZN => n193);
   U59 : XNOR2_X1 port map( A => n244, B => B(10), ZN => DIFF_10_port);
   U60 : NOR2_X1 port map( A1 => n190, A2 => B(9), ZN => n244);
   U61 : XNOR2_X1 port map( A => n248, B => B(6), ZN => DIFF_6_port);
   U62 : NOR2_X1 port map( A1 => n194, A2 => B(5), ZN => n248);
   U63 : NOR2_X1 port map( A1 => B(19), A2 => n241, ZN => n242);
   U64 : XNOR2_X1 port map( A => B(16), B => n246, ZN => DIFF_16_port);
   U65 : NOR2_X1 port map( A1 => B(15), A2 => n245, ZN => n246);
   U66 : XNOR2_X1 port map( A => B(12), B => n250, ZN => DIFF_12_port);
   U67 : NOR2_X1 port map( A1 => B(11), A2 => n249, ZN => n250);
   U68 : XNOR2_X1 port map( A => B(8), B => n191, ZN => DIFF_8_port);
   U69 : NOR2_X1 port map( A1 => B(7), A2 => n192, ZN => n191);
   U70 : XNOR2_X1 port map( A => B(2), B => n232, ZN => DIFF_2_port);
   U71 : NOR2_X1 port map( A1 => B(0), A2 => B(1), ZN => n232);
   U72 : XNOR2_X1 port map( A => B(4), B => n210, ZN => DIFF_4_port);
   U73 : NOR2_X1 port map( A1 => B(3), A2 => n211, ZN => n210);
   U74 : OR3_X1 port map( A1 => B(5), A2 => B(6), A3 => n194, ZN => n192);
   U75 : OR3_X1 port map( A1 => B(10), A2 => B(9), A3 => n190, ZN => n249);
   U76 : OR3_X1 port map( A1 => B(13), A2 => B(14), A3 => n247, ZN => n245);
   U77 : OR3_X1 port map( A1 => B(17), A2 => B(18), A3 => n243, ZN => n241);
   U78 : OR3_X1 port map( A1 => B(7), A2 => B(8), A3 => n192, ZN => n190);
   U79 : OR3_X1 port map( A1 => B(11), A2 => B(12), A3 => n249, ZN => n247);
   U80 : OR3_X1 port map( A1 => B(15), A2 => B(16), A3 => n245, ZN => n243);
   U83 : OR3_X1 port map( A1 => B(19), A2 => B(20), A3 => n241, ZN => n239);
   U120 : OR3_X1 port map( A1 => B(3), A2 => B(4), A3 => n211, ZN => n194);
   U123 : OR3_X1 port map( A1 => B(1), A2 => B(2), A3 => B(0), ZN => n211);
   U126 : INV_X1 port map( A => B(61), ZN => n251);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_12_DW01_sub_0 is

   port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (63 downto 0);  CO : out std_logic);

end complementer_N64_12_DW01_sub_0;

architecture SYN_rpl of complementer_N64_12_DW01_sub_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal DIFF_62_port, DIFF_61_port, DIFF_60_port, DIFF_59_port, DIFF_58_port,
      DIFF_57_port, DIFF_56_port, DIFF_55_port, DIFF_54_port, DIFF_53_port, 
      DIFF_52_port, DIFF_51_port, DIFF_50_port, DIFF_49_port, DIFF_48_port, 
      DIFF_47_port, DIFF_46_port, DIFF_45_port, DIFF_44_port, DIFF_43_port, 
      DIFF_42_port, DIFF_41_port, DIFF_40_port, DIFF_39_port, DIFF_38_port, 
      DIFF_37_port, DIFF_36_port, DIFF_35_port, DIFF_34_port, DIFF_33_port, 
      DIFF_32_port, DIFF_31_port, DIFF_30_port, DIFF_29_port, DIFF_28_port, 
      DIFF_27_port, DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, 
      DIFF_22_port, DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, 
      DIFF_17_port, DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, 
      DIFF_12_port, DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, 
      DIFF_7_port, DIFF_6_port, DIFF_5_port, DIFF_4_port, DIFF_3_port, 
      DIFF_2_port, DIFF_1_port, DIFF_63_port, n190, n191, n192, n193, n194, 
      n196, n197, n198, n199, n200, n202, n203, n204, n206, n207, n208, n210, 
      n211, n212, n213, n214, n216, n217, n218, n220, n221, n222, n224, n225, 
      n226, n228, n229, n230, n232, n233, n234, n235, n237, n238, n239, n241, 
      n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n189, n195, 
      n201, n205, n209, n215, n219, n223, n227, n231, n236, n240 : std_logic;

begin
   DIFF <= ( DIFF_63_port, DIFF_62_port, DIFF_61_port, DIFF_60_port, 
      DIFF_59_port, DIFF_58_port, DIFF_57_port, DIFF_56_port, DIFF_55_port, 
      DIFF_54_port, DIFF_53_port, DIFF_52_port, DIFF_51_port, DIFF_50_port, 
      DIFF_49_port, DIFF_48_port, DIFF_47_port, DIFF_46_port, DIFF_45_port, 
      DIFF_44_port, DIFF_43_port, DIFF_42_port, DIFF_41_port, DIFF_40_port, 
      DIFF_39_port, DIFF_38_port, DIFF_37_port, DIFF_36_port, DIFF_35_port, 
      DIFF_34_port, DIFF_33_port, DIFF_32_port, DIFF_31_port, DIFF_30_port, 
      DIFF_29_port, DIFF_28_port, DIFF_27_port, DIFF_26_port, DIFF_25_port, 
      DIFF_24_port, DIFF_23_port, DIFF_22_port, DIFF_21_port, DIFF_20_port, 
      DIFF_19_port, DIFF_18_port, DIFF_17_port, DIFF_16_port, DIFF_15_port, 
      DIFF_14_port, DIFF_13_port, DIFF_12_port, DIFF_11_port, DIFF_10_port, 
      DIFF_9_port, DIFF_8_port, DIFF_7_port, DIFF_6_port, DIFF_5_port, 
      DIFF_4_port, DIFF_3_port, DIFF_2_port, DIFF_1_port, B(0) );
   
   U81 : XOR2_X1 port map( A => n190, B => B(9), Z => DIFF_9_port);
   U82 : XOR2_X1 port map( A => n192, B => B(7), Z => DIFF_7_port);
   U83 : XOR2_X1 port map( A => n193, B => B(6), Z => DIFF_6_port);
   U85 : XOR2_X1 port map( A => n196, B => B(62), Z => DIFF_62_port);
   U86 : XOR2_X1 port map( A => n194, B => B(5), Z => DIFF_5_port);
   U87 : XOR2_X1 port map( A => n198, B => B(59), Z => DIFF_59_port);
   U89 : XOR2_X1 port map( A => n200, B => B(57), Z => DIFF_57_port);
   U90 : XOR2_X1 port map( A => n202, B => B(55), Z => DIFF_55_port);
   U92 : XOR2_X1 port map( A => n204, B => B(53), Z => DIFF_53_port);
   U93 : XOR2_X1 port map( A => n206, B => B(51), Z => DIFF_51_port);
   U95 : XOR2_X1 port map( A => n208, B => B(49), Z => DIFF_49_port);
   U96 : XOR2_X1 port map( A => n212, B => B(47), Z => DIFF_47_port);
   U98 : XOR2_X1 port map( A => n214, B => B(45), Z => DIFF_45_port);
   U99 : XOR2_X1 port map( A => n216, B => B(43), Z => DIFF_43_port);
   U101 : XOR2_X1 port map( A => n218, B => B(41), Z => DIFF_41_port);
   U102 : XOR2_X1 port map( A => n211, B => B(3), Z => DIFF_3_port);
   U103 : XOR2_X1 port map( A => n220, B => B(39), Z => DIFF_39_port);
   U105 : XOR2_X1 port map( A => n222, B => B(37), Z => DIFF_37_port);
   U106 : XOR2_X1 port map( A => n224, B => B(35), Z => DIFF_35_port);
   U108 : XOR2_X1 port map( A => n226, B => B(33), Z => DIFF_33_port);
   U109 : XOR2_X1 port map( A => n228, B => B(31), Z => DIFF_31_port);
   U111 : XOR2_X1 port map( A => n230, B => B(29), Z => DIFF_29_port);
   U112 : XOR2_X1 port map( A => n233, B => B(27), Z => DIFF_27_port);
   U114 : XOR2_X1 port map( A => n235, B => B(25), Z => DIFF_25_port);
   U115 : XOR2_X1 port map( A => n237, B => B(23), Z => DIFF_23_port);
   U117 : XOR2_X1 port map( A => n239, B => B(21), Z => DIFF_21_port);
   U118 : XOR2_X1 port map( A => B(1), B => B(0), Z => DIFF_1_port);
   U119 : XOR2_X1 port map( A => n241, B => B(19), Z => DIFF_19_port);
   U120 : XOR2_X1 port map( A => n244, B => B(18), Z => DIFF_18_port);
   U121 : XOR2_X1 port map( A => n243, B => B(17), Z => DIFF_17_port);
   U122 : XOR2_X1 port map( A => n245, B => B(15), Z => DIFF_15_port);
   U123 : XOR2_X1 port map( A => n248, B => B(14), Z => DIFF_14_port);
   U124 : XOR2_X1 port map( A => n247, B => B(13), Z => DIFF_13_port);
   U125 : XOR2_X1 port map( A => n249, B => B(11), Z => DIFF_11_port);
   U126 : XOR2_X1 port map( A => n251, B => B(10), Z => DIFF_10_port);
   U1 : XOR2_X1 port map( A => n197, B => n240, Z => DIFF_61_port);
   U2 : NAND2_X1 port map( A1 => n197, A2 => n240, ZN => n196);
   U3 : OR3_X1 port map( A1 => B(57), A2 => B(58), A3 => n200, ZN => n198);
   U4 : XNOR2_X1 port map( A => n189, B => B(58), ZN => DIFF_58_port);
   U5 : NOR2_X1 port map( A1 => n200, A2 => B(57), ZN => n189);
   U6 : XNOR2_X1 port map( A => B(36), B => n225, ZN => DIFF_36_port);
   U7 : NOR2_X1 port map( A1 => B(35), A2 => n224, ZN => n225);
   U8 : XNOR2_X1 port map( A => B(32), B => n229, ZN => DIFF_32_port);
   U9 : NOR2_X1 port map( A1 => B(31), A2 => n228, ZN => n229);
   U10 : XNOR2_X1 port map( A => B(28), B => n234, ZN => DIFF_28_port);
   U11 : NOR2_X1 port map( A1 => B(27), A2 => n233, ZN => n234);
   U12 : OR3_X1 port map( A1 => B(29), A2 => B(30), A3 => n230, ZN => n228);
   U13 : OR3_X1 port map( A1 => B(33), A2 => B(34), A3 => n226, ZN => n224);
   U14 : OR3_X1 port map( A1 => B(27), A2 => B(28), A3 => n233, ZN => n230);
   U15 : OR3_X1 port map( A1 => B(31), A2 => B(32), A3 => n228, ZN => n226);
   U16 : OR3_X1 port map( A1 => B(35), A2 => B(36), A3 => n224, ZN => n222);
   U17 : XNOR2_X1 port map( A => n195, B => B(34), ZN => DIFF_34_port);
   U18 : NOR2_X1 port map( A1 => n226, A2 => B(33), ZN => n195);
   U19 : XNOR2_X1 port map( A => n201, B => B(30), ZN => DIFF_30_port);
   U20 : NOR2_X1 port map( A1 => n230, A2 => B(29), ZN => n201);
   U21 : NOR3_X1 port map( A1 => B(59), A2 => B(60), A3 => n198, ZN => n197);
   U22 : XNOR2_X1 port map( A => n205, B => B(46), ZN => DIFF_46_port);
   U23 : NOR2_X1 port map( A1 => n214, A2 => B(45), ZN => n205);
   U24 : XNOR2_X1 port map( A => n209, B => B(42), ZN => DIFF_42_port);
   U25 : NOR2_X1 port map( A1 => n218, A2 => B(41), ZN => n209);
   U26 : XNOR2_X1 port map( A => n215, B => B(38), ZN => DIFF_38_port);
   U27 : NOR2_X1 port map( A1 => n222, A2 => B(37), ZN => n215);
   U28 : XNOR2_X1 port map( A => n219, B => B(50), ZN => DIFF_50_port);
   U29 : NOR2_X1 port map( A1 => n208, A2 => B(49), ZN => n219);
   U30 : XNOR2_X1 port map( A => n223, B => B(54), ZN => DIFF_54_port);
   U31 : NOR2_X1 port map( A1 => n204, A2 => B(53), ZN => n223);
   U32 : XNOR2_X1 port map( A => B(40), B => n221, ZN => DIFF_40_port);
   U33 : NOR2_X1 port map( A1 => B(39), A2 => n220, ZN => n221);
   U34 : XNOR2_X1 port map( A => B(48), B => n213, ZN => DIFF_48_port);
   U35 : NOR2_X1 port map( A1 => B(47), A2 => n212, ZN => n213);
   U36 : XNOR2_X1 port map( A => B(44), B => n217, ZN => DIFF_44_port);
   U37 : NOR2_X1 port map( A1 => B(43), A2 => n216, ZN => n217);
   U38 : XNOR2_X1 port map( A => B(52), B => n207, ZN => DIFF_52_port);
   U39 : NOR2_X1 port map( A1 => B(51), A2 => n206, ZN => n207);
   U40 : XNOR2_X1 port map( A => B(60), B => n199, ZN => DIFF_60_port);
   U41 : NOR2_X1 port map( A1 => B(59), A2 => n198, ZN => n199);
   U42 : XNOR2_X1 port map( A => B(56), B => n203, ZN => DIFF_56_port);
   U43 : NOR2_X1 port map( A1 => B(55), A2 => n202, ZN => n203);
   U44 : OR3_X1 port map( A1 => B(37), A2 => B(38), A3 => n222, ZN => n220);
   U45 : OR3_X1 port map( A1 => B(41), A2 => B(42), A3 => n218, ZN => n216);
   U46 : OR3_X1 port map( A1 => B(45), A2 => B(46), A3 => n214, ZN => n212);
   U47 : OR3_X1 port map( A1 => B(53), A2 => B(54), A3 => n204, ZN => n202);
   U48 : OR3_X1 port map( A1 => B(49), A2 => B(50), A3 => n208, ZN => n206);
   U49 : OR3_X1 port map( A1 => B(51), A2 => B(52), A3 => n206, ZN => n204);
   U50 : OR3_X1 port map( A1 => B(39), A2 => B(40), A3 => n220, ZN => n218);
   U51 : OR3_X1 port map( A1 => B(43), A2 => B(44), A3 => n216, ZN => n214);
   U52 : OR3_X1 port map( A1 => B(47), A2 => B(48), A3 => n212, ZN => n208);
   U53 : OR3_X1 port map( A1 => B(55), A2 => B(56), A3 => n202, ZN => n200);
   U54 : OR3_X1 port map( A1 => B(25), A2 => B(26), A3 => n235, ZN => n233);
   U55 : XNOR2_X1 port map( A => n227, B => B(26), ZN => DIFF_26_port);
   U56 : NOR2_X1 port map( A1 => n235, A2 => B(25), ZN => n227);
   U57 : XNOR2_X1 port map( A => n231, B => B(63), ZN => DIFF_63_port);
   U58 : NOR2_X1 port map( A1 => n196, A2 => B(62), ZN => n231);
   U59 : XNOR2_X1 port map( A => B(24), B => n238, ZN => DIFF_24_port);
   U60 : NOR2_X1 port map( A1 => B(23), A2 => n237, ZN => n238);
   U61 : OR3_X1 port map( A1 => B(23), A2 => B(24), A3 => n237, ZN => n235);
   U62 : XNOR2_X1 port map( A => n236, B => B(22), ZN => DIFF_22_port);
   U63 : NOR2_X1 port map( A1 => n239, A2 => B(21), ZN => n236);
   U64 : OR3_X1 port map( A1 => B(21), A2 => B(22), A3 => n239, ZN => n237);
   U65 : OR3_X1 port map( A1 => B(19), A2 => B(20), A3 => n241, ZN => n239);
   U66 : XNOR2_X1 port map( A => B(20), B => n242, ZN => DIFF_20_port);
   U67 : NOR2_X1 port map( A1 => B(19), A2 => n241, ZN => n242);
   U68 : NOR2_X1 port map( A1 => B(15), A2 => n245, ZN => n246);
   U69 : NOR2_X1 port map( A1 => B(11), A2 => n249, ZN => n250);
   U70 : NOR2_X1 port map( A1 => B(7), A2 => n192, ZN => n191);
   U71 : NOR2_X1 port map( A1 => B(3), A2 => n211, ZN => n210);
   U72 : OR3_X1 port map( A1 => B(17), A2 => B(18), A3 => n243, ZN => n241);
   U73 : OR3_X1 port map( A1 => B(13), A2 => B(14), A3 => n247, ZN => n245);
   U74 : OR3_X1 port map( A1 => B(10), A2 => B(9), A3 => n190, ZN => n249);
   U75 : OR3_X1 port map( A1 => B(5), A2 => B(6), A3 => n194, ZN => n192);
   U76 : OR3_X1 port map( A1 => B(15), A2 => B(16), A3 => n245, ZN => n243);
   U77 : OR3_X1 port map( A1 => B(11), A2 => B(12), A3 => n249, ZN => n247);
   U78 : OR3_X1 port map( A1 => B(7), A2 => B(8), A3 => n192, ZN => n190);
   U79 : OR3_X1 port map( A1 => B(3), A2 => B(4), A3 => n211, ZN => n194);
   U80 : XNOR2_X1 port map( A => B(16), B => n246, ZN => DIFF_16_port);
   U84 : XNOR2_X1 port map( A => B(12), B => n250, ZN => DIFF_12_port);
   U88 : XNOR2_X1 port map( A => B(8), B => n191, ZN => DIFF_8_port);
   U91 : XNOR2_X1 port map( A => B(4), B => n210, ZN => DIFF_4_port);
   U94 : XNOR2_X1 port map( A => B(2), B => n232, ZN => DIFF_2_port);
   U97 : OR2_X1 port map( A1 => n243, A2 => B(17), ZN => n244);
   U100 : OR2_X1 port map( A1 => n247, A2 => B(13), ZN => n248);
   U104 : OR2_X1 port map( A1 => n190, A2 => B(9), ZN => n251);
   U107 : OR2_X1 port map( A1 => n194, A2 => B(5), ZN => n193);
   U110 : OR3_X1 port map( A1 => B(1), A2 => B(2), A3 => B(0), ZN => n211);
   U113 : NOR2_X1 port map( A1 => B(0), A2 => B(1), ZN => n232);
   U116 : INV_X1 port map( A => B(61), ZN => n240);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_13_DW01_sub_0 is

   port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (63 downto 0);  CO : out std_logic);

end complementer_N64_13_DW01_sub_0;

architecture SYN_rpl of complementer_N64_13_DW01_sub_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal DIFF_62_port, DIFF_63_port, DIFF_19_port, DIFF_20_port, DIFF_21_port,
      DIFF_22_port, DIFF_23_port, DIFF_24_port, DIFF_25_port, DIFF_26_port, 
      DIFF_27_port, DIFF_28_port, DIFF_29_port, DIFF_30_port, DIFF_31_port, 
      DIFF_32_port, DIFF_33_port, DIFF_34_port, DIFF_35_port, DIFF_36_port, 
      DIFF_37_port, DIFF_38_port, DIFF_39_port, DIFF_40_port, DIFF_41_port, 
      DIFF_42_port, DIFF_43_port, DIFF_44_port, DIFF_45_port, DIFF_46_port, 
      DIFF_47_port, DIFF_48_port, DIFF_49_port, DIFF_50_port, DIFF_51_port, 
      DIFF_52_port, DIFF_53_port, DIFF_54_port, DIFF_55_port, DIFF_56_port, 
      DIFF_57_port, DIFF_58_port, DIFF_59_port, DIFF_60_port, DIFF_61_port, 
      DIFF_3_port, DIFF_4_port, DIFF_5_port, DIFF_6_port, DIFF_7_port, 
      DIFF_8_port, DIFF_9_port, DIFF_10_port, DIFF_11_port, DIFF_12_port, 
      DIFF_13_port, DIFF_14_port, DIFF_15_port, DIFF_16_port, DIFF_17_port, 
      DIFF_18_port, DIFF_2_port, DIFF_1_port, n190, n191, n192, n194, n195, 
      n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, 
      n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, 
      n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, 
      n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, 
      n244, n245, n246, n247, n249, n250, n189, n193, n248, n251 : std_logic;

begin
   DIFF <= ( DIFF_63_port, DIFF_62_port, DIFF_61_port, DIFF_60_port, 
      DIFF_59_port, DIFF_58_port, DIFF_57_port, DIFF_56_port, DIFF_55_port, 
      DIFF_54_port, DIFF_53_port, DIFF_52_port, DIFF_51_port, DIFF_50_port, 
      DIFF_49_port, DIFF_48_port, DIFF_47_port, DIFF_46_port, DIFF_45_port, 
      DIFF_44_port, DIFF_43_port, DIFF_42_port, DIFF_41_port, DIFF_40_port, 
      DIFF_39_port, DIFF_38_port, DIFF_37_port, DIFF_36_port, DIFF_35_port, 
      DIFF_34_port, DIFF_33_port, DIFF_32_port, DIFF_31_port, DIFF_30_port, 
      DIFF_29_port, DIFF_28_port, DIFF_27_port, DIFF_26_port, DIFF_25_port, 
      DIFF_24_port, DIFF_23_port, DIFF_22_port, DIFF_21_port, DIFF_20_port, 
      DIFF_19_port, DIFF_18_port, DIFF_17_port, DIFF_16_port, DIFF_15_port, 
      DIFF_14_port, DIFF_13_port, DIFF_12_port, DIFF_11_port, DIFF_10_port, 
      DIFF_9_port, DIFF_8_port, DIFF_7_port, DIFF_6_port, DIFF_5_port, 
      DIFF_4_port, DIFF_3_port, DIFF_2_port, DIFF_1_port, B(0) );
   
   U81 : XOR2_X1 port map( A => n190, B => B(9), Z => DIFF_9_port);
   U82 : XOR2_X1 port map( A => n192, B => B(7), Z => DIFF_7_port);
   U84 : XOR2_X1 port map( A => n195, B => B(63), Z => DIFF_63_port);
   U85 : XOR2_X1 port map( A => n196, B => B(62), Z => DIFF_62_port);
   U86 : XOR2_X1 port map( A => n194, B => B(5), Z => DIFF_5_port);
   U87 : XOR2_X1 port map( A => n198, B => B(59), Z => DIFF_59_port);
   U88 : XOR2_X1 port map( A => n201, B => B(58), Z => DIFF_58_port);
   U89 : XOR2_X1 port map( A => n200, B => B(57), Z => DIFF_57_port);
   U90 : XOR2_X1 port map( A => n202, B => B(55), Z => DIFF_55_port);
   U91 : XOR2_X1 port map( A => n205, B => B(54), Z => DIFF_54_port);
   U92 : XOR2_X1 port map( A => n204, B => B(53), Z => DIFF_53_port);
   U93 : XOR2_X1 port map( A => n206, B => B(51), Z => DIFF_51_port);
   U94 : XOR2_X1 port map( A => n209, B => B(50), Z => DIFF_50_port);
   U95 : XOR2_X1 port map( A => n208, B => B(49), Z => DIFF_49_port);
   U96 : XOR2_X1 port map( A => n212, B => B(47), Z => DIFF_47_port);
   U97 : XOR2_X1 port map( A => n215, B => B(46), Z => DIFF_46_port);
   U98 : XOR2_X1 port map( A => n214, B => B(45), Z => DIFF_45_port);
   U99 : XOR2_X1 port map( A => n216, B => B(43), Z => DIFF_43_port);
   U100 : XOR2_X1 port map( A => n219, B => B(42), Z => DIFF_42_port);
   U101 : XOR2_X1 port map( A => n218, B => B(41), Z => DIFF_41_port);
   U102 : XOR2_X1 port map( A => n211, B => B(3), Z => DIFF_3_port);
   U103 : XOR2_X1 port map( A => n220, B => B(39), Z => DIFF_39_port);
   U104 : XOR2_X1 port map( A => n223, B => B(38), Z => DIFF_38_port);
   U105 : XOR2_X1 port map( A => n222, B => B(37), Z => DIFF_37_port);
   U106 : XOR2_X1 port map( A => n224, B => B(35), Z => DIFF_35_port);
   U107 : XOR2_X1 port map( A => n227, B => B(34), Z => DIFF_34_port);
   U108 : XOR2_X1 port map( A => n226, B => B(33), Z => DIFF_33_port);
   U109 : XOR2_X1 port map( A => n228, B => B(31), Z => DIFF_31_port);
   U110 : XOR2_X1 port map( A => n231, B => B(30), Z => DIFF_30_port);
   U111 : XOR2_X1 port map( A => n230, B => B(29), Z => DIFF_29_port);
   U112 : XOR2_X1 port map( A => n233, B => B(27), Z => DIFF_27_port);
   U113 : XOR2_X1 port map( A => n236, B => B(26), Z => DIFF_26_port);
   U114 : XOR2_X1 port map( A => n235, B => B(25), Z => DIFF_25_port);
   U115 : XOR2_X1 port map( A => n237, B => B(23), Z => DIFF_23_port);
   U116 : XOR2_X1 port map( A => n240, B => B(22), Z => DIFF_22_port);
   U117 : XOR2_X1 port map( A => n239, B => B(21), Z => DIFF_21_port);
   U118 : XOR2_X1 port map( A => B(1), B => B(0), Z => DIFF_1_port);
   U119 : XOR2_X1 port map( A => n241, B => B(19), Z => DIFF_19_port);
   U120 : XOR2_X1 port map( A => n244, B => B(18), Z => DIFF_18_port);
   U121 : XOR2_X1 port map( A => n243, B => B(17), Z => DIFF_17_port);
   U122 : XOR2_X1 port map( A => n245, B => B(15), Z => DIFF_15_port);
   U124 : XOR2_X1 port map( A => n247, B => B(13), Z => DIFF_13_port);
   U125 : XOR2_X1 port map( A => n249, B => B(11), Z => DIFF_11_port);
   U1 : NAND2_X1 port map( A1 => n197, A2 => n251, ZN => n196);
   U2 : NOR2_X1 port map( A1 => B(39), A2 => n220, ZN => n221);
   U3 : NOR2_X1 port map( A1 => B(35), A2 => n224, ZN => n225);
   U4 : NOR2_X1 port map( A1 => B(31), A2 => n228, ZN => n229);
   U5 : NOR2_X1 port map( A1 => B(27), A2 => n233, ZN => n234);
   U6 : OR3_X1 port map( A1 => B(37), A2 => B(38), A3 => n222, ZN => n220);
   U7 : OR3_X1 port map( A1 => B(33), A2 => B(34), A3 => n226, ZN => n224);
   U8 : OR3_X1 port map( A1 => B(29), A2 => B(30), A3 => n230, ZN => n228);
   U9 : OR3_X1 port map( A1 => B(25), A2 => B(26), A3 => n235, ZN => n233);
   U10 : OR3_X1 port map( A1 => B(39), A2 => B(40), A3 => n220, ZN => n218);
   U11 : OR3_X1 port map( A1 => B(35), A2 => B(36), A3 => n224, ZN => n222);
   U12 : OR3_X1 port map( A1 => B(31), A2 => B(32), A3 => n228, ZN => n226);
   U13 : OR3_X1 port map( A1 => B(27), A2 => B(28), A3 => n233, ZN => n230);
   U14 : OR2_X1 port map( A1 => n222, A2 => B(37), ZN => n223);
   U15 : OR2_X1 port map( A1 => n226, A2 => B(33), ZN => n227);
   U16 : OR2_X1 port map( A1 => n230, A2 => B(29), ZN => n231);
   U17 : OR2_X1 port map( A1 => n235, A2 => B(25), ZN => n236);
   U18 : NOR3_X1 port map( A1 => B(59), A2 => B(60), A3 => n198, ZN => n197);
   U19 : NOR2_X1 port map( A1 => B(47), A2 => n212, ZN => n213);
   U20 : NOR2_X1 port map( A1 => B(43), A2 => n216, ZN => n217);
   U21 : NOR2_X1 port map( A1 => B(51), A2 => n206, ZN => n207);
   U22 : NOR2_X1 port map( A1 => B(59), A2 => n198, ZN => n199);
   U23 : NOR2_X1 port map( A1 => B(55), A2 => n202, ZN => n203);
   U24 : OR3_X1 port map( A1 => B(57), A2 => B(58), A3 => n200, ZN => n198);
   U25 : OR3_X1 port map( A1 => B(45), A2 => B(46), A3 => n214, ZN => n212);
   U26 : OR3_X1 port map( A1 => B(41), A2 => B(42), A3 => n218, ZN => n216);
   U27 : OR3_X1 port map( A1 => B(49), A2 => B(50), A3 => n208, ZN => n206);
   U28 : OR3_X1 port map( A1 => B(53), A2 => B(54), A3 => n204, ZN => n202);
   U29 : OR3_X1 port map( A1 => B(47), A2 => B(48), A3 => n212, ZN => n208);
   U30 : OR3_X1 port map( A1 => B(43), A2 => B(44), A3 => n216, ZN => n214);
   U31 : OR3_X1 port map( A1 => B(51), A2 => B(52), A3 => n206, ZN => n204);
   U32 : OR3_X1 port map( A1 => B(55), A2 => B(56), A3 => n202, ZN => n200);
   U33 : OR2_X1 port map( A1 => n214, A2 => B(45), ZN => n215);
   U34 : OR2_X1 port map( A1 => n218, A2 => B(41), ZN => n219);
   U35 : OR2_X1 port map( A1 => n208, A2 => B(49), ZN => n209);
   U36 : OR2_X1 port map( A1 => n200, A2 => B(57), ZN => n201);
   U37 : OR2_X1 port map( A1 => n204, A2 => B(53), ZN => n205);
   U38 : NOR2_X1 port map( A1 => B(23), A2 => n237, ZN => n238);
   U39 : XNOR2_X1 port map( A => B(44), B => n217, ZN => DIFF_44_port);
   U40 : OR3_X1 port map( A1 => B(23), A2 => B(24), A3 => n237, ZN => n235);
   U41 : XNOR2_X1 port map( A => B(40), B => n221, ZN => DIFF_40_port);
   U42 : XNOR2_X1 port map( A => B(36), B => n225, ZN => DIFF_36_port);
   U43 : XNOR2_X1 port map( A => B(32), B => n229, ZN => DIFF_32_port);
   U44 : XNOR2_X1 port map( A => B(28), B => n234, ZN => DIFF_28_port);
   U45 : XNOR2_X1 port map( A => B(24), B => n238, ZN => DIFF_24_port);
   U46 : XNOR2_X1 port map( A => n197, B => B(61), ZN => DIFF_61_port);
   U47 : XNOR2_X1 port map( A => B(60), B => n199, ZN => DIFF_60_port);
   U48 : XNOR2_X1 port map( A => B(56), B => n203, ZN => DIFF_56_port);
   U49 : XNOR2_X1 port map( A => B(52), B => n207, ZN => DIFF_52_port);
   U50 : XNOR2_X1 port map( A => B(48), B => n213, ZN => DIFF_48_port);
   U51 : OR2_X1 port map( A1 => n196, A2 => B(62), ZN => n195);
   U52 : OR3_X1 port map( A1 => B(21), A2 => B(22), A3 => n239, ZN => n237);
   U53 : XNOR2_X1 port map( A => B(20), B => n242, ZN => DIFF_20_port);
   U54 : OR2_X1 port map( A1 => n239, A2 => B(21), ZN => n240);
   U55 : NOR2_X1 port map( A1 => B(19), A2 => n241, ZN => n242);
   U56 : OR3_X1 port map( A1 => B(19), A2 => B(20), A3 => n241, ZN => n239);
   U57 : XNOR2_X1 port map( A => n189, B => B(14), ZN => DIFF_14_port);
   U58 : NOR2_X1 port map( A1 => n247, A2 => B(13), ZN => n189);
   U59 : XNOR2_X1 port map( A => n193, B => B(6), ZN => DIFF_6_port);
   U60 : NOR2_X1 port map( A1 => n194, A2 => B(5), ZN => n193);
   U61 : XNOR2_X1 port map( A => n248, B => B(10), ZN => DIFF_10_port);
   U62 : NOR2_X1 port map( A1 => n190, A2 => B(9), ZN => n248);
   U63 : XNOR2_X1 port map( A => B(16), B => n246, ZN => DIFF_16_port);
   U64 : NOR2_X1 port map( A1 => B(15), A2 => n245, ZN => n246);
   U65 : XNOR2_X1 port map( A => B(12), B => n250, ZN => DIFF_12_port);
   U66 : NOR2_X1 port map( A1 => B(11), A2 => n249, ZN => n250);
   U67 : XNOR2_X1 port map( A => B(8), B => n191, ZN => DIFF_8_port);
   U68 : NOR2_X1 port map( A1 => B(7), A2 => n192, ZN => n191);
   U69 : XNOR2_X1 port map( A => B(2), B => n232, ZN => DIFF_2_port);
   U70 : NOR2_X1 port map( A1 => B(0), A2 => B(1), ZN => n232);
   U71 : XNOR2_X1 port map( A => B(4), B => n210, ZN => DIFF_4_port);
   U72 : NOR2_X1 port map( A1 => B(3), A2 => n211, ZN => n210);
   U73 : OR3_X1 port map( A1 => B(5), A2 => B(6), A3 => n194, ZN => n192);
   U74 : OR3_X1 port map( A1 => B(10), A2 => B(9), A3 => n190, ZN => n249);
   U75 : OR3_X1 port map( A1 => B(13), A2 => B(14), A3 => n247, ZN => n245);
   U76 : OR3_X1 port map( A1 => B(17), A2 => B(18), A3 => n243, ZN => n241);
   U77 : OR3_X1 port map( A1 => B(7), A2 => B(8), A3 => n192, ZN => n190);
   U78 : OR3_X1 port map( A1 => B(11), A2 => B(12), A3 => n249, ZN => n247);
   U79 : OR3_X1 port map( A1 => B(15), A2 => B(16), A3 => n245, ZN => n243);
   U80 : OR3_X1 port map( A1 => B(3), A2 => B(4), A3 => n211, ZN => n194);
   U83 : OR2_X1 port map( A1 => n243, A2 => B(17), ZN => n244);
   U123 : OR3_X1 port map( A1 => B(1), A2 => B(2), A3 => B(0), ZN => n211);
   U126 : INV_X1 port map( A => B(61), ZN => n251);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_14_DW01_sub_0 is

   port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (63 downto 0);  CO : out std_logic);

end complementer_N64_14_DW01_sub_0;

architecture SYN_rpl of complementer_N64_14_DW01_sub_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal DIFF_62_port, DIFF_61_port, DIFF_60_port, DIFF_59_port, DIFF_58_port,
      DIFF_57_port, DIFF_56_port, DIFF_55_port, DIFF_54_port, DIFF_53_port, 
      DIFF_52_port, DIFF_51_port, DIFF_50_port, DIFF_49_port, DIFF_48_port, 
      DIFF_47_port, DIFF_46_port, DIFF_45_port, DIFF_44_port, DIFF_43_port, 
      DIFF_42_port, DIFF_41_port, DIFF_40_port, DIFF_39_port, DIFF_38_port, 
      DIFF_37_port, DIFF_36_port, DIFF_35_port, DIFF_34_port, DIFF_33_port, 
      DIFF_32_port, DIFF_31_port, DIFF_30_port, DIFF_29_port, DIFF_28_port, 
      DIFF_27_port, DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, 
      DIFF_22_port, DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, 
      DIFF_17_port, DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, 
      DIFF_12_port, DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, 
      DIFF_7_port, DIFF_6_port, DIFF_5_port, DIFF_4_port, DIFF_3_port, 
      DIFF_2_port, DIFF_1_port, DIFF_63_port, n190, n191, n192, n193, n194, 
      n196, n197, n198, n199, n200, n202, n203, n204, n206, n207, n208, n210, 
      n211, n212, n213, n214, n216, n217, n218, n220, n221, n222, n224, n225, 
      n226, n228, n229, n230, n232, n233, n234, n235, n237, n238, n239, n241, 
      n242, n243, n245, n246, n247, n248, n249, n250, n251, n189, n195, n201, 
      n205, n209, n215, n219, n223, n227, n231, n236, n240, n244 : std_logic;

begin
   DIFF <= ( DIFF_63_port, DIFF_62_port, DIFF_61_port, DIFF_60_port, 
      DIFF_59_port, DIFF_58_port, DIFF_57_port, DIFF_56_port, DIFF_55_port, 
      DIFF_54_port, DIFF_53_port, DIFF_52_port, DIFF_51_port, DIFF_50_port, 
      DIFF_49_port, DIFF_48_port, DIFF_47_port, DIFF_46_port, DIFF_45_port, 
      DIFF_44_port, DIFF_43_port, DIFF_42_port, DIFF_41_port, DIFF_40_port, 
      DIFF_39_port, DIFF_38_port, DIFF_37_port, DIFF_36_port, DIFF_35_port, 
      DIFF_34_port, DIFF_33_port, DIFF_32_port, DIFF_31_port, DIFF_30_port, 
      DIFF_29_port, DIFF_28_port, DIFF_27_port, DIFF_26_port, DIFF_25_port, 
      DIFF_24_port, DIFF_23_port, DIFF_22_port, DIFF_21_port, DIFF_20_port, 
      DIFF_19_port, DIFF_18_port, DIFF_17_port, DIFF_16_port, DIFF_15_port, 
      DIFF_14_port, DIFF_13_port, DIFF_12_port, DIFF_11_port, DIFF_10_port, 
      DIFF_9_port, DIFF_8_port, DIFF_7_port, DIFF_6_port, DIFF_5_port, 
      DIFF_4_port, DIFF_3_port, DIFF_2_port, DIFF_1_port, B(0) );
   
   U81 : XOR2_X1 port map( A => n190, B => B(9), Z => DIFF_9_port);
   U82 : XOR2_X1 port map( A => n192, B => B(7), Z => DIFF_7_port);
   U83 : XOR2_X1 port map( A => n193, B => B(6), Z => DIFF_6_port);
   U85 : XOR2_X1 port map( A => n196, B => B(62), Z => DIFF_62_port);
   U86 : XOR2_X1 port map( A => n194, B => B(5), Z => DIFF_5_port);
   U87 : XOR2_X1 port map( A => n198, B => B(59), Z => DIFF_59_port);
   U89 : XOR2_X1 port map( A => n200, B => B(57), Z => DIFF_57_port);
   U90 : XOR2_X1 port map( A => n202, B => B(55), Z => DIFF_55_port);
   U92 : XOR2_X1 port map( A => n204, B => B(53), Z => DIFF_53_port);
   U93 : XOR2_X1 port map( A => n206, B => B(51), Z => DIFF_51_port);
   U95 : XOR2_X1 port map( A => n208, B => B(49), Z => DIFF_49_port);
   U96 : XOR2_X1 port map( A => n212, B => B(47), Z => DIFF_47_port);
   U98 : XOR2_X1 port map( A => n214, B => B(45), Z => DIFF_45_port);
   U99 : XOR2_X1 port map( A => n216, B => B(43), Z => DIFF_43_port);
   U101 : XOR2_X1 port map( A => n218, B => B(41), Z => DIFF_41_port);
   U102 : XOR2_X1 port map( A => n211, B => B(3), Z => DIFF_3_port);
   U103 : XOR2_X1 port map( A => n220, B => B(39), Z => DIFF_39_port);
   U105 : XOR2_X1 port map( A => n222, B => B(37), Z => DIFF_37_port);
   U106 : XOR2_X1 port map( A => n224, B => B(35), Z => DIFF_35_port);
   U108 : XOR2_X1 port map( A => n226, B => B(33), Z => DIFF_33_port);
   U109 : XOR2_X1 port map( A => n228, B => B(31), Z => DIFF_31_port);
   U111 : XOR2_X1 port map( A => n230, B => B(29), Z => DIFF_29_port);
   U112 : XOR2_X1 port map( A => n233, B => B(27), Z => DIFF_27_port);
   U114 : XOR2_X1 port map( A => n235, B => B(25), Z => DIFF_25_port);
   U115 : XOR2_X1 port map( A => n237, B => B(23), Z => DIFF_23_port);
   U117 : XOR2_X1 port map( A => n239, B => B(21), Z => DIFF_21_port);
   U118 : XOR2_X1 port map( A => B(1), B => B(0), Z => DIFF_1_port);
   U119 : XOR2_X1 port map( A => n241, B => B(19), Z => DIFF_19_port);
   U121 : XOR2_X1 port map( A => n243, B => B(17), Z => DIFF_17_port);
   U122 : XOR2_X1 port map( A => n245, B => B(15), Z => DIFF_15_port);
   U123 : XOR2_X1 port map( A => n248, B => B(14), Z => DIFF_14_port);
   U124 : XOR2_X1 port map( A => n247, B => B(13), Z => DIFF_13_port);
   U125 : XOR2_X1 port map( A => n249, B => B(11), Z => DIFF_11_port);
   U126 : XOR2_X1 port map( A => n251, B => B(10), Z => DIFF_10_port);
   U1 : XNOR2_X1 port map( A => B(44), B => n217, ZN => DIFF_44_port);
   U2 : NOR2_X1 port map( A1 => B(43), A2 => n216, ZN => n217);
   U3 : XNOR2_X1 port map( A => B(40), B => n221, ZN => DIFF_40_port);
   U4 : NOR2_X1 port map( A1 => B(39), A2 => n220, ZN => n221);
   U5 : XNOR2_X1 port map( A => B(36), B => n225, ZN => DIFF_36_port);
   U6 : NOR2_X1 port map( A1 => B(35), A2 => n224, ZN => n225);
   U7 : XNOR2_X1 port map( A => B(32), B => n229, ZN => DIFF_32_port);
   U8 : NOR2_X1 port map( A1 => B(31), A2 => n228, ZN => n229);
   U9 : XNOR2_X1 port map( A => B(28), B => n234, ZN => DIFF_28_port);
   U10 : NOR2_X1 port map( A1 => B(27), A2 => n233, ZN => n234);
   U11 : OR3_X1 port map( A1 => B(25), A2 => B(26), A3 => n235, ZN => n233);
   U12 : OR3_X1 port map( A1 => B(29), A2 => B(30), A3 => n230, ZN => n228);
   U13 : OR3_X1 port map( A1 => B(33), A2 => B(34), A3 => n226, ZN => n224);
   U14 : OR3_X1 port map( A1 => B(37), A2 => B(38), A3 => n222, ZN => n220);
   U15 : OR3_X1 port map( A1 => B(41), A2 => B(42), A3 => n218, ZN => n216);
   U16 : OR3_X1 port map( A1 => B(27), A2 => B(28), A3 => n233, ZN => n230);
   U17 : OR3_X1 port map( A1 => B(31), A2 => B(32), A3 => n228, ZN => n226);
   U18 : OR3_X1 port map( A1 => B(35), A2 => B(36), A3 => n224, ZN => n222);
   U19 : OR3_X1 port map( A1 => B(39), A2 => B(40), A3 => n220, ZN => n218);
   U20 : XNOR2_X1 port map( A => n189, B => B(42), ZN => DIFF_42_port);
   U21 : NOR2_X1 port map( A1 => n218, A2 => B(41), ZN => n189);
   U22 : XNOR2_X1 port map( A => n195, B => B(38), ZN => DIFF_38_port);
   U23 : NOR2_X1 port map( A1 => n222, A2 => B(37), ZN => n195);
   U24 : XNOR2_X1 port map( A => n201, B => B(34), ZN => DIFF_34_port);
   U25 : NOR2_X1 port map( A1 => n226, A2 => B(33), ZN => n201);
   U26 : XNOR2_X1 port map( A => n205, B => B(30), ZN => DIFF_30_port);
   U27 : NOR2_X1 port map( A1 => n230, A2 => B(29), ZN => n205);
   U28 : XNOR2_X1 port map( A => n209, B => B(26), ZN => DIFF_26_port);
   U29 : NOR2_X1 port map( A1 => n235, A2 => B(25), ZN => n209);
   U30 : NOR3_X1 port map( A1 => B(59), A2 => B(60), A3 => n198, ZN => n197);
   U31 : XNOR2_X1 port map( A => n215, B => B(46), ZN => DIFF_46_port);
   U32 : NOR2_X1 port map( A1 => n214, A2 => B(45), ZN => n215);
   U33 : XNOR2_X1 port map( A => n219, B => B(50), ZN => DIFF_50_port);
   U34 : NOR2_X1 port map( A1 => n208, A2 => B(49), ZN => n219);
   U35 : XNOR2_X1 port map( A => n223, B => B(54), ZN => DIFF_54_port);
   U36 : NOR2_X1 port map( A1 => n204, A2 => B(53), ZN => n223);
   U37 : XNOR2_X1 port map( A => B(48), B => n213, ZN => DIFF_48_port);
   U38 : NOR2_X1 port map( A1 => B(47), A2 => n212, ZN => n213);
   U39 : XNOR2_X1 port map( A => B(60), B => n199, ZN => DIFF_60_port);
   U40 : NOR2_X1 port map( A1 => B(59), A2 => n198, ZN => n199);
   U41 : XNOR2_X1 port map( A => B(56), B => n203, ZN => DIFF_56_port);
   U42 : NOR2_X1 port map( A1 => B(55), A2 => n202, ZN => n203);
   U43 : XOR2_X1 port map( A => n197, B => n244, Z => DIFF_61_port);
   U44 : NAND2_X1 port map( A1 => n197, A2 => n244, ZN => n196);
   U45 : OR3_X1 port map( A1 => B(57), A2 => B(58), A3 => n200, ZN => n198);
   U46 : OR3_X1 port map( A1 => B(49), A2 => B(50), A3 => n208, ZN => n206);
   U47 : OR3_X1 port map( A1 => B(45), A2 => B(46), A3 => n214, ZN => n212);
   U48 : OR3_X1 port map( A1 => B(53), A2 => B(54), A3 => n204, ZN => n202);
   U49 : OR3_X1 port map( A1 => B(43), A2 => B(44), A3 => n216, ZN => n214);
   U50 : OR3_X1 port map( A1 => B(55), A2 => B(56), A3 => n202, ZN => n200);
   U51 : OR3_X1 port map( A1 => B(47), A2 => B(48), A3 => n212, ZN => n208);
   U52 : XNOR2_X1 port map( A => n227, B => B(58), ZN => DIFF_58_port);
   U53 : NOR2_X1 port map( A1 => n200, A2 => B(57), ZN => n227);
   U54 : XNOR2_X1 port map( A => B(24), B => n238, ZN => DIFF_24_port);
   U55 : NOR2_X1 port map( A1 => B(23), A2 => n237, ZN => n238);
   U56 : OR3_X1 port map( A1 => B(23), A2 => B(24), A3 => n237, ZN => n235);
   U57 : XNOR2_X1 port map( A => n231, B => B(63), ZN => DIFF_63_port);
   U58 : NOR2_X1 port map( A1 => n196, A2 => B(62), ZN => n231);
   U59 : XNOR2_X1 port map( A => B(52), B => n207, ZN => DIFF_52_port);
   U60 : NOR2_X1 port map( A1 => B(51), A2 => n206, ZN => n207);
   U61 : OR3_X1 port map( A1 => B(51), A2 => B(52), A3 => n206, ZN => n204);
   U62 : XNOR2_X1 port map( A => n236, B => B(22), ZN => DIFF_22_port);
   U63 : NOR2_X1 port map( A1 => n239, A2 => B(21), ZN => n236);
   U64 : OR3_X1 port map( A1 => B(21), A2 => B(22), A3 => n239, ZN => n237);
   U65 : XNOR2_X1 port map( A => B(20), B => n242, ZN => DIFF_20_port);
   U66 : NOR2_X1 port map( A1 => B(19), A2 => n241, ZN => n242);
   U67 : OR3_X1 port map( A1 => B(19), A2 => B(20), A3 => n241, ZN => n239);
   U68 : XNOR2_X1 port map( A => n240, B => B(18), ZN => DIFF_18_port);
   U69 : NOR2_X1 port map( A1 => n243, A2 => B(17), ZN => n240);
   U70 : OR3_X1 port map( A1 => B(17), A2 => B(18), A3 => n243, ZN => n241);
   U71 : NOR2_X1 port map( A1 => B(15), A2 => n245, ZN => n246);
   U72 : NOR2_X1 port map( A1 => B(11), A2 => n249, ZN => n250);
   U73 : NOR2_X1 port map( A1 => B(7), A2 => n192, ZN => n191);
   U74 : NOR2_X1 port map( A1 => B(3), A2 => n211, ZN => n210);
   U75 : OR3_X1 port map( A1 => B(13), A2 => B(14), A3 => n247, ZN => n245);
   U76 : OR3_X1 port map( A1 => B(10), A2 => B(9), A3 => n190, ZN => n249);
   U77 : OR3_X1 port map( A1 => B(5), A2 => B(6), A3 => n194, ZN => n192);
   U78 : OR3_X1 port map( A1 => B(15), A2 => B(16), A3 => n245, ZN => n243);
   U79 : OR3_X1 port map( A1 => B(11), A2 => B(12), A3 => n249, ZN => n247);
   U80 : OR3_X1 port map( A1 => B(7), A2 => B(8), A3 => n192, ZN => n190);
   U84 : OR3_X1 port map( A1 => B(3), A2 => B(4), A3 => n211, ZN => n194);
   U88 : XNOR2_X1 port map( A => B(16), B => n246, ZN => DIFF_16_port);
   U91 : XNOR2_X1 port map( A => B(12), B => n250, ZN => DIFF_12_port);
   U94 : XNOR2_X1 port map( A => B(8), B => n191, ZN => DIFF_8_port);
   U97 : XNOR2_X1 port map( A => B(4), B => n210, ZN => DIFF_4_port);
   U100 : XNOR2_X1 port map( A => B(2), B => n232, ZN => DIFF_2_port);
   U104 : OR2_X1 port map( A1 => n247, A2 => B(13), ZN => n248);
   U107 : OR2_X1 port map( A1 => n190, A2 => B(9), ZN => n251);
   U110 : OR2_X1 port map( A1 => n194, A2 => B(5), ZN => n193);
   U113 : OR3_X1 port map( A1 => B(1), A2 => B(2), A3 => B(0), ZN => n211);
   U116 : NOR2_X1 port map( A1 => B(0), A2 => B(1), ZN => n232);
   U120 : INV_X1 port map( A => B(61), ZN => n244);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_15_DW01_sub_0 is

   port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (63 downto 0);  CO : out std_logic);

end complementer_N64_15_DW01_sub_0;

architecture SYN_rpl of complementer_N64_15_DW01_sub_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal DIFF_62_port, DIFF_63_port, DIFF_17_port, DIFF_18_port, DIFF_19_port,
      DIFF_20_port, DIFF_21_port, DIFF_22_port, DIFF_23_port, DIFF_24_port, 
      DIFF_25_port, DIFF_26_port, DIFF_27_port, DIFF_28_port, DIFF_29_port, 
      DIFF_30_port, DIFF_31_port, DIFF_32_port, DIFF_33_port, DIFF_34_port, 
      DIFF_35_port, DIFF_36_port, DIFF_37_port, DIFF_38_port, DIFF_39_port, 
      DIFF_40_port, DIFF_41_port, DIFF_42_port, DIFF_43_port, DIFF_44_port, 
      DIFF_45_port, DIFF_46_port, DIFF_47_port, DIFF_48_port, DIFF_49_port, 
      DIFF_50_port, DIFF_51_port, DIFF_52_port, DIFF_53_port, DIFF_54_port, 
      DIFF_55_port, DIFF_56_port, DIFF_57_port, DIFF_58_port, DIFF_59_port, 
      DIFF_60_port, DIFF_61_port, DIFF_3_port, DIFF_4_port, DIFF_5_port, 
      DIFF_6_port, DIFF_7_port, DIFF_8_port, DIFF_9_port, DIFF_10_port, 
      DIFF_11_port, DIFF_12_port, DIFF_13_port, DIFF_14_port, DIFF_15_port, 
      DIFF_16_port, DIFF_2_port, DIFF_1_port, n190, n191, n192, n194, n196, 
      n197, n198, n199, n200, n202, n203, n204, n206, n207, n208, n210, n211, 
      n212, n213, n214, n216, n217, n218, n220, n221, n222, n224, n225, n226, 
      n228, n229, n230, n232, n233, n234, n235, n237, n238, n239, n241, n242, 
      n243, n245, n246, n247, n249, n250, n189, n193, n195, n201, n205, n209, 
      n215, n219, n223, n227, n231, n236, n240, n244, n248, n251 : std_logic;

begin
   DIFF <= ( DIFF_63_port, DIFF_62_port, DIFF_61_port, DIFF_60_port, 
      DIFF_59_port, DIFF_58_port, DIFF_57_port, DIFF_56_port, DIFF_55_port, 
      DIFF_54_port, DIFF_53_port, DIFF_52_port, DIFF_51_port, DIFF_50_port, 
      DIFF_49_port, DIFF_48_port, DIFF_47_port, DIFF_46_port, DIFF_45_port, 
      DIFF_44_port, DIFF_43_port, DIFF_42_port, DIFF_41_port, DIFF_40_port, 
      DIFF_39_port, DIFF_38_port, DIFF_37_port, DIFF_36_port, DIFF_35_port, 
      DIFF_34_port, DIFF_33_port, DIFF_32_port, DIFF_31_port, DIFF_30_port, 
      DIFF_29_port, DIFF_28_port, DIFF_27_port, DIFF_26_port, DIFF_25_port, 
      DIFF_24_port, DIFF_23_port, DIFF_22_port, DIFF_21_port, DIFF_20_port, 
      DIFF_19_port, DIFF_18_port, DIFF_17_port, DIFF_16_port, DIFF_15_port, 
      DIFF_14_port, DIFF_13_port, DIFF_12_port, DIFF_11_port, DIFF_10_port, 
      DIFF_9_port, DIFF_8_port, DIFF_7_port, DIFF_6_port, DIFF_5_port, 
      DIFF_4_port, DIFF_3_port, DIFF_2_port, DIFF_1_port, B(0) );
   
   U81 : XOR2_X1 port map( A => n190, B => B(9), Z => DIFF_9_port);
   U82 : XOR2_X1 port map( A => n192, B => B(7), Z => DIFF_7_port);
   U85 : XOR2_X1 port map( A => n196, B => B(62), Z => DIFF_62_port);
   U86 : XOR2_X1 port map( A => n194, B => B(5), Z => DIFF_5_port);
   U87 : XOR2_X1 port map( A => n198, B => B(59), Z => DIFF_59_port);
   U89 : XOR2_X1 port map( A => n200, B => B(57), Z => DIFF_57_port);
   U90 : XOR2_X1 port map( A => n202, B => B(55), Z => DIFF_55_port);
   U92 : XOR2_X1 port map( A => n204, B => B(53), Z => DIFF_53_port);
   U93 : XOR2_X1 port map( A => n206, B => B(51), Z => DIFF_51_port);
   U95 : XOR2_X1 port map( A => n208, B => B(49), Z => DIFF_49_port);
   U96 : XOR2_X1 port map( A => n212, B => B(47), Z => DIFF_47_port);
   U98 : XOR2_X1 port map( A => n214, B => B(45), Z => DIFF_45_port);
   U99 : XOR2_X1 port map( A => n216, B => B(43), Z => DIFF_43_port);
   U101 : XOR2_X1 port map( A => n218, B => B(41), Z => DIFF_41_port);
   U102 : XOR2_X1 port map( A => n211, B => B(3), Z => DIFF_3_port);
   U103 : XOR2_X1 port map( A => n220, B => B(39), Z => DIFF_39_port);
   U105 : XOR2_X1 port map( A => n222, B => B(37), Z => DIFF_37_port);
   U106 : XOR2_X1 port map( A => n224, B => B(35), Z => DIFF_35_port);
   U108 : XOR2_X1 port map( A => n226, B => B(33), Z => DIFF_33_port);
   U109 : XOR2_X1 port map( A => n228, B => B(31), Z => DIFF_31_port);
   U111 : XOR2_X1 port map( A => n230, B => B(29), Z => DIFF_29_port);
   U112 : XOR2_X1 port map( A => n233, B => B(27), Z => DIFF_27_port);
   U114 : XOR2_X1 port map( A => n235, B => B(25), Z => DIFF_25_port);
   U115 : XOR2_X1 port map( A => n237, B => B(23), Z => DIFF_23_port);
   U117 : XOR2_X1 port map( A => n239, B => B(21), Z => DIFF_21_port);
   U118 : XOR2_X1 port map( A => B(1), B => B(0), Z => DIFF_1_port);
   U119 : XOR2_X1 port map( A => n241, B => B(19), Z => DIFF_19_port);
   U121 : XOR2_X1 port map( A => n243, B => B(17), Z => DIFF_17_port);
   U122 : XOR2_X1 port map( A => n245, B => B(15), Z => DIFF_15_port);
   U124 : XOR2_X1 port map( A => n247, B => B(13), Z => DIFF_13_port);
   U125 : XOR2_X1 port map( A => n249, B => B(11), Z => DIFF_11_port);
   U1 : XNOR2_X1 port map( A => n189, B => B(46), ZN => DIFF_46_port);
   U2 : NOR2_X1 port map( A1 => n214, A2 => B(45), ZN => n189);
   U3 : XNOR2_X1 port map( A => B(44), B => n217, ZN => DIFF_44_port);
   U4 : NOR2_X1 port map( A1 => B(43), A2 => n216, ZN => n217);
   U5 : XNOR2_X1 port map( A => B(40), B => n221, ZN => DIFF_40_port);
   U6 : NOR2_X1 port map( A1 => B(39), A2 => n220, ZN => n221);
   U7 : XNOR2_X1 port map( A => B(36), B => n225, ZN => DIFF_36_port);
   U8 : NOR2_X1 port map( A1 => B(35), A2 => n224, ZN => n225);
   U9 : XNOR2_X1 port map( A => B(32), B => n229, ZN => DIFF_32_port);
   U10 : NOR2_X1 port map( A1 => B(31), A2 => n228, ZN => n229);
   U11 : XNOR2_X1 port map( A => B(28), B => n234, ZN => DIFF_28_port);
   U12 : NOR2_X1 port map( A1 => B(27), A2 => n233, ZN => n234);
   U13 : XNOR2_X1 port map( A => B(48), B => n213, ZN => DIFF_48_port);
   U14 : NOR2_X1 port map( A1 => B(47), A2 => n212, ZN => n213);
   U15 : XNOR2_X1 port map( A => B(24), B => n238, ZN => DIFF_24_port);
   U16 : NOR2_X1 port map( A1 => B(23), A2 => n237, ZN => n238);
   U17 : OR3_X1 port map( A1 => B(25), A2 => B(26), A3 => n235, ZN => n233);
   U18 : OR3_X1 port map( A1 => B(29), A2 => B(30), A3 => n230, ZN => n228);
   U19 : OR3_X1 port map( A1 => B(33), A2 => B(34), A3 => n226, ZN => n224);
   U20 : OR3_X1 port map( A1 => B(37), A2 => B(38), A3 => n222, ZN => n220);
   U21 : OR3_X1 port map( A1 => B(41), A2 => B(42), A3 => n218, ZN => n216);
   U22 : OR3_X1 port map( A1 => B(45), A2 => B(46), A3 => n214, ZN => n212);
   U23 : OR3_X1 port map( A1 => B(23), A2 => B(24), A3 => n237, ZN => n235);
   U24 : OR3_X1 port map( A1 => B(27), A2 => B(28), A3 => n233, ZN => n230);
   U25 : OR3_X1 port map( A1 => B(31), A2 => B(32), A3 => n228, ZN => n226);
   U26 : OR3_X1 port map( A1 => B(35), A2 => B(36), A3 => n224, ZN => n222);
   U27 : OR3_X1 port map( A1 => B(39), A2 => B(40), A3 => n220, ZN => n218);
   U28 : OR3_X1 port map( A1 => B(43), A2 => B(44), A3 => n216, ZN => n214);
   U29 : OR3_X1 port map( A1 => B(47), A2 => B(48), A3 => n212, ZN => n208);
   U30 : XNOR2_X1 port map( A => n193, B => B(42), ZN => DIFF_42_port);
   U31 : NOR2_X1 port map( A1 => n218, A2 => B(41), ZN => n193);
   U32 : XNOR2_X1 port map( A => n195, B => B(38), ZN => DIFF_38_port);
   U33 : NOR2_X1 port map( A1 => n222, A2 => B(37), ZN => n195);
   U34 : XNOR2_X1 port map( A => n201, B => B(34), ZN => DIFF_34_port);
   U35 : NOR2_X1 port map( A1 => n226, A2 => B(33), ZN => n201);
   U36 : XNOR2_X1 port map( A => n205, B => B(30), ZN => DIFF_30_port);
   U37 : NOR2_X1 port map( A1 => n230, A2 => B(29), ZN => n205);
   U38 : XNOR2_X1 port map( A => n209, B => B(26), ZN => DIFF_26_port);
   U39 : NOR2_X1 port map( A1 => n235, A2 => B(25), ZN => n209);
   U40 : XOR2_X1 port map( A => n197, B => n251, Z => DIFF_61_port);
   U41 : NAND2_X1 port map( A1 => n197, A2 => n251, ZN => n196);
   U42 : OR3_X1 port map( A1 => B(53), A2 => B(54), A3 => n204, ZN => n202);
   U43 : XNOR2_X1 port map( A => n215, B => B(54), ZN => DIFF_54_port);
   U44 : NOR2_X1 port map( A1 => n204, A2 => B(53), ZN => n215);
   U45 : XNOR2_X1 port map( A => n219, B => B(22), ZN => DIFF_22_port);
   U46 : NOR2_X1 port map( A1 => n239, A2 => B(21), ZN => n219);
   U47 : OR3_X1 port map( A1 => B(21), A2 => B(22), A3 => n239, ZN => n237);
   U48 : NOR3_X1 port map( A1 => B(59), A2 => B(60), A3 => n198, ZN => n197);
   U49 : XNOR2_X1 port map( A => n223, B => B(63), ZN => DIFF_63_port);
   U50 : NOR2_X1 port map( A1 => n196, A2 => B(62), ZN => n223);
   U51 : XNOR2_X1 port map( A => B(60), B => n199, ZN => DIFF_60_port);
   U52 : NOR2_X1 port map( A1 => B(59), A2 => n198, ZN => n199);
   U53 : XNOR2_X1 port map( A => B(56), B => n203, ZN => DIFF_56_port);
   U54 : NOR2_X1 port map( A1 => B(55), A2 => n202, ZN => n203);
   U55 : XNOR2_X1 port map( A => B(52), B => n207, ZN => DIFF_52_port);
   U56 : NOR2_X1 port map( A1 => B(51), A2 => n206, ZN => n207);
   U57 : OR3_X1 port map( A1 => B(57), A2 => B(58), A3 => n200, ZN => n198);
   U58 : OR3_X1 port map( A1 => B(49), A2 => B(50), A3 => n208, ZN => n206);
   U59 : OR3_X1 port map( A1 => B(51), A2 => B(52), A3 => n206, ZN => n204);
   U60 : OR3_X1 port map( A1 => B(55), A2 => B(56), A3 => n202, ZN => n200);
   U61 : XNOR2_X1 port map( A => n227, B => B(50), ZN => DIFF_50_port);
   U62 : NOR2_X1 port map( A1 => n208, A2 => B(49), ZN => n227);
   U63 : XNOR2_X1 port map( A => n231, B => B(58), ZN => DIFF_58_port);
   U64 : NOR2_X1 port map( A1 => n200, A2 => B(57), ZN => n231);
   U65 : XNOR2_X1 port map( A => B(20), B => n242, ZN => DIFF_20_port);
   U66 : NOR2_X1 port map( A1 => B(19), A2 => n241, ZN => n242);
   U67 : OR3_X1 port map( A1 => B(19), A2 => B(20), A3 => n241, ZN => n239);
   U68 : XNOR2_X1 port map( A => n236, B => B(18), ZN => DIFF_18_port);
   U69 : NOR2_X1 port map( A1 => n243, A2 => B(17), ZN => n236);
   U70 : OR3_X1 port map( A1 => B(17), A2 => B(18), A3 => n243, ZN => n241);
   U71 : XNOR2_X1 port map( A => B(16), B => n246, ZN => DIFF_16_port);
   U72 : XNOR2_X1 port map( A => n240, B => B(14), ZN => DIFF_14_port);
   U73 : NOR2_X1 port map( A1 => n247, A2 => B(13), ZN => n240);
   U74 : XNOR2_X1 port map( A => n244, B => B(10), ZN => DIFF_10_port);
   U75 : NOR2_X1 port map( A1 => n190, A2 => B(9), ZN => n244);
   U76 : XNOR2_X1 port map( A => n248, B => B(6), ZN => DIFF_6_port);
   U77 : NOR2_X1 port map( A1 => n194, A2 => B(5), ZN => n248);
   U78 : NOR2_X1 port map( A1 => B(15), A2 => n245, ZN => n246);
   U79 : XNOR2_X1 port map( A => B(12), B => n250, ZN => DIFF_12_port);
   U80 : NOR2_X1 port map( A1 => B(11), A2 => n249, ZN => n250);
   U83 : XNOR2_X1 port map( A => B(8), B => n191, ZN => DIFF_8_port);
   U84 : NOR2_X1 port map( A1 => B(7), A2 => n192, ZN => n191);
   U88 : XNOR2_X1 port map( A => B(2), B => n232, ZN => DIFF_2_port);
   U91 : NOR2_X1 port map( A1 => B(0), A2 => B(1), ZN => n232);
   U94 : XNOR2_X1 port map( A => B(4), B => n210, ZN => DIFF_4_port);
   U97 : NOR2_X1 port map( A1 => B(3), A2 => n211, ZN => n210);
   U100 : OR3_X1 port map( A1 => B(5), A2 => B(6), A3 => n194, ZN => n192);
   U104 : OR3_X1 port map( A1 => B(10), A2 => B(9), A3 => n190, ZN => n249);
   U107 : OR3_X1 port map( A1 => B(13), A2 => B(14), A3 => n247, ZN => n245);
   U110 : OR3_X1 port map( A1 => B(7), A2 => B(8), A3 => n192, ZN => n190);
   U113 : OR3_X1 port map( A1 => B(11), A2 => B(12), A3 => n249, ZN => n247);
   U116 : OR3_X1 port map( A1 => B(15), A2 => B(16), A3 => n245, ZN => n243);
   U120 : OR3_X1 port map( A1 => B(3), A2 => B(4), A3 => n211, ZN => n194);
   U123 : OR3_X1 port map( A1 => B(1), A2 => B(2), A3 => B(0), ZN => n211);
   U126 : INV_X1 port map( A => B(61), ZN => n251);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_16_DW01_sub_0 is

   port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (63 downto 0);  CO : out std_logic);

end complementer_N64_16_DW01_sub_0;

architecture SYN_rpl of complementer_N64_16_DW01_sub_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal DIFF_62_port, DIFF_61_port, DIFF_60_port, DIFF_59_port, DIFF_58_port,
      DIFF_57_port, DIFF_56_port, DIFF_55_port, DIFF_54_port, DIFF_53_port, 
      DIFF_52_port, DIFF_51_port, DIFF_50_port, DIFF_49_port, DIFF_48_port, 
      DIFF_47_port, DIFF_46_port, DIFF_45_port, DIFF_44_port, DIFF_43_port, 
      DIFF_42_port, DIFF_41_port, DIFF_40_port, DIFF_39_port, DIFF_38_port, 
      DIFF_37_port, DIFF_36_port, DIFF_35_port, DIFF_34_port, DIFF_33_port, 
      DIFF_32_port, DIFF_31_port, DIFF_30_port, DIFF_29_port, DIFF_28_port, 
      DIFF_27_port, DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, 
      DIFF_22_port, DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, 
      DIFF_17_port, DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, 
      DIFF_12_port, DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, 
      DIFF_7_port, DIFF_6_port, DIFF_5_port, DIFF_4_port, DIFF_3_port, 
      DIFF_2_port, DIFF_1_port, DIFF_63_port, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, 
      n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, 
      n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, 
      n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, 
      n243, n244, n245, n246, n247, n248, n249, n250, n251, n189 : std_logic;

begin
   DIFF <= ( DIFF_63_port, DIFF_62_port, DIFF_61_port, DIFF_60_port, 
      DIFF_59_port, DIFF_58_port, DIFF_57_port, DIFF_56_port, DIFF_55_port, 
      DIFF_54_port, DIFF_53_port, DIFF_52_port, DIFF_51_port, DIFF_50_port, 
      DIFF_49_port, DIFF_48_port, DIFF_47_port, DIFF_46_port, DIFF_45_port, 
      DIFF_44_port, DIFF_43_port, DIFF_42_port, DIFF_41_port, DIFF_40_port, 
      DIFF_39_port, DIFF_38_port, DIFF_37_port, DIFF_36_port, DIFF_35_port, 
      DIFF_34_port, DIFF_33_port, DIFF_32_port, DIFF_31_port, DIFF_30_port, 
      DIFF_29_port, DIFF_28_port, DIFF_27_port, DIFF_26_port, DIFF_25_port, 
      DIFF_24_port, DIFF_23_port, DIFF_22_port, DIFF_21_port, DIFF_20_port, 
      DIFF_19_port, DIFF_18_port, DIFF_17_port, DIFF_16_port, DIFF_15_port, 
      DIFF_14_port, DIFF_13_port, DIFF_12_port, DIFF_11_port, DIFF_10_port, 
      DIFF_9_port, DIFF_8_port, DIFF_7_port, DIFF_6_port, DIFF_5_port, 
      DIFF_4_port, DIFF_3_port, DIFF_2_port, DIFF_1_port, B(0) );
   
   U81 : XOR2_X1 port map( A => n190, B => B(9), Z => DIFF_9_port);
   U82 : XOR2_X1 port map( A => n192, B => B(7), Z => DIFF_7_port);
   U83 : XOR2_X1 port map( A => n193, B => B(6), Z => DIFF_6_port);
   U84 : XOR2_X1 port map( A => n195, B => B(63), Z => DIFF_63_port);
   U85 : XOR2_X1 port map( A => n196, B => B(62), Z => DIFF_62_port);
   U86 : XOR2_X1 port map( A => n194, B => B(5), Z => DIFF_5_port);
   U87 : XOR2_X1 port map( A => n198, B => B(59), Z => DIFF_59_port);
   U88 : XOR2_X1 port map( A => n201, B => B(58), Z => DIFF_58_port);
   U89 : XOR2_X1 port map( A => n200, B => B(57), Z => DIFF_57_port);
   U90 : XOR2_X1 port map( A => n202, B => B(55), Z => DIFF_55_port);
   U91 : XOR2_X1 port map( A => n205, B => B(54), Z => DIFF_54_port);
   U92 : XOR2_X1 port map( A => n204, B => B(53), Z => DIFF_53_port);
   U93 : XOR2_X1 port map( A => n206, B => B(51), Z => DIFF_51_port);
   U94 : XOR2_X1 port map( A => n209, B => B(50), Z => DIFF_50_port);
   U95 : XOR2_X1 port map( A => n208, B => B(49), Z => DIFF_49_port);
   U96 : XOR2_X1 port map( A => n212, B => B(47), Z => DIFF_47_port);
   U97 : XOR2_X1 port map( A => n215, B => B(46), Z => DIFF_46_port);
   U98 : XOR2_X1 port map( A => n214, B => B(45), Z => DIFF_45_port);
   U99 : XOR2_X1 port map( A => n216, B => B(43), Z => DIFF_43_port);
   U100 : XOR2_X1 port map( A => n219, B => B(42), Z => DIFF_42_port);
   U101 : XOR2_X1 port map( A => n218, B => B(41), Z => DIFF_41_port);
   U102 : XOR2_X1 port map( A => n211, B => B(3), Z => DIFF_3_port);
   U103 : XOR2_X1 port map( A => n220, B => B(39), Z => DIFF_39_port);
   U104 : XOR2_X1 port map( A => n223, B => B(38), Z => DIFF_38_port);
   U105 : XOR2_X1 port map( A => n222, B => B(37), Z => DIFF_37_port);
   U106 : XOR2_X1 port map( A => n224, B => B(35), Z => DIFF_35_port);
   U107 : XOR2_X1 port map( A => n227, B => B(34), Z => DIFF_34_port);
   U108 : XOR2_X1 port map( A => n226, B => B(33), Z => DIFF_33_port);
   U109 : XOR2_X1 port map( A => n228, B => B(31), Z => DIFF_31_port);
   U110 : XOR2_X1 port map( A => n231, B => B(30), Z => DIFF_30_port);
   U111 : XOR2_X1 port map( A => n230, B => B(29), Z => DIFF_29_port);
   U112 : XOR2_X1 port map( A => n233, B => B(27), Z => DIFF_27_port);
   U113 : XOR2_X1 port map( A => n236, B => B(26), Z => DIFF_26_port);
   U114 : XOR2_X1 port map( A => n235, B => B(25), Z => DIFF_25_port);
   U115 : XOR2_X1 port map( A => n237, B => B(23), Z => DIFF_23_port);
   U116 : XOR2_X1 port map( A => n240, B => B(22), Z => DIFF_22_port);
   U117 : XOR2_X1 port map( A => n239, B => B(21), Z => DIFF_21_port);
   U118 : XOR2_X1 port map( A => B(1), B => B(0), Z => DIFF_1_port);
   U119 : XOR2_X1 port map( A => n241, B => B(19), Z => DIFF_19_port);
   U120 : XOR2_X1 port map( A => n244, B => B(18), Z => DIFF_18_port);
   U121 : XOR2_X1 port map( A => n243, B => B(17), Z => DIFF_17_port);
   U122 : XOR2_X1 port map( A => n245, B => B(15), Z => DIFF_15_port);
   U123 : XOR2_X1 port map( A => n248, B => B(14), Z => DIFF_14_port);
   U124 : XOR2_X1 port map( A => n247, B => B(13), Z => DIFF_13_port);
   U125 : XOR2_X1 port map( A => n249, B => B(11), Z => DIFF_11_port);
   U126 : XOR2_X1 port map( A => n251, B => B(10), Z => DIFF_10_port);
   U1 : NOR2_X1 port map( A1 => B(47), A2 => n212, ZN => n213);
   U2 : NAND2_X1 port map( A1 => n197, A2 => n189, ZN => n196);
   U3 : OR3_X1 port map( A1 => B(57), A2 => B(58), A3 => n200, ZN => n198);
   U4 : OR3_X1 port map( A1 => B(53), A2 => B(54), A3 => n204, ZN => n202);
   U5 : OR3_X1 port map( A1 => B(47), A2 => B(48), A3 => n212, ZN => n208);
   U6 : OR2_X1 port map( A1 => n200, A2 => B(57), ZN => n201);
   U7 : OR2_X1 port map( A1 => n204, A2 => B(53), ZN => n205);
   U8 : XNOR2_X1 port map( A => B(20), B => n242, ZN => DIFF_20_port);
   U9 : NOR2_X1 port map( A1 => B(43), A2 => n216, ZN => n217);
   U10 : NOR2_X1 port map( A1 => B(39), A2 => n220, ZN => n221);
   U11 : NOR2_X1 port map( A1 => B(35), A2 => n224, ZN => n225);
   U12 : NOR2_X1 port map( A1 => B(31), A2 => n228, ZN => n229);
   U13 : NOR2_X1 port map( A1 => B(27), A2 => n233, ZN => n234);
   U14 : NOR2_X1 port map( A1 => B(23), A2 => n237, ZN => n238);
   U15 : XNOR2_X1 port map( A => B(48), B => n213, ZN => DIFF_48_port);
   U16 : OR3_X1 port map( A1 => B(45), A2 => B(46), A3 => n214, ZN => n212);
   U17 : OR3_X1 port map( A1 => B(41), A2 => B(42), A3 => n218, ZN => n216);
   U18 : OR3_X1 port map( A1 => B(37), A2 => B(38), A3 => n222, ZN => n220);
   U19 : OR3_X1 port map( A1 => B(33), A2 => B(34), A3 => n226, ZN => n224);
   U20 : OR3_X1 port map( A1 => B(29), A2 => B(30), A3 => n230, ZN => n228);
   U21 : OR3_X1 port map( A1 => B(25), A2 => B(26), A3 => n235, ZN => n233);
   U22 : OR3_X1 port map( A1 => B(21), A2 => B(22), A3 => n239, ZN => n237);
   U23 : OR3_X1 port map( A1 => B(43), A2 => B(44), A3 => n216, ZN => n214);
   U24 : OR3_X1 port map( A1 => B(39), A2 => B(40), A3 => n220, ZN => n218);
   U25 : OR3_X1 port map( A1 => B(35), A2 => B(36), A3 => n224, ZN => n222);
   U26 : OR3_X1 port map( A1 => B(31), A2 => B(32), A3 => n228, ZN => n226);
   U27 : OR3_X1 port map( A1 => B(27), A2 => B(28), A3 => n233, ZN => n230);
   U28 : OR3_X1 port map( A1 => B(23), A2 => B(24), A3 => n237, ZN => n235);
   U29 : XNOR2_X1 port map( A => B(44), B => n217, ZN => DIFF_44_port);
   U30 : XNOR2_X1 port map( A => B(40), B => n221, ZN => DIFF_40_port);
   U31 : XNOR2_X1 port map( A => B(36), B => n225, ZN => DIFF_36_port);
   U32 : XNOR2_X1 port map( A => B(32), B => n229, ZN => DIFF_32_port);
   U33 : XNOR2_X1 port map( A => B(28), B => n234, ZN => DIFF_28_port);
   U34 : XNOR2_X1 port map( A => B(24), B => n238, ZN => DIFF_24_port);
   U35 : OR2_X1 port map( A1 => n214, A2 => B(45), ZN => n215);
   U36 : OR2_X1 port map( A1 => n218, A2 => B(41), ZN => n219);
   U37 : OR2_X1 port map( A1 => n222, A2 => B(37), ZN => n223);
   U38 : OR2_X1 port map( A1 => n226, A2 => B(33), ZN => n227);
   U39 : OR2_X1 port map( A1 => n230, A2 => B(29), ZN => n231);
   U40 : OR2_X1 port map( A1 => n235, A2 => B(25), ZN => n236);
   U41 : OR2_X1 port map( A1 => n239, A2 => B(21), ZN => n240);
   U42 : NOR3_X1 port map( A1 => B(59), A2 => B(60), A3 => n198, ZN => n197);
   U43 : XNOR2_X1 port map( A => n197, B => B(61), ZN => DIFF_61_port);
   U44 : XNOR2_X1 port map( A => B(60), B => n199, ZN => DIFF_60_port);
   U45 : NOR2_X1 port map( A1 => B(59), A2 => n198, ZN => n199);
   U46 : NOR2_X1 port map( A1 => B(51), A2 => n206, ZN => n207);
   U47 : XNOR2_X1 port map( A => B(56), B => n203, ZN => DIFF_56_port);
   U48 : XNOR2_X1 port map( A => B(52), B => n207, ZN => DIFF_52_port);
   U49 : NOR2_X1 port map( A1 => B(55), A2 => n202, ZN => n203);
   U50 : OR3_X1 port map( A1 => B(49), A2 => B(50), A3 => n208, ZN => n206);
   U51 : OR3_X1 port map( A1 => B(51), A2 => B(52), A3 => n206, ZN => n204);
   U52 : OR3_X1 port map( A1 => B(55), A2 => B(56), A3 => n202, ZN => n200);
   U53 : OR2_X1 port map( A1 => n208, A2 => B(49), ZN => n209);
   U54 : OR2_X1 port map( A1 => n196, A2 => B(62), ZN => n195);
   U55 : NOR2_X1 port map( A1 => B(19), A2 => n241, ZN => n242);
   U56 : OR3_X1 port map( A1 => B(19), A2 => B(20), A3 => n241, ZN => n239);
   U57 : OR3_X1 port map( A1 => B(17), A2 => B(18), A3 => n243, ZN => n241);
   U58 : OR2_X1 port map( A1 => n243, A2 => B(17), ZN => n244);
   U59 : OR3_X1 port map( A1 => B(15), A2 => B(16), A3 => n245, ZN => n243);
   U60 : XNOR2_X1 port map( A => B(16), B => n246, ZN => DIFF_16_port);
   U61 : NOR2_X1 port map( A1 => B(15), A2 => n245, ZN => n246);
   U62 : NOR2_X1 port map( A1 => B(11), A2 => n249, ZN => n250);
   U63 : NOR2_X1 port map( A1 => B(7), A2 => n192, ZN => n191);
   U64 : NOR2_X1 port map( A1 => B(3), A2 => n211, ZN => n210);
   U65 : OR3_X1 port map( A1 => B(13), A2 => B(14), A3 => n247, ZN => n245);
   U66 : OR3_X1 port map( A1 => B(10), A2 => B(9), A3 => n190, ZN => n249);
   U67 : OR3_X1 port map( A1 => B(5), A2 => B(6), A3 => n194, ZN => n192);
   U68 : OR3_X1 port map( A1 => B(11), A2 => B(12), A3 => n249, ZN => n247);
   U69 : OR3_X1 port map( A1 => B(7), A2 => B(8), A3 => n192, ZN => n190);
   U70 : OR3_X1 port map( A1 => B(3), A2 => B(4), A3 => n211, ZN => n194);
   U71 : XNOR2_X1 port map( A => B(12), B => n250, ZN => DIFF_12_port);
   U72 : XNOR2_X1 port map( A => B(8), B => n191, ZN => DIFF_8_port);
   U73 : XNOR2_X1 port map( A => B(4), B => n210, ZN => DIFF_4_port);
   U74 : XNOR2_X1 port map( A => B(2), B => n232, ZN => DIFF_2_port);
   U75 : OR2_X1 port map( A1 => n247, A2 => B(13), ZN => n248);
   U76 : OR2_X1 port map( A1 => n190, A2 => B(9), ZN => n251);
   U77 : OR2_X1 port map( A1 => n194, A2 => B(5), ZN => n193);
   U78 : OR3_X1 port map( A1 => B(1), A2 => B(2), A3 => B(0), ZN => n211);
   U79 : NOR2_X1 port map( A1 => B(0), A2 => B(1), ZN => n232);
   U80 : INV_X1 port map( A => B(61), ZN => n189);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_17_DW01_sub_0 is

   port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (63 downto 0);  CO : out std_logic);

end complementer_N64_17_DW01_sub_0;

architecture SYN_rpl of complementer_N64_17_DW01_sub_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal DIFF_62_port, DIFF_63_port, DIFF_15_port, DIFF_16_port, DIFF_17_port,
      DIFF_18_port, DIFF_19_port, DIFF_20_port, DIFF_21_port, DIFF_22_port, 
      DIFF_23_port, DIFF_24_port, DIFF_25_port, DIFF_26_port, DIFF_27_port, 
      DIFF_28_port, DIFF_29_port, DIFF_30_port, DIFF_31_port, DIFF_32_port, 
      DIFF_33_port, DIFF_34_port, DIFF_35_port, DIFF_36_port, DIFF_37_port, 
      DIFF_38_port, DIFF_39_port, DIFF_40_port, DIFF_41_port, DIFF_42_port, 
      DIFF_43_port, DIFF_44_port, DIFF_45_port, DIFF_46_port, DIFF_47_port, 
      DIFF_48_port, DIFF_49_port, DIFF_50_port, DIFF_51_port, DIFF_52_port, 
      DIFF_53_port, DIFF_54_port, DIFF_55_port, DIFF_56_port, DIFF_57_port, 
      DIFF_58_port, DIFF_59_port, DIFF_60_port, DIFF_61_port, DIFF_3_port, 
      DIFF_4_port, DIFF_5_port, DIFF_6_port, DIFF_7_port, DIFF_8_port, 
      DIFF_9_port, DIFF_10_port, DIFF_11_port, DIFF_12_port, DIFF_13_port, 
      DIFF_14_port, DIFF_2_port, DIFF_1_port, n190, n191, n192, n194, n195, 
      n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, 
      n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, 
      n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, 
      n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, 
      n244, n245, n246, n247, n248, n249, n250, n189, n193, n251 : std_logic;

begin
   DIFF <= ( DIFF_63_port, DIFF_62_port, DIFF_61_port, DIFF_60_port, 
      DIFF_59_port, DIFF_58_port, DIFF_57_port, DIFF_56_port, DIFF_55_port, 
      DIFF_54_port, DIFF_53_port, DIFF_52_port, DIFF_51_port, DIFF_50_port, 
      DIFF_49_port, DIFF_48_port, DIFF_47_port, DIFF_46_port, DIFF_45_port, 
      DIFF_44_port, DIFF_43_port, DIFF_42_port, DIFF_41_port, DIFF_40_port, 
      DIFF_39_port, DIFF_38_port, DIFF_37_port, DIFF_36_port, DIFF_35_port, 
      DIFF_34_port, DIFF_33_port, DIFF_32_port, DIFF_31_port, DIFF_30_port, 
      DIFF_29_port, DIFF_28_port, DIFF_27_port, DIFF_26_port, DIFF_25_port, 
      DIFF_24_port, DIFF_23_port, DIFF_22_port, DIFF_21_port, DIFF_20_port, 
      DIFF_19_port, DIFF_18_port, DIFF_17_port, DIFF_16_port, DIFF_15_port, 
      DIFF_14_port, DIFF_13_port, DIFF_12_port, DIFF_11_port, DIFF_10_port, 
      DIFF_9_port, DIFF_8_port, DIFF_7_port, DIFF_6_port, DIFF_5_port, 
      DIFF_4_port, DIFF_3_port, DIFF_2_port, DIFF_1_port, B(0) );
   
   U81 : XOR2_X1 port map( A => n190, B => B(9), Z => DIFF_9_port);
   U82 : XOR2_X1 port map( A => n192, B => B(7), Z => DIFF_7_port);
   U84 : XOR2_X1 port map( A => n195, B => B(63), Z => DIFF_63_port);
   U85 : XOR2_X1 port map( A => n196, B => B(62), Z => DIFF_62_port);
   U86 : XOR2_X1 port map( A => n194, B => B(5), Z => DIFF_5_port);
   U87 : XOR2_X1 port map( A => n198, B => B(59), Z => DIFF_59_port);
   U88 : XOR2_X1 port map( A => n201, B => B(58), Z => DIFF_58_port);
   U89 : XOR2_X1 port map( A => n200, B => B(57), Z => DIFF_57_port);
   U90 : XOR2_X1 port map( A => n202, B => B(55), Z => DIFF_55_port);
   U91 : XOR2_X1 port map( A => n205, B => B(54), Z => DIFF_54_port);
   U92 : XOR2_X1 port map( A => n204, B => B(53), Z => DIFF_53_port);
   U93 : XOR2_X1 port map( A => n206, B => B(51), Z => DIFF_51_port);
   U94 : XOR2_X1 port map( A => n209, B => B(50), Z => DIFF_50_port);
   U95 : XOR2_X1 port map( A => n208, B => B(49), Z => DIFF_49_port);
   U96 : XOR2_X1 port map( A => n212, B => B(47), Z => DIFF_47_port);
   U97 : XOR2_X1 port map( A => n215, B => B(46), Z => DIFF_46_port);
   U98 : XOR2_X1 port map( A => n214, B => B(45), Z => DIFF_45_port);
   U99 : XOR2_X1 port map( A => n216, B => B(43), Z => DIFF_43_port);
   U100 : XOR2_X1 port map( A => n219, B => B(42), Z => DIFF_42_port);
   U101 : XOR2_X1 port map( A => n218, B => B(41), Z => DIFF_41_port);
   U102 : XOR2_X1 port map( A => n211, B => B(3), Z => DIFF_3_port);
   U103 : XOR2_X1 port map( A => n220, B => B(39), Z => DIFF_39_port);
   U104 : XOR2_X1 port map( A => n223, B => B(38), Z => DIFF_38_port);
   U105 : XOR2_X1 port map( A => n222, B => B(37), Z => DIFF_37_port);
   U106 : XOR2_X1 port map( A => n224, B => B(35), Z => DIFF_35_port);
   U107 : XOR2_X1 port map( A => n227, B => B(34), Z => DIFF_34_port);
   U108 : XOR2_X1 port map( A => n226, B => B(33), Z => DIFF_33_port);
   U109 : XOR2_X1 port map( A => n228, B => B(31), Z => DIFF_31_port);
   U110 : XOR2_X1 port map( A => n231, B => B(30), Z => DIFF_30_port);
   U111 : XOR2_X1 port map( A => n230, B => B(29), Z => DIFF_29_port);
   U112 : XOR2_X1 port map( A => n233, B => B(27), Z => DIFF_27_port);
   U113 : XOR2_X1 port map( A => n236, B => B(26), Z => DIFF_26_port);
   U114 : XOR2_X1 port map( A => n235, B => B(25), Z => DIFF_25_port);
   U115 : XOR2_X1 port map( A => n237, B => B(23), Z => DIFF_23_port);
   U116 : XOR2_X1 port map( A => n240, B => B(22), Z => DIFF_22_port);
   U117 : XOR2_X1 port map( A => n239, B => B(21), Z => DIFF_21_port);
   U118 : XOR2_X1 port map( A => B(1), B => B(0), Z => DIFF_1_port);
   U119 : XOR2_X1 port map( A => n241, B => B(19), Z => DIFF_19_port);
   U120 : XOR2_X1 port map( A => n244, B => B(18), Z => DIFF_18_port);
   U121 : XOR2_X1 port map( A => n243, B => B(17), Z => DIFF_17_port);
   U122 : XOR2_X1 port map( A => n245, B => B(15), Z => DIFF_15_port);
   U123 : XOR2_X1 port map( A => n248, B => B(14), Z => DIFF_14_port);
   U124 : XOR2_X1 port map( A => n247, B => B(13), Z => DIFF_13_port);
   U125 : XOR2_X1 port map( A => n249, B => B(11), Z => DIFF_11_port);
   U1 : NAND2_X1 port map( A1 => n197, A2 => n251, ZN => n196);
   U2 : OR2_X1 port map( A1 => n204, A2 => B(53), ZN => n205);
   U3 : NOR2_X1 port map( A1 => B(23), A2 => n237, ZN => n238);
   U4 : NOR2_X1 port map( A1 => B(19), A2 => n241, ZN => n242);
   U5 : OR3_X1 port map( A1 => B(21), A2 => B(22), A3 => n239, ZN => n237);
   U6 : OR3_X1 port map( A1 => B(23), A2 => B(24), A3 => n237, ZN => n235);
   U7 : OR3_X1 port map( A1 => B(19), A2 => B(20), A3 => n241, ZN => n239);
   U8 : XNOR2_X1 port map( A => B(28), B => n234, ZN => DIFF_28_port);
   U9 : XNOR2_X1 port map( A => B(24), B => n238, ZN => DIFF_24_port);
   U10 : XNOR2_X1 port map( A => B(20), B => n242, ZN => DIFF_20_port);
   U11 : OR2_X1 port map( A1 => n235, A2 => B(25), ZN => n236);
   U12 : OR2_X1 port map( A1 => n239, A2 => B(21), ZN => n240);
   U13 : NOR2_X1 port map( A1 => B(47), A2 => n212, ZN => n213);
   U14 : NOR2_X1 port map( A1 => B(51), A2 => n206, ZN => n207);
   U15 : NOR2_X1 port map( A1 => B(43), A2 => n216, ZN => n217);
   U16 : NOR2_X1 port map( A1 => B(39), A2 => n220, ZN => n221);
   U17 : NOR2_X1 port map( A1 => B(35), A2 => n224, ZN => n225);
   U18 : NOR2_X1 port map( A1 => B(31), A2 => n228, ZN => n229);
   U19 : NOR2_X1 port map( A1 => B(27), A2 => n233, ZN => n234);
   U20 : XNOR2_X1 port map( A => B(52), B => n207, ZN => DIFF_52_port);
   U21 : XNOR2_X1 port map( A => B(48), B => n213, ZN => DIFF_48_port);
   U22 : OR3_X1 port map( A1 => B(49), A2 => B(50), A3 => n208, ZN => n206);
   U23 : OR3_X1 port map( A1 => B(41), A2 => B(42), A3 => n218, ZN => n216);
   U24 : OR3_X1 port map( A1 => B(37), A2 => B(38), A3 => n222, ZN => n220);
   U25 : OR3_X1 port map( A1 => B(33), A2 => B(34), A3 => n226, ZN => n224);
   U26 : OR3_X1 port map( A1 => B(29), A2 => B(30), A3 => n230, ZN => n228);
   U27 : OR3_X1 port map( A1 => B(25), A2 => B(26), A3 => n235, ZN => n233);
   U28 : OR3_X1 port map( A1 => B(45), A2 => B(46), A3 => n214, ZN => n212);
   U29 : OR3_X1 port map( A1 => B(47), A2 => B(48), A3 => n212, ZN => n208);
   U30 : OR3_X1 port map( A1 => B(43), A2 => B(44), A3 => n216, ZN => n214);
   U31 : OR3_X1 port map( A1 => B(39), A2 => B(40), A3 => n220, ZN => n218);
   U32 : OR3_X1 port map( A1 => B(35), A2 => B(36), A3 => n224, ZN => n222);
   U33 : OR3_X1 port map( A1 => B(31), A2 => B(32), A3 => n228, ZN => n226);
   U34 : OR3_X1 port map( A1 => B(27), A2 => B(28), A3 => n233, ZN => n230);
   U35 : XNOR2_X1 port map( A => B(44), B => n217, ZN => DIFF_44_port);
   U36 : XNOR2_X1 port map( A => B(40), B => n221, ZN => DIFF_40_port);
   U37 : XNOR2_X1 port map( A => B(36), B => n225, ZN => DIFF_36_port);
   U38 : XNOR2_X1 port map( A => B(32), B => n229, ZN => DIFF_32_port);
   U39 : OR2_X1 port map( A1 => n214, A2 => B(45), ZN => n215);
   U40 : OR2_X1 port map( A1 => n208, A2 => B(49), ZN => n209);
   U41 : OR2_X1 port map( A1 => n218, A2 => B(41), ZN => n219);
   U42 : OR2_X1 port map( A1 => n222, A2 => B(37), ZN => n223);
   U43 : OR2_X1 port map( A1 => n226, A2 => B(33), ZN => n227);
   U44 : OR2_X1 port map( A1 => n230, A2 => B(29), ZN => n231);
   U45 : NOR3_X1 port map( A1 => B(59), A2 => B(60), A3 => n198, ZN => n197);
   U46 : XNOR2_X1 port map( A => n197, B => B(61), ZN => DIFF_61_port);
   U47 : XNOR2_X1 port map( A => B(60), B => n199, ZN => DIFF_60_port);
   U48 : NOR2_X1 port map( A1 => B(59), A2 => n198, ZN => n199);
   U49 : NOR2_X1 port map( A1 => B(55), A2 => n202, ZN => n203);
   U50 : OR3_X1 port map( A1 => B(57), A2 => B(58), A3 => n200, ZN => n198);
   U51 : OR3_X1 port map( A1 => B(53), A2 => B(54), A3 => n204, ZN => n202);
   U52 : OR3_X1 port map( A1 => B(51), A2 => B(52), A3 => n206, ZN => n204);
   U53 : OR3_X1 port map( A1 => B(55), A2 => B(56), A3 => n202, ZN => n200);
   U54 : XNOR2_X1 port map( A => B(56), B => n203, ZN => DIFF_56_port);
   U55 : OR2_X1 port map( A1 => n196, A2 => B(62), ZN => n195);
   U56 : OR2_X1 port map( A1 => n200, A2 => B(57), ZN => n201);
   U57 : OR3_X1 port map( A1 => B(17), A2 => B(18), A3 => n243, ZN => n241);
   U58 : XNOR2_X1 port map( A => B(16), B => n246, ZN => DIFF_16_port);
   U59 : OR2_X1 port map( A1 => n243, A2 => B(17), ZN => n244);
   U60 : NOR2_X1 port map( A1 => B(15), A2 => n245, ZN => n246);
   U61 : OR3_X1 port map( A1 => B(15), A2 => B(16), A3 => n245, ZN => n243);
   U62 : XNOR2_X1 port map( A => n189, B => B(10), ZN => DIFF_10_port);
   U63 : NOR2_X1 port map( A1 => n190, A2 => B(9), ZN => n189);
   U64 : XNOR2_X1 port map( A => n193, B => B(6), ZN => DIFF_6_port);
   U65 : NOR2_X1 port map( A1 => n194, A2 => B(5), ZN => n193);
   U66 : XNOR2_X1 port map( A => B(12), B => n250, ZN => DIFF_12_port);
   U67 : NOR2_X1 port map( A1 => B(11), A2 => n249, ZN => n250);
   U68 : XNOR2_X1 port map( A => B(8), B => n191, ZN => DIFF_8_port);
   U69 : NOR2_X1 port map( A1 => B(7), A2 => n192, ZN => n191);
   U70 : XNOR2_X1 port map( A => B(2), B => n232, ZN => DIFF_2_port);
   U71 : NOR2_X1 port map( A1 => B(0), A2 => B(1), ZN => n232);
   U72 : XNOR2_X1 port map( A => B(4), B => n210, ZN => DIFF_4_port);
   U73 : NOR2_X1 port map( A1 => B(3), A2 => n211, ZN => n210);
   U74 : OR3_X1 port map( A1 => B(5), A2 => B(6), A3 => n194, ZN => n192);
   U75 : OR3_X1 port map( A1 => B(10), A2 => B(9), A3 => n190, ZN => n249);
   U76 : OR3_X1 port map( A1 => B(13), A2 => B(14), A3 => n247, ZN => n245);
   U77 : OR3_X1 port map( A1 => B(7), A2 => B(8), A3 => n192, ZN => n190);
   U78 : OR3_X1 port map( A1 => B(11), A2 => B(12), A3 => n249, ZN => n247);
   U79 : OR3_X1 port map( A1 => B(3), A2 => B(4), A3 => n211, ZN => n194);
   U80 : OR2_X1 port map( A1 => n247, A2 => B(13), ZN => n248);
   U83 : OR3_X1 port map( A1 => B(1), A2 => B(2), A3 => B(0), ZN => n211);
   U126 : INV_X1 port map( A => B(61), ZN => n251);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_18_DW01_sub_0 is

   port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (63 downto 0);  CO : out std_logic);

end complementer_N64_18_DW01_sub_0;

architecture SYN_rpl of complementer_N64_18_DW01_sub_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal DIFF_62_port, DIFF_61_port, DIFF_60_port, DIFF_59_port, DIFF_58_port,
      DIFF_57_port, DIFF_56_port, DIFF_55_port, DIFF_54_port, DIFF_53_port, 
      DIFF_52_port, DIFF_51_port, DIFF_50_port, DIFF_49_port, DIFF_48_port, 
      DIFF_47_port, DIFF_46_port, DIFF_45_port, DIFF_44_port, DIFF_43_port, 
      DIFF_42_port, DIFF_41_port, DIFF_40_port, DIFF_39_port, DIFF_38_port, 
      DIFF_37_port, DIFF_36_port, DIFF_35_port, DIFF_34_port, DIFF_33_port, 
      DIFF_32_port, DIFF_31_port, DIFF_30_port, DIFF_29_port, DIFF_28_port, 
      DIFF_27_port, DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, 
      DIFF_22_port, DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, 
      DIFF_17_port, DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, 
      DIFF_12_port, DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, 
      DIFF_7_port, DIFF_6_port, DIFF_5_port, DIFF_4_port, DIFF_3_port, 
      DIFF_2_port, DIFF_1_port, DIFF_63_port, n190, n191, n192, n193, n194, 
      n196, n197, n198, n199, n200, n202, n203, n204, n206, n207, n208, n210, 
      n211, n212, n213, n214, n216, n217, n218, n220, n221, n222, n224, n225, 
      n226, n228, n229, n230, n232, n233, n234, n235, n237, n238, n239, n241, 
      n242, n243, n245, n246, n247, n249, n250, n251, n189, n195, n201, n205, 
      n209, n215, n219, n223, n227, n231, n236, n240, n244, n248 : std_logic;

begin
   DIFF <= ( DIFF_63_port, DIFF_62_port, DIFF_61_port, DIFF_60_port, 
      DIFF_59_port, DIFF_58_port, DIFF_57_port, DIFF_56_port, DIFF_55_port, 
      DIFF_54_port, DIFF_53_port, DIFF_52_port, DIFF_51_port, DIFF_50_port, 
      DIFF_49_port, DIFF_48_port, DIFF_47_port, DIFF_46_port, DIFF_45_port, 
      DIFF_44_port, DIFF_43_port, DIFF_42_port, DIFF_41_port, DIFF_40_port, 
      DIFF_39_port, DIFF_38_port, DIFF_37_port, DIFF_36_port, DIFF_35_port, 
      DIFF_34_port, DIFF_33_port, DIFF_32_port, DIFF_31_port, DIFF_30_port, 
      DIFF_29_port, DIFF_28_port, DIFF_27_port, DIFF_26_port, DIFF_25_port, 
      DIFF_24_port, DIFF_23_port, DIFF_22_port, DIFF_21_port, DIFF_20_port, 
      DIFF_19_port, DIFF_18_port, DIFF_17_port, DIFF_16_port, DIFF_15_port, 
      DIFF_14_port, DIFF_13_port, DIFF_12_port, DIFF_11_port, DIFF_10_port, 
      DIFF_9_port, DIFF_8_port, DIFF_7_port, DIFF_6_port, DIFF_5_port, 
      DIFF_4_port, DIFF_3_port, DIFF_2_port, DIFF_1_port, B(0) );
   
   U81 : XOR2_X1 port map( A => n190, B => B(9), Z => DIFF_9_port);
   U82 : XOR2_X1 port map( A => n192, B => B(7), Z => DIFF_7_port);
   U83 : XOR2_X1 port map( A => n193, B => B(6), Z => DIFF_6_port);
   U85 : XOR2_X1 port map( A => n196, B => B(62), Z => DIFF_62_port);
   U86 : XOR2_X1 port map( A => n194, B => B(5), Z => DIFF_5_port);
   U87 : XOR2_X1 port map( A => n198, B => B(59), Z => DIFF_59_port);
   U89 : XOR2_X1 port map( A => n200, B => B(57), Z => DIFF_57_port);
   U90 : XOR2_X1 port map( A => n202, B => B(55), Z => DIFF_55_port);
   U92 : XOR2_X1 port map( A => n204, B => B(53), Z => DIFF_53_port);
   U93 : XOR2_X1 port map( A => n206, B => B(51), Z => DIFF_51_port);
   U95 : XOR2_X1 port map( A => n208, B => B(49), Z => DIFF_49_port);
   U96 : XOR2_X1 port map( A => n212, B => B(47), Z => DIFF_47_port);
   U98 : XOR2_X1 port map( A => n214, B => B(45), Z => DIFF_45_port);
   U99 : XOR2_X1 port map( A => n216, B => B(43), Z => DIFF_43_port);
   U101 : XOR2_X1 port map( A => n218, B => B(41), Z => DIFF_41_port);
   U102 : XOR2_X1 port map( A => n211, B => B(3), Z => DIFF_3_port);
   U103 : XOR2_X1 port map( A => n220, B => B(39), Z => DIFF_39_port);
   U105 : XOR2_X1 port map( A => n222, B => B(37), Z => DIFF_37_port);
   U106 : XOR2_X1 port map( A => n224, B => B(35), Z => DIFF_35_port);
   U108 : XOR2_X1 port map( A => n226, B => B(33), Z => DIFF_33_port);
   U109 : XOR2_X1 port map( A => n228, B => B(31), Z => DIFF_31_port);
   U111 : XOR2_X1 port map( A => n230, B => B(29), Z => DIFF_29_port);
   U112 : XOR2_X1 port map( A => n233, B => B(27), Z => DIFF_27_port);
   U114 : XOR2_X1 port map( A => n235, B => B(25), Z => DIFF_25_port);
   U115 : XOR2_X1 port map( A => n237, B => B(23), Z => DIFF_23_port);
   U117 : XOR2_X1 port map( A => n239, B => B(21), Z => DIFF_21_port);
   U118 : XOR2_X1 port map( A => B(1), B => B(0), Z => DIFF_1_port);
   U119 : XOR2_X1 port map( A => n241, B => B(19), Z => DIFF_19_port);
   U121 : XOR2_X1 port map( A => n243, B => B(17), Z => DIFF_17_port);
   U122 : XOR2_X1 port map( A => n245, B => B(15), Z => DIFF_15_port);
   U124 : XOR2_X1 port map( A => n247, B => B(13), Z => DIFF_13_port);
   U125 : XOR2_X1 port map( A => n249, B => B(11), Z => DIFF_11_port);
   U126 : XOR2_X1 port map( A => n251, B => B(10), Z => DIFF_10_port);
   U1 : XOR2_X1 port map( A => n197, B => n248, Z => DIFF_61_port);
   U2 : NAND2_X1 port map( A1 => n197, A2 => n248, ZN => n196);
   U3 : XNOR2_X1 port map( A => n189, B => B(26), ZN => DIFF_26_port);
   U4 : NOR2_X1 port map( A1 => n235, A2 => B(25), ZN => n189);
   U5 : XNOR2_X1 port map( A => n195, B => B(22), ZN => DIFF_22_port);
   U6 : NOR2_X1 port map( A1 => n239, A2 => B(21), ZN => n195);
   U7 : XNOR2_X1 port map( A => B(28), B => n234, ZN => DIFF_28_port);
   U8 : NOR2_X1 port map( A1 => B(27), A2 => n233, ZN => n234);
   U9 : XNOR2_X1 port map( A => B(24), B => n238, ZN => DIFF_24_port);
   U10 : NOR2_X1 port map( A1 => B(23), A2 => n237, ZN => n238);
   U11 : XNOR2_X1 port map( A => B(20), B => n242, ZN => DIFF_20_port);
   U12 : NOR2_X1 port map( A1 => B(19), A2 => n241, ZN => n242);
   U13 : OR3_X1 port map( A1 => B(21), A2 => B(22), A3 => n239, ZN => n237);
   U14 : OR3_X1 port map( A1 => B(25), A2 => B(26), A3 => n235, ZN => n233);
   U15 : OR3_X1 port map( A1 => B(19), A2 => B(20), A3 => n241, ZN => n239);
   U16 : OR3_X1 port map( A1 => B(23), A2 => B(24), A3 => n237, ZN => n235);
   U17 : OR3_X1 port map( A1 => B(27), A2 => B(28), A3 => n233, ZN => n230);
   U18 : XNOR2_X1 port map( A => n201, B => B(46), ZN => DIFF_46_port);
   U19 : NOR2_X1 port map( A1 => n214, A2 => B(45), ZN => n201);
   U20 : XNOR2_X1 port map( A => n205, B => B(50), ZN => DIFF_50_port);
   U21 : NOR2_X1 port map( A1 => n208, A2 => B(49), ZN => n205);
   U22 : XNOR2_X1 port map( A => n209, B => B(54), ZN => DIFF_54_port);
   U23 : NOR2_X1 port map( A1 => n204, A2 => B(53), ZN => n209);
   U24 : XNOR2_X1 port map( A => B(40), B => n221, ZN => DIFF_40_port);
   U25 : NOR2_X1 port map( A1 => B(39), A2 => n220, ZN => n221);
   U26 : XNOR2_X1 port map( A => B(36), B => n225, ZN => DIFF_36_port);
   U27 : NOR2_X1 port map( A1 => B(35), A2 => n224, ZN => n225);
   U28 : XNOR2_X1 port map( A => B(32), B => n229, ZN => DIFF_32_port);
   U29 : NOR2_X1 port map( A1 => B(31), A2 => n228, ZN => n229);
   U30 : XNOR2_X1 port map( A => B(44), B => n217, ZN => DIFF_44_port);
   U31 : NOR2_X1 port map( A1 => B(43), A2 => n216, ZN => n217);
   U32 : XNOR2_X1 port map( A => B(52), B => n207, ZN => DIFF_52_port);
   U33 : NOR2_X1 port map( A1 => B(51), A2 => n206, ZN => n207);
   U34 : XNOR2_X1 port map( A => B(48), B => n213, ZN => DIFF_48_port);
   U35 : NOR2_X1 port map( A1 => B(47), A2 => n212, ZN => n213);
   U36 : OR3_X1 port map( A1 => B(29), A2 => B(30), A3 => n230, ZN => n228);
   U37 : OR3_X1 port map( A1 => B(33), A2 => B(34), A3 => n226, ZN => n224);
   U38 : OR3_X1 port map( A1 => B(37), A2 => B(38), A3 => n222, ZN => n220);
   U39 : OR3_X1 port map( A1 => B(41), A2 => B(42), A3 => n218, ZN => n216);
   U40 : OR3_X1 port map( A1 => B(49), A2 => B(50), A3 => n208, ZN => n206);
   U41 : OR3_X1 port map( A1 => B(45), A2 => B(46), A3 => n214, ZN => n212);
   U42 : OR3_X1 port map( A1 => B(53), A2 => B(54), A3 => n204, ZN => n202);
   U43 : OR3_X1 port map( A1 => B(47), A2 => B(48), A3 => n212, ZN => n208);
   U44 : OR3_X1 port map( A1 => B(51), A2 => B(52), A3 => n206, ZN => n204);
   U45 : OR3_X1 port map( A1 => B(31), A2 => B(32), A3 => n228, ZN => n226);
   U46 : OR3_X1 port map( A1 => B(35), A2 => B(36), A3 => n224, ZN => n222);
   U47 : OR3_X1 port map( A1 => B(39), A2 => B(40), A3 => n220, ZN => n218);
   U48 : OR3_X1 port map( A1 => B(43), A2 => B(44), A3 => n216, ZN => n214);
   U49 : XNOR2_X1 port map( A => n215, B => B(42), ZN => DIFF_42_port);
   U50 : NOR2_X1 port map( A1 => n218, A2 => B(41), ZN => n215);
   U51 : XNOR2_X1 port map( A => n219, B => B(38), ZN => DIFF_38_port);
   U52 : NOR2_X1 port map( A1 => n222, A2 => B(37), ZN => n219);
   U53 : XNOR2_X1 port map( A => n223, B => B(34), ZN => DIFF_34_port);
   U54 : NOR2_X1 port map( A1 => n226, A2 => B(33), ZN => n223);
   U55 : XNOR2_X1 port map( A => n227, B => B(30), ZN => DIFF_30_port);
   U56 : NOR2_X1 port map( A1 => n230, A2 => B(29), ZN => n227);
   U57 : NOR3_X1 port map( A1 => B(59), A2 => B(60), A3 => n198, ZN => n197);
   U58 : XNOR2_X1 port map( A => B(60), B => n199, ZN => DIFF_60_port);
   U59 : NOR2_X1 port map( A1 => B(59), A2 => n198, ZN => n199);
   U60 : XNOR2_X1 port map( A => B(56), B => n203, ZN => DIFF_56_port);
   U61 : NOR2_X1 port map( A1 => B(55), A2 => n202, ZN => n203);
   U62 : OR3_X1 port map( A1 => B(57), A2 => B(58), A3 => n200, ZN => n198);
   U63 : OR3_X1 port map( A1 => B(55), A2 => B(56), A3 => n202, ZN => n200);
   U64 : XNOR2_X1 port map( A => n231, B => B(58), ZN => DIFF_58_port);
   U65 : NOR2_X1 port map( A1 => n200, A2 => B(57), ZN => n231);
   U66 : XNOR2_X1 port map( A => n236, B => B(18), ZN => DIFF_18_port);
   U67 : NOR2_X1 port map( A1 => n243, A2 => B(17), ZN => n236);
   U68 : OR3_X1 port map( A1 => B(17), A2 => B(18), A3 => n243, ZN => n241);
   U69 : XNOR2_X1 port map( A => n240, B => B(63), ZN => DIFF_63_port);
   U70 : NOR2_X1 port map( A1 => n196, A2 => B(62), ZN => n240);
   U71 : XNOR2_X1 port map( A => B(16), B => n246, ZN => DIFF_16_port);
   U72 : NOR2_X1 port map( A1 => B(15), A2 => n245, ZN => n246);
   U73 : OR3_X1 port map( A1 => B(15), A2 => B(16), A3 => n245, ZN => n243);
   U74 : XNOR2_X1 port map( A => n244, B => B(14), ZN => DIFF_14_port);
   U75 : NOR2_X1 port map( A1 => n247, A2 => B(13), ZN => n244);
   U76 : OR3_X1 port map( A1 => B(13), A2 => B(14), A3 => n247, ZN => n245);
   U77 : NOR2_X1 port map( A1 => B(11), A2 => n249, ZN => n250);
   U78 : NOR2_X1 port map( A1 => B(7), A2 => n192, ZN => n191);
   U79 : NOR2_X1 port map( A1 => B(3), A2 => n211, ZN => n210);
   U80 : OR3_X1 port map( A1 => B(10), A2 => B(9), A3 => n190, ZN => n249);
   U84 : OR3_X1 port map( A1 => B(5), A2 => B(6), A3 => n194, ZN => n192);
   U88 : OR3_X1 port map( A1 => B(11), A2 => B(12), A3 => n249, ZN => n247);
   U91 : OR3_X1 port map( A1 => B(7), A2 => B(8), A3 => n192, ZN => n190);
   U94 : OR3_X1 port map( A1 => B(3), A2 => B(4), A3 => n211, ZN => n194);
   U97 : XNOR2_X1 port map( A => B(12), B => n250, ZN => DIFF_12_port);
   U100 : XNOR2_X1 port map( A => B(8), B => n191, ZN => DIFF_8_port);
   U104 : XNOR2_X1 port map( A => B(4), B => n210, ZN => DIFF_4_port);
   U107 : XNOR2_X1 port map( A => B(2), B => n232, ZN => DIFF_2_port);
   U110 : OR2_X1 port map( A1 => n190, A2 => B(9), ZN => n251);
   U113 : OR2_X1 port map( A1 => n194, A2 => B(5), ZN => n193);
   U116 : OR3_X1 port map( A1 => B(1), A2 => B(2), A3 => B(0), ZN => n211);
   U120 : NOR2_X1 port map( A1 => B(0), A2 => B(1), ZN => n232);
   U123 : INV_X1 port map( A => B(61), ZN => n248);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_19_DW01_sub_0 is

   port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (63 downto 0);  CO : out std_logic);

end complementer_N64_19_DW01_sub_0;

architecture SYN_rpl of complementer_N64_19_DW01_sub_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal DIFF_62_port, DIFF_63_port, DIFF_13_port, DIFF_14_port, DIFF_15_port,
      DIFF_16_port, DIFF_17_port, DIFF_18_port, DIFF_19_port, DIFF_20_port, 
      DIFF_21_port, DIFF_22_port, DIFF_23_port, DIFF_24_port, DIFF_25_port, 
      DIFF_26_port, DIFF_27_port, DIFF_28_port, DIFF_29_port, DIFF_30_port, 
      DIFF_31_port, DIFF_32_port, DIFF_33_port, DIFF_34_port, DIFF_35_port, 
      DIFF_36_port, DIFF_37_port, DIFF_38_port, DIFF_39_port, DIFF_40_port, 
      DIFF_41_port, DIFF_42_port, DIFF_43_port, DIFF_44_port, DIFF_45_port, 
      DIFF_46_port, DIFF_47_port, DIFF_48_port, DIFF_49_port, DIFF_50_port, 
      DIFF_51_port, DIFF_52_port, DIFF_53_port, DIFF_54_port, DIFF_55_port, 
      DIFF_56_port, DIFF_57_port, DIFF_58_port, DIFF_59_port, DIFF_60_port, 
      DIFF_61_port, DIFF_3_port, DIFF_4_port, DIFF_5_port, DIFF_6_port, 
      DIFF_7_port, DIFF_8_port, DIFF_9_port, DIFF_10_port, DIFF_11_port, 
      DIFF_12_port, DIFF_2_port, DIFF_1_port, n190, n191, n192, n194, n195, 
      n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, 
      n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, 
      n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, 
      n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, 
      n244, n245, n246, n247, n248, n249, n250, n189, n193, n251 : std_logic;

begin
   DIFF <= ( DIFF_63_port, DIFF_62_port, DIFF_61_port, DIFF_60_port, 
      DIFF_59_port, DIFF_58_port, DIFF_57_port, DIFF_56_port, DIFF_55_port, 
      DIFF_54_port, DIFF_53_port, DIFF_52_port, DIFF_51_port, DIFF_50_port, 
      DIFF_49_port, DIFF_48_port, DIFF_47_port, DIFF_46_port, DIFF_45_port, 
      DIFF_44_port, DIFF_43_port, DIFF_42_port, DIFF_41_port, DIFF_40_port, 
      DIFF_39_port, DIFF_38_port, DIFF_37_port, DIFF_36_port, DIFF_35_port, 
      DIFF_34_port, DIFF_33_port, DIFF_32_port, DIFF_31_port, DIFF_30_port, 
      DIFF_29_port, DIFF_28_port, DIFF_27_port, DIFF_26_port, DIFF_25_port, 
      DIFF_24_port, DIFF_23_port, DIFF_22_port, DIFF_21_port, DIFF_20_port, 
      DIFF_19_port, DIFF_18_port, DIFF_17_port, DIFF_16_port, DIFF_15_port, 
      DIFF_14_port, DIFF_13_port, DIFF_12_port, DIFF_11_port, DIFF_10_port, 
      DIFF_9_port, DIFF_8_port, DIFF_7_port, DIFF_6_port, DIFF_5_port, 
      DIFF_4_port, DIFF_3_port, DIFF_2_port, DIFF_1_port, B(0) );
   
   U81 : XOR2_X1 port map( A => n190, B => B(9), Z => DIFF_9_port);
   U82 : XOR2_X1 port map( A => n192, B => B(7), Z => DIFF_7_port);
   U84 : XOR2_X1 port map( A => n195, B => B(63), Z => DIFF_63_port);
   U85 : XOR2_X1 port map( A => n196, B => B(62), Z => DIFF_62_port);
   U86 : XOR2_X1 port map( A => n194, B => B(5), Z => DIFF_5_port);
   U87 : XOR2_X1 port map( A => n198, B => B(59), Z => DIFF_59_port);
   U88 : XOR2_X1 port map( A => n201, B => B(58), Z => DIFF_58_port);
   U89 : XOR2_X1 port map( A => n200, B => B(57), Z => DIFF_57_port);
   U90 : XOR2_X1 port map( A => n202, B => B(55), Z => DIFF_55_port);
   U91 : XOR2_X1 port map( A => n205, B => B(54), Z => DIFF_54_port);
   U92 : XOR2_X1 port map( A => n204, B => B(53), Z => DIFF_53_port);
   U93 : XOR2_X1 port map( A => n206, B => B(51), Z => DIFF_51_port);
   U94 : XOR2_X1 port map( A => n209, B => B(50), Z => DIFF_50_port);
   U95 : XOR2_X1 port map( A => n208, B => B(49), Z => DIFF_49_port);
   U96 : XOR2_X1 port map( A => n212, B => B(47), Z => DIFF_47_port);
   U97 : XOR2_X1 port map( A => n215, B => B(46), Z => DIFF_46_port);
   U98 : XOR2_X1 port map( A => n214, B => B(45), Z => DIFF_45_port);
   U99 : XOR2_X1 port map( A => n216, B => B(43), Z => DIFF_43_port);
   U100 : XOR2_X1 port map( A => n219, B => B(42), Z => DIFF_42_port);
   U101 : XOR2_X1 port map( A => n218, B => B(41), Z => DIFF_41_port);
   U102 : XOR2_X1 port map( A => n211, B => B(3), Z => DIFF_3_port);
   U103 : XOR2_X1 port map( A => n220, B => B(39), Z => DIFF_39_port);
   U104 : XOR2_X1 port map( A => n223, B => B(38), Z => DIFF_38_port);
   U105 : XOR2_X1 port map( A => n222, B => B(37), Z => DIFF_37_port);
   U106 : XOR2_X1 port map( A => n224, B => B(35), Z => DIFF_35_port);
   U107 : XOR2_X1 port map( A => n227, B => B(34), Z => DIFF_34_port);
   U108 : XOR2_X1 port map( A => n226, B => B(33), Z => DIFF_33_port);
   U109 : XOR2_X1 port map( A => n228, B => B(31), Z => DIFF_31_port);
   U110 : XOR2_X1 port map( A => n231, B => B(30), Z => DIFF_30_port);
   U111 : XOR2_X1 port map( A => n230, B => B(29), Z => DIFF_29_port);
   U112 : XOR2_X1 port map( A => n233, B => B(27), Z => DIFF_27_port);
   U113 : XOR2_X1 port map( A => n236, B => B(26), Z => DIFF_26_port);
   U114 : XOR2_X1 port map( A => n235, B => B(25), Z => DIFF_25_port);
   U115 : XOR2_X1 port map( A => n237, B => B(23), Z => DIFF_23_port);
   U116 : XOR2_X1 port map( A => n240, B => B(22), Z => DIFF_22_port);
   U117 : XOR2_X1 port map( A => n239, B => B(21), Z => DIFF_21_port);
   U118 : XOR2_X1 port map( A => B(1), B => B(0), Z => DIFF_1_port);
   U119 : XOR2_X1 port map( A => n241, B => B(19), Z => DIFF_19_port);
   U120 : XOR2_X1 port map( A => n244, B => B(18), Z => DIFF_18_port);
   U121 : XOR2_X1 port map( A => n243, B => B(17), Z => DIFF_17_port);
   U122 : XOR2_X1 port map( A => n245, B => B(15), Z => DIFF_15_port);
   U123 : XOR2_X1 port map( A => n248, B => B(14), Z => DIFF_14_port);
   U124 : XOR2_X1 port map( A => n247, B => B(13), Z => DIFF_13_port);
   U125 : XOR2_X1 port map( A => n249, B => B(11), Z => DIFF_11_port);
   U1 : NAND2_X1 port map( A1 => n197, A2 => n251, ZN => n196);
   U2 : NOR2_X1 port map( A1 => B(31), A2 => n228, ZN => n229);
   U3 : NOR2_X1 port map( A1 => B(27), A2 => n233, ZN => n234);
   U4 : NOR2_X1 port map( A1 => B(23), A2 => n237, ZN => n238);
   U5 : NOR2_X1 port map( A1 => B(19), A2 => n241, ZN => n242);
   U6 : OR3_X1 port map( A1 => B(29), A2 => B(30), A3 => n230, ZN => n228);
   U7 : OR3_X1 port map( A1 => B(25), A2 => B(26), A3 => n235, ZN => n233);
   U8 : OR3_X1 port map( A1 => B(21), A2 => B(22), A3 => n239, ZN => n237);
   U9 : OR3_X1 port map( A1 => B(17), A2 => B(18), A3 => n243, ZN => n241);
   U10 : OR3_X1 port map( A1 => B(31), A2 => B(32), A3 => n228, ZN => n226);
   U11 : OR3_X1 port map( A1 => B(27), A2 => B(28), A3 => n233, ZN => n230);
   U12 : OR3_X1 port map( A1 => B(23), A2 => B(24), A3 => n237, ZN => n235);
   U13 : OR3_X1 port map( A1 => B(19), A2 => B(20), A3 => n241, ZN => n239);
   U14 : XNOR2_X1 port map( A => B(36), B => n225, ZN => DIFF_36_port);
   U15 : XNOR2_X1 port map( A => B(32), B => n229, ZN => DIFF_32_port);
   U16 : XNOR2_X1 port map( A => B(28), B => n234, ZN => DIFF_28_port);
   U17 : XNOR2_X1 port map( A => B(24), B => n238, ZN => DIFF_24_port);
   U18 : XNOR2_X1 port map( A => B(20), B => n242, ZN => DIFF_20_port);
   U19 : XNOR2_X1 port map( A => B(16), B => n246, ZN => DIFF_16_port);
   U20 : OR2_X1 port map( A1 => n230, A2 => B(29), ZN => n231);
   U21 : OR2_X1 port map( A1 => n235, A2 => B(25), ZN => n236);
   U22 : OR2_X1 port map( A1 => n239, A2 => B(21), ZN => n240);
   U23 : OR2_X1 port map( A1 => n243, A2 => B(17), ZN => n244);
   U24 : XNOR2_X1 port map( A => B(60), B => n199, ZN => DIFF_60_port);
   U25 : NOR2_X1 port map( A1 => B(43), A2 => n216, ZN => n217);
   U26 : NOR2_X1 port map( A1 => B(51), A2 => n206, ZN => n207);
   U27 : NOR2_X1 port map( A1 => B(39), A2 => n220, ZN => n221);
   U28 : NOR2_X1 port map( A1 => B(35), A2 => n224, ZN => n225);
   U29 : NOR2_X1 port map( A1 => B(59), A2 => n198, ZN => n199);
   U30 : NOR2_X1 port map( A1 => B(55), A2 => n202, ZN => n203);
   U31 : OR3_X1 port map( A1 => B(49), A2 => B(50), A3 => n208, ZN => n206);
   U32 : OR3_X1 port map( A1 => B(41), A2 => B(42), A3 => n218, ZN => n216);
   U33 : OR3_X1 port map( A1 => B(37), A2 => B(38), A3 => n222, ZN => n220);
   U34 : OR3_X1 port map( A1 => B(33), A2 => B(34), A3 => n226, ZN => n224);
   U35 : OR3_X1 port map( A1 => B(53), A2 => B(54), A3 => n204, ZN => n202);
   U36 : OR3_X1 port map( A1 => B(39), A2 => B(40), A3 => n220, ZN => n218);
   U37 : OR3_X1 port map( A1 => B(35), A2 => B(36), A3 => n224, ZN => n222);
   U38 : OR3_X1 port map( A1 => B(43), A2 => B(44), A3 => n216, ZN => n214);
   U39 : OR3_X1 port map( A1 => B(51), A2 => B(52), A3 => n206, ZN => n204);
   U40 : XNOR2_X1 port map( A => B(48), B => n213, ZN => DIFF_48_port);
   U41 : XNOR2_X1 port map( A => B(40), B => n221, ZN => DIFF_40_port);
   U42 : XNOR2_X1 port map( A => B(44), B => n217, ZN => DIFF_44_port);
   U43 : OR2_X1 port map( A1 => n214, A2 => B(45), ZN => n215);
   U44 : OR2_X1 port map( A1 => n208, A2 => B(49), ZN => n209);
   U45 : OR2_X1 port map( A1 => n218, A2 => B(41), ZN => n219);
   U46 : OR2_X1 port map( A1 => n222, A2 => B(37), ZN => n223);
   U47 : OR2_X1 port map( A1 => n226, A2 => B(33), ZN => n227);
   U48 : OR2_X1 port map( A1 => n204, A2 => B(53), ZN => n205);
   U49 : NOR3_X1 port map( A1 => B(59), A2 => B(60), A3 => n198, ZN => n197);
   U50 : NOR2_X1 port map( A1 => B(15), A2 => n245, ZN => n246);
   U51 : OR3_X1 port map( A1 => B(15), A2 => B(16), A3 => n245, ZN => n243);
   U52 : XNOR2_X1 port map( A => n197, B => B(61), ZN => DIFF_61_port);
   U53 : NOR2_X1 port map( A1 => B(47), A2 => n212, ZN => n213);
   U54 : XNOR2_X1 port map( A => B(52), B => n207, ZN => DIFF_52_port);
   U55 : OR3_X1 port map( A1 => B(57), A2 => B(58), A3 => n200, ZN => n198);
   U56 : OR3_X1 port map( A1 => B(45), A2 => B(46), A3 => n214, ZN => n212);
   U57 : OR3_X1 port map( A1 => B(47), A2 => B(48), A3 => n212, ZN => n208);
   U58 : OR3_X1 port map( A1 => B(55), A2 => B(56), A3 => n202, ZN => n200);
   U59 : XNOR2_X1 port map( A => B(56), B => n203, ZN => DIFF_56_port);
   U60 : OR2_X1 port map( A1 => n200, A2 => B(57), ZN => n201);
   U61 : OR2_X1 port map( A1 => n196, A2 => B(62), ZN => n195);
   U62 : OR3_X1 port map( A1 => B(13), A2 => B(14), A3 => n247, ZN => n245);
   U63 : OR2_X1 port map( A1 => n247, A2 => B(13), ZN => n248);
   U64 : XNOR2_X1 port map( A => B(12), B => n250, ZN => DIFF_12_port);
   U65 : XNOR2_X1 port map( A => n189, B => B(10), ZN => DIFF_10_port);
   U66 : NOR2_X1 port map( A1 => n190, A2 => B(9), ZN => n189);
   U67 : XNOR2_X1 port map( A => n193, B => B(6), ZN => DIFF_6_port);
   U68 : NOR2_X1 port map( A1 => n194, A2 => B(5), ZN => n193);
   U69 : NOR2_X1 port map( A1 => B(11), A2 => n249, ZN => n250);
   U70 : XNOR2_X1 port map( A => B(8), B => n191, ZN => DIFF_8_port);
   U71 : NOR2_X1 port map( A1 => B(7), A2 => n192, ZN => n191);
   U72 : XNOR2_X1 port map( A => B(2), B => n232, ZN => DIFF_2_port);
   U73 : NOR2_X1 port map( A1 => B(0), A2 => B(1), ZN => n232);
   U74 : XNOR2_X1 port map( A => B(4), B => n210, ZN => DIFF_4_port);
   U75 : NOR2_X1 port map( A1 => B(3), A2 => n211, ZN => n210);
   U76 : OR3_X1 port map( A1 => B(5), A2 => B(6), A3 => n194, ZN => n192);
   U77 : OR3_X1 port map( A1 => B(10), A2 => B(9), A3 => n190, ZN => n249);
   U78 : OR3_X1 port map( A1 => B(7), A2 => B(8), A3 => n192, ZN => n190);
   U79 : OR3_X1 port map( A1 => B(11), A2 => B(12), A3 => n249, ZN => n247);
   U80 : OR3_X1 port map( A1 => B(3), A2 => B(4), A3 => n211, ZN => n194);
   U83 : OR3_X1 port map( A1 => B(1), A2 => B(2), A3 => B(0), ZN => n211);
   U126 : INV_X1 port map( A => B(61), ZN => n251);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_20_DW01_sub_0 is

   port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (63 downto 0);  CO : out std_logic);

end complementer_N64_20_DW01_sub_0;

architecture SYN_rpl of complementer_N64_20_DW01_sub_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal DIFF_62_port, DIFF_61_port, DIFF_60_port, DIFF_59_port, DIFF_58_port,
      DIFF_57_port, DIFF_56_port, DIFF_55_port, DIFF_54_port, DIFF_53_port, 
      DIFF_52_port, DIFF_51_port, DIFF_50_port, DIFF_49_port, DIFF_48_port, 
      DIFF_47_port, DIFF_46_port, DIFF_45_port, DIFF_44_port, DIFF_43_port, 
      DIFF_42_port, DIFF_41_port, DIFF_40_port, DIFF_39_port, DIFF_38_port, 
      DIFF_37_port, DIFF_36_port, DIFF_35_port, DIFF_34_port, DIFF_33_port, 
      DIFF_32_port, DIFF_31_port, DIFF_30_port, DIFF_29_port, DIFF_28_port, 
      DIFF_27_port, DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, 
      DIFF_22_port, DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, 
      DIFF_17_port, DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, 
      DIFF_12_port, DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, 
      DIFF_7_port, DIFF_6_port, DIFF_5_port, DIFF_4_port, DIFF_3_port, 
      DIFF_2_port, DIFF_1_port, DIFF_63_port, n190, n191, n192, n193, n194, 
      n196, n197, n198, n199, n200, n202, n203, n204, n206, n207, n208, n210, 
      n211, n212, n213, n214, n216, n217, n218, n220, n221, n222, n224, n225, 
      n226, n228, n229, n230, n232, n233, n234, n235, n237, n238, n239, n241, 
      n242, n243, n245, n246, n247, n249, n250, n251, n189, n195, n201, n205, 
      n209, n215, n219, n223, n227, n231, n236, n240, n244, n248 : std_logic;

begin
   DIFF <= ( DIFF_63_port, DIFF_62_port, DIFF_61_port, DIFF_60_port, 
      DIFF_59_port, DIFF_58_port, DIFF_57_port, DIFF_56_port, DIFF_55_port, 
      DIFF_54_port, DIFF_53_port, DIFF_52_port, DIFF_51_port, DIFF_50_port, 
      DIFF_49_port, DIFF_48_port, DIFF_47_port, DIFF_46_port, DIFF_45_port, 
      DIFF_44_port, DIFF_43_port, DIFF_42_port, DIFF_41_port, DIFF_40_port, 
      DIFF_39_port, DIFF_38_port, DIFF_37_port, DIFF_36_port, DIFF_35_port, 
      DIFF_34_port, DIFF_33_port, DIFF_32_port, DIFF_31_port, DIFF_30_port, 
      DIFF_29_port, DIFF_28_port, DIFF_27_port, DIFF_26_port, DIFF_25_port, 
      DIFF_24_port, DIFF_23_port, DIFF_22_port, DIFF_21_port, DIFF_20_port, 
      DIFF_19_port, DIFF_18_port, DIFF_17_port, DIFF_16_port, DIFF_15_port, 
      DIFF_14_port, DIFF_13_port, DIFF_12_port, DIFF_11_port, DIFF_10_port, 
      DIFF_9_port, DIFF_8_port, DIFF_7_port, DIFF_6_port, DIFF_5_port, 
      DIFF_4_port, DIFF_3_port, DIFF_2_port, DIFF_1_port, B(0) );
   
   U81 : XOR2_X1 port map( A => n190, B => B(9), Z => DIFF_9_port);
   U82 : XOR2_X1 port map( A => n192, B => B(7), Z => DIFF_7_port);
   U83 : XOR2_X1 port map( A => n193, B => B(6), Z => DIFF_6_port);
   U85 : XOR2_X1 port map( A => n196, B => B(62), Z => DIFF_62_port);
   U86 : XOR2_X1 port map( A => n194, B => B(5), Z => DIFF_5_port);
   U87 : XOR2_X1 port map( A => n198, B => B(59), Z => DIFF_59_port);
   U89 : XOR2_X1 port map( A => n200, B => B(57), Z => DIFF_57_port);
   U90 : XOR2_X1 port map( A => n202, B => B(55), Z => DIFF_55_port);
   U92 : XOR2_X1 port map( A => n204, B => B(53), Z => DIFF_53_port);
   U93 : XOR2_X1 port map( A => n206, B => B(51), Z => DIFF_51_port);
   U95 : XOR2_X1 port map( A => n208, B => B(49), Z => DIFF_49_port);
   U96 : XOR2_X1 port map( A => n212, B => B(47), Z => DIFF_47_port);
   U98 : XOR2_X1 port map( A => n214, B => B(45), Z => DIFF_45_port);
   U99 : XOR2_X1 port map( A => n216, B => B(43), Z => DIFF_43_port);
   U101 : XOR2_X1 port map( A => n218, B => B(41), Z => DIFF_41_port);
   U102 : XOR2_X1 port map( A => n211, B => B(3), Z => DIFF_3_port);
   U103 : XOR2_X1 port map( A => n220, B => B(39), Z => DIFF_39_port);
   U105 : XOR2_X1 port map( A => n222, B => B(37), Z => DIFF_37_port);
   U106 : XOR2_X1 port map( A => n224, B => B(35), Z => DIFF_35_port);
   U108 : XOR2_X1 port map( A => n226, B => B(33), Z => DIFF_33_port);
   U109 : XOR2_X1 port map( A => n228, B => B(31), Z => DIFF_31_port);
   U111 : XOR2_X1 port map( A => n230, B => B(29), Z => DIFF_29_port);
   U112 : XOR2_X1 port map( A => n233, B => B(27), Z => DIFF_27_port);
   U114 : XOR2_X1 port map( A => n235, B => B(25), Z => DIFF_25_port);
   U115 : XOR2_X1 port map( A => n237, B => B(23), Z => DIFF_23_port);
   U117 : XOR2_X1 port map( A => n239, B => B(21), Z => DIFF_21_port);
   U118 : XOR2_X1 port map( A => B(1), B => B(0), Z => DIFF_1_port);
   U119 : XOR2_X1 port map( A => n241, B => B(19), Z => DIFF_19_port);
   U121 : XOR2_X1 port map( A => n243, B => B(17), Z => DIFF_17_port);
   U122 : XOR2_X1 port map( A => n245, B => B(15), Z => DIFF_15_port);
   U124 : XOR2_X1 port map( A => n247, B => B(13), Z => DIFF_13_port);
   U125 : XOR2_X1 port map( A => n249, B => B(11), Z => DIFF_11_port);
   U126 : XOR2_X1 port map( A => n251, B => B(10), Z => DIFF_10_port);
   U1 : XNOR2_X1 port map( A => n189, B => B(34), ZN => DIFF_34_port);
   U2 : NOR2_X1 port map( A1 => n226, A2 => B(33), ZN => n189);
   U3 : XNOR2_X1 port map( A => n195, B => B(30), ZN => DIFF_30_port);
   U4 : NOR2_X1 port map( A1 => n230, A2 => B(29), ZN => n195);
   U5 : XNOR2_X1 port map( A => n201, B => B(26), ZN => DIFF_26_port);
   U6 : NOR2_X1 port map( A1 => n235, A2 => B(25), ZN => n201);
   U7 : XNOR2_X1 port map( A => n205, B => B(22), ZN => DIFF_22_port);
   U8 : NOR2_X1 port map( A1 => n239, A2 => B(21), ZN => n205);
   U9 : XNOR2_X1 port map( A => n209, B => B(18), ZN => DIFF_18_port);
   U10 : NOR2_X1 port map( A1 => n243, A2 => B(17), ZN => n209);
   U11 : XNOR2_X1 port map( A => B(36), B => n225, ZN => DIFF_36_port);
   U12 : NOR2_X1 port map( A1 => B(35), A2 => n224, ZN => n225);
   U13 : XNOR2_X1 port map( A => B(32), B => n229, ZN => DIFF_32_port);
   U14 : NOR2_X1 port map( A1 => B(31), A2 => n228, ZN => n229);
   U15 : XNOR2_X1 port map( A => B(28), B => n234, ZN => DIFF_28_port);
   U16 : NOR2_X1 port map( A1 => B(27), A2 => n233, ZN => n234);
   U17 : XNOR2_X1 port map( A => B(24), B => n238, ZN => DIFF_24_port);
   U18 : NOR2_X1 port map( A1 => B(23), A2 => n237, ZN => n238);
   U19 : XNOR2_X1 port map( A => B(20), B => n242, ZN => DIFF_20_port);
   U20 : NOR2_X1 port map( A1 => B(19), A2 => n241, ZN => n242);
   U21 : OR3_X1 port map( A1 => B(17), A2 => B(18), A3 => n243, ZN => n241);
   U22 : OR3_X1 port map( A1 => B(21), A2 => B(22), A3 => n239, ZN => n237);
   U23 : OR3_X1 port map( A1 => B(25), A2 => B(26), A3 => n235, ZN => n233);
   U24 : OR3_X1 port map( A1 => B(29), A2 => B(30), A3 => n230, ZN => n228);
   U25 : OR3_X1 port map( A1 => B(33), A2 => B(34), A3 => n226, ZN => n224);
   U26 : OR3_X1 port map( A1 => B(19), A2 => B(20), A3 => n241, ZN => n239);
   U27 : OR3_X1 port map( A1 => B(23), A2 => B(24), A3 => n237, ZN => n235);
   U28 : OR3_X1 port map( A1 => B(27), A2 => B(28), A3 => n233, ZN => n230);
   U29 : OR3_X1 port map( A1 => B(31), A2 => B(32), A3 => n228, ZN => n226);
   U30 : NOR3_X1 port map( A1 => B(59), A2 => B(60), A3 => n198, ZN => n197);
   U31 : XNOR2_X1 port map( A => n215, B => B(42), ZN => DIFF_42_port);
   U32 : NOR2_X1 port map( A1 => n218, A2 => B(41), ZN => n215);
   U33 : XNOR2_X1 port map( A => n219, B => B(50), ZN => DIFF_50_port);
   U34 : NOR2_X1 port map( A1 => n208, A2 => B(49), ZN => n219);
   U35 : XNOR2_X1 port map( A => n223, B => B(38), ZN => DIFF_38_port);
   U36 : NOR2_X1 port map( A1 => n222, A2 => B(37), ZN => n223);
   U37 : XNOR2_X1 port map( A => n227, B => B(54), ZN => DIFF_54_port);
   U38 : NOR2_X1 port map( A1 => n204, A2 => B(53), ZN => n227);
   U39 : XNOR2_X1 port map( A => B(40), B => n221, ZN => DIFF_40_port);
   U40 : NOR2_X1 port map( A1 => B(39), A2 => n220, ZN => n221);
   U41 : XNOR2_X1 port map( A => B(44), B => n217, ZN => DIFF_44_port);
   U42 : NOR2_X1 port map( A1 => B(43), A2 => n216, ZN => n217);
   U43 : XNOR2_X1 port map( A => B(48), B => n213, ZN => DIFF_48_port);
   U44 : NOR2_X1 port map( A1 => B(47), A2 => n212, ZN => n213);
   U45 : XNOR2_X1 port map( A => B(60), B => n199, ZN => DIFF_60_port);
   U46 : NOR2_X1 port map( A1 => B(59), A2 => n198, ZN => n199);
   U47 : XOR2_X1 port map( A => n197, B => n248, Z => DIFF_61_port);
   U48 : NAND2_X1 port map( A1 => n197, A2 => n248, ZN => n196);
   U49 : OR3_X1 port map( A1 => B(57), A2 => B(58), A3 => n200, ZN => n198);
   U50 : OR3_X1 port map( A1 => B(49), A2 => B(50), A3 => n208, ZN => n206);
   U51 : OR3_X1 port map( A1 => B(37), A2 => B(38), A3 => n222, ZN => n220);
   U52 : OR3_X1 port map( A1 => B(41), A2 => B(42), A3 => n218, ZN => n216);
   U53 : OR3_X1 port map( A1 => B(53), A2 => B(54), A3 => n204, ZN => n202);
   U54 : OR3_X1 port map( A1 => B(35), A2 => B(36), A3 => n224, ZN => n222);
   U55 : OR3_X1 port map( A1 => B(39), A2 => B(40), A3 => n220, ZN => n218);
   U56 : OR3_X1 port map( A1 => B(47), A2 => B(48), A3 => n212, ZN => n208);
   U57 : OR3_X1 port map( A1 => B(43), A2 => B(44), A3 => n216, ZN => n214);
   U58 : XNOR2_X1 port map( A => n231, B => B(58), ZN => DIFF_58_port);
   U59 : NOR2_X1 port map( A1 => n200, A2 => B(57), ZN => n231);
   U60 : XNOR2_X1 port map( A => B(16), B => n246, ZN => DIFF_16_port);
   U61 : NOR2_X1 port map( A1 => B(15), A2 => n245, ZN => n246);
   U62 : OR3_X1 port map( A1 => B(15), A2 => B(16), A3 => n245, ZN => n243);
   U63 : XNOR2_X1 port map( A => n236, B => B(63), ZN => DIFF_63_port);
   U64 : NOR2_X1 port map( A1 => n196, A2 => B(62), ZN => n236);
   U65 : XNOR2_X1 port map( A => n240, B => B(46), ZN => DIFF_46_port);
   U66 : NOR2_X1 port map( A1 => n214, A2 => B(45), ZN => n240);
   U67 : XNOR2_X1 port map( A => B(52), B => n207, ZN => DIFF_52_port);
   U68 : NOR2_X1 port map( A1 => B(51), A2 => n206, ZN => n207);
   U69 : XNOR2_X1 port map( A => B(56), B => n203, ZN => DIFF_56_port);
   U70 : NOR2_X1 port map( A1 => B(55), A2 => n202, ZN => n203);
   U71 : OR3_X1 port map( A1 => B(45), A2 => B(46), A3 => n214, ZN => n212);
   U72 : OR3_X1 port map( A1 => B(51), A2 => B(52), A3 => n206, ZN => n204);
   U73 : OR3_X1 port map( A1 => B(55), A2 => B(56), A3 => n202, ZN => n200);
   U74 : XNOR2_X1 port map( A => n244, B => B(14), ZN => DIFF_14_port);
   U75 : NOR2_X1 port map( A1 => n247, A2 => B(13), ZN => n244);
   U76 : OR3_X1 port map( A1 => B(13), A2 => B(14), A3 => n247, ZN => n245);
   U77 : OR3_X1 port map( A1 => B(11), A2 => B(12), A3 => n249, ZN => n247);
   U78 : XNOR2_X1 port map( A => B(12), B => n250, ZN => DIFF_12_port);
   U79 : NOR2_X1 port map( A1 => B(11), A2 => n249, ZN => n250);
   U80 : NOR2_X1 port map( A1 => B(7), A2 => n192, ZN => n191);
   U84 : NOR2_X1 port map( A1 => B(3), A2 => n211, ZN => n210);
   U88 : OR3_X1 port map( A1 => B(10), A2 => B(9), A3 => n190, ZN => n249);
   U91 : OR3_X1 port map( A1 => B(5), A2 => B(6), A3 => n194, ZN => n192);
   U94 : OR3_X1 port map( A1 => B(7), A2 => B(8), A3 => n192, ZN => n190);
   U97 : OR3_X1 port map( A1 => B(3), A2 => B(4), A3 => n211, ZN => n194);
   U100 : XNOR2_X1 port map( A => B(8), B => n191, ZN => DIFF_8_port);
   U104 : XNOR2_X1 port map( A => B(4), B => n210, ZN => DIFF_4_port);
   U107 : XNOR2_X1 port map( A => B(2), B => n232, ZN => DIFF_2_port);
   U110 : OR2_X1 port map( A1 => n190, A2 => B(9), ZN => n251);
   U113 : OR2_X1 port map( A1 => n194, A2 => B(5), ZN => n193);
   U116 : OR3_X1 port map( A1 => B(1), A2 => B(2), A3 => B(0), ZN => n211);
   U120 : NOR2_X1 port map( A1 => B(0), A2 => B(1), ZN => n232);
   U123 : INV_X1 port map( A => B(61), ZN => n248);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_21_DW01_sub_0 is

   port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (63 downto 0);  CO : out std_logic);

end complementer_N64_21_DW01_sub_0;

architecture SYN_rpl of complementer_N64_21_DW01_sub_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal DIFF_62_port, DIFF_63_port, DIFF_11_port, DIFF_12_port, DIFF_13_port,
      DIFF_14_port, DIFF_15_port, DIFF_16_port, DIFF_17_port, DIFF_18_port, 
      DIFF_19_port, DIFF_20_port, DIFF_21_port, DIFF_22_port, DIFF_23_port, 
      DIFF_24_port, DIFF_25_port, DIFF_26_port, DIFF_27_port, DIFF_28_port, 
      DIFF_29_port, DIFF_30_port, DIFF_31_port, DIFF_32_port, DIFF_33_port, 
      DIFF_34_port, DIFF_35_port, DIFF_36_port, DIFF_37_port, DIFF_38_port, 
      DIFF_39_port, DIFF_40_port, DIFF_41_port, DIFF_42_port, DIFF_43_port, 
      DIFF_44_port, DIFF_45_port, DIFF_46_port, DIFF_47_port, DIFF_48_port, 
      DIFF_49_port, DIFF_50_port, DIFF_51_port, DIFF_52_port, DIFF_53_port, 
      DIFF_54_port, DIFF_55_port, DIFF_56_port, DIFF_57_port, DIFF_58_port, 
      DIFF_59_port, DIFF_60_port, DIFF_61_port, DIFF_3_port, DIFF_4_port, 
      DIFF_5_port, DIFF_6_port, DIFF_7_port, DIFF_8_port, DIFF_9_port, 
      DIFF_10_port, DIFF_2_port, DIFF_1_port, n190, n191, n192, n194, n195, 
      n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, 
      n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, 
      n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, 
      n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, 
      n244, n245, n246, n247, n248, n249, n250, n251, n189, n193 : std_logic;

begin
   DIFF <= ( DIFF_63_port, DIFF_62_port, DIFF_61_port, DIFF_60_port, 
      DIFF_59_port, DIFF_58_port, DIFF_57_port, DIFF_56_port, DIFF_55_port, 
      DIFF_54_port, DIFF_53_port, DIFF_52_port, DIFF_51_port, DIFF_50_port, 
      DIFF_49_port, DIFF_48_port, DIFF_47_port, DIFF_46_port, DIFF_45_port, 
      DIFF_44_port, DIFF_43_port, DIFF_42_port, DIFF_41_port, DIFF_40_port, 
      DIFF_39_port, DIFF_38_port, DIFF_37_port, DIFF_36_port, DIFF_35_port, 
      DIFF_34_port, DIFF_33_port, DIFF_32_port, DIFF_31_port, DIFF_30_port, 
      DIFF_29_port, DIFF_28_port, DIFF_27_port, DIFF_26_port, DIFF_25_port, 
      DIFF_24_port, DIFF_23_port, DIFF_22_port, DIFF_21_port, DIFF_20_port, 
      DIFF_19_port, DIFF_18_port, DIFF_17_port, DIFF_16_port, DIFF_15_port, 
      DIFF_14_port, DIFF_13_port, DIFF_12_port, DIFF_11_port, DIFF_10_port, 
      DIFF_9_port, DIFF_8_port, DIFF_7_port, DIFF_6_port, DIFF_5_port, 
      DIFF_4_port, DIFF_3_port, DIFF_2_port, DIFF_1_port, B(0) );
   
   U81 : XOR2_X1 port map( A => n190, B => B(9), Z => DIFF_9_port);
   U82 : XOR2_X1 port map( A => n192, B => B(7), Z => DIFF_7_port);
   U84 : XOR2_X1 port map( A => n195, B => B(63), Z => DIFF_63_port);
   U85 : XOR2_X1 port map( A => n196, B => B(62), Z => DIFF_62_port);
   U86 : XOR2_X1 port map( A => n194, B => B(5), Z => DIFF_5_port);
   U87 : XOR2_X1 port map( A => n198, B => B(59), Z => DIFF_59_port);
   U88 : XOR2_X1 port map( A => n201, B => B(58), Z => DIFF_58_port);
   U89 : XOR2_X1 port map( A => n200, B => B(57), Z => DIFF_57_port);
   U90 : XOR2_X1 port map( A => n202, B => B(55), Z => DIFF_55_port);
   U91 : XOR2_X1 port map( A => n205, B => B(54), Z => DIFF_54_port);
   U92 : XOR2_X1 port map( A => n204, B => B(53), Z => DIFF_53_port);
   U93 : XOR2_X1 port map( A => n206, B => B(51), Z => DIFF_51_port);
   U94 : XOR2_X1 port map( A => n209, B => B(50), Z => DIFF_50_port);
   U95 : XOR2_X1 port map( A => n208, B => B(49), Z => DIFF_49_port);
   U96 : XOR2_X1 port map( A => n212, B => B(47), Z => DIFF_47_port);
   U97 : XOR2_X1 port map( A => n215, B => B(46), Z => DIFF_46_port);
   U98 : XOR2_X1 port map( A => n214, B => B(45), Z => DIFF_45_port);
   U99 : XOR2_X1 port map( A => n216, B => B(43), Z => DIFF_43_port);
   U100 : XOR2_X1 port map( A => n219, B => B(42), Z => DIFF_42_port);
   U101 : XOR2_X1 port map( A => n218, B => B(41), Z => DIFF_41_port);
   U102 : XOR2_X1 port map( A => n211, B => B(3), Z => DIFF_3_port);
   U103 : XOR2_X1 port map( A => n220, B => B(39), Z => DIFF_39_port);
   U104 : XOR2_X1 port map( A => n223, B => B(38), Z => DIFF_38_port);
   U105 : XOR2_X1 port map( A => n222, B => B(37), Z => DIFF_37_port);
   U106 : XOR2_X1 port map( A => n224, B => B(35), Z => DIFF_35_port);
   U107 : XOR2_X1 port map( A => n227, B => B(34), Z => DIFF_34_port);
   U108 : XOR2_X1 port map( A => n226, B => B(33), Z => DIFF_33_port);
   U109 : XOR2_X1 port map( A => n228, B => B(31), Z => DIFF_31_port);
   U110 : XOR2_X1 port map( A => n231, B => B(30), Z => DIFF_30_port);
   U111 : XOR2_X1 port map( A => n230, B => B(29), Z => DIFF_29_port);
   U112 : XOR2_X1 port map( A => n233, B => B(27), Z => DIFF_27_port);
   U113 : XOR2_X1 port map( A => n236, B => B(26), Z => DIFF_26_port);
   U114 : XOR2_X1 port map( A => n235, B => B(25), Z => DIFF_25_port);
   U115 : XOR2_X1 port map( A => n237, B => B(23), Z => DIFF_23_port);
   U116 : XOR2_X1 port map( A => n240, B => B(22), Z => DIFF_22_port);
   U117 : XOR2_X1 port map( A => n239, B => B(21), Z => DIFF_21_port);
   U118 : XOR2_X1 port map( A => B(1), B => B(0), Z => DIFF_1_port);
   U119 : XOR2_X1 port map( A => n241, B => B(19), Z => DIFF_19_port);
   U120 : XOR2_X1 port map( A => n244, B => B(18), Z => DIFF_18_port);
   U121 : XOR2_X1 port map( A => n243, B => B(17), Z => DIFF_17_port);
   U122 : XOR2_X1 port map( A => n245, B => B(15), Z => DIFF_15_port);
   U123 : XOR2_X1 port map( A => n248, B => B(14), Z => DIFF_14_port);
   U124 : XOR2_X1 port map( A => n247, B => B(13), Z => DIFF_13_port);
   U125 : XOR2_X1 port map( A => n249, B => B(11), Z => DIFF_11_port);
   U126 : XOR2_X1 port map( A => n251, B => B(10), Z => DIFF_10_port);
   U1 : NOR2_X1 port map( A1 => B(43), A2 => n216, ZN => n217);
   U2 : NOR2_X1 port map( A1 => B(59), A2 => n198, ZN => n199);
   U3 : NAND2_X1 port map( A1 => n197, A2 => n193, ZN => n196);
   U4 : OR3_X1 port map( A1 => B(41), A2 => B(42), A3 => n218, ZN => n216);
   U5 : XNOR2_X1 port map( A => B(48), B => n213, ZN => DIFF_48_port);
   U6 : OR2_X1 port map( A1 => n218, A2 => B(41), ZN => n219);
   U7 : OR2_X1 port map( A1 => n208, A2 => B(49), ZN => n209);
   U8 : OR2_X1 port map( A1 => n204, A2 => B(53), ZN => n205);
   U9 : NOR2_X1 port map( A1 => B(35), A2 => n224, ZN => n225);
   U10 : NOR2_X1 port map( A1 => B(31), A2 => n228, ZN => n229);
   U11 : NOR2_X1 port map( A1 => B(27), A2 => n233, ZN => n234);
   U12 : NOR2_X1 port map( A1 => B(23), A2 => n237, ZN => n238);
   U13 : NOR2_X1 port map( A1 => B(19), A2 => n241, ZN => n242);
   U14 : NOR2_X1 port map( A1 => B(15), A2 => n245, ZN => n246);
   U15 : OR3_X1 port map( A1 => B(13), A2 => B(14), A3 => n247, ZN => n245);
   U16 : OR3_X1 port map( A1 => B(33), A2 => B(34), A3 => n226, ZN => n224);
   U17 : OR3_X1 port map( A1 => B(29), A2 => B(30), A3 => n230, ZN => n228);
   U18 : OR3_X1 port map( A1 => B(25), A2 => B(26), A3 => n235, ZN => n233);
   U19 : OR3_X1 port map( A1 => B(21), A2 => B(22), A3 => n239, ZN => n237);
   U20 : OR3_X1 port map( A1 => B(17), A2 => B(18), A3 => n243, ZN => n241);
   U21 : OR3_X1 port map( A1 => B(35), A2 => B(36), A3 => n224, ZN => n222);
   U22 : OR3_X1 port map( A1 => B(31), A2 => B(32), A3 => n228, ZN => n226);
   U23 : OR3_X1 port map( A1 => B(27), A2 => B(28), A3 => n233, ZN => n230);
   U24 : OR3_X1 port map( A1 => B(23), A2 => B(24), A3 => n237, ZN => n235);
   U25 : OR3_X1 port map( A1 => B(19), A2 => B(20), A3 => n241, ZN => n239);
   U26 : OR3_X1 port map( A1 => B(15), A2 => B(16), A3 => n245, ZN => n243);
   U27 : XNOR2_X1 port map( A => B(16), B => n246, ZN => DIFF_16_port);
   U28 : XNOR2_X1 port map( A => B(12), B => n250, ZN => DIFF_12_port);
   U29 : XNOR2_X1 port map( A => B(36), B => n225, ZN => DIFF_36_port);
   U30 : XNOR2_X1 port map( A => B(32), B => n229, ZN => DIFF_32_port);
   U31 : XNOR2_X1 port map( A => B(28), B => n234, ZN => DIFF_28_port);
   U32 : XNOR2_X1 port map( A => B(24), B => n238, ZN => DIFF_24_port);
   U33 : XNOR2_X1 port map( A => B(20), B => n242, ZN => DIFF_20_port);
   U34 : OR2_X1 port map( A1 => n247, A2 => B(13), ZN => n248);
   U35 : OR2_X1 port map( A1 => n226, A2 => B(33), ZN => n227);
   U36 : OR2_X1 port map( A1 => n230, A2 => B(29), ZN => n231);
   U37 : OR2_X1 port map( A1 => n235, A2 => B(25), ZN => n236);
   U38 : OR2_X1 port map( A1 => n239, A2 => B(21), ZN => n240);
   U39 : OR2_X1 port map( A1 => n243, A2 => B(17), ZN => n244);
   U40 : NOR3_X1 port map( A1 => B(59), A2 => B(60), A3 => n198, ZN => n197);
   U41 : XNOR2_X1 port map( A => n197, B => B(61), ZN => DIFF_61_port);
   U42 : XNOR2_X1 port map( A => B(60), B => n199, ZN => DIFF_60_port);
   U43 : NOR2_X1 port map( A1 => B(47), A2 => n212, ZN => n213);
   U44 : NOR2_X1 port map( A1 => B(39), A2 => n220, ZN => n221);
   U45 : NOR2_X1 port map( A1 => B(51), A2 => n206, ZN => n207);
   U46 : XNOR2_X1 port map( A => B(52), B => n207, ZN => DIFF_52_port);
   U47 : NOR2_X1 port map( A1 => B(55), A2 => n202, ZN => n203);
   U48 : OR3_X1 port map( A1 => B(57), A2 => B(58), A3 => n200, ZN => n198);
   U49 : OR3_X1 port map( A1 => B(45), A2 => B(46), A3 => n214, ZN => n212);
   U50 : OR3_X1 port map( A1 => B(49), A2 => B(50), A3 => n208, ZN => n206);
   U51 : OR3_X1 port map( A1 => B(37), A2 => B(38), A3 => n222, ZN => n220);
   U52 : OR3_X1 port map( A1 => B(53), A2 => B(54), A3 => n204, ZN => n202);
   U53 : OR3_X1 port map( A1 => B(47), A2 => B(48), A3 => n212, ZN => n208);
   U54 : OR3_X1 port map( A1 => B(43), A2 => B(44), A3 => n216, ZN => n214);
   U55 : OR3_X1 port map( A1 => B(39), A2 => B(40), A3 => n220, ZN => n218);
   U56 : OR3_X1 port map( A1 => B(51), A2 => B(52), A3 => n206, ZN => n204);
   U57 : OR3_X1 port map( A1 => B(55), A2 => B(56), A3 => n202, ZN => n200);
   U58 : XNOR2_X1 port map( A => B(56), B => n203, ZN => DIFF_56_port);
   U59 : XNOR2_X1 port map( A => B(40), B => n221, ZN => DIFF_40_port);
   U60 : XNOR2_X1 port map( A => B(44), B => n217, ZN => DIFF_44_port);
   U61 : OR2_X1 port map( A1 => n196, A2 => B(62), ZN => n195);
   U62 : OR2_X1 port map( A1 => n214, A2 => B(45), ZN => n215);
   U63 : OR2_X1 port map( A1 => n222, A2 => B(37), ZN => n223);
   U64 : OR2_X1 port map( A1 => n200, A2 => B(57), ZN => n201);
   U65 : NOR2_X1 port map( A1 => B(11), A2 => n249, ZN => n250);
   U66 : OR3_X1 port map( A1 => B(11), A2 => B(12), A3 => n249, ZN => n247);
   U67 : XNOR2_X1 port map( A => n189, B => B(6), ZN => DIFF_6_port);
   U68 : NOR2_X1 port map( A1 => n194, A2 => B(5), ZN => n189);
   U69 : XNOR2_X1 port map( A => B(8), B => n191, ZN => DIFF_8_port);
   U70 : NOR2_X1 port map( A1 => B(7), A2 => n192, ZN => n191);
   U71 : XNOR2_X1 port map( A => B(2), B => n232, ZN => DIFF_2_port);
   U72 : NOR2_X1 port map( A1 => B(0), A2 => B(1), ZN => n232);
   U73 : XNOR2_X1 port map( A => B(4), B => n210, ZN => DIFF_4_port);
   U74 : NOR2_X1 port map( A1 => B(3), A2 => n211, ZN => n210);
   U75 : OR3_X1 port map( A1 => B(5), A2 => B(6), A3 => n194, ZN => n192);
   U76 : OR3_X1 port map( A1 => B(10), A2 => B(9), A3 => n190, ZN => n249);
   U77 : OR3_X1 port map( A1 => B(7), A2 => B(8), A3 => n192, ZN => n190);
   U78 : OR3_X1 port map( A1 => B(3), A2 => B(4), A3 => n211, ZN => n194);
   U79 : OR2_X1 port map( A1 => n190, A2 => B(9), ZN => n251);
   U80 : OR3_X1 port map( A1 => B(1), A2 => B(2), A3 => B(0), ZN => n211);
   U83 : INV_X1 port map( A => B(61), ZN => n193);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_22_DW01_sub_0 is

   port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (63 downto 0);  CO : out std_logic);

end complementer_N64_22_DW01_sub_0;

architecture SYN_rpl of complementer_N64_22_DW01_sub_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal DIFF_62_port, DIFF_61_port, DIFF_60_port, DIFF_59_port, DIFF_58_port,
      DIFF_57_port, DIFF_56_port, DIFF_55_port, DIFF_54_port, DIFF_53_port, 
      DIFF_52_port, DIFF_51_port, DIFF_50_port, DIFF_49_port, DIFF_48_port, 
      DIFF_47_port, DIFF_46_port, DIFF_45_port, DIFF_44_port, DIFF_43_port, 
      DIFF_42_port, DIFF_41_port, DIFF_40_port, DIFF_39_port, DIFF_38_port, 
      DIFF_37_port, DIFF_36_port, DIFF_35_port, DIFF_34_port, DIFF_33_port, 
      DIFF_32_port, DIFF_31_port, DIFF_30_port, DIFF_29_port, DIFF_28_port, 
      DIFF_27_port, DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, 
      DIFF_22_port, DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, 
      DIFF_17_port, DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, 
      DIFF_12_port, DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, 
      DIFF_7_port, DIFF_6_port, DIFF_5_port, DIFF_4_port, DIFF_3_port, 
      DIFF_2_port, DIFF_1_port, DIFF_63_port, n190, n191, n192, n193, n194, 
      n196, n197, n198, n199, n200, n202, n203, n204, n206, n207, n208, n210, 
      n211, n212, n213, n214, n216, n217, n218, n220, n221, n222, n224, n225, 
      n226, n228, n229, n230, n232, n233, n234, n235, n237, n238, n239, n241, 
      n242, n243, n245, n246, n247, n249, n250, n189, n195, n201, n205, n209, 
      n215, n219, n223, n227, n231, n236, n240, n244, n248, n251 : std_logic;

begin
   DIFF <= ( DIFF_63_port, DIFF_62_port, DIFF_61_port, DIFF_60_port, 
      DIFF_59_port, DIFF_58_port, DIFF_57_port, DIFF_56_port, DIFF_55_port, 
      DIFF_54_port, DIFF_53_port, DIFF_52_port, DIFF_51_port, DIFF_50_port, 
      DIFF_49_port, DIFF_48_port, DIFF_47_port, DIFF_46_port, DIFF_45_port, 
      DIFF_44_port, DIFF_43_port, DIFF_42_port, DIFF_41_port, DIFF_40_port, 
      DIFF_39_port, DIFF_38_port, DIFF_37_port, DIFF_36_port, DIFF_35_port, 
      DIFF_34_port, DIFF_33_port, DIFF_32_port, DIFF_31_port, DIFF_30_port, 
      DIFF_29_port, DIFF_28_port, DIFF_27_port, DIFF_26_port, DIFF_25_port, 
      DIFF_24_port, DIFF_23_port, DIFF_22_port, DIFF_21_port, DIFF_20_port, 
      DIFF_19_port, DIFF_18_port, DIFF_17_port, DIFF_16_port, DIFF_15_port, 
      DIFF_14_port, DIFF_13_port, DIFF_12_port, DIFF_11_port, DIFF_10_port, 
      DIFF_9_port, DIFF_8_port, DIFF_7_port, DIFF_6_port, DIFF_5_port, 
      DIFF_4_port, DIFF_3_port, DIFF_2_port, DIFF_1_port, B(0) );
   
   U81 : XOR2_X1 port map( A => n190, B => B(9), Z => DIFF_9_port);
   U82 : XOR2_X1 port map( A => n192, B => B(7), Z => DIFF_7_port);
   U83 : XOR2_X1 port map( A => n193, B => B(6), Z => DIFF_6_port);
   U85 : XOR2_X1 port map( A => n196, B => B(62), Z => DIFF_62_port);
   U86 : XOR2_X1 port map( A => n194, B => B(5), Z => DIFF_5_port);
   U87 : XOR2_X1 port map( A => n198, B => B(59), Z => DIFF_59_port);
   U89 : XOR2_X1 port map( A => n200, B => B(57), Z => DIFF_57_port);
   U90 : XOR2_X1 port map( A => n202, B => B(55), Z => DIFF_55_port);
   U92 : XOR2_X1 port map( A => n204, B => B(53), Z => DIFF_53_port);
   U93 : XOR2_X1 port map( A => n206, B => B(51), Z => DIFF_51_port);
   U95 : XOR2_X1 port map( A => n208, B => B(49), Z => DIFF_49_port);
   U96 : XOR2_X1 port map( A => n212, B => B(47), Z => DIFF_47_port);
   U98 : XOR2_X1 port map( A => n214, B => B(45), Z => DIFF_45_port);
   U99 : XOR2_X1 port map( A => n216, B => B(43), Z => DIFF_43_port);
   U101 : XOR2_X1 port map( A => n218, B => B(41), Z => DIFF_41_port);
   U102 : XOR2_X1 port map( A => n211, B => B(3), Z => DIFF_3_port);
   U103 : XOR2_X1 port map( A => n220, B => B(39), Z => DIFF_39_port);
   U105 : XOR2_X1 port map( A => n222, B => B(37), Z => DIFF_37_port);
   U106 : XOR2_X1 port map( A => n224, B => B(35), Z => DIFF_35_port);
   U108 : XOR2_X1 port map( A => n226, B => B(33), Z => DIFF_33_port);
   U109 : XOR2_X1 port map( A => n228, B => B(31), Z => DIFF_31_port);
   U111 : XOR2_X1 port map( A => n230, B => B(29), Z => DIFF_29_port);
   U112 : XOR2_X1 port map( A => n233, B => B(27), Z => DIFF_27_port);
   U114 : XOR2_X1 port map( A => n235, B => B(25), Z => DIFF_25_port);
   U115 : XOR2_X1 port map( A => n237, B => B(23), Z => DIFF_23_port);
   U117 : XOR2_X1 port map( A => n239, B => B(21), Z => DIFF_21_port);
   U118 : XOR2_X1 port map( A => B(1), B => B(0), Z => DIFF_1_port);
   U119 : XOR2_X1 port map( A => n241, B => B(19), Z => DIFF_19_port);
   U121 : XOR2_X1 port map( A => n243, B => B(17), Z => DIFF_17_port);
   U122 : XOR2_X1 port map( A => n245, B => B(15), Z => DIFF_15_port);
   U124 : XOR2_X1 port map( A => n247, B => B(13), Z => DIFF_13_port);
   U125 : XOR2_X1 port map( A => n249, B => B(11), Z => DIFF_11_port);
   U1 : XNOR2_X1 port map( A => B(48), B => n213, ZN => DIFF_48_port);
   U2 : NOR2_X1 port map( A1 => B(47), A2 => n212, ZN => n213);
   U3 : XOR2_X1 port map( A => n197, B => n251, Z => DIFF_61_port);
   U4 : NAND2_X1 port map( A1 => n197, A2 => n251, ZN => n196);
   U5 : OR3_X1 port map( A1 => B(57), A2 => B(58), A3 => n200, ZN => n198);
   U6 : OR3_X1 port map( A1 => B(47), A2 => B(48), A3 => n212, ZN => n208);
   U7 : XNOR2_X1 port map( A => n189, B => B(58), ZN => DIFF_58_port);
   U8 : NOR2_X1 port map( A1 => n200, A2 => B(57), ZN => n189);
   U9 : XNOR2_X1 port map( A => n195, B => B(18), ZN => DIFF_18_port);
   U10 : NOR2_X1 port map( A1 => n243, A2 => B(17), ZN => n195);
   U11 : XNOR2_X1 port map( A => n201, B => B(14), ZN => DIFF_14_port);
   U12 : NOR2_X1 port map( A1 => n247, A2 => B(13), ZN => n201);
   U13 : XNOR2_X1 port map( A => n205, B => B(30), ZN => DIFF_30_port);
   U14 : NOR2_X1 port map( A1 => n230, A2 => B(29), ZN => n205);
   U15 : XNOR2_X1 port map( A => n209, B => B(26), ZN => DIFF_26_port);
   U16 : NOR2_X1 port map( A1 => n235, A2 => B(25), ZN => n209);
   U17 : XNOR2_X1 port map( A => n215, B => B(22), ZN => DIFF_22_port);
   U18 : NOR2_X1 port map( A1 => n239, A2 => B(21), ZN => n215);
   U19 : XNOR2_X1 port map( A => B(36), B => n225, ZN => DIFF_36_port);
   U20 : NOR2_X1 port map( A1 => B(35), A2 => n224, ZN => n225);
   U21 : XNOR2_X1 port map( A => B(32), B => n229, ZN => DIFF_32_port);
   U22 : NOR2_X1 port map( A1 => B(31), A2 => n228, ZN => n229);
   U23 : XNOR2_X1 port map( A => B(16), B => n246, ZN => DIFF_16_port);
   U24 : NOR2_X1 port map( A1 => B(15), A2 => n245, ZN => n246);
   U25 : XNOR2_X1 port map( A => B(28), B => n234, ZN => DIFF_28_port);
   U26 : NOR2_X1 port map( A1 => B(27), A2 => n233, ZN => n234);
   U27 : XNOR2_X1 port map( A => B(24), B => n238, ZN => DIFF_24_port);
   U28 : NOR2_X1 port map( A1 => B(23), A2 => n237, ZN => n238);
   U29 : XNOR2_X1 port map( A => B(20), B => n242, ZN => DIFF_20_port);
   U30 : NOR2_X1 port map( A1 => B(19), A2 => n241, ZN => n242);
   U31 : OR3_X1 port map( A1 => B(13), A2 => B(14), A3 => n247, ZN => n245);
   U32 : OR3_X1 port map( A1 => B(17), A2 => B(18), A3 => n243, ZN => n241);
   U33 : OR3_X1 port map( A1 => B(21), A2 => B(22), A3 => n239, ZN => n237);
   U34 : OR3_X1 port map( A1 => B(25), A2 => B(26), A3 => n235, ZN => n233);
   U35 : OR3_X1 port map( A1 => B(29), A2 => B(30), A3 => n230, ZN => n228);
   U36 : OR3_X1 port map( A1 => B(33), A2 => B(34), A3 => n226, ZN => n224);
   U37 : OR3_X1 port map( A1 => B(37), A2 => B(38), A3 => n222, ZN => n220);
   U38 : OR3_X1 port map( A1 => B(15), A2 => B(16), A3 => n245, ZN => n243);
   U39 : OR3_X1 port map( A1 => B(19), A2 => B(20), A3 => n241, ZN => n239);
   U40 : OR3_X1 port map( A1 => B(23), A2 => B(24), A3 => n237, ZN => n235);
   U41 : OR3_X1 port map( A1 => B(27), A2 => B(28), A3 => n233, ZN => n230);
   U42 : OR3_X1 port map( A1 => B(31), A2 => B(32), A3 => n228, ZN => n226);
   U43 : OR3_X1 port map( A1 => B(35), A2 => B(36), A3 => n224, ZN => n222);
   U44 : XNOR2_X1 port map( A => n219, B => B(38), ZN => DIFF_38_port);
   U45 : NOR2_X1 port map( A1 => n222, A2 => B(37), ZN => n219);
   U46 : XNOR2_X1 port map( A => n223, B => B(34), ZN => DIFF_34_port);
   U47 : NOR2_X1 port map( A1 => n226, A2 => B(33), ZN => n223);
   U48 : NOR3_X1 port map( A1 => B(59), A2 => B(60), A3 => n198, ZN => n197);
   U49 : XNOR2_X1 port map( A => n227, B => B(46), ZN => DIFF_46_port);
   U50 : NOR2_X1 port map( A1 => n214, A2 => B(45), ZN => n227);
   U51 : XNOR2_X1 port map( A => n231, B => B(50), ZN => DIFF_50_port);
   U52 : NOR2_X1 port map( A1 => n208, A2 => B(49), ZN => n231);
   U53 : XNOR2_X1 port map( A => n236, B => B(42), ZN => DIFF_42_port);
   U54 : NOR2_X1 port map( A1 => n218, A2 => B(41), ZN => n236);
   U55 : XNOR2_X1 port map( A => n240, B => B(54), ZN => DIFF_54_port);
   U56 : NOR2_X1 port map( A1 => n204, A2 => B(53), ZN => n240);
   U57 : XNOR2_X1 port map( A => B(52), B => n207, ZN => DIFF_52_port);
   U58 : NOR2_X1 port map( A1 => B(51), A2 => n206, ZN => n207);
   U59 : XNOR2_X1 port map( A => B(40), B => n221, ZN => DIFF_40_port);
   U60 : NOR2_X1 port map( A1 => B(39), A2 => n220, ZN => n221);
   U61 : XNOR2_X1 port map( A => B(44), B => n217, ZN => DIFF_44_port);
   U62 : NOR2_X1 port map( A1 => B(43), A2 => n216, ZN => n217);
   U63 : XNOR2_X1 port map( A => B(60), B => n199, ZN => DIFF_60_port);
   U64 : NOR2_X1 port map( A1 => B(59), A2 => n198, ZN => n199);
   U65 : XNOR2_X1 port map( A => B(56), B => n203, ZN => DIFF_56_port);
   U66 : NOR2_X1 port map( A1 => B(55), A2 => n202, ZN => n203);
   U67 : OR3_X1 port map( A1 => B(49), A2 => B(50), A3 => n208, ZN => n206);
   U68 : OR3_X1 port map( A1 => B(45), A2 => B(46), A3 => n214, ZN => n212);
   U69 : OR3_X1 port map( A1 => B(41), A2 => B(42), A3 => n218, ZN => n216);
   U70 : OR3_X1 port map( A1 => B(53), A2 => B(54), A3 => n204, ZN => n202);
   U71 : OR3_X1 port map( A1 => B(51), A2 => B(52), A3 => n206, ZN => n204);
   U72 : OR3_X1 port map( A1 => B(43), A2 => B(44), A3 => n216, ZN => n214);
   U73 : OR3_X1 port map( A1 => B(39), A2 => B(40), A3 => n220, ZN => n218);
   U74 : OR3_X1 port map( A1 => B(55), A2 => B(56), A3 => n202, ZN => n200);
   U75 : XNOR2_X1 port map( A => B(12), B => n250, ZN => DIFF_12_port);
   U76 : NOR2_X1 port map( A1 => B(11), A2 => n249, ZN => n250);
   U77 : OR3_X1 port map( A1 => B(11), A2 => B(12), A3 => n249, ZN => n247);
   U78 : XNOR2_X1 port map( A => n244, B => B(63), ZN => DIFF_63_port);
   U79 : NOR2_X1 port map( A1 => n196, A2 => B(62), ZN => n244);
   U80 : XNOR2_X1 port map( A => n248, B => B(10), ZN => DIFF_10_port);
   U84 : NOR2_X1 port map( A1 => n190, A2 => B(9), ZN => n248);
   U88 : OR3_X1 port map( A1 => B(10), A2 => B(9), A3 => n190, ZN => n249);
   U91 : NOR2_X1 port map( A1 => B(7), A2 => n192, ZN => n191);
   U94 : NOR2_X1 port map( A1 => B(3), A2 => n211, ZN => n210);
   U97 : OR3_X1 port map( A1 => B(5), A2 => B(6), A3 => n194, ZN => n192);
   U100 : OR3_X1 port map( A1 => B(7), A2 => B(8), A3 => n192, ZN => n190);
   U104 : OR3_X1 port map( A1 => B(3), A2 => B(4), A3 => n211, ZN => n194);
   U107 : XNOR2_X1 port map( A => B(8), B => n191, ZN => DIFF_8_port);
   U110 : XNOR2_X1 port map( A => B(4), B => n210, ZN => DIFF_4_port);
   U113 : XNOR2_X1 port map( A => B(2), B => n232, ZN => DIFF_2_port);
   U116 : OR2_X1 port map( A1 => n194, A2 => B(5), ZN => n193);
   U120 : OR3_X1 port map( A1 => B(1), A2 => B(2), A3 => B(0), ZN => n211);
   U123 : NOR2_X1 port map( A1 => B(0), A2 => B(1), ZN => n232);
   U126 : INV_X1 port map( A => B(61), ZN => n251);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_23_DW01_sub_0 is

   port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (63 downto 0);  CO : out std_logic);

end complementer_N64_23_DW01_sub_0;

architecture SYN_rpl of complementer_N64_23_DW01_sub_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal DIFF_62_port, DIFF_63_port, DIFF_9_port, DIFF_10_port, DIFF_11_port, 
      DIFF_12_port, DIFF_13_port, DIFF_14_port, DIFF_15_port, DIFF_16_port, 
      DIFF_17_port, DIFF_18_port, DIFF_19_port, DIFF_20_port, DIFF_21_port, 
      DIFF_22_port, DIFF_23_port, DIFF_24_port, DIFF_25_port, DIFF_26_port, 
      DIFF_27_port, DIFF_28_port, DIFF_29_port, DIFF_30_port, DIFF_31_port, 
      DIFF_32_port, DIFF_33_port, DIFF_34_port, DIFF_35_port, DIFF_36_port, 
      DIFF_37_port, DIFF_38_port, DIFF_39_port, DIFF_40_port, DIFF_41_port, 
      DIFF_42_port, DIFF_43_port, DIFF_44_port, DIFF_45_port, DIFF_46_port, 
      DIFF_47_port, DIFF_48_port, DIFF_49_port, DIFF_50_port, DIFF_51_port, 
      DIFF_52_port, DIFF_53_port, DIFF_54_port, DIFF_55_port, DIFF_56_port, 
      DIFF_57_port, DIFF_58_port, DIFF_59_port, DIFF_60_port, DIFF_61_port, 
      DIFF_3_port, DIFF_4_port, DIFF_5_port, DIFF_6_port, DIFF_7_port, 
      DIFF_8_port, DIFF_2_port, DIFF_1_port, n190, n191, n192, n194, n195, n196
      , n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
      n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, 
      n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, 
      n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, 
      n245, n246, n247, n248, n249, n250, n251, n189, n193 : std_logic;

begin
   DIFF <= ( DIFF_63_port, DIFF_62_port, DIFF_61_port, DIFF_60_port, 
      DIFF_59_port, DIFF_58_port, DIFF_57_port, DIFF_56_port, DIFF_55_port, 
      DIFF_54_port, DIFF_53_port, DIFF_52_port, DIFF_51_port, DIFF_50_port, 
      DIFF_49_port, DIFF_48_port, DIFF_47_port, DIFF_46_port, DIFF_45_port, 
      DIFF_44_port, DIFF_43_port, DIFF_42_port, DIFF_41_port, DIFF_40_port, 
      DIFF_39_port, DIFF_38_port, DIFF_37_port, DIFF_36_port, DIFF_35_port, 
      DIFF_34_port, DIFF_33_port, DIFF_32_port, DIFF_31_port, DIFF_30_port, 
      DIFF_29_port, DIFF_28_port, DIFF_27_port, DIFF_26_port, DIFF_25_port, 
      DIFF_24_port, DIFF_23_port, DIFF_22_port, DIFF_21_port, DIFF_20_port, 
      DIFF_19_port, DIFF_18_port, DIFF_17_port, DIFF_16_port, DIFF_15_port, 
      DIFF_14_port, DIFF_13_port, DIFF_12_port, DIFF_11_port, DIFF_10_port, 
      DIFF_9_port, DIFF_8_port, DIFF_7_port, DIFF_6_port, DIFF_5_port, 
      DIFF_4_port, DIFF_3_port, DIFF_2_port, DIFF_1_port, B(0) );
   
   U81 : XOR2_X1 port map( A => n190, B => B(9), Z => DIFF_9_port);
   U82 : XOR2_X1 port map( A => n192, B => B(7), Z => DIFF_7_port);
   U84 : XOR2_X1 port map( A => n195, B => B(63), Z => DIFF_63_port);
   U85 : XOR2_X1 port map( A => n196, B => B(62), Z => DIFF_62_port);
   U86 : XOR2_X1 port map( A => n194, B => B(5), Z => DIFF_5_port);
   U87 : XOR2_X1 port map( A => n198, B => B(59), Z => DIFF_59_port);
   U88 : XOR2_X1 port map( A => n201, B => B(58), Z => DIFF_58_port);
   U89 : XOR2_X1 port map( A => n200, B => B(57), Z => DIFF_57_port);
   U90 : XOR2_X1 port map( A => n202, B => B(55), Z => DIFF_55_port);
   U91 : XOR2_X1 port map( A => n205, B => B(54), Z => DIFF_54_port);
   U92 : XOR2_X1 port map( A => n204, B => B(53), Z => DIFF_53_port);
   U93 : XOR2_X1 port map( A => n206, B => B(51), Z => DIFF_51_port);
   U94 : XOR2_X1 port map( A => n209, B => B(50), Z => DIFF_50_port);
   U95 : XOR2_X1 port map( A => n208, B => B(49), Z => DIFF_49_port);
   U96 : XOR2_X1 port map( A => n212, B => B(47), Z => DIFF_47_port);
   U97 : XOR2_X1 port map( A => n215, B => B(46), Z => DIFF_46_port);
   U98 : XOR2_X1 port map( A => n214, B => B(45), Z => DIFF_45_port);
   U99 : XOR2_X1 port map( A => n216, B => B(43), Z => DIFF_43_port);
   U100 : XOR2_X1 port map( A => n219, B => B(42), Z => DIFF_42_port);
   U101 : XOR2_X1 port map( A => n218, B => B(41), Z => DIFF_41_port);
   U102 : XOR2_X1 port map( A => n211, B => B(3), Z => DIFF_3_port);
   U103 : XOR2_X1 port map( A => n220, B => B(39), Z => DIFF_39_port);
   U104 : XOR2_X1 port map( A => n223, B => B(38), Z => DIFF_38_port);
   U105 : XOR2_X1 port map( A => n222, B => B(37), Z => DIFF_37_port);
   U106 : XOR2_X1 port map( A => n224, B => B(35), Z => DIFF_35_port);
   U107 : XOR2_X1 port map( A => n227, B => B(34), Z => DIFF_34_port);
   U108 : XOR2_X1 port map( A => n226, B => B(33), Z => DIFF_33_port);
   U109 : XOR2_X1 port map( A => n228, B => B(31), Z => DIFF_31_port);
   U110 : XOR2_X1 port map( A => n231, B => B(30), Z => DIFF_30_port);
   U111 : XOR2_X1 port map( A => n230, B => B(29), Z => DIFF_29_port);
   U112 : XOR2_X1 port map( A => n233, B => B(27), Z => DIFF_27_port);
   U113 : XOR2_X1 port map( A => n236, B => B(26), Z => DIFF_26_port);
   U114 : XOR2_X1 port map( A => n235, B => B(25), Z => DIFF_25_port);
   U115 : XOR2_X1 port map( A => n237, B => B(23), Z => DIFF_23_port);
   U116 : XOR2_X1 port map( A => n240, B => B(22), Z => DIFF_22_port);
   U117 : XOR2_X1 port map( A => n239, B => B(21), Z => DIFF_21_port);
   U118 : XOR2_X1 port map( A => B(1), B => B(0), Z => DIFF_1_port);
   U119 : XOR2_X1 port map( A => n241, B => B(19), Z => DIFF_19_port);
   U120 : XOR2_X1 port map( A => n244, B => B(18), Z => DIFF_18_port);
   U121 : XOR2_X1 port map( A => n243, B => B(17), Z => DIFF_17_port);
   U122 : XOR2_X1 port map( A => n245, B => B(15), Z => DIFF_15_port);
   U123 : XOR2_X1 port map( A => n248, B => B(14), Z => DIFF_14_port);
   U124 : XOR2_X1 port map( A => n247, B => B(13), Z => DIFF_13_port);
   U125 : XOR2_X1 port map( A => n249, B => B(11), Z => DIFF_11_port);
   U126 : XOR2_X1 port map( A => n251, B => B(10), Z => DIFF_10_port);
   U1 : NAND2_X1 port map( A1 => n197, A2 => n193, ZN => n196);
   U2 : NOR2_X1 port map( A1 => B(43), A2 => n216, ZN => n217);
   U3 : NOR2_X1 port map( A1 => B(19), A2 => n241, ZN => n242);
   U4 : NOR2_X1 port map( A1 => B(11), A2 => n249, ZN => n250);
   U5 : NOR2_X1 port map( A1 => B(15), A2 => n245, ZN => n246);
   U6 : NOR2_X1 port map( A1 => B(35), A2 => n224, ZN => n225);
   U7 : NOR2_X1 port map( A1 => B(31), A2 => n228, ZN => n229);
   U8 : NOR2_X1 port map( A1 => B(27), A2 => n233, ZN => n234);
   U9 : NOR2_X1 port map( A1 => B(23), A2 => n237, ZN => n238);
   U10 : NOR2_X1 port map( A1 => B(39), A2 => n220, ZN => n221);
   U11 : XNOR2_X1 port map( A => B(36), B => n225, ZN => DIFF_36_port);
   U12 : XNOR2_X1 port map( A => B(32), B => n229, ZN => DIFF_32_port);
   U13 : OR3_X1 port map( A1 => B(17), A2 => B(18), A3 => n243, ZN => n241);
   U14 : OR3_X1 port map( A1 => B(21), A2 => B(22), A3 => n239, ZN => n237);
   U15 : OR3_X1 port map( A1 => B(13), A2 => B(14), A3 => n247, ZN => n245);
   U16 : OR3_X1 port map( A1 => B(37), A2 => B(38), A3 => n222, ZN => n220);
   U17 : OR3_X1 port map( A1 => B(33), A2 => B(34), A3 => n226, ZN => n224);
   U18 : OR3_X1 port map( A1 => B(29), A2 => B(30), A3 => n230, ZN => n228);
   U19 : OR3_X1 port map( A1 => B(25), A2 => B(26), A3 => n235, ZN => n233);
   U20 : OR3_X1 port map( A1 => B(41), A2 => B(42), A3 => n218, ZN => n216);
   U21 : OR3_X1 port map( A1 => B(19), A2 => B(20), A3 => n241, ZN => n239);
   U22 : OR3_X1 port map( A1 => B(11), A2 => B(12), A3 => n249, ZN => n247);
   U23 : OR3_X1 port map( A1 => B(15), A2 => B(16), A3 => n245, ZN => n243);
   U24 : OR3_X1 port map( A1 => B(35), A2 => B(36), A3 => n224, ZN => n222);
   U25 : OR3_X1 port map( A1 => B(31), A2 => B(32), A3 => n228, ZN => n226);
   U26 : OR3_X1 port map( A1 => B(27), A2 => B(28), A3 => n233, ZN => n230);
   U27 : OR3_X1 port map( A1 => B(23), A2 => B(24), A3 => n237, ZN => n235);
   U28 : OR3_X1 port map( A1 => B(39), A2 => B(40), A3 => n220, ZN => n218);
   U29 : XNOR2_X1 port map( A => B(40), B => n221, ZN => DIFF_40_port);
   U30 : XNOR2_X1 port map( A => B(12), B => n250, ZN => DIFF_12_port);
   U31 : XNOR2_X1 port map( A => B(24), B => n238, ZN => DIFF_24_port);
   U32 : XNOR2_X1 port map( A => B(16), B => n246, ZN => DIFF_16_port);
   U33 : XNOR2_X1 port map( A => B(20), B => n242, ZN => DIFF_20_port);
   U34 : XNOR2_X1 port map( A => B(44), B => n217, ZN => DIFF_44_port);
   U35 : XNOR2_X1 port map( A => B(28), B => n234, ZN => DIFF_28_port);
   U36 : OR2_X1 port map( A1 => n239, A2 => B(21), ZN => n240);
   U37 : OR2_X1 port map( A1 => n243, A2 => B(17), ZN => n244);
   U38 : OR2_X1 port map( A1 => n247, A2 => B(13), ZN => n248);
   U39 : OR2_X1 port map( A1 => n222, A2 => B(37), ZN => n223);
   U40 : OR2_X1 port map( A1 => n226, A2 => B(33), ZN => n227);
   U41 : OR2_X1 port map( A1 => n230, A2 => B(29), ZN => n231);
   U42 : OR2_X1 port map( A1 => n235, A2 => B(25), ZN => n236);
   U43 : OR2_X1 port map( A1 => n218, A2 => B(41), ZN => n219);
   U44 : NOR3_X1 port map( A1 => B(59), A2 => B(60), A3 => n198, ZN => n197);
   U45 : XNOR2_X1 port map( A => B(60), B => n199, ZN => DIFF_60_port);
   U46 : NOR2_X1 port map( A1 => B(47), A2 => n212, ZN => n213);
   U47 : NOR2_X1 port map( A1 => B(51), A2 => n206, ZN => n207);
   U48 : NOR2_X1 port map( A1 => B(59), A2 => n198, ZN => n199);
   U49 : NOR2_X1 port map( A1 => B(55), A2 => n202, ZN => n203);
   U50 : OR3_X1 port map( A1 => B(57), A2 => B(58), A3 => n200, ZN => n198);
   U51 : OR3_X1 port map( A1 => B(45), A2 => B(46), A3 => n214, ZN => n212);
   U52 : OR3_X1 port map( A1 => B(49), A2 => B(50), A3 => n208, ZN => n206);
   U53 : OR3_X1 port map( A1 => B(53), A2 => B(54), A3 => n204, ZN => n202);
   U54 : OR3_X1 port map( A1 => B(47), A2 => B(48), A3 => n212, ZN => n208);
   U55 : OR3_X1 port map( A1 => B(43), A2 => B(44), A3 => n216, ZN => n214);
   U56 : OR3_X1 port map( A1 => B(51), A2 => B(52), A3 => n206, ZN => n204);
   U57 : OR3_X1 port map( A1 => B(55), A2 => B(56), A3 => n202, ZN => n200);
   U58 : XNOR2_X1 port map( A => B(48), B => n213, ZN => DIFF_48_port);
   U59 : XNOR2_X1 port map( A => B(56), B => n203, ZN => DIFF_56_port);
   U60 : OR2_X1 port map( A1 => n214, A2 => B(45), ZN => n215);
   U61 : OR2_X1 port map( A1 => n208, A2 => B(49), ZN => n209);
   U62 : OR2_X1 port map( A1 => n200, A2 => B(57), ZN => n201);
   U63 : OR2_X1 port map( A1 => n204, A2 => B(53), ZN => n205);
   U64 : OR3_X1 port map( A1 => B(10), A2 => B(9), A3 => n190, ZN => n249);
   U65 : OR2_X1 port map( A1 => n190, A2 => B(9), ZN => n251);
   U66 : XNOR2_X1 port map( A => n197, B => B(61), ZN => DIFF_61_port);
   U67 : XNOR2_X1 port map( A => B(52), B => n207, ZN => DIFF_52_port);
   U68 : OR2_X1 port map( A1 => n196, A2 => B(62), ZN => n195);
   U69 : XNOR2_X1 port map( A => B(8), B => n191, ZN => DIFF_8_port);
   U70 : XNOR2_X1 port map( A => n189, B => B(6), ZN => DIFF_6_port);
   U71 : NOR2_X1 port map( A1 => n194, A2 => B(5), ZN => n189);
   U72 : NOR2_X1 port map( A1 => B(7), A2 => n192, ZN => n191);
   U73 : XNOR2_X1 port map( A => B(2), B => n232, ZN => DIFF_2_port);
   U74 : NOR2_X1 port map( A1 => B(0), A2 => B(1), ZN => n232);
   U75 : XNOR2_X1 port map( A => B(4), B => n210, ZN => DIFF_4_port);
   U76 : NOR2_X1 port map( A1 => B(3), A2 => n211, ZN => n210);
   U77 : OR3_X1 port map( A1 => B(5), A2 => B(6), A3 => n194, ZN => n192);
   U78 : OR3_X1 port map( A1 => B(7), A2 => B(8), A3 => n192, ZN => n190);
   U79 : OR3_X1 port map( A1 => B(3), A2 => B(4), A3 => n211, ZN => n194);
   U80 : OR3_X1 port map( A1 => B(1), A2 => B(2), A3 => B(0), ZN => n211);
   U83 : INV_X1 port map( A => B(61), ZN => n193);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_24_DW01_sub_0 is

   port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (63 downto 0);  CO : out std_logic);

end complementer_N64_24_DW01_sub_0;

architecture SYN_rpl of complementer_N64_24_DW01_sub_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal DIFF_62_port, DIFF_61_port, DIFF_60_port, DIFF_59_port, DIFF_58_port,
      DIFF_57_port, DIFF_56_port, DIFF_55_port, DIFF_54_port, DIFF_53_port, 
      DIFF_52_port, DIFF_51_port, DIFF_50_port, DIFF_49_port, DIFF_48_port, 
      DIFF_47_port, DIFF_46_port, DIFF_45_port, DIFF_44_port, DIFF_43_port, 
      DIFF_42_port, DIFF_41_port, DIFF_40_port, DIFF_39_port, DIFF_38_port, 
      DIFF_37_port, DIFF_36_port, DIFF_35_port, DIFF_34_port, DIFF_33_port, 
      DIFF_32_port, DIFF_31_port, DIFF_30_port, DIFF_29_port, DIFF_28_port, 
      DIFF_27_port, DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, 
      DIFF_22_port, DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, 
      DIFF_17_port, DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, 
      DIFF_12_port, DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, 
      DIFF_7_port, DIFF_6_port, DIFF_5_port, DIFF_4_port, DIFF_3_port, 
      DIFF_2_port, DIFF_1_port, DIFF_63_port, n190, n191, n192, n193, n194, 
      n196, n197, n198, n199, n200, n202, n203, n204, n206, n207, n208, n210, 
      n211, n212, n213, n214, n216, n217, n218, n220, n221, n222, n224, n225, 
      n226, n228, n229, n230, n232, n233, n234, n235, n237, n238, n239, n241, 
      n242, n243, n245, n246, n247, n249, n250, n189, n195, n201, n205, n209, 
      n215, n219, n223, n227, n231, n236, n240, n244, n248, n251 : std_logic;

begin
   DIFF <= ( DIFF_63_port, DIFF_62_port, DIFF_61_port, DIFF_60_port, 
      DIFF_59_port, DIFF_58_port, DIFF_57_port, DIFF_56_port, DIFF_55_port, 
      DIFF_54_port, DIFF_53_port, DIFF_52_port, DIFF_51_port, DIFF_50_port, 
      DIFF_49_port, DIFF_48_port, DIFF_47_port, DIFF_46_port, DIFF_45_port, 
      DIFF_44_port, DIFF_43_port, DIFF_42_port, DIFF_41_port, DIFF_40_port, 
      DIFF_39_port, DIFF_38_port, DIFF_37_port, DIFF_36_port, DIFF_35_port, 
      DIFF_34_port, DIFF_33_port, DIFF_32_port, DIFF_31_port, DIFF_30_port, 
      DIFF_29_port, DIFF_28_port, DIFF_27_port, DIFF_26_port, DIFF_25_port, 
      DIFF_24_port, DIFF_23_port, DIFF_22_port, DIFF_21_port, DIFF_20_port, 
      DIFF_19_port, DIFF_18_port, DIFF_17_port, DIFF_16_port, DIFF_15_port, 
      DIFF_14_port, DIFF_13_port, DIFF_12_port, DIFF_11_port, DIFF_10_port, 
      DIFF_9_port, DIFF_8_port, DIFF_7_port, DIFF_6_port, DIFF_5_port, 
      DIFF_4_port, DIFF_3_port, DIFF_2_port, DIFF_1_port, B(0) );
   
   U81 : XOR2_X1 port map( A => n190, B => B(9), Z => DIFF_9_port);
   U82 : XOR2_X1 port map( A => n192, B => B(7), Z => DIFF_7_port);
   U83 : XOR2_X1 port map( A => n193, B => B(6), Z => DIFF_6_port);
   U85 : XOR2_X1 port map( A => n196, B => B(62), Z => DIFF_62_port);
   U86 : XOR2_X1 port map( A => n194, B => B(5), Z => DIFF_5_port);
   U87 : XOR2_X1 port map( A => n198, B => B(59), Z => DIFF_59_port);
   U89 : XOR2_X1 port map( A => n200, B => B(57), Z => DIFF_57_port);
   U90 : XOR2_X1 port map( A => n202, B => B(55), Z => DIFF_55_port);
   U92 : XOR2_X1 port map( A => n204, B => B(53), Z => DIFF_53_port);
   U93 : XOR2_X1 port map( A => n206, B => B(51), Z => DIFF_51_port);
   U95 : XOR2_X1 port map( A => n208, B => B(49), Z => DIFF_49_port);
   U96 : XOR2_X1 port map( A => n212, B => B(47), Z => DIFF_47_port);
   U98 : XOR2_X1 port map( A => n214, B => B(45), Z => DIFF_45_port);
   U99 : XOR2_X1 port map( A => n216, B => B(43), Z => DIFF_43_port);
   U101 : XOR2_X1 port map( A => n218, B => B(41), Z => DIFF_41_port);
   U102 : XOR2_X1 port map( A => n211, B => B(3), Z => DIFF_3_port);
   U103 : XOR2_X1 port map( A => n220, B => B(39), Z => DIFF_39_port);
   U105 : XOR2_X1 port map( A => n222, B => B(37), Z => DIFF_37_port);
   U106 : XOR2_X1 port map( A => n224, B => B(35), Z => DIFF_35_port);
   U108 : XOR2_X1 port map( A => n226, B => B(33), Z => DIFF_33_port);
   U109 : XOR2_X1 port map( A => n228, B => B(31), Z => DIFF_31_port);
   U111 : XOR2_X1 port map( A => n230, B => B(29), Z => DIFF_29_port);
   U112 : XOR2_X1 port map( A => n233, B => B(27), Z => DIFF_27_port);
   U114 : XOR2_X1 port map( A => n235, B => B(25), Z => DIFF_25_port);
   U115 : XOR2_X1 port map( A => n237, B => B(23), Z => DIFF_23_port);
   U117 : XOR2_X1 port map( A => n239, B => B(21), Z => DIFF_21_port);
   U118 : XOR2_X1 port map( A => B(1), B => B(0), Z => DIFF_1_port);
   U119 : XOR2_X1 port map( A => n241, B => B(19), Z => DIFF_19_port);
   U121 : XOR2_X1 port map( A => n243, B => B(17), Z => DIFF_17_port);
   U122 : XOR2_X1 port map( A => n245, B => B(15), Z => DIFF_15_port);
   U124 : XOR2_X1 port map( A => n247, B => B(13), Z => DIFF_13_port);
   U125 : XOR2_X1 port map( A => n249, B => B(11), Z => DIFF_11_port);
   U1 : XNOR2_X1 port map( A => n189, B => B(46), ZN => DIFF_46_port);
   U2 : NOR2_X1 port map( A1 => n214, A2 => B(45), ZN => n189);
   U3 : XNOR2_X1 port map( A => n195, B => B(26), ZN => DIFF_26_port);
   U4 : NOR2_X1 port map( A1 => n235, A2 => B(25), ZN => n195);
   U5 : XNOR2_X1 port map( A => n201, B => B(22), ZN => DIFF_22_port);
   U6 : NOR2_X1 port map( A1 => n239, A2 => B(21), ZN => n201);
   U7 : XNOR2_X1 port map( A => n205, B => B(14), ZN => DIFF_14_port);
   U8 : NOR2_X1 port map( A1 => n247, A2 => B(13), ZN => n205);
   U9 : XNOR2_X1 port map( A => n209, B => B(18), ZN => DIFF_18_port);
   U10 : NOR2_X1 port map( A1 => n243, A2 => B(17), ZN => n209);
   U11 : XNOR2_X1 port map( A => n215, B => B(30), ZN => DIFF_30_port);
   U12 : NOR2_X1 port map( A1 => n230, A2 => B(29), ZN => n215);
   U13 : XNOR2_X1 port map( A => B(12), B => n250, ZN => DIFF_12_port);
   U14 : NOR2_X1 port map( A1 => B(11), A2 => n249, ZN => n250);
   U15 : XNOR2_X1 port map( A => B(24), B => n238, ZN => DIFF_24_port);
   U16 : NOR2_X1 port map( A1 => B(23), A2 => n237, ZN => n238);
   U17 : XNOR2_X1 port map( A => B(16), B => n246, ZN => DIFF_16_port);
   U18 : NOR2_X1 port map( A1 => B(15), A2 => n245, ZN => n246);
   U19 : XNOR2_X1 port map( A => B(20), B => n242, ZN => DIFF_20_port);
   U20 : NOR2_X1 port map( A1 => B(19), A2 => n241, ZN => n242);
   U21 : XNOR2_X1 port map( A => B(44), B => n217, ZN => DIFF_44_port);
   U22 : NOR2_X1 port map( A1 => B(43), A2 => n216, ZN => n217);
   U23 : XNOR2_X1 port map( A => B(28), B => n234, ZN => DIFF_28_port);
   U24 : NOR2_X1 port map( A1 => B(27), A2 => n233, ZN => n234);
   U25 : XNOR2_X1 port map( A => B(36), B => n225, ZN => DIFF_36_port);
   U26 : NOR2_X1 port map( A1 => B(35), A2 => n224, ZN => n225);
   U27 : XNOR2_X1 port map( A => B(32), B => n229, ZN => DIFF_32_port);
   U28 : NOR2_X1 port map( A1 => B(31), A2 => n228, ZN => n229);
   U29 : XNOR2_X1 port map( A => B(40), B => n221, ZN => DIFF_40_port);
   U30 : NOR2_X1 port map( A1 => B(39), A2 => n220, ZN => n221);
   U31 : OR3_X1 port map( A1 => B(45), A2 => B(46), A3 => n214, ZN => n212);
   U32 : OR3_X1 port map( A1 => B(17), A2 => B(18), A3 => n243, ZN => n241);
   U33 : OR3_X1 port map( A1 => B(21), A2 => B(22), A3 => n239, ZN => n237);
   U34 : OR3_X1 port map( A1 => B(13), A2 => B(14), A3 => n247, ZN => n245);
   U35 : OR3_X1 port map( A1 => B(25), A2 => B(26), A3 => n235, ZN => n233);
   U36 : OR3_X1 port map( A1 => B(29), A2 => B(30), A3 => n230, ZN => n228);
   U37 : OR3_X1 port map( A1 => B(33), A2 => B(34), A3 => n226, ZN => n224);
   U38 : OR3_X1 port map( A1 => B(37), A2 => B(38), A3 => n222, ZN => n220);
   U39 : OR3_X1 port map( A1 => B(19), A2 => B(20), A3 => n241, ZN => n239);
   U40 : OR3_X1 port map( A1 => B(15), A2 => B(16), A3 => n245, ZN => n243);
   U41 : OR3_X1 port map( A1 => B(11), A2 => B(12), A3 => n249, ZN => n247);
   U42 : OR3_X1 port map( A1 => B(23), A2 => B(24), A3 => n237, ZN => n235);
   U43 : OR3_X1 port map( A1 => B(27), A2 => B(28), A3 => n233, ZN => n230);
   U44 : OR3_X1 port map( A1 => B(31), A2 => B(32), A3 => n228, ZN => n226);
   U45 : OR3_X1 port map( A1 => B(35), A2 => B(36), A3 => n224, ZN => n222);
   U46 : OR3_X1 port map( A1 => B(43), A2 => B(44), A3 => n216, ZN => n214);
   U47 : OR3_X1 port map( A1 => B(39), A2 => B(40), A3 => n220, ZN => n218);
   U48 : XNOR2_X1 port map( A => n219, B => B(38), ZN => DIFF_38_port);
   U49 : NOR2_X1 port map( A1 => n222, A2 => B(37), ZN => n219);
   U50 : XNOR2_X1 port map( A => n223, B => B(34), ZN => DIFF_34_port);
   U51 : NOR2_X1 port map( A1 => n226, A2 => B(33), ZN => n223);
   U52 : NOR3_X1 port map( A1 => B(59), A2 => B(60), A3 => n198, ZN => n197);
   U53 : XNOR2_X1 port map( A => n227, B => B(50), ZN => DIFF_50_port);
   U54 : NOR2_X1 port map( A1 => n208, A2 => B(49), ZN => n227);
   U55 : XNOR2_X1 port map( A => n231, B => B(54), ZN => DIFF_54_port);
   U56 : NOR2_X1 port map( A1 => n204, A2 => B(53), ZN => n231);
   U57 : XNOR2_X1 port map( A => B(48), B => n213, ZN => DIFF_48_port);
   U58 : NOR2_X1 port map( A1 => B(47), A2 => n212, ZN => n213);
   U59 : XNOR2_X1 port map( A => B(60), B => n199, ZN => DIFF_60_port);
   U60 : NOR2_X1 port map( A1 => B(59), A2 => n198, ZN => n199);
   U61 : XNOR2_X1 port map( A => B(56), B => n203, ZN => DIFF_56_port);
   U62 : NOR2_X1 port map( A1 => B(55), A2 => n202, ZN => n203);
   U63 : XOR2_X1 port map( A => n197, B => n251, Z => DIFF_61_port);
   U64 : NAND2_X1 port map( A1 => n197, A2 => n251, ZN => n196);
   U65 : OR3_X1 port map( A1 => B(57), A2 => B(58), A3 => n200, ZN => n198);
   U66 : OR3_X1 port map( A1 => B(49), A2 => B(50), A3 => n208, ZN => n206);
   U67 : OR3_X1 port map( A1 => B(53), A2 => B(54), A3 => n204, ZN => n202);
   U68 : OR3_X1 port map( A1 => B(47), A2 => B(48), A3 => n212, ZN => n208);
   U69 : OR3_X1 port map( A1 => B(55), A2 => B(56), A3 => n202, ZN => n200);
   U70 : XNOR2_X1 port map( A => n236, B => B(58), ZN => DIFF_58_port);
   U71 : NOR2_X1 port map( A1 => n200, A2 => B(57), ZN => n236);
   U72 : XNOR2_X1 port map( A => n240, B => B(10), ZN => DIFF_10_port);
   U73 : NOR2_X1 port map( A1 => n190, A2 => B(9), ZN => n240);
   U74 : XNOR2_X1 port map( A => n244, B => B(42), ZN => DIFF_42_port);
   U75 : NOR2_X1 port map( A1 => n218, A2 => B(41), ZN => n244);
   U76 : OR3_X1 port map( A1 => B(10), A2 => B(9), A3 => n190, ZN => n249);
   U77 : OR3_X1 port map( A1 => B(41), A2 => B(42), A3 => n218, ZN => n216);
   U78 : XNOR2_X1 port map( A => n248, B => B(63), ZN => DIFF_63_port);
   U79 : NOR2_X1 port map( A1 => n196, A2 => B(62), ZN => n248);
   U80 : XNOR2_X1 port map( A => B(52), B => n207, ZN => DIFF_52_port);
   U84 : NOR2_X1 port map( A1 => B(51), A2 => n206, ZN => n207);
   U88 : OR3_X1 port map( A1 => B(51), A2 => B(52), A3 => n206, ZN => n204);
   U91 : OR3_X1 port map( A1 => B(7), A2 => B(8), A3 => n192, ZN => n190);
   U94 : XNOR2_X1 port map( A => B(8), B => n191, ZN => DIFF_8_port);
   U97 : NOR2_X1 port map( A1 => B(7), A2 => n192, ZN => n191);
   U100 : NOR2_X1 port map( A1 => B(3), A2 => n211, ZN => n210);
   U104 : OR3_X1 port map( A1 => B(5), A2 => B(6), A3 => n194, ZN => n192);
   U107 : OR3_X1 port map( A1 => B(3), A2 => B(4), A3 => n211, ZN => n194);
   U110 : XNOR2_X1 port map( A => B(4), B => n210, ZN => DIFF_4_port);
   U113 : XNOR2_X1 port map( A => B(2), B => n232, ZN => DIFF_2_port);
   U116 : OR2_X1 port map( A1 => n194, A2 => B(5), ZN => n193);
   U120 : OR3_X1 port map( A1 => B(1), A2 => B(2), A3 => B(0), ZN => n211);
   U123 : NOR2_X1 port map( A1 => B(0), A2 => B(1), ZN => n232);
   U126 : INV_X1 port map( A => B(61), ZN => n251);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_25_DW01_sub_0 is

   port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (63 downto 0);  CO : out std_logic);

end complementer_N64_25_DW01_sub_0;

architecture SYN_rpl of complementer_N64_25_DW01_sub_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal DIFF_62_port, DIFF_63_port, DIFF_7_port, DIFF_8_port, DIFF_9_port, 
      DIFF_10_port, DIFF_11_port, DIFF_12_port, DIFF_13_port, DIFF_14_port, 
      DIFF_15_port, DIFF_16_port, DIFF_17_port, DIFF_18_port, DIFF_19_port, 
      DIFF_20_port, DIFF_21_port, DIFF_22_port, DIFF_23_port, DIFF_24_port, 
      DIFF_25_port, DIFF_26_port, DIFF_27_port, DIFF_28_port, DIFF_29_port, 
      DIFF_30_port, DIFF_31_port, DIFF_32_port, DIFF_33_port, DIFF_34_port, 
      DIFF_35_port, DIFF_36_port, DIFF_37_port, DIFF_38_port, DIFF_39_port, 
      DIFF_40_port, DIFF_41_port, DIFF_42_port, DIFF_43_port, DIFF_44_port, 
      DIFF_45_port, DIFF_46_port, DIFF_47_port, DIFF_48_port, DIFF_49_port, 
      DIFF_50_port, DIFF_51_port, DIFF_52_port, DIFF_53_port, DIFF_54_port, 
      DIFF_55_port, DIFF_56_port, DIFF_57_port, DIFF_58_port, DIFF_59_port, 
      DIFF_60_port, DIFF_61_port, DIFF_3_port, DIFF_4_port, DIFF_5_port, 
      DIFF_6_port, DIFF_2_port, DIFF_1_port, n190, n191, n192, n193, n194, n196
      , n197, n198, n199, n200, n202, n203, n204, n206, n207, n208, n210, n211,
      n212, n213, n214, n216, n217, n218, n220, n221, n222, n224, n225, n226, 
      n228, n229, n230, n232, n233, n234, n235, n237, n238, n239, n241, n242, 
      n243, n245, n246, n247, n249, n250, n189, n195, n201, n205, n209, n215, 
      n219, n223, n227, n231, n236, n240, n244, n248, n251 : std_logic;

begin
   DIFF <= ( DIFF_63_port, DIFF_62_port, DIFF_61_port, DIFF_60_port, 
      DIFF_59_port, DIFF_58_port, DIFF_57_port, DIFF_56_port, DIFF_55_port, 
      DIFF_54_port, DIFF_53_port, DIFF_52_port, DIFF_51_port, DIFF_50_port, 
      DIFF_49_port, DIFF_48_port, DIFF_47_port, DIFF_46_port, DIFF_45_port, 
      DIFF_44_port, DIFF_43_port, DIFF_42_port, DIFF_41_port, DIFF_40_port, 
      DIFF_39_port, DIFF_38_port, DIFF_37_port, DIFF_36_port, DIFF_35_port, 
      DIFF_34_port, DIFF_33_port, DIFF_32_port, DIFF_31_port, DIFF_30_port, 
      DIFF_29_port, DIFF_28_port, DIFF_27_port, DIFF_26_port, DIFF_25_port, 
      DIFF_24_port, DIFF_23_port, DIFF_22_port, DIFF_21_port, DIFF_20_port, 
      DIFF_19_port, DIFF_18_port, DIFF_17_port, DIFF_16_port, DIFF_15_port, 
      DIFF_14_port, DIFF_13_port, DIFF_12_port, DIFF_11_port, DIFF_10_port, 
      DIFF_9_port, DIFF_8_port, DIFF_7_port, DIFF_6_port, DIFF_5_port, 
      DIFF_4_port, DIFF_3_port, DIFF_2_port, DIFF_1_port, B(0) );
   
   U81 : XOR2_X1 port map( A => n190, B => B(9), Z => DIFF_9_port);
   U82 : XOR2_X1 port map( A => n192, B => B(7), Z => DIFF_7_port);
   U83 : XOR2_X1 port map( A => n193, B => B(6), Z => DIFF_6_port);
   U85 : XOR2_X1 port map( A => n196, B => B(62), Z => DIFF_62_port);
   U86 : XOR2_X1 port map( A => n194, B => B(5), Z => DIFF_5_port);
   U87 : XOR2_X1 port map( A => n198, B => B(59), Z => DIFF_59_port);
   U89 : XOR2_X1 port map( A => n200, B => B(57), Z => DIFF_57_port);
   U90 : XOR2_X1 port map( A => n202, B => B(55), Z => DIFF_55_port);
   U92 : XOR2_X1 port map( A => n204, B => B(53), Z => DIFF_53_port);
   U93 : XOR2_X1 port map( A => n206, B => B(51), Z => DIFF_51_port);
   U95 : XOR2_X1 port map( A => n208, B => B(49), Z => DIFF_49_port);
   U96 : XOR2_X1 port map( A => n212, B => B(47), Z => DIFF_47_port);
   U98 : XOR2_X1 port map( A => n214, B => B(45), Z => DIFF_45_port);
   U99 : XOR2_X1 port map( A => n216, B => B(43), Z => DIFF_43_port);
   U101 : XOR2_X1 port map( A => n218, B => B(41), Z => DIFF_41_port);
   U102 : XOR2_X1 port map( A => n211, B => B(3), Z => DIFF_3_port);
   U103 : XOR2_X1 port map( A => n220, B => B(39), Z => DIFF_39_port);
   U105 : XOR2_X1 port map( A => n222, B => B(37), Z => DIFF_37_port);
   U106 : XOR2_X1 port map( A => n224, B => B(35), Z => DIFF_35_port);
   U108 : XOR2_X1 port map( A => n226, B => B(33), Z => DIFF_33_port);
   U109 : XOR2_X1 port map( A => n228, B => B(31), Z => DIFF_31_port);
   U111 : XOR2_X1 port map( A => n230, B => B(29), Z => DIFF_29_port);
   U112 : XOR2_X1 port map( A => n233, B => B(27), Z => DIFF_27_port);
   U114 : XOR2_X1 port map( A => n235, B => B(25), Z => DIFF_25_port);
   U115 : XOR2_X1 port map( A => n237, B => B(23), Z => DIFF_23_port);
   U117 : XOR2_X1 port map( A => n239, B => B(21), Z => DIFF_21_port);
   U118 : XOR2_X1 port map( A => B(1), B => B(0), Z => DIFF_1_port);
   U119 : XOR2_X1 port map( A => n241, B => B(19), Z => DIFF_19_port);
   U121 : XOR2_X1 port map( A => n243, B => B(17), Z => DIFF_17_port);
   U122 : XOR2_X1 port map( A => n245, B => B(15), Z => DIFF_15_port);
   U124 : XOR2_X1 port map( A => n247, B => B(13), Z => DIFF_13_port);
   U125 : XOR2_X1 port map( A => n249, B => B(11), Z => DIFF_11_port);
   U1 : XNOR2_X1 port map( A => n189, B => B(10), ZN => DIFF_10_port);
   U2 : NOR2_X1 port map( A1 => n190, A2 => B(9), ZN => n189);
   U3 : XNOR2_X1 port map( A => n195, B => B(30), ZN => DIFF_30_port);
   U4 : NOR2_X1 port map( A1 => n230, A2 => B(29), ZN => n195);
   U5 : XNOR2_X1 port map( A => n201, B => B(26), ZN => DIFF_26_port);
   U6 : NOR2_X1 port map( A1 => n235, A2 => B(25), ZN => n201);
   U7 : XNOR2_X1 port map( A => n205, B => B(18), ZN => DIFF_18_port);
   U8 : NOR2_X1 port map( A1 => n243, A2 => B(17), ZN => n205);
   U9 : XNOR2_X1 port map( A => n209, B => B(22), ZN => DIFF_22_port);
   U10 : NOR2_X1 port map( A1 => n239, A2 => B(21), ZN => n209);
   U11 : XNOR2_X1 port map( A => B(36), B => n225, ZN => DIFF_36_port);
   U12 : NOR2_X1 port map( A1 => B(35), A2 => n224, ZN => n225);
   U13 : XNOR2_X1 port map( A => B(12), B => n250, ZN => DIFF_12_port);
   U14 : NOR2_X1 port map( A1 => B(11), A2 => n249, ZN => n250);
   U15 : XNOR2_X1 port map( A => B(16), B => n246, ZN => DIFF_16_port);
   U16 : NOR2_X1 port map( A1 => B(15), A2 => n245, ZN => n246);
   U17 : XNOR2_X1 port map( A => B(28), B => n234, ZN => DIFF_28_port);
   U18 : NOR2_X1 port map( A1 => B(27), A2 => n233, ZN => n234);
   U19 : XNOR2_X1 port map( A => B(20), B => n242, ZN => DIFF_20_port);
   U20 : NOR2_X1 port map( A1 => B(19), A2 => n241, ZN => n242);
   U21 : XNOR2_X1 port map( A => B(24), B => n238, ZN => DIFF_24_port);
   U22 : NOR2_X1 port map( A1 => B(23), A2 => n237, ZN => n238);
   U23 : XNOR2_X1 port map( A => B(32), B => n229, ZN => DIFF_32_port);
   U24 : NOR2_X1 port map( A1 => B(31), A2 => n228, ZN => n229);
   U25 : XNOR2_X1 port map( A => B(44), B => n217, ZN => DIFF_44_port);
   U26 : NOR2_X1 port map( A1 => B(43), A2 => n216, ZN => n217);
   U27 : OR3_X1 port map( A1 => B(17), A2 => B(18), A3 => n243, ZN => n241);
   U28 : OR3_X1 port map( A1 => B(21), A2 => B(22), A3 => n239, ZN => n237);
   U29 : OR3_X1 port map( A1 => B(13), A2 => B(14), A3 => n247, ZN => n245);
   U30 : OR3_X1 port map( A1 => B(25), A2 => B(26), A3 => n235, ZN => n233);
   U31 : OR3_X1 port map( A1 => B(29), A2 => B(30), A3 => n230, ZN => n228);
   U32 : OR3_X1 port map( A1 => B(33), A2 => B(34), A3 => n226, ZN => n224);
   U33 : OR3_X1 port map( A1 => B(37), A2 => B(38), A3 => n222, ZN => n220);
   U34 : OR3_X1 port map( A1 => B(10), A2 => B(9), A3 => n190, ZN => n249);
   U35 : OR3_X1 port map( A1 => B(15), A2 => B(16), A3 => n245, ZN => n243);
   U36 : OR3_X1 port map( A1 => B(19), A2 => B(20), A3 => n241, ZN => n239);
   U37 : OR3_X1 port map( A1 => B(11), A2 => B(12), A3 => n249, ZN => n247);
   U38 : OR3_X1 port map( A1 => B(23), A2 => B(24), A3 => n237, ZN => n235);
   U39 : OR3_X1 port map( A1 => B(27), A2 => B(28), A3 => n233, ZN => n230);
   U40 : OR3_X1 port map( A1 => B(31), A2 => B(32), A3 => n228, ZN => n226);
   U41 : OR3_X1 port map( A1 => B(35), A2 => B(36), A3 => n224, ZN => n222);
   U42 : OR3_X1 port map( A1 => B(43), A2 => B(44), A3 => n216, ZN => n214);
   U43 : XNOR2_X1 port map( A => n215, B => B(14), ZN => DIFF_14_port);
   U44 : NOR2_X1 port map( A1 => n247, A2 => B(13), ZN => n215);
   U45 : XNOR2_X1 port map( A => n219, B => B(34), ZN => DIFF_34_port);
   U46 : NOR2_X1 port map( A1 => n226, A2 => B(33), ZN => n219);
   U47 : XNOR2_X1 port map( A => n223, B => B(38), ZN => DIFF_38_port);
   U48 : NOR2_X1 port map( A1 => n222, A2 => B(37), ZN => n223);
   U49 : XNOR2_X1 port map( A => n227, B => B(54), ZN => DIFF_54_port);
   U50 : NOR2_X1 port map( A1 => n204, A2 => B(53), ZN => n227);
   U51 : XOR2_X1 port map( A => n197, B => n251, Z => DIFF_61_port);
   U52 : NAND2_X1 port map( A1 => n197, A2 => n251, ZN => n196);
   U53 : OR3_X1 port map( A1 => B(53), A2 => B(54), A3 => n204, ZN => n202);
   U54 : XNOR2_X1 port map( A => n231, B => B(50), ZN => DIFF_50_port);
   U55 : NOR2_X1 port map( A1 => n208, A2 => B(49), ZN => n231);
   U56 : XNOR2_X1 port map( A => n236, B => B(42), ZN => DIFF_42_port);
   U57 : NOR2_X1 port map( A1 => n218, A2 => B(41), ZN => n236);
   U58 : XNOR2_X1 port map( A => n240, B => B(46), ZN => DIFF_46_port);
   U59 : NOR2_X1 port map( A1 => n214, A2 => B(45), ZN => n240);
   U60 : XNOR2_X1 port map( A => B(48), B => n213, ZN => DIFF_48_port);
   U61 : NOR2_X1 port map( A1 => B(47), A2 => n212, ZN => n213);
   U62 : XNOR2_X1 port map( A => B(40), B => n221, ZN => DIFF_40_port);
   U63 : NOR2_X1 port map( A1 => B(39), A2 => n220, ZN => n221);
   U64 : XNOR2_X1 port map( A => B(8), B => n191, ZN => DIFF_8_port);
   U65 : NOR2_X1 port map( A1 => B(7), A2 => n192, ZN => n191);
   U66 : XNOR2_X1 port map( A => B(52), B => n207, ZN => DIFF_52_port);
   U67 : NOR2_X1 port map( A1 => B(51), A2 => n206, ZN => n207);
   U68 : OR3_X1 port map( A1 => B(45), A2 => B(46), A3 => n214, ZN => n212);
   U69 : OR3_X1 port map( A1 => B(49), A2 => B(50), A3 => n208, ZN => n206);
   U70 : OR3_X1 port map( A1 => B(41), A2 => B(42), A3 => n218, ZN => n216);
   U71 : OR3_X1 port map( A1 => B(7), A2 => B(8), A3 => n192, ZN => n190);
   U72 : OR3_X1 port map( A1 => B(47), A2 => B(48), A3 => n212, ZN => n208);
   U73 : OR3_X1 port map( A1 => B(39), A2 => B(40), A3 => n220, ZN => n218);
   U74 : NOR3_X1 port map( A1 => B(59), A2 => B(60), A3 => n198, ZN => n197);
   U75 : XNOR2_X1 port map( A => n244, B => B(58), ZN => DIFF_58_port);
   U76 : NOR2_X1 port map( A1 => n200, A2 => B(57), ZN => n244);
   U77 : XNOR2_X1 port map( A => n248, B => B(63), ZN => DIFF_63_port);
   U78 : NOR2_X1 port map( A1 => n196, A2 => B(62), ZN => n248);
   U79 : XNOR2_X1 port map( A => B(60), B => n199, ZN => DIFF_60_port);
   U80 : NOR2_X1 port map( A1 => B(59), A2 => n198, ZN => n199);
   U84 : XNOR2_X1 port map( A => B(56), B => n203, ZN => DIFF_56_port);
   U88 : NOR2_X1 port map( A1 => B(55), A2 => n202, ZN => n203);
   U91 : OR3_X1 port map( A1 => B(57), A2 => B(58), A3 => n200, ZN => n198);
   U94 : OR3_X1 port map( A1 => B(51), A2 => B(52), A3 => n206, ZN => n204);
   U97 : OR3_X1 port map( A1 => B(55), A2 => B(56), A3 => n202, ZN => n200);
   U100 : XNOR2_X1 port map( A => B(2), B => n232, ZN => DIFF_2_port);
   U104 : NOR2_X1 port map( A1 => B(0), A2 => B(1), ZN => n232);
   U107 : XNOR2_X1 port map( A => B(4), B => n210, ZN => DIFF_4_port);
   U110 : NOR2_X1 port map( A1 => B(3), A2 => n211, ZN => n210);
   U113 : OR3_X1 port map( A1 => B(5), A2 => B(6), A3 => n194, ZN => n192);
   U116 : OR3_X1 port map( A1 => B(3), A2 => B(4), A3 => n211, ZN => n194);
   U120 : OR2_X1 port map( A1 => n194, A2 => B(5), ZN => n193);
   U123 : OR3_X1 port map( A1 => B(1), A2 => B(2), A3 => B(0), ZN => n211);
   U126 : INV_X1 port map( A => B(61), ZN => n251);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_26_DW01_sub_0 is

   port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (63 downto 0);  CO : out std_logic);

end complementer_N64_26_DW01_sub_0;

architecture SYN_rpl of complementer_N64_26_DW01_sub_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal DIFF_62_port, DIFF_61_port, DIFF_60_port, DIFF_59_port, DIFF_58_port,
      DIFF_57_port, DIFF_56_port, DIFF_55_port, DIFF_54_port, DIFF_53_port, 
      DIFF_52_port, DIFF_51_port, DIFF_50_port, DIFF_49_port, DIFF_48_port, 
      DIFF_47_port, DIFF_46_port, DIFF_45_port, DIFF_44_port, DIFF_43_port, 
      DIFF_42_port, DIFF_41_port, DIFF_40_port, DIFF_39_port, DIFF_38_port, 
      DIFF_37_port, DIFF_36_port, DIFF_35_port, DIFF_34_port, DIFF_33_port, 
      DIFF_32_port, DIFF_31_port, DIFF_30_port, DIFF_29_port, DIFF_28_port, 
      DIFF_27_port, DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, 
      DIFF_22_port, DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, 
      DIFF_17_port, DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, 
      DIFF_12_port, DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, 
      DIFF_7_port, DIFF_6_port, DIFF_5_port, DIFF_4_port, DIFF_3_port, 
      DIFF_2_port, DIFF_1_port, DIFF_63_port, n190, n191, n192, n194, n195, 
      n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, 
      n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, 
      n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, 
      n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, 
      n244, n245, n246, n247, n248, n249, n250, n251, n189, n193 : std_logic;

begin
   DIFF <= ( DIFF_63_port, DIFF_62_port, DIFF_61_port, DIFF_60_port, 
      DIFF_59_port, DIFF_58_port, DIFF_57_port, DIFF_56_port, DIFF_55_port, 
      DIFF_54_port, DIFF_53_port, DIFF_52_port, DIFF_51_port, DIFF_50_port, 
      DIFF_49_port, DIFF_48_port, DIFF_47_port, DIFF_46_port, DIFF_45_port, 
      DIFF_44_port, DIFF_43_port, DIFF_42_port, DIFF_41_port, DIFF_40_port, 
      DIFF_39_port, DIFF_38_port, DIFF_37_port, DIFF_36_port, DIFF_35_port, 
      DIFF_34_port, DIFF_33_port, DIFF_32_port, DIFF_31_port, DIFF_30_port, 
      DIFF_29_port, DIFF_28_port, DIFF_27_port, DIFF_26_port, DIFF_25_port, 
      DIFF_24_port, DIFF_23_port, DIFF_22_port, DIFF_21_port, DIFF_20_port, 
      DIFF_19_port, DIFF_18_port, DIFF_17_port, DIFF_16_port, DIFF_15_port, 
      DIFF_14_port, DIFF_13_port, DIFF_12_port, DIFF_11_port, DIFF_10_port, 
      DIFF_9_port, DIFF_8_port, DIFF_7_port, DIFF_6_port, DIFF_5_port, 
      DIFF_4_port, DIFF_3_port, DIFF_2_port, DIFF_1_port, B(0) );
   
   U81 : XOR2_X1 port map( A => n190, B => B(9), Z => DIFF_9_port);
   U82 : XOR2_X1 port map( A => n192, B => B(7), Z => DIFF_7_port);
   U84 : XOR2_X1 port map( A => n195, B => B(63), Z => DIFF_63_port);
   U85 : XOR2_X1 port map( A => n196, B => B(62), Z => DIFF_62_port);
   U86 : XOR2_X1 port map( A => n194, B => B(5), Z => DIFF_5_port);
   U87 : XOR2_X1 port map( A => n198, B => B(59), Z => DIFF_59_port);
   U88 : XOR2_X1 port map( A => n201, B => B(58), Z => DIFF_58_port);
   U89 : XOR2_X1 port map( A => n200, B => B(57), Z => DIFF_57_port);
   U90 : XOR2_X1 port map( A => n202, B => B(55), Z => DIFF_55_port);
   U91 : XOR2_X1 port map( A => n205, B => B(54), Z => DIFF_54_port);
   U92 : XOR2_X1 port map( A => n204, B => B(53), Z => DIFF_53_port);
   U93 : XOR2_X1 port map( A => n206, B => B(51), Z => DIFF_51_port);
   U94 : XOR2_X1 port map( A => n209, B => B(50), Z => DIFF_50_port);
   U95 : XOR2_X1 port map( A => n208, B => B(49), Z => DIFF_49_port);
   U96 : XOR2_X1 port map( A => n212, B => B(47), Z => DIFF_47_port);
   U97 : XOR2_X1 port map( A => n215, B => B(46), Z => DIFF_46_port);
   U98 : XOR2_X1 port map( A => n214, B => B(45), Z => DIFF_45_port);
   U99 : XOR2_X1 port map( A => n216, B => B(43), Z => DIFF_43_port);
   U100 : XOR2_X1 port map( A => n219, B => B(42), Z => DIFF_42_port);
   U101 : XOR2_X1 port map( A => n218, B => B(41), Z => DIFF_41_port);
   U102 : XOR2_X1 port map( A => n211, B => B(3), Z => DIFF_3_port);
   U103 : XOR2_X1 port map( A => n220, B => B(39), Z => DIFF_39_port);
   U104 : XOR2_X1 port map( A => n223, B => B(38), Z => DIFF_38_port);
   U105 : XOR2_X1 port map( A => n222, B => B(37), Z => DIFF_37_port);
   U106 : XOR2_X1 port map( A => n224, B => B(35), Z => DIFF_35_port);
   U107 : XOR2_X1 port map( A => n227, B => B(34), Z => DIFF_34_port);
   U108 : XOR2_X1 port map( A => n226, B => B(33), Z => DIFF_33_port);
   U109 : XOR2_X1 port map( A => n228, B => B(31), Z => DIFF_31_port);
   U110 : XOR2_X1 port map( A => n231, B => B(30), Z => DIFF_30_port);
   U111 : XOR2_X1 port map( A => n230, B => B(29), Z => DIFF_29_port);
   U112 : XOR2_X1 port map( A => n233, B => B(27), Z => DIFF_27_port);
   U113 : XOR2_X1 port map( A => n236, B => B(26), Z => DIFF_26_port);
   U114 : XOR2_X1 port map( A => n235, B => B(25), Z => DIFF_25_port);
   U115 : XOR2_X1 port map( A => n237, B => B(23), Z => DIFF_23_port);
   U116 : XOR2_X1 port map( A => n240, B => B(22), Z => DIFF_22_port);
   U117 : XOR2_X1 port map( A => n239, B => B(21), Z => DIFF_21_port);
   U118 : XOR2_X1 port map( A => B(1), B => B(0), Z => DIFF_1_port);
   U119 : XOR2_X1 port map( A => n241, B => B(19), Z => DIFF_19_port);
   U120 : XOR2_X1 port map( A => n244, B => B(18), Z => DIFF_18_port);
   U121 : XOR2_X1 port map( A => n243, B => B(17), Z => DIFF_17_port);
   U122 : XOR2_X1 port map( A => n245, B => B(15), Z => DIFF_15_port);
   U123 : XOR2_X1 port map( A => n248, B => B(14), Z => DIFF_14_port);
   U124 : XOR2_X1 port map( A => n247, B => B(13), Z => DIFF_13_port);
   U125 : XOR2_X1 port map( A => n249, B => B(11), Z => DIFF_11_port);
   U126 : XOR2_X1 port map( A => n251, B => B(10), Z => DIFF_10_port);
   U1 : NOR2_X1 port map( A1 => B(47), A2 => n212, ZN => n213);
   U2 : NOR2_X1 port map( A1 => B(43), A2 => n216, ZN => n217);
   U3 : OR3_X1 port map( A1 => B(37), A2 => B(38), A3 => n222, ZN => n220);
   U4 : OR3_X1 port map( A1 => B(47), A2 => B(48), A3 => n212, ZN => n208);
   U5 : OR3_X1 port map( A1 => B(43), A2 => B(44), A3 => n216, ZN => n214);
   U6 : XNOR2_X1 port map( A => B(48), B => n213, ZN => DIFF_48_port);
   U7 : XNOR2_X1 port map( A => B(36), B => n225, ZN => DIFF_36_port);
   U8 : XNOR2_X1 port map( A => B(44), B => n217, ZN => DIFF_44_port);
   U9 : OR2_X1 port map( A1 => n222, A2 => B(37), ZN => n223);
   U10 : NAND2_X1 port map( A1 => n197, A2 => n193, ZN => n196);
   U11 : OR3_X1 port map( A1 => B(57), A2 => B(58), A3 => n200, ZN => n198);
   U12 : OR3_X1 port map( A1 => B(53), A2 => B(54), A3 => n204, ZN => n202);
   U13 : OR2_X1 port map( A1 => n200, A2 => B(57), ZN => n201);
   U14 : OR2_X1 port map( A1 => n204, A2 => B(53), ZN => n205);
   U15 : NOR2_X1 port map( A1 => B(7), A2 => n192, ZN => n191);
   U16 : NOR2_X1 port map( A1 => B(11), A2 => n249, ZN => n250);
   U17 : NOR2_X1 port map( A1 => B(15), A2 => n245, ZN => n246);
   U18 : NOR2_X1 port map( A1 => B(27), A2 => n233, ZN => n234);
   U19 : NOR2_X1 port map( A1 => B(19), A2 => n241, ZN => n242);
   U20 : NOR2_X1 port map( A1 => B(23), A2 => n237, ZN => n238);
   U21 : NOR2_X1 port map( A1 => B(35), A2 => n224, ZN => n225);
   U22 : NOR2_X1 port map( A1 => B(31), A2 => n228, ZN => n229);
   U23 : NOR2_X1 port map( A1 => B(39), A2 => n220, ZN => n221);
   U24 : XNOR2_X1 port map( A => B(8), B => n191, ZN => DIFF_8_port);
   U25 : OR3_X1 port map( A1 => B(49), A2 => B(50), A3 => n208, ZN => n206);
   U26 : OR3_X1 port map( A1 => B(45), A2 => B(46), A3 => n214, ZN => n212);
   U27 : OR3_X1 port map( A1 => B(25), A2 => B(26), A3 => n235, ZN => n233);
   U28 : OR3_X1 port map( A1 => B(13), A2 => B(14), A3 => n247, ZN => n245);
   U29 : OR3_X1 port map( A1 => B(17), A2 => B(18), A3 => n243, ZN => n241);
   U30 : OR3_X1 port map( A1 => B(21), A2 => B(22), A3 => n239, ZN => n237);
   U31 : OR3_X1 port map( A1 => B(41), A2 => B(42), A3 => n218, ZN => n216);
   U32 : OR3_X1 port map( A1 => B(33), A2 => B(34), A3 => n226, ZN => n224);
   U33 : OR3_X1 port map( A1 => B(29), A2 => B(30), A3 => n230, ZN => n228);
   U34 : OR3_X1 port map( A1 => B(10), A2 => B(9), A3 => n190, ZN => n249);
   U35 : OR3_X1 port map( A1 => B(7), A2 => B(8), A3 => n192, ZN => n190);
   U36 : OR3_X1 port map( A1 => B(11), A2 => B(12), A3 => n249, ZN => n247);
   U37 : OR3_X1 port map( A1 => B(15), A2 => B(16), A3 => n245, ZN => n243);
   U38 : OR3_X1 port map( A1 => B(19), A2 => B(20), A3 => n241, ZN => n239);
   U39 : OR3_X1 port map( A1 => B(23), A2 => B(24), A3 => n237, ZN => n235);
   U40 : OR3_X1 port map( A1 => B(27), A2 => B(28), A3 => n233, ZN => n230);
   U41 : OR3_X1 port map( A1 => B(35), A2 => B(36), A3 => n224, ZN => n222);
   U42 : OR3_X1 port map( A1 => B(31), A2 => B(32), A3 => n228, ZN => n226);
   U43 : OR3_X1 port map( A1 => B(39), A2 => B(40), A3 => n220, ZN => n218);
   U44 : XNOR2_X1 port map( A => B(40), B => n221, ZN => DIFF_40_port);
   U45 : XNOR2_X1 port map( A => B(12), B => n250, ZN => DIFF_12_port);
   U46 : XNOR2_X1 port map( A => B(16), B => n246, ZN => DIFF_16_port);
   U47 : XNOR2_X1 port map( A => B(28), B => n234, ZN => DIFF_28_port);
   U48 : XNOR2_X1 port map( A => B(20), B => n242, ZN => DIFF_20_port);
   U49 : XNOR2_X1 port map( A => B(24), B => n238, ZN => DIFF_24_port);
   U50 : XNOR2_X1 port map( A => B(52), B => n207, ZN => DIFF_52_port);
   U51 : XNOR2_X1 port map( A => B(32), B => n229, ZN => DIFF_32_port);
   U52 : OR2_X1 port map( A1 => n208, A2 => B(49), ZN => n209);
   U53 : OR2_X1 port map( A1 => n190, A2 => B(9), ZN => n251);
   U54 : OR2_X1 port map( A1 => n247, A2 => B(13), ZN => n248);
   U55 : OR2_X1 port map( A1 => n230, A2 => B(29), ZN => n231);
   U56 : OR2_X1 port map( A1 => n235, A2 => B(25), ZN => n236);
   U57 : OR2_X1 port map( A1 => n243, A2 => B(17), ZN => n244);
   U58 : OR2_X1 port map( A1 => n239, A2 => B(21), ZN => n240);
   U59 : OR2_X1 port map( A1 => n218, A2 => B(41), ZN => n219);
   U60 : OR2_X1 port map( A1 => n226, A2 => B(33), ZN => n227);
   U61 : OR2_X1 port map( A1 => n214, A2 => B(45), ZN => n215);
   U62 : NOR3_X1 port map( A1 => B(59), A2 => B(60), A3 => n198, ZN => n197);
   U63 : XNOR2_X1 port map( A => n197, B => B(61), ZN => DIFF_61_port);
   U64 : XNOR2_X1 port map( A => B(60), B => n199, ZN => DIFF_60_port);
   U65 : NOR2_X1 port map( A1 => B(59), A2 => n198, ZN => n199);
   U66 : NOR2_X1 port map( A1 => B(51), A2 => n206, ZN => n207);
   U67 : XNOR2_X1 port map( A => B(56), B => n203, ZN => DIFF_56_port);
   U68 : NOR2_X1 port map( A1 => B(55), A2 => n202, ZN => n203);
   U69 : OR3_X1 port map( A1 => B(51), A2 => B(52), A3 => n206, ZN => n204);
   U70 : OR3_X1 port map( A1 => B(55), A2 => B(56), A3 => n202, ZN => n200);
   U71 : OR2_X1 port map( A1 => n196, A2 => B(62), ZN => n195);
   U72 : XNOR2_X1 port map( A => n189, B => B(6), ZN => DIFF_6_port);
   U73 : NOR2_X1 port map( A1 => n194, A2 => B(5), ZN => n189);
   U74 : OR3_X1 port map( A1 => B(5), A2 => B(6), A3 => n194, ZN => n192);
   U75 : NOR2_X1 port map( A1 => B(3), A2 => n211, ZN => n210);
   U76 : OR3_X1 port map( A1 => B(3), A2 => B(4), A3 => n211, ZN => n194);
   U77 : XNOR2_X1 port map( A => B(4), B => n210, ZN => DIFF_4_port);
   U78 : XNOR2_X1 port map( A => B(2), B => n232, ZN => DIFF_2_port);
   U79 : OR3_X1 port map( A1 => B(1), A2 => B(2), A3 => B(0), ZN => n211);
   U80 : NOR2_X1 port map( A1 => B(0), A2 => B(1), ZN => n232);
   U83 : INV_X1 port map( A => B(61), ZN => n193);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_27_DW01_sub_0 is

   port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (63 downto 0);  CO : out std_logic);

end complementer_N64_27_DW01_sub_0;

architecture SYN_rpl of complementer_N64_27_DW01_sub_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal DIFF_62_port, DIFF_63_port, DIFF_5_port, DIFF_6_port, DIFF_7_port, 
      DIFF_8_port, DIFF_9_port, DIFF_10_port, DIFF_11_port, DIFF_12_port, 
      DIFF_13_port, DIFF_14_port, DIFF_15_port, DIFF_16_port, DIFF_17_port, 
      DIFF_18_port, DIFF_19_port, DIFF_20_port, DIFF_21_port, DIFF_22_port, 
      DIFF_23_port, DIFF_24_port, DIFF_25_port, DIFF_26_port, DIFF_27_port, 
      DIFF_28_port, DIFF_29_port, DIFF_30_port, DIFF_31_port, DIFF_32_port, 
      DIFF_33_port, DIFF_34_port, DIFF_35_port, DIFF_36_port, DIFF_37_port, 
      DIFF_38_port, DIFF_39_port, DIFF_40_port, DIFF_41_port, DIFF_42_port, 
      DIFF_43_port, DIFF_44_port, DIFF_45_port, DIFF_46_port, DIFF_47_port, 
      DIFF_48_port, DIFF_49_port, DIFF_50_port, DIFF_51_port, DIFF_52_port, 
      DIFF_53_port, DIFF_54_port, DIFF_55_port, DIFF_56_port, DIFF_57_port, 
      DIFF_58_port, DIFF_59_port, DIFF_60_port, DIFF_61_port, DIFF_3_port, 
      DIFF_4_port, DIFF_2_port, DIFF_1_port, n190, n191, n192, n193, n194, n195
      , n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
      n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, 
      n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, 
      n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, 
      n244, n245, n246, n247, n248, n249, n250, n251, n189 : std_logic;

begin
   DIFF <= ( DIFF_63_port, DIFF_62_port, DIFF_61_port, DIFF_60_port, 
      DIFF_59_port, DIFF_58_port, DIFF_57_port, DIFF_56_port, DIFF_55_port, 
      DIFF_54_port, DIFF_53_port, DIFF_52_port, DIFF_51_port, DIFF_50_port, 
      DIFF_49_port, DIFF_48_port, DIFF_47_port, DIFF_46_port, DIFF_45_port, 
      DIFF_44_port, DIFF_43_port, DIFF_42_port, DIFF_41_port, DIFF_40_port, 
      DIFF_39_port, DIFF_38_port, DIFF_37_port, DIFF_36_port, DIFF_35_port, 
      DIFF_34_port, DIFF_33_port, DIFF_32_port, DIFF_31_port, DIFF_30_port, 
      DIFF_29_port, DIFF_28_port, DIFF_27_port, DIFF_26_port, DIFF_25_port, 
      DIFF_24_port, DIFF_23_port, DIFF_22_port, DIFF_21_port, DIFF_20_port, 
      DIFF_19_port, DIFF_18_port, DIFF_17_port, DIFF_16_port, DIFF_15_port, 
      DIFF_14_port, DIFF_13_port, DIFF_12_port, DIFF_11_port, DIFF_10_port, 
      DIFF_9_port, DIFF_8_port, DIFF_7_port, DIFF_6_port, DIFF_5_port, 
      DIFF_4_port, DIFF_3_port, DIFF_2_port, DIFF_1_port, B(0) );
   
   U81 : XOR2_X1 port map( A => n190, B => B(9), Z => DIFF_9_port);
   U82 : XOR2_X1 port map( A => n192, B => B(7), Z => DIFF_7_port);
   U83 : XOR2_X1 port map( A => n193, B => B(6), Z => DIFF_6_port);
   U84 : XOR2_X1 port map( A => n195, B => B(63), Z => DIFF_63_port);
   U85 : XOR2_X1 port map( A => n196, B => B(62), Z => DIFF_62_port);
   U86 : XOR2_X1 port map( A => n194, B => B(5), Z => DIFF_5_port);
   U87 : XOR2_X1 port map( A => n198, B => B(59), Z => DIFF_59_port);
   U88 : XOR2_X1 port map( A => n201, B => B(58), Z => DIFF_58_port);
   U89 : XOR2_X1 port map( A => n200, B => B(57), Z => DIFF_57_port);
   U90 : XOR2_X1 port map( A => n202, B => B(55), Z => DIFF_55_port);
   U91 : XOR2_X1 port map( A => n205, B => B(54), Z => DIFF_54_port);
   U92 : XOR2_X1 port map( A => n204, B => B(53), Z => DIFF_53_port);
   U93 : XOR2_X1 port map( A => n206, B => B(51), Z => DIFF_51_port);
   U94 : XOR2_X1 port map( A => n209, B => B(50), Z => DIFF_50_port);
   U95 : XOR2_X1 port map( A => n208, B => B(49), Z => DIFF_49_port);
   U96 : XOR2_X1 port map( A => n212, B => B(47), Z => DIFF_47_port);
   U97 : XOR2_X1 port map( A => n215, B => B(46), Z => DIFF_46_port);
   U98 : XOR2_X1 port map( A => n214, B => B(45), Z => DIFF_45_port);
   U99 : XOR2_X1 port map( A => n216, B => B(43), Z => DIFF_43_port);
   U100 : XOR2_X1 port map( A => n219, B => B(42), Z => DIFF_42_port);
   U101 : XOR2_X1 port map( A => n218, B => B(41), Z => DIFF_41_port);
   U102 : XOR2_X1 port map( A => n211, B => B(3), Z => DIFF_3_port);
   U103 : XOR2_X1 port map( A => n220, B => B(39), Z => DIFF_39_port);
   U104 : XOR2_X1 port map( A => n223, B => B(38), Z => DIFF_38_port);
   U105 : XOR2_X1 port map( A => n222, B => B(37), Z => DIFF_37_port);
   U106 : XOR2_X1 port map( A => n224, B => B(35), Z => DIFF_35_port);
   U107 : XOR2_X1 port map( A => n227, B => B(34), Z => DIFF_34_port);
   U108 : XOR2_X1 port map( A => n226, B => B(33), Z => DIFF_33_port);
   U109 : XOR2_X1 port map( A => n228, B => B(31), Z => DIFF_31_port);
   U110 : XOR2_X1 port map( A => n231, B => B(30), Z => DIFF_30_port);
   U111 : XOR2_X1 port map( A => n230, B => B(29), Z => DIFF_29_port);
   U112 : XOR2_X1 port map( A => n233, B => B(27), Z => DIFF_27_port);
   U113 : XOR2_X1 port map( A => n236, B => B(26), Z => DIFF_26_port);
   U114 : XOR2_X1 port map( A => n235, B => B(25), Z => DIFF_25_port);
   U115 : XOR2_X1 port map( A => n237, B => B(23), Z => DIFF_23_port);
   U116 : XOR2_X1 port map( A => n240, B => B(22), Z => DIFF_22_port);
   U117 : XOR2_X1 port map( A => n239, B => B(21), Z => DIFF_21_port);
   U118 : XOR2_X1 port map( A => B(1), B => B(0), Z => DIFF_1_port);
   U119 : XOR2_X1 port map( A => n241, B => B(19), Z => DIFF_19_port);
   U120 : XOR2_X1 port map( A => n244, B => B(18), Z => DIFF_18_port);
   U121 : XOR2_X1 port map( A => n243, B => B(17), Z => DIFF_17_port);
   U122 : XOR2_X1 port map( A => n245, B => B(15), Z => DIFF_15_port);
   U123 : XOR2_X1 port map( A => n248, B => B(14), Z => DIFF_14_port);
   U124 : XOR2_X1 port map( A => n247, B => B(13), Z => DIFF_13_port);
   U125 : XOR2_X1 port map( A => n249, B => B(11), Z => DIFF_11_port);
   U126 : XOR2_X1 port map( A => n251, B => B(10), Z => DIFF_10_port);
   U1 : NOR2_X1 port map( A1 => B(43), A2 => n216, ZN => n217);
   U2 : OR2_X1 port map( A1 => n204, A2 => B(53), ZN => n205);
   U3 : NAND2_X1 port map( A1 => n197, A2 => n189, ZN => n196);
   U4 : NOR2_X1 port map( A1 => B(47), A2 => n212, ZN => n213);
   U5 : NOR2_X1 port map( A1 => B(35), A2 => n224, ZN => n225);
   U6 : NOR2_X1 port map( A1 => B(7), A2 => n192, ZN => n191);
   U7 : NOR2_X1 port map( A1 => B(11), A2 => n249, ZN => n250);
   U8 : NOR2_X1 port map( A1 => B(15), A2 => n245, ZN => n246);
   U9 : NOR2_X1 port map( A1 => B(19), A2 => n241, ZN => n242);
   U10 : NOR2_X1 port map( A1 => B(31), A2 => n228, ZN => n229);
   U11 : NOR2_X1 port map( A1 => B(23), A2 => n237, ZN => n238);
   U12 : NOR2_X1 port map( A1 => B(27), A2 => n233, ZN => n234);
   U13 : NOR2_X1 port map( A1 => B(51), A2 => n206, ZN => n207);
   U14 : NOR2_X1 port map( A1 => B(39), A2 => n220, ZN => n221);
   U15 : NOR2_X1 port map( A1 => B(55), A2 => n202, ZN => n203);
   U16 : OR3_X1 port map( A1 => B(10), A2 => B(9), A3 => n190, ZN => n249);
   U17 : OR3_X1 port map( A1 => B(45), A2 => B(46), A3 => n214, ZN => n212);
   U18 : OR3_X1 port map( A1 => B(5), A2 => B(6), A3 => n194, ZN => n192);
   U19 : OR3_X1 port map( A1 => B(25), A2 => B(26), A3 => n235, ZN => n233);
   U20 : OR3_X1 port map( A1 => B(13), A2 => B(14), A3 => n247, ZN => n245);
   U21 : OR3_X1 port map( A1 => B(29), A2 => B(30), A3 => n230, ZN => n228);
   U22 : OR3_X1 port map( A1 => B(17), A2 => B(18), A3 => n243, ZN => n241);
   U23 : OR3_X1 port map( A1 => B(21), A2 => B(22), A3 => n239, ZN => n237);
   U24 : OR3_X1 port map( A1 => B(49), A2 => B(50), A3 => n208, ZN => n206);
   U25 : OR3_X1 port map( A1 => B(33), A2 => B(34), A3 => n226, ZN => n224);
   U26 : OR3_X1 port map( A1 => B(37), A2 => B(38), A3 => n222, ZN => n220);
   U27 : OR3_X1 port map( A1 => B(53), A2 => B(54), A3 => n204, ZN => n202);
   U28 : OR3_X1 port map( A1 => B(41), A2 => B(42), A3 => n218, ZN => n216);
   U29 : OR3_X1 port map( A1 => B(43), A2 => B(44), A3 => n216, ZN => n214);
   U30 : OR3_X1 port map( A1 => B(47), A2 => B(48), A3 => n212, ZN => n208);
   U31 : OR3_X1 port map( A1 => B(35), A2 => B(36), A3 => n224, ZN => n222);
   U32 : OR3_X1 port map( A1 => B(7), A2 => B(8), A3 => n192, ZN => n190);
   U33 : OR3_X1 port map( A1 => B(11), A2 => B(12), A3 => n249, ZN => n247);
   U34 : OR3_X1 port map( A1 => B(27), A2 => B(28), A3 => n233, ZN => n230);
   U35 : OR3_X1 port map( A1 => B(15), A2 => B(16), A3 => n245, ZN => n243);
   U36 : OR3_X1 port map( A1 => B(23), A2 => B(24), A3 => n237, ZN => n235);
   U37 : OR3_X1 port map( A1 => B(19), A2 => B(20), A3 => n241, ZN => n239);
   U38 : OR3_X1 port map( A1 => B(31), A2 => B(32), A3 => n228, ZN => n226);
   U39 : OR3_X1 port map( A1 => B(39), A2 => B(40), A3 => n220, ZN => n218);
   U40 : OR3_X1 port map( A1 => B(51), A2 => B(52), A3 => n206, ZN => n204);
   U41 : XNOR2_X1 port map( A => B(48), B => n213, ZN => DIFF_48_port);
   U42 : XNOR2_X1 port map( A => B(8), B => n191, ZN => DIFF_8_port);
   U43 : XNOR2_X1 port map( A => B(12), B => n250, ZN => DIFF_12_port);
   U44 : XNOR2_X1 port map( A => B(16), B => n246, ZN => DIFF_16_port);
   U45 : XNOR2_X1 port map( A => B(20), B => n242, ZN => DIFF_20_port);
   U46 : XNOR2_X1 port map( A => B(24), B => n238, ZN => DIFF_24_port);
   U47 : XNOR2_X1 port map( A => B(28), B => n234, ZN => DIFF_28_port);
   U48 : XNOR2_X1 port map( A => B(32), B => n229, ZN => DIFF_32_port);
   U49 : XNOR2_X1 port map( A => B(40), B => n221, ZN => DIFF_40_port);
   U50 : XNOR2_X1 port map( A => B(52), B => n207, ZN => DIFF_52_port);
   U51 : XNOR2_X1 port map( A => B(36), B => n225, ZN => DIFF_36_port);
   U52 : XNOR2_X1 port map( A => B(56), B => n203, ZN => DIFF_56_port);
   U53 : XNOR2_X1 port map( A => B(44), B => n217, ZN => DIFF_44_port);
   U54 : OR2_X1 port map( A1 => n214, A2 => B(45), ZN => n215);
   U55 : OR2_X1 port map( A1 => n222, A2 => B(37), ZN => n223);
   U56 : OR2_X1 port map( A1 => n194, A2 => B(5), ZN => n193);
   U57 : OR2_X1 port map( A1 => n208, A2 => B(49), ZN => n209);
   U58 : OR2_X1 port map( A1 => n190, A2 => B(9), ZN => n251);
   U59 : OR2_X1 port map( A1 => n247, A2 => B(13), ZN => n248);
   U60 : OR2_X1 port map( A1 => n243, A2 => B(17), ZN => n244);
   U61 : OR2_X1 port map( A1 => n226, A2 => B(33), ZN => n227);
   U62 : OR2_X1 port map( A1 => n230, A2 => B(29), ZN => n231);
   U63 : OR2_X1 port map( A1 => n239, A2 => B(21), ZN => n240);
   U64 : OR2_X1 port map( A1 => n235, A2 => B(25), ZN => n236);
   U65 : OR2_X1 port map( A1 => n218, A2 => B(41), ZN => n219);
   U66 : NOR3_X1 port map( A1 => B(59), A2 => B(60), A3 => n198, ZN => n197);
   U67 : XNOR2_X1 port map( A => n197, B => B(61), ZN => DIFF_61_port);
   U68 : XNOR2_X1 port map( A => B(60), B => n199, ZN => DIFF_60_port);
   U69 : NOR2_X1 port map( A1 => B(59), A2 => n198, ZN => n199);
   U70 : OR3_X1 port map( A1 => B(57), A2 => B(58), A3 => n200, ZN => n198);
   U71 : OR3_X1 port map( A1 => B(55), A2 => B(56), A3 => n202, ZN => n200);
   U72 : OR2_X1 port map( A1 => n196, A2 => B(62), ZN => n195);
   U73 : OR2_X1 port map( A1 => n200, A2 => B(57), ZN => n201);
   U74 : XNOR2_X1 port map( A => B(4), B => n210, ZN => DIFF_4_port);
   U75 : NOR2_X1 port map( A1 => B(3), A2 => n211, ZN => n210);
   U76 : XNOR2_X1 port map( A => B(2), B => n232, ZN => DIFF_2_port);
   U77 : NOR2_X1 port map( A1 => B(0), A2 => B(1), ZN => n232);
   U78 : OR3_X1 port map( A1 => B(3), A2 => B(4), A3 => n211, ZN => n194);
   U79 : OR3_X1 port map( A1 => B(1), A2 => B(2), A3 => B(0), ZN => n211);
   U80 : INV_X1 port map( A => B(61), ZN => n189);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_28_DW01_sub_0 is

   port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (63 downto 0);  CO : out std_logic);

end complementer_N64_28_DW01_sub_0;

architecture SYN_rpl of complementer_N64_28_DW01_sub_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal DIFF_62_port, DIFF_61_port, DIFF_60_port, DIFF_59_port, DIFF_58_port,
      DIFF_57_port, DIFF_56_port, DIFF_55_port, DIFF_54_port, DIFF_53_port, 
      DIFF_52_port, DIFF_51_port, DIFF_50_port, DIFF_49_port, DIFF_48_port, 
      DIFF_47_port, DIFF_46_port, DIFF_45_port, DIFF_44_port, DIFF_43_port, 
      DIFF_42_port, DIFF_41_port, DIFF_40_port, DIFF_39_port, DIFF_38_port, 
      DIFF_37_port, DIFF_36_port, DIFF_35_port, DIFF_34_port, DIFF_33_port, 
      DIFF_32_port, DIFF_31_port, DIFF_30_port, DIFF_29_port, DIFF_28_port, 
      DIFF_27_port, DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, 
      DIFF_22_port, DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, 
      DIFF_17_port, DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, 
      DIFF_12_port, DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, 
      DIFF_7_port, DIFF_6_port, DIFF_5_port, DIFF_4_port, DIFF_3_port, 
      DIFF_2_port, DIFF_1_port, DIFF_63_port, n190, n191, n192, n194, n196, 
      n197, n198, n199, n200, n202, n203, n204, n206, n207, n208, n210, n211, 
      n212, n213, n214, n216, n217, n218, n220, n221, n222, n224, n225, n226, 
      n228, n229, n230, n232, n233, n234, n235, n237, n238, n239, n241, n242, 
      n243, n245, n246, n247, n249, n250, n189, n193, n195, n201, n205, n209, 
      n215, n219, n223, n227, n231, n236, n240, n244, n248, n251 : std_logic;

begin
   DIFF <= ( DIFF_63_port, DIFF_62_port, DIFF_61_port, DIFF_60_port, 
      DIFF_59_port, DIFF_58_port, DIFF_57_port, DIFF_56_port, DIFF_55_port, 
      DIFF_54_port, DIFF_53_port, DIFF_52_port, DIFF_51_port, DIFF_50_port, 
      DIFF_49_port, DIFF_48_port, DIFF_47_port, DIFF_46_port, DIFF_45_port, 
      DIFF_44_port, DIFF_43_port, DIFF_42_port, DIFF_41_port, DIFF_40_port, 
      DIFF_39_port, DIFF_38_port, DIFF_37_port, DIFF_36_port, DIFF_35_port, 
      DIFF_34_port, DIFF_33_port, DIFF_32_port, DIFF_31_port, DIFF_30_port, 
      DIFF_29_port, DIFF_28_port, DIFF_27_port, DIFF_26_port, DIFF_25_port, 
      DIFF_24_port, DIFF_23_port, DIFF_22_port, DIFF_21_port, DIFF_20_port, 
      DIFF_19_port, DIFF_18_port, DIFF_17_port, DIFF_16_port, DIFF_15_port, 
      DIFF_14_port, DIFF_13_port, DIFF_12_port, DIFF_11_port, DIFF_10_port, 
      DIFF_9_port, DIFF_8_port, DIFF_7_port, DIFF_6_port, DIFF_5_port, 
      DIFF_4_port, DIFF_3_port, DIFF_2_port, DIFF_1_port, B(0) );
   
   U81 : XOR2_X1 port map( A => n190, B => B(9), Z => DIFF_9_port);
   U82 : XOR2_X1 port map( A => n192, B => B(7), Z => DIFF_7_port);
   U85 : XOR2_X1 port map( A => n196, B => B(62), Z => DIFF_62_port);
   U86 : XOR2_X1 port map( A => n194, B => B(5), Z => DIFF_5_port);
   U87 : XOR2_X1 port map( A => n198, B => B(59), Z => DIFF_59_port);
   U89 : XOR2_X1 port map( A => n200, B => B(57), Z => DIFF_57_port);
   U90 : XOR2_X1 port map( A => n202, B => B(55), Z => DIFF_55_port);
   U92 : XOR2_X1 port map( A => n204, B => B(53), Z => DIFF_53_port);
   U93 : XOR2_X1 port map( A => n206, B => B(51), Z => DIFF_51_port);
   U95 : XOR2_X1 port map( A => n208, B => B(49), Z => DIFF_49_port);
   U96 : XOR2_X1 port map( A => n212, B => B(47), Z => DIFF_47_port);
   U98 : XOR2_X1 port map( A => n214, B => B(45), Z => DIFF_45_port);
   U99 : XOR2_X1 port map( A => n216, B => B(43), Z => DIFF_43_port);
   U101 : XOR2_X1 port map( A => n218, B => B(41), Z => DIFF_41_port);
   U102 : XOR2_X1 port map( A => n211, B => B(3), Z => DIFF_3_port);
   U103 : XOR2_X1 port map( A => n220, B => B(39), Z => DIFF_39_port);
   U105 : XOR2_X1 port map( A => n222, B => B(37), Z => DIFF_37_port);
   U106 : XOR2_X1 port map( A => n224, B => B(35), Z => DIFF_35_port);
   U108 : XOR2_X1 port map( A => n226, B => B(33), Z => DIFF_33_port);
   U109 : XOR2_X1 port map( A => n228, B => B(31), Z => DIFF_31_port);
   U111 : XOR2_X1 port map( A => n230, B => B(29), Z => DIFF_29_port);
   U112 : XOR2_X1 port map( A => n233, B => B(27), Z => DIFF_27_port);
   U114 : XOR2_X1 port map( A => n235, B => B(25), Z => DIFF_25_port);
   U115 : XOR2_X1 port map( A => n237, B => B(23), Z => DIFF_23_port);
   U117 : XOR2_X1 port map( A => n239, B => B(21), Z => DIFF_21_port);
   U118 : XOR2_X1 port map( A => B(1), B => B(0), Z => DIFF_1_port);
   U119 : XOR2_X1 port map( A => n241, B => B(19), Z => DIFF_19_port);
   U121 : XOR2_X1 port map( A => n243, B => B(17), Z => DIFF_17_port);
   U122 : XOR2_X1 port map( A => n245, B => B(15), Z => DIFF_15_port);
   U124 : XOR2_X1 port map( A => n247, B => B(13), Z => DIFF_13_port);
   U125 : XOR2_X1 port map( A => n249, B => B(11), Z => DIFF_11_port);
   U1 : XOR2_X1 port map( A => n197, B => n251, Z => DIFF_61_port);
   U2 : NAND2_X1 port map( A1 => n197, A2 => n251, ZN => n196);
   U3 : XNOR2_X1 port map( A => n189, B => B(34), ZN => DIFF_34_port);
   U4 : NOR2_X1 port map( A1 => n226, A2 => B(33), ZN => n189);
   U5 : XNOR2_X1 port map( A => n193, B => B(46), ZN => DIFF_46_port);
   U6 : NOR2_X1 port map( A1 => n214, A2 => B(45), ZN => n193);
   U7 : XNOR2_X1 port map( A => n195, B => B(6), ZN => DIFF_6_port);
   U8 : NOR2_X1 port map( A1 => n194, A2 => B(5), ZN => n195);
   U9 : XNOR2_X1 port map( A => n201, B => B(10), ZN => DIFF_10_port);
   U10 : NOR2_X1 port map( A1 => n190, A2 => B(9), ZN => n201);
   U11 : XNOR2_X1 port map( A => n205, B => B(14), ZN => DIFF_14_port);
   U12 : NOR2_X1 port map( A1 => n247, A2 => B(13), ZN => n205);
   U13 : XNOR2_X1 port map( A => n209, B => B(18), ZN => DIFF_18_port);
   U14 : NOR2_X1 port map( A1 => n243, A2 => B(17), ZN => n209);
   U15 : XNOR2_X1 port map( A => n215, B => B(26), ZN => DIFF_26_port);
   U16 : NOR2_X1 port map( A1 => n235, A2 => B(25), ZN => n215);
   U17 : XNOR2_X1 port map( A => n219, B => B(30), ZN => DIFF_30_port);
   U18 : NOR2_X1 port map( A1 => n230, A2 => B(29), ZN => n219);
   U19 : XNOR2_X1 port map( A => n223, B => B(50), ZN => DIFF_50_port);
   U20 : NOR2_X1 port map( A1 => n208, A2 => B(49), ZN => n223);
   U21 : XNOR2_X1 port map( A => n227, B => B(42), ZN => DIFF_42_port);
   U22 : NOR2_X1 port map( A1 => n218, A2 => B(41), ZN => n227);
   U23 : XNOR2_X1 port map( A => n231, B => B(38), ZN => DIFF_38_port);
   U24 : NOR2_X1 port map( A1 => n222, A2 => B(37), ZN => n231);
   U25 : XNOR2_X1 port map( A => n236, B => B(58), ZN => DIFF_58_port);
   U26 : NOR2_X1 port map( A1 => n200, A2 => B(57), ZN => n236);
   U27 : XNOR2_X1 port map( A => n240, B => B(54), ZN => DIFF_54_port);
   U28 : NOR2_X1 port map( A1 => n204, A2 => B(53), ZN => n240);
   U29 : XNOR2_X1 port map( A => B(20), B => n242, ZN => DIFF_20_port);
   U30 : NOR2_X1 port map( A1 => B(19), A2 => n241, ZN => n242);
   U31 : XNOR2_X1 port map( A => B(24), B => n238, ZN => DIFF_24_port);
   U32 : NOR2_X1 port map( A1 => B(23), A2 => n237, ZN => n238);
   U33 : XNOR2_X1 port map( A => B(36), B => n225, ZN => DIFF_36_port);
   U34 : NOR2_X1 port map( A1 => B(35), A2 => n224, ZN => n225);
   U35 : XNOR2_X1 port map( A => B(44), B => n217, ZN => DIFF_44_port);
   U36 : NOR2_X1 port map( A1 => B(43), A2 => n216, ZN => n217);
   U37 : XNOR2_X1 port map( A => B(52), B => n207, ZN => DIFF_52_port);
   U38 : NOR2_X1 port map( A1 => B(51), A2 => n206, ZN => n207);
   U39 : XNOR2_X1 port map( A => B(48), B => n213, ZN => DIFF_48_port);
   U40 : NOR2_X1 port map( A1 => B(47), A2 => n212, ZN => n213);
   U41 : XNOR2_X1 port map( A => B(8), B => n191, ZN => DIFF_8_port);
   U42 : NOR2_X1 port map( A1 => B(7), A2 => n192, ZN => n191);
   U43 : XNOR2_X1 port map( A => B(12), B => n250, ZN => DIFF_12_port);
   U44 : NOR2_X1 port map( A1 => B(11), A2 => n249, ZN => n250);
   U45 : XNOR2_X1 port map( A => B(16), B => n246, ZN => DIFF_16_port);
   U46 : NOR2_X1 port map( A1 => B(15), A2 => n245, ZN => n246);
   U47 : XNOR2_X1 port map( A => B(28), B => n234, ZN => DIFF_28_port);
   U48 : NOR2_X1 port map( A1 => B(27), A2 => n233, ZN => n234);
   U49 : XNOR2_X1 port map( A => B(32), B => n229, ZN => DIFF_32_port);
   U50 : NOR2_X1 port map( A1 => B(31), A2 => n228, ZN => n229);
   U51 : XNOR2_X1 port map( A => B(40), B => n221, ZN => DIFF_40_port);
   U52 : NOR2_X1 port map( A1 => B(39), A2 => n220, ZN => n221);
   U53 : XNOR2_X1 port map( A => B(56), B => n203, ZN => DIFF_56_port);
   U54 : NOR2_X1 port map( A1 => B(55), A2 => n202, ZN => n203);
   U55 : OR3_X1 port map( A1 => B(57), A2 => B(58), A3 => n200, ZN => n198);
   U56 : OR3_X1 port map( A1 => B(25), A2 => B(26), A3 => n235, ZN => n233);
   U57 : OR3_X1 port map( A1 => B(5), A2 => B(6), A3 => n194, ZN => n192);
   U58 : OR3_X1 port map( A1 => B(13), A2 => B(14), A3 => n247, ZN => n245);
   U59 : OR3_X1 port map( A1 => B(17), A2 => B(18), A3 => n243, ZN => n241);
   U60 : OR3_X1 port map( A1 => B(29), A2 => B(30), A3 => n230, ZN => n228);
   U61 : OR3_X1 port map( A1 => B(21), A2 => B(22), A3 => n239, ZN => n237);
   U62 : OR3_X1 port map( A1 => B(33), A2 => B(34), A3 => n226, ZN => n224);
   U63 : OR3_X1 port map( A1 => B(49), A2 => B(50), A3 => n208, ZN => n206);
   U64 : OR3_X1 port map( A1 => B(10), A2 => B(9), A3 => n190, ZN => n249);
   U65 : OR3_X1 port map( A1 => B(45), A2 => B(46), A3 => n214, ZN => n212);
   U66 : OR3_X1 port map( A1 => B(37), A2 => B(38), A3 => n222, ZN => n220);
   U67 : OR3_X1 port map( A1 => B(41), A2 => B(42), A3 => n218, ZN => n216);
   U68 : OR3_X1 port map( A1 => B(53), A2 => B(54), A3 => n204, ZN => n202);
   U69 : OR3_X1 port map( A1 => B(47), A2 => B(48), A3 => n212, ZN => n208);
   U70 : OR3_X1 port map( A1 => B(51), A2 => B(52), A3 => n206, ZN => n204);
   U71 : OR3_X1 port map( A1 => B(43), A2 => B(44), A3 => n216, ZN => n214);
   U72 : OR3_X1 port map( A1 => B(23), A2 => B(24), A3 => n237, ZN => n235);
   U73 : OR3_X1 port map( A1 => B(7), A2 => B(8), A3 => n192, ZN => n190);
   U74 : OR3_X1 port map( A1 => B(15), A2 => B(16), A3 => n245, ZN => n243);
   U75 : OR3_X1 port map( A1 => B(11), A2 => B(12), A3 => n249, ZN => n247);
   U76 : OR3_X1 port map( A1 => B(27), A2 => B(28), A3 => n233, ZN => n230);
   U77 : OR3_X1 port map( A1 => B(31), A2 => B(32), A3 => n228, ZN => n226);
   U78 : OR3_X1 port map( A1 => B(19), A2 => B(20), A3 => n241, ZN => n239);
   U79 : OR3_X1 port map( A1 => B(39), A2 => B(40), A3 => n220, ZN => n218);
   U80 : OR3_X1 port map( A1 => B(35), A2 => B(36), A3 => n224, ZN => n222);
   U83 : OR3_X1 port map( A1 => B(55), A2 => B(56), A3 => n202, ZN => n200);
   U84 : XNOR2_X1 port map( A => n244, B => B(22), ZN => DIFF_22_port);
   U88 : NOR2_X1 port map( A1 => n239, A2 => B(21), ZN => n244);
   U91 : NOR3_X1 port map( A1 => B(59), A2 => B(60), A3 => n198, ZN => n197);
   U94 : XNOR2_X1 port map( A => B(60), B => n199, ZN => DIFF_60_port);
   U97 : NOR2_X1 port map( A1 => B(59), A2 => n198, ZN => n199);
   U100 : OR3_X1 port map( A1 => B(3), A2 => B(4), A3 => n211, ZN => n194);
   U104 : XNOR2_X1 port map( A => B(4), B => n210, ZN => DIFF_4_port);
   U107 : NOR2_X1 port map( A1 => B(3), A2 => n211, ZN => n210);
   U110 : XNOR2_X1 port map( A => n248, B => B(63), ZN => DIFF_63_port);
   U113 : NOR2_X1 port map( A1 => n196, A2 => B(62), ZN => n248);
   U116 : XNOR2_X1 port map( A => B(2), B => n232, ZN => DIFF_2_port);
   U120 : OR3_X1 port map( A1 => B(1), A2 => B(2), A3 => B(0), ZN => n211);
   U123 : NOR2_X1 port map( A1 => B(0), A2 => B(1), ZN => n232);
   U126 : INV_X1 port map( A => B(61), ZN => n251);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_29_DW01_sub_0 is

   port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (63 downto 0);  CO : out std_logic);

end complementer_N64_29_DW01_sub_0;

architecture SYN_rpl of complementer_N64_29_DW01_sub_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal DIFF_62_port, DIFF_63_port, DIFF_3_port, DIFF_4_port, DIFF_5_port, 
      DIFF_6_port, DIFF_7_port, DIFF_8_port, DIFF_9_port, DIFF_10_port, 
      DIFF_11_port, DIFF_12_port, DIFF_13_port, DIFF_14_port, DIFF_15_port, 
      DIFF_16_port, DIFF_17_port, DIFF_18_port, DIFF_19_port, DIFF_20_port, 
      DIFF_21_port, DIFF_22_port, DIFF_23_port, DIFF_24_port, DIFF_25_port, 
      DIFF_26_port, DIFF_27_port, DIFF_28_port, DIFF_29_port, DIFF_30_port, 
      DIFF_31_port, DIFF_32_port, DIFF_33_port, DIFF_34_port, DIFF_35_port, 
      DIFF_36_port, DIFF_37_port, DIFF_38_port, DIFF_39_port, DIFF_40_port, 
      DIFF_41_port, DIFF_42_port, DIFF_43_port, DIFF_44_port, DIFF_45_port, 
      DIFF_46_port, DIFF_47_port, DIFF_48_port, DIFF_49_port, DIFF_50_port, 
      DIFF_51_port, DIFF_52_port, DIFF_53_port, DIFF_54_port, DIFF_55_port, 
      DIFF_56_port, DIFF_57_port, DIFF_58_port, DIFF_59_port, DIFF_60_port, 
      DIFF_61_port, DIFF_2_port, DIFF_1_port, n190, n191, n192, n194, n195, 
      n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, 
      n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, 
      n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, 
      n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, 
      n244, n245, n246, n247, n248, n249, n250, n251, n189, n193 : std_logic;

begin
   DIFF <= ( DIFF_63_port, DIFF_62_port, DIFF_61_port, DIFF_60_port, 
      DIFF_59_port, DIFF_58_port, DIFF_57_port, DIFF_56_port, DIFF_55_port, 
      DIFF_54_port, DIFF_53_port, DIFF_52_port, DIFF_51_port, DIFF_50_port, 
      DIFF_49_port, DIFF_48_port, DIFF_47_port, DIFF_46_port, DIFF_45_port, 
      DIFF_44_port, DIFF_43_port, DIFF_42_port, DIFF_41_port, DIFF_40_port, 
      DIFF_39_port, DIFF_38_port, DIFF_37_port, DIFF_36_port, DIFF_35_port, 
      DIFF_34_port, DIFF_33_port, DIFF_32_port, DIFF_31_port, DIFF_30_port, 
      DIFF_29_port, DIFF_28_port, DIFF_27_port, DIFF_26_port, DIFF_25_port, 
      DIFF_24_port, DIFF_23_port, DIFF_22_port, DIFF_21_port, DIFF_20_port, 
      DIFF_19_port, DIFF_18_port, DIFF_17_port, DIFF_16_port, DIFF_15_port, 
      DIFF_14_port, DIFF_13_port, DIFF_12_port, DIFF_11_port, DIFF_10_port, 
      DIFF_9_port, DIFF_8_port, DIFF_7_port, DIFF_6_port, DIFF_5_port, 
      DIFF_4_port, DIFF_3_port, DIFF_2_port, DIFF_1_port, B(0) );
   
   U81 : XOR2_X1 port map( A => n190, B => B(9), Z => DIFF_9_port);
   U82 : XOR2_X1 port map( A => n192, B => B(7), Z => DIFF_7_port);
   U84 : XOR2_X1 port map( A => n195, B => B(63), Z => DIFF_63_port);
   U85 : XOR2_X1 port map( A => n196, B => B(62), Z => DIFF_62_port);
   U86 : XOR2_X1 port map( A => n194, B => B(5), Z => DIFF_5_port);
   U87 : XOR2_X1 port map( A => n198, B => B(59), Z => DIFF_59_port);
   U88 : XOR2_X1 port map( A => n201, B => B(58), Z => DIFF_58_port);
   U89 : XOR2_X1 port map( A => n200, B => B(57), Z => DIFF_57_port);
   U90 : XOR2_X1 port map( A => n202, B => B(55), Z => DIFF_55_port);
   U91 : XOR2_X1 port map( A => n205, B => B(54), Z => DIFF_54_port);
   U92 : XOR2_X1 port map( A => n204, B => B(53), Z => DIFF_53_port);
   U93 : XOR2_X1 port map( A => n206, B => B(51), Z => DIFF_51_port);
   U94 : XOR2_X1 port map( A => n209, B => B(50), Z => DIFF_50_port);
   U95 : XOR2_X1 port map( A => n208, B => B(49), Z => DIFF_49_port);
   U96 : XOR2_X1 port map( A => n212, B => B(47), Z => DIFF_47_port);
   U97 : XOR2_X1 port map( A => n215, B => B(46), Z => DIFF_46_port);
   U98 : XOR2_X1 port map( A => n214, B => B(45), Z => DIFF_45_port);
   U99 : XOR2_X1 port map( A => n216, B => B(43), Z => DIFF_43_port);
   U100 : XOR2_X1 port map( A => n219, B => B(42), Z => DIFF_42_port);
   U101 : XOR2_X1 port map( A => n218, B => B(41), Z => DIFF_41_port);
   U102 : XOR2_X1 port map( A => n211, B => B(3), Z => DIFF_3_port);
   U103 : XOR2_X1 port map( A => n220, B => B(39), Z => DIFF_39_port);
   U104 : XOR2_X1 port map( A => n223, B => B(38), Z => DIFF_38_port);
   U105 : XOR2_X1 port map( A => n222, B => B(37), Z => DIFF_37_port);
   U106 : XOR2_X1 port map( A => n224, B => B(35), Z => DIFF_35_port);
   U107 : XOR2_X1 port map( A => n227, B => B(34), Z => DIFF_34_port);
   U108 : XOR2_X1 port map( A => n226, B => B(33), Z => DIFF_33_port);
   U109 : XOR2_X1 port map( A => n228, B => B(31), Z => DIFF_31_port);
   U110 : XOR2_X1 port map( A => n231, B => B(30), Z => DIFF_30_port);
   U111 : XOR2_X1 port map( A => n230, B => B(29), Z => DIFF_29_port);
   U112 : XOR2_X1 port map( A => n233, B => B(27), Z => DIFF_27_port);
   U113 : XOR2_X1 port map( A => n236, B => B(26), Z => DIFF_26_port);
   U114 : XOR2_X1 port map( A => n235, B => B(25), Z => DIFF_25_port);
   U115 : XOR2_X1 port map( A => n237, B => B(23), Z => DIFF_23_port);
   U116 : XOR2_X1 port map( A => n240, B => B(22), Z => DIFF_22_port);
   U117 : XOR2_X1 port map( A => n239, B => B(21), Z => DIFF_21_port);
   U118 : XOR2_X1 port map( A => B(1), B => B(0), Z => DIFF_1_port);
   U119 : XOR2_X1 port map( A => n241, B => B(19), Z => DIFF_19_port);
   U120 : XOR2_X1 port map( A => n244, B => B(18), Z => DIFF_18_port);
   U121 : XOR2_X1 port map( A => n243, B => B(17), Z => DIFF_17_port);
   U122 : XOR2_X1 port map( A => n245, B => B(15), Z => DIFF_15_port);
   U123 : XOR2_X1 port map( A => n248, B => B(14), Z => DIFF_14_port);
   U124 : XOR2_X1 port map( A => n247, B => B(13), Z => DIFF_13_port);
   U125 : XOR2_X1 port map( A => n249, B => B(11), Z => DIFF_11_port);
   U126 : XOR2_X1 port map( A => n251, B => B(10), Z => DIFF_10_port);
   U1 : XNOR2_X1 port map( A => n189, B => B(6), ZN => DIFF_6_port);
   U2 : NOR2_X1 port map( A1 => n194, A2 => B(5), ZN => n189);
   U3 : NOR2_X1 port map( A1 => B(3), A2 => n211, ZN => n210);
   U4 : NOR2_X1 port map( A1 => B(7), A2 => n192, ZN => n191);
   U5 : XNOR2_X1 port map( A => B(8), B => n191, ZN => DIFF_8_port);
   U6 : OR3_X1 port map( A1 => B(5), A2 => B(6), A3 => n194, ZN => n192);
   U7 : OR3_X1 port map( A1 => B(7), A2 => B(8), A3 => n192, ZN => n190);
   U8 : OR3_X1 port map( A1 => B(3), A2 => B(4), A3 => n211, ZN => n194);
   U9 : XNOR2_X1 port map( A => B(4), B => n210, ZN => DIFF_4_port);
   U10 : XNOR2_X1 port map( A => B(12), B => n250, ZN => DIFF_12_port);
   U11 : NOR3_X1 port map( A1 => B(59), A2 => B(60), A3 => n198, ZN => n197);
   U12 : NOR2_X1 port map( A1 => B(43), A2 => n216, ZN => n217);
   U13 : NOR2_X1 port map( A1 => B(35), A2 => n224, ZN => n225);
   U14 : NOR2_X1 port map( A1 => B(51), A2 => n206, ZN => n207);
   U15 : NOR2_X1 port map( A1 => B(11), A2 => n249, ZN => n250);
   U16 : NOR2_X1 port map( A1 => B(15), A2 => n245, ZN => n246);
   U17 : NOR2_X1 port map( A1 => B(19), A2 => n241, ZN => n242);
   U18 : NOR2_X1 port map( A1 => B(23), A2 => n237, ZN => n238);
   U19 : NOR2_X1 port map( A1 => B(27), A2 => n233, ZN => n234);
   U20 : NOR2_X1 port map( A1 => B(39), A2 => n220, ZN => n221);
   U21 : NOR2_X1 port map( A1 => B(31), A2 => n228, ZN => n229);
   U22 : NOR2_X1 port map( A1 => B(59), A2 => n198, ZN => n199);
   U23 : NOR2_X1 port map( A1 => B(55), A2 => n202, ZN => n203);
   U24 : NAND2_X1 port map( A1 => n197, A2 => n193, ZN => n196);
   U25 : OR3_X1 port map( A1 => B(33), A2 => B(34), A3 => n226, ZN => n224);
   U26 : OR3_X1 port map( A1 => B(49), A2 => B(50), A3 => n208, ZN => n206);
   U27 : OR3_X1 port map( A1 => B(10), A2 => B(9), A3 => n190, ZN => n249);
   U28 : OR3_X1 port map( A1 => B(21), A2 => B(22), A3 => n239, ZN => n237);
   U29 : OR3_X1 port map( A1 => B(25), A2 => B(26), A3 => n235, ZN => n233);
   U30 : OR3_X1 port map( A1 => B(17), A2 => B(18), A3 => n243, ZN => n241);
   U31 : OR3_X1 port map( A1 => B(29), A2 => B(30), A3 => n230, ZN => n228);
   U32 : OR3_X1 port map( A1 => B(13), A2 => B(14), A3 => n247, ZN => n245);
   U33 : OR3_X1 port map( A1 => B(53), A2 => B(54), A3 => n204, ZN => n202);
   U34 : OR3_X1 port map( A1 => B(41), A2 => B(42), A3 => n218, ZN => n216);
   U35 : OR3_X1 port map( A1 => B(43), A2 => B(44), A3 => n216, ZN => n214);
   U36 : OR3_X1 port map( A1 => B(23), A2 => B(24), A3 => n237, ZN => n235);
   U37 : OR3_X1 port map( A1 => B(27), A2 => B(28), A3 => n233, ZN => n230);
   U38 : OR3_X1 port map( A1 => B(19), A2 => B(20), A3 => n241, ZN => n239);
   U39 : OR3_X1 port map( A1 => B(15), A2 => B(16), A3 => n245, ZN => n243);
   U40 : OR3_X1 port map( A1 => B(11), A2 => B(12), A3 => n249, ZN => n247);
   U41 : OR3_X1 port map( A1 => B(31), A2 => B(32), A3 => n228, ZN => n226);
   U42 : OR3_X1 port map( A1 => B(39), A2 => B(40), A3 => n220, ZN => n218);
   U43 : OR3_X1 port map( A1 => B(51), A2 => B(52), A3 => n206, ZN => n204);
   U44 : XNOR2_X1 port map( A => B(16), B => n246, ZN => DIFF_16_port);
   U45 : XNOR2_X1 port map( A => B(20), B => n242, ZN => DIFF_20_port);
   U46 : XNOR2_X1 port map( A => B(24), B => n238, ZN => DIFF_24_port);
   U47 : XNOR2_X1 port map( A => B(28), B => n234, ZN => DIFF_28_port);
   U48 : XNOR2_X1 port map( A => B(32), B => n229, ZN => DIFF_32_port);
   U49 : XNOR2_X1 port map( A => B(48), B => n213, ZN => DIFF_48_port);
   U50 : XNOR2_X1 port map( A => B(40), B => n221, ZN => DIFF_40_port);
   U51 : XNOR2_X1 port map( A => B(44), B => n217, ZN => DIFF_44_port);
   U52 : OR2_X1 port map( A1 => n226, A2 => B(33), ZN => n227);
   U53 : OR2_X1 port map( A1 => n214, A2 => B(45), ZN => n215);
   U54 : OR2_X1 port map( A1 => n190, A2 => B(9), ZN => n251);
   U55 : OR2_X1 port map( A1 => n247, A2 => B(13), ZN => n248);
   U56 : OR2_X1 port map( A1 => n230, A2 => B(29), ZN => n231);
   U57 : OR2_X1 port map( A1 => n243, A2 => B(17), ZN => n244);
   U58 : OR2_X1 port map( A1 => n239, A2 => B(21), ZN => n240);
   U59 : OR2_X1 port map( A1 => n235, A2 => B(25), ZN => n236);
   U60 : OR2_X1 port map( A1 => n208, A2 => B(49), ZN => n209);
   U61 : OR2_X1 port map( A1 => n218, A2 => B(41), ZN => n219);
   U62 : OR2_X1 port map( A1 => n204, A2 => B(53), ZN => n205);
   U63 : XNOR2_X1 port map( A => B(2), B => n232, ZN => DIFF_2_port);
   U64 : XNOR2_X1 port map( A => B(36), B => n225, ZN => DIFF_36_port);
   U65 : NOR2_X1 port map( A1 => B(47), A2 => n212, ZN => n213);
   U66 : XNOR2_X1 port map( A => B(60), B => n199, ZN => DIFF_60_port);
   U67 : XNOR2_X1 port map( A => B(52), B => n207, ZN => DIFF_52_port);
   U68 : OR3_X1 port map( A1 => B(57), A2 => B(58), A3 => n200, ZN => n198);
   U69 : OR3_X1 port map( A1 => B(45), A2 => B(46), A3 => n214, ZN => n212);
   U70 : OR3_X1 port map( A1 => B(37), A2 => B(38), A3 => n222, ZN => n220);
   U71 : OR3_X1 port map( A1 => B(47), A2 => B(48), A3 => n212, ZN => n208);
   U72 : OR3_X1 port map( A1 => B(35), A2 => B(36), A3 => n224, ZN => n222);
   U73 : OR3_X1 port map( A1 => B(55), A2 => B(56), A3 => n202, ZN => n200);
   U74 : XNOR2_X1 port map( A => n197, B => B(61), ZN => DIFF_61_port);
   U75 : XNOR2_X1 port map( A => B(56), B => n203, ZN => DIFF_56_port);
   U76 : OR2_X1 port map( A1 => n196, A2 => B(62), ZN => n195);
   U77 : OR2_X1 port map( A1 => n222, A2 => B(37), ZN => n223);
   U78 : OR2_X1 port map( A1 => n200, A2 => B(57), ZN => n201);
   U79 : OR3_X1 port map( A1 => B(1), A2 => B(2), A3 => B(0), ZN => n211);
   U80 : NOR2_X1 port map( A1 => B(0), A2 => B(1), ZN => n232);
   U83 : INV_X1 port map( A => B(61), ZN => n193);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_30_DW01_sub_0 is

   port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (63 downto 0);  CO : out std_logic);

end complementer_N64_30_DW01_sub_0;

architecture SYN_rpl of complementer_N64_30_DW01_sub_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal DIFF_62_port, DIFF_61_port, DIFF_60_port, DIFF_59_port, DIFF_58_port,
      DIFF_57_port, DIFF_56_port, DIFF_55_port, DIFF_54_port, DIFF_53_port, 
      DIFF_52_port, DIFF_51_port, DIFF_50_port, DIFF_49_port, DIFF_48_port, 
      DIFF_47_port, DIFF_46_port, DIFF_45_port, DIFF_44_port, DIFF_43_port, 
      DIFF_42_port, DIFF_41_port, DIFF_40_port, DIFF_39_port, DIFF_38_port, 
      DIFF_37_port, DIFF_36_port, DIFF_35_port, DIFF_34_port, DIFF_33_port, 
      DIFF_32_port, DIFF_31_port, DIFF_30_port, DIFF_29_port, DIFF_28_port, 
      DIFF_27_port, DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, 
      DIFF_22_port, DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, 
      DIFF_17_port, DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, 
      DIFF_12_port, DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, 
      DIFF_7_port, DIFF_6_port, DIFF_5_port, DIFF_4_port, DIFF_3_port, 
      DIFF_2_port, DIFF_1_port, DIFF_63_port, n190, n191, n192, n194, n196, 
      n197, n198, n199, n200, n202, n203, n204, n206, n207, n208, n210, n211, 
      n212, n213, n214, n216, n217, n218, n220, n221, n222, n224, n225, n226, 
      n228, n229, n230, n232, n233, n234, n235, n237, n238, n239, n241, n242, 
      n243, n245, n246, n247, n249, n250, n189, n193, n195, n201, n205, n209, 
      n215, n219, n223, n227, n231, n236, n240, n244, n248, n251 : std_logic;

begin
   DIFF <= ( DIFF_63_port, DIFF_62_port, DIFF_61_port, DIFF_60_port, 
      DIFF_59_port, DIFF_58_port, DIFF_57_port, DIFF_56_port, DIFF_55_port, 
      DIFF_54_port, DIFF_53_port, DIFF_52_port, DIFF_51_port, DIFF_50_port, 
      DIFF_49_port, DIFF_48_port, DIFF_47_port, DIFF_46_port, DIFF_45_port, 
      DIFF_44_port, DIFF_43_port, DIFF_42_port, DIFF_41_port, DIFF_40_port, 
      DIFF_39_port, DIFF_38_port, DIFF_37_port, DIFF_36_port, DIFF_35_port, 
      DIFF_34_port, DIFF_33_port, DIFF_32_port, DIFF_31_port, DIFF_30_port, 
      DIFF_29_port, DIFF_28_port, DIFF_27_port, DIFF_26_port, DIFF_25_port, 
      DIFF_24_port, DIFF_23_port, DIFF_22_port, DIFF_21_port, DIFF_20_port, 
      DIFF_19_port, DIFF_18_port, DIFF_17_port, DIFF_16_port, DIFF_15_port, 
      DIFF_14_port, DIFF_13_port, DIFF_12_port, DIFF_11_port, DIFF_10_port, 
      DIFF_9_port, DIFF_8_port, DIFF_7_port, DIFF_6_port, DIFF_5_port, 
      DIFF_4_port, DIFF_3_port, DIFF_2_port, DIFF_1_port, B(0) );
   
   U81 : XOR2_X1 port map( A => n190, B => B(9), Z => DIFF_9_port);
   U82 : XOR2_X1 port map( A => n192, B => B(7), Z => DIFF_7_port);
   U85 : XOR2_X1 port map( A => n196, B => B(62), Z => DIFF_62_port);
   U86 : XOR2_X1 port map( A => n194, B => B(5), Z => DIFF_5_port);
   U87 : XOR2_X1 port map( A => n198, B => B(59), Z => DIFF_59_port);
   U89 : XOR2_X1 port map( A => n200, B => B(57), Z => DIFF_57_port);
   U90 : XOR2_X1 port map( A => n202, B => B(55), Z => DIFF_55_port);
   U92 : XOR2_X1 port map( A => n204, B => B(53), Z => DIFF_53_port);
   U93 : XOR2_X1 port map( A => n206, B => B(51), Z => DIFF_51_port);
   U95 : XOR2_X1 port map( A => n208, B => B(49), Z => DIFF_49_port);
   U96 : XOR2_X1 port map( A => n212, B => B(47), Z => DIFF_47_port);
   U98 : XOR2_X1 port map( A => n214, B => B(45), Z => DIFF_45_port);
   U99 : XOR2_X1 port map( A => n216, B => B(43), Z => DIFF_43_port);
   U101 : XOR2_X1 port map( A => n218, B => B(41), Z => DIFF_41_port);
   U102 : XOR2_X1 port map( A => n211, B => B(3), Z => DIFF_3_port);
   U103 : XOR2_X1 port map( A => n220, B => B(39), Z => DIFF_39_port);
   U105 : XOR2_X1 port map( A => n222, B => B(37), Z => DIFF_37_port);
   U106 : XOR2_X1 port map( A => n224, B => B(35), Z => DIFF_35_port);
   U108 : XOR2_X1 port map( A => n226, B => B(33), Z => DIFF_33_port);
   U109 : XOR2_X1 port map( A => n228, B => B(31), Z => DIFF_31_port);
   U111 : XOR2_X1 port map( A => n230, B => B(29), Z => DIFF_29_port);
   U112 : XOR2_X1 port map( A => n233, B => B(27), Z => DIFF_27_port);
   U114 : XOR2_X1 port map( A => n235, B => B(25), Z => DIFF_25_port);
   U115 : XOR2_X1 port map( A => n237, B => B(23), Z => DIFF_23_port);
   U117 : XOR2_X1 port map( A => n239, B => B(21), Z => DIFF_21_port);
   U118 : XOR2_X1 port map( A => B(1), B => B(0), Z => DIFF_1_port);
   U119 : XOR2_X1 port map( A => n241, B => B(19), Z => DIFF_19_port);
   U121 : XOR2_X1 port map( A => n243, B => B(17), Z => DIFF_17_port);
   U122 : XOR2_X1 port map( A => n245, B => B(15), Z => DIFF_15_port);
   U124 : XOR2_X1 port map( A => n247, B => B(13), Z => DIFF_13_port);
   U125 : XOR2_X1 port map( A => n249, B => B(11), Z => DIFF_11_port);
   U1 : OR3_X1 port map( A1 => B(1), A2 => B(2), A3 => B(0), ZN => n211);
   U2 : XNOR2_X1 port map( A => n189, B => B(6), ZN => DIFF_6_port);
   U3 : NOR2_X1 port map( A1 => n194, A2 => B(5), ZN => n189);
   U4 : XNOR2_X1 port map( A => n193, B => B(10), ZN => DIFF_10_port);
   U5 : NOR2_X1 port map( A1 => n190, A2 => B(9), ZN => n193);
   U6 : XNOR2_X1 port map( A => B(12), B => n250, ZN => DIFF_12_port);
   U7 : NOR2_X1 port map( A1 => B(11), A2 => n249, ZN => n250);
   U8 : XNOR2_X1 port map( A => B(4), B => n210, ZN => DIFF_4_port);
   U9 : NOR2_X1 port map( A1 => B(3), A2 => n211, ZN => n210);
   U10 : XNOR2_X1 port map( A => B(8), B => n191, ZN => DIFF_8_port);
   U11 : NOR2_X1 port map( A1 => B(7), A2 => n192, ZN => n191);
   U12 : OR3_X1 port map( A1 => B(5), A2 => B(6), A3 => n194, ZN => n192);
   U13 : OR3_X1 port map( A1 => B(10), A2 => B(9), A3 => n190, ZN => n249);
   U14 : OR3_X1 port map( A1 => B(7), A2 => B(8), A3 => n192, ZN => n190);
   U15 : OR3_X1 port map( A1 => B(3), A2 => B(4), A3 => n211, ZN => n194);
   U16 : XNOR2_X1 port map( A => n195, B => B(50), ZN => DIFF_50_port);
   U17 : NOR2_X1 port map( A1 => n208, A2 => B(49), ZN => n195);
   U18 : XNOR2_X1 port map( A => n201, B => B(14), ZN => DIFF_14_port);
   U19 : NOR2_X1 port map( A1 => n247, A2 => B(13), ZN => n201);
   U20 : XNOR2_X1 port map( A => n205, B => B(30), ZN => DIFF_30_port);
   U21 : NOR2_X1 port map( A1 => n230, A2 => B(29), ZN => n205);
   U22 : XNOR2_X1 port map( A => n209, B => B(18), ZN => DIFF_18_port);
   U23 : NOR2_X1 port map( A1 => n243, A2 => B(17), ZN => n209);
   U24 : XNOR2_X1 port map( A => n215, B => B(22), ZN => DIFF_22_port);
   U25 : NOR2_X1 port map( A1 => n239, A2 => B(21), ZN => n215);
   U26 : XNOR2_X1 port map( A => n219, B => B(26), ZN => DIFF_26_port);
   U27 : NOR2_X1 port map( A1 => n235, A2 => B(25), ZN => n219);
   U28 : XNOR2_X1 port map( A => n223, B => B(38), ZN => DIFF_38_port);
   U29 : NOR2_X1 port map( A1 => n222, A2 => B(37), ZN => n223);
   U30 : XNOR2_X1 port map( A => n227, B => B(58), ZN => DIFF_58_port);
   U31 : NOR2_X1 port map( A1 => n200, A2 => B(57), ZN => n227);
   U32 : XNOR2_X1 port map( A => n231, B => B(54), ZN => DIFF_54_port);
   U33 : NOR2_X1 port map( A1 => n204, A2 => B(53), ZN => n231);
   U34 : XNOR2_X1 port map( A => B(20), B => n242, ZN => DIFF_20_port);
   U35 : NOR2_X1 port map( A1 => B(19), A2 => n241, ZN => n242);
   U36 : XNOR2_X1 port map( A => B(24), B => n238, ZN => DIFF_24_port);
   U37 : NOR2_X1 port map( A1 => B(23), A2 => n237, ZN => n238);
   U38 : XNOR2_X1 port map( A => B(44), B => n217, ZN => DIFF_44_port);
   U39 : NOR2_X1 port map( A1 => B(43), A2 => n216, ZN => n217);
   U40 : XNOR2_X1 port map( A => B(32), B => n229, ZN => DIFF_32_port);
   U41 : NOR2_X1 port map( A1 => B(31), A2 => n228, ZN => n229);
   U42 : XNOR2_X1 port map( A => B(16), B => n246, ZN => DIFF_16_port);
   U43 : NOR2_X1 port map( A1 => B(15), A2 => n245, ZN => n246);
   U44 : XNOR2_X1 port map( A => B(28), B => n234, ZN => DIFF_28_port);
   U45 : NOR2_X1 port map( A1 => B(27), A2 => n233, ZN => n234);
   U46 : XNOR2_X1 port map( A => B(48), B => n213, ZN => DIFF_48_port);
   U47 : NOR2_X1 port map( A1 => B(47), A2 => n212, ZN => n213);
   U48 : XNOR2_X1 port map( A => B(40), B => n221, ZN => DIFF_40_port);
   U49 : NOR2_X1 port map( A1 => B(39), A2 => n220, ZN => n221);
   U50 : XOR2_X1 port map( A => n197, B => n251, Z => DIFF_61_port);
   U51 : NAND2_X1 port map( A1 => n197, A2 => n251, ZN => n196);
   U52 : OR3_X1 port map( A1 => B(57), A2 => B(58), A3 => n200, ZN => n198);
   U53 : OR3_X1 port map( A1 => B(49), A2 => B(50), A3 => n208, ZN => n206);
   U54 : OR3_X1 port map( A1 => B(21), A2 => B(22), A3 => n239, ZN => n237);
   U55 : OR3_X1 port map( A1 => B(25), A2 => B(26), A3 => n235, ZN => n233);
   U56 : OR3_X1 port map( A1 => B(13), A2 => B(14), A3 => n247, ZN => n245);
   U57 : OR3_X1 port map( A1 => B(17), A2 => B(18), A3 => n243, ZN => n241);
   U58 : OR3_X1 port map( A1 => B(29), A2 => B(30), A3 => n230, ZN => n228);
   U59 : OR3_X1 port map( A1 => B(37), A2 => B(38), A3 => n222, ZN => n220);
   U60 : OR3_X1 port map( A1 => B(33), A2 => B(34), A3 => n226, ZN => n224);
   U61 : OR3_X1 port map( A1 => B(53), A2 => B(54), A3 => n204, ZN => n202);
   U62 : OR3_X1 port map( A1 => B(23), A2 => B(24), A3 => n237, ZN => n235);
   U63 : OR3_X1 port map( A1 => B(19), A2 => B(20), A3 => n241, ZN => n239);
   U64 : OR3_X1 port map( A1 => B(15), A2 => B(16), A3 => n245, ZN => n243);
   U65 : OR3_X1 port map( A1 => B(27), A2 => B(28), A3 => n233, ZN => n230);
   U66 : OR3_X1 port map( A1 => B(11), A2 => B(12), A3 => n249, ZN => n247);
   U67 : OR3_X1 port map( A1 => B(31), A2 => B(32), A3 => n228, ZN => n226);
   U68 : OR3_X1 port map( A1 => B(47), A2 => B(48), A3 => n212, ZN => n208);
   U69 : OR3_X1 port map( A1 => B(43), A2 => B(44), A3 => n216, ZN => n214);
   U70 : OR3_X1 port map( A1 => B(39), A2 => B(40), A3 => n220, ZN => n218);
   U71 : XNOR2_X1 port map( A => n236, B => B(34), ZN => DIFF_34_port);
   U72 : NOR2_X1 port map( A1 => n226, A2 => B(33), ZN => n236);
   U73 : XNOR2_X1 port map( A => B(2), B => n232, ZN => DIFF_2_port);
   U74 : NOR2_X1 port map( A1 => B(0), A2 => B(1), ZN => n232);
   U75 : NOR3_X1 port map( A1 => B(59), A2 => B(60), A3 => n198, ZN => n197);
   U76 : XNOR2_X1 port map( A => n240, B => B(42), ZN => DIFF_42_port);
   U77 : NOR2_X1 port map( A1 => n218, A2 => B(41), ZN => n240);
   U78 : XNOR2_X1 port map( A => n244, B => B(63), ZN => DIFF_63_port);
   U79 : NOR2_X1 port map( A1 => n196, A2 => B(62), ZN => n244);
   U80 : XNOR2_X1 port map( A => n248, B => B(46), ZN => DIFF_46_port);
   U83 : NOR2_X1 port map( A1 => n214, A2 => B(45), ZN => n248);
   U84 : XNOR2_X1 port map( A => B(60), B => n199, ZN => DIFF_60_port);
   U88 : NOR2_X1 port map( A1 => B(59), A2 => n198, ZN => n199);
   U91 : XNOR2_X1 port map( A => B(36), B => n225, ZN => DIFF_36_port);
   U94 : NOR2_X1 port map( A1 => B(35), A2 => n224, ZN => n225);
   U97 : XNOR2_X1 port map( A => B(56), B => n203, ZN => DIFF_56_port);
   U100 : NOR2_X1 port map( A1 => B(55), A2 => n202, ZN => n203);
   U104 : XNOR2_X1 port map( A => B(52), B => n207, ZN => DIFF_52_port);
   U107 : NOR2_X1 port map( A1 => B(51), A2 => n206, ZN => n207);
   U110 : OR3_X1 port map( A1 => B(41), A2 => B(42), A3 => n218, ZN => n216);
   U113 : OR3_X1 port map( A1 => B(45), A2 => B(46), A3 => n214, ZN => n212);
   U116 : OR3_X1 port map( A1 => B(35), A2 => B(36), A3 => n224, ZN => n222);
   U120 : OR3_X1 port map( A1 => B(51), A2 => B(52), A3 => n206, ZN => n204);
   U123 : OR3_X1 port map( A1 => B(55), A2 => B(56), A3 => n202, ZN => n200);
   U126 : INV_X1 port map( A => B(61), ZN => n251);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_31_DW01_sub_0 is

   port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (63 downto 0);  CO : out std_logic);

end complementer_N64_31_DW01_sub_0;

architecture SYN_rpl of complementer_N64_31_DW01_sub_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal DIFF_62_port, DIFF_63_port, DIFF_1_port, DIFF_2_port, DIFF_3_port, 
      DIFF_4_port, DIFF_5_port, DIFF_6_port, DIFF_7_port, DIFF_8_port, 
      DIFF_9_port, DIFF_10_port, DIFF_11_port, DIFF_12_port, DIFF_13_port, 
      DIFF_14_port, DIFF_15_port, DIFF_16_port, DIFF_17_port, DIFF_18_port, 
      DIFF_19_port, DIFF_20_port, DIFF_21_port, DIFF_22_port, DIFF_23_port, 
      DIFF_24_port, DIFF_25_port, DIFF_26_port, DIFF_27_port, DIFF_28_port, 
      DIFF_29_port, DIFF_30_port, DIFF_31_port, DIFF_32_port, DIFF_33_port, 
      DIFF_34_port, DIFF_35_port, DIFF_36_port, DIFF_37_port, DIFF_38_port, 
      DIFF_39_port, DIFF_40_port, DIFF_41_port, DIFF_42_port, DIFF_43_port, 
      DIFF_44_port, DIFF_45_port, DIFF_46_port, DIFF_47_port, DIFF_48_port, 
      DIFF_49_port, DIFF_50_port, DIFF_51_port, DIFF_52_port, DIFF_53_port, 
      DIFF_54_port, DIFF_55_port, DIFF_56_port, DIFF_57_port, DIFF_58_port, 
      DIFF_59_port, DIFF_60_port, DIFF_61_port, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, 
      n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, 
      n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, 
      n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, 
      n243, n244, n245, n246, n247, n248, n249, n250, n251, n189 : std_logic;

begin
   DIFF <= ( DIFF_63_port, DIFF_62_port, DIFF_61_port, DIFF_60_port, 
      DIFF_59_port, DIFF_58_port, DIFF_57_port, DIFF_56_port, DIFF_55_port, 
      DIFF_54_port, DIFF_53_port, DIFF_52_port, DIFF_51_port, DIFF_50_port, 
      DIFF_49_port, DIFF_48_port, DIFF_47_port, DIFF_46_port, DIFF_45_port, 
      DIFF_44_port, DIFF_43_port, DIFF_42_port, DIFF_41_port, DIFF_40_port, 
      DIFF_39_port, DIFF_38_port, DIFF_37_port, DIFF_36_port, DIFF_35_port, 
      DIFF_34_port, DIFF_33_port, DIFF_32_port, DIFF_31_port, DIFF_30_port, 
      DIFF_29_port, DIFF_28_port, DIFF_27_port, DIFF_26_port, DIFF_25_port, 
      DIFF_24_port, DIFF_23_port, DIFF_22_port, DIFF_21_port, DIFF_20_port, 
      DIFF_19_port, DIFF_18_port, DIFF_17_port, DIFF_16_port, DIFF_15_port, 
      DIFF_14_port, DIFF_13_port, DIFF_12_port, DIFF_11_port, DIFF_10_port, 
      DIFF_9_port, DIFF_8_port, DIFF_7_port, DIFF_6_port, DIFF_5_port, 
      DIFF_4_port, DIFF_3_port, DIFF_2_port, DIFF_1_port, B(0) );
   
   U81 : XOR2_X1 port map( A => n190, B => B(9), Z => DIFF_9_port);
   U82 : XOR2_X1 port map( A => n192, B => B(7), Z => DIFF_7_port);
   U83 : XOR2_X1 port map( A => n193, B => B(6), Z => DIFF_6_port);
   U84 : XOR2_X1 port map( A => n195, B => B(63), Z => DIFF_63_port);
   U85 : XOR2_X1 port map( A => n196, B => B(62), Z => DIFF_62_port);
   U86 : XOR2_X1 port map( A => n194, B => B(5), Z => DIFF_5_port);
   U87 : XOR2_X1 port map( A => n198, B => B(59), Z => DIFF_59_port);
   U88 : XOR2_X1 port map( A => n201, B => B(58), Z => DIFF_58_port);
   U89 : XOR2_X1 port map( A => n200, B => B(57), Z => DIFF_57_port);
   U90 : XOR2_X1 port map( A => n202, B => B(55), Z => DIFF_55_port);
   U91 : XOR2_X1 port map( A => n205, B => B(54), Z => DIFF_54_port);
   U92 : XOR2_X1 port map( A => n204, B => B(53), Z => DIFF_53_port);
   U93 : XOR2_X1 port map( A => n206, B => B(51), Z => DIFF_51_port);
   U94 : XOR2_X1 port map( A => n209, B => B(50), Z => DIFF_50_port);
   U95 : XOR2_X1 port map( A => n208, B => B(49), Z => DIFF_49_port);
   U96 : XOR2_X1 port map( A => n212, B => B(47), Z => DIFF_47_port);
   U97 : XOR2_X1 port map( A => n215, B => B(46), Z => DIFF_46_port);
   U98 : XOR2_X1 port map( A => n214, B => B(45), Z => DIFF_45_port);
   U99 : XOR2_X1 port map( A => n216, B => B(43), Z => DIFF_43_port);
   U100 : XOR2_X1 port map( A => n219, B => B(42), Z => DIFF_42_port);
   U101 : XOR2_X1 port map( A => n218, B => B(41), Z => DIFF_41_port);
   U102 : XOR2_X1 port map( A => n211, B => B(3), Z => DIFF_3_port);
   U103 : XOR2_X1 port map( A => n220, B => B(39), Z => DIFF_39_port);
   U104 : XOR2_X1 port map( A => n223, B => B(38), Z => DIFF_38_port);
   U105 : XOR2_X1 port map( A => n222, B => B(37), Z => DIFF_37_port);
   U106 : XOR2_X1 port map( A => n224, B => B(35), Z => DIFF_35_port);
   U107 : XOR2_X1 port map( A => n227, B => B(34), Z => DIFF_34_port);
   U108 : XOR2_X1 port map( A => n226, B => B(33), Z => DIFF_33_port);
   U109 : XOR2_X1 port map( A => n228, B => B(31), Z => DIFF_31_port);
   U110 : XOR2_X1 port map( A => n231, B => B(30), Z => DIFF_30_port);
   U111 : XOR2_X1 port map( A => n230, B => B(29), Z => DIFF_29_port);
   U112 : XOR2_X1 port map( A => n233, B => B(27), Z => DIFF_27_port);
   U113 : XOR2_X1 port map( A => n236, B => B(26), Z => DIFF_26_port);
   U114 : XOR2_X1 port map( A => n235, B => B(25), Z => DIFF_25_port);
   U115 : XOR2_X1 port map( A => n237, B => B(23), Z => DIFF_23_port);
   U116 : XOR2_X1 port map( A => n240, B => B(22), Z => DIFF_22_port);
   U117 : XOR2_X1 port map( A => n239, B => B(21), Z => DIFF_21_port);
   U118 : XOR2_X1 port map( A => B(1), B => B(0), Z => DIFF_1_port);
   U119 : XOR2_X1 port map( A => n241, B => B(19), Z => DIFF_19_port);
   U120 : XOR2_X1 port map( A => n244, B => B(18), Z => DIFF_18_port);
   U121 : XOR2_X1 port map( A => n243, B => B(17), Z => DIFF_17_port);
   U122 : XOR2_X1 port map( A => n245, B => B(15), Z => DIFF_15_port);
   U123 : XOR2_X1 port map( A => n248, B => B(14), Z => DIFF_14_port);
   U124 : XOR2_X1 port map( A => n247, B => B(13), Z => DIFF_13_port);
   U125 : XOR2_X1 port map( A => n249, B => B(11), Z => DIFF_11_port);
   U126 : XOR2_X1 port map( A => n251, B => B(10), Z => DIFF_10_port);
   U1 : NOR2_X1 port map( A1 => B(31), A2 => n228, ZN => n229);
   U2 : NOR2_X1 port map( A1 => B(43), A2 => n216, ZN => n217);
   U3 : NOR2_X1 port map( A1 => B(39), A2 => n220, ZN => n221);
   U4 : NAND2_X1 port map( A1 => n197, A2 => n189, ZN => n196);
   U5 : OR3_X1 port map( A1 => B(31), A2 => B(32), A3 => n228, ZN => n226);
   U6 : XNOR2_X1 port map( A => B(48), B => n213, ZN => DIFF_48_port);
   U7 : OR2_X1 port map( A1 => n226, A2 => B(33), ZN => n227);
   U8 : OR2_X1 port map( A1 => n208, A2 => B(49), ZN => n209);
   U9 : OR2_X1 port map( A1 => n204, A2 => B(53), ZN => n205);
   U10 : XNOR2_X1 port map( A => B(4), B => n210, ZN => DIFF_4_port);
   U11 : NOR2_X1 port map( A1 => B(3), A2 => n211, ZN => n210);
   U12 : NOR2_X1 port map( A1 => B(7), A2 => n192, ZN => n191);
   U13 : NOR2_X1 port map( A1 => B(0), A2 => B(1), ZN => n232);
   U14 : OR3_X1 port map( A1 => B(5), A2 => B(6), A3 => n194, ZN => n192);
   U15 : OR3_X1 port map( A1 => B(1), A2 => B(2), A3 => B(0), ZN => n211);
   U16 : OR3_X1 port map( A1 => B(7), A2 => B(8), A3 => n192, ZN => n190);
   U17 : OR3_X1 port map( A1 => B(3), A2 => B(4), A3 => n211, ZN => n194);
   U18 : XNOR2_X1 port map( A => B(2), B => n232, ZN => DIFF_2_port);
   U19 : XNOR2_X1 port map( A => B(8), B => n191, ZN => DIFF_8_port);
   U20 : OR2_X1 port map( A1 => n194, A2 => B(5), ZN => n193);
   U21 : NOR3_X1 port map( A1 => B(59), A2 => B(60), A3 => n198, ZN => n197);
   U22 : XNOR2_X1 port map( A => n197, B => B(61), ZN => DIFF_61_port);
   U23 : XNOR2_X1 port map( A => B(60), B => n199, ZN => DIFF_60_port);
   U24 : XNOR2_X1 port map( A => B(12), B => n250, ZN => DIFF_12_port);
   U25 : NOR2_X1 port map( A1 => B(59), A2 => n198, ZN => n199);
   U26 : NOR2_X1 port map( A1 => B(11), A2 => n249, ZN => n250);
   U27 : NOR2_X1 port map( A1 => B(15), A2 => n245, ZN => n246);
   U28 : NOR2_X1 port map( A1 => B(19), A2 => n241, ZN => n242);
   U29 : NOR2_X1 port map( A1 => B(23), A2 => n237, ZN => n238);
   U30 : NOR2_X1 port map( A1 => B(27), A2 => n233, ZN => n234);
   U31 : NOR2_X1 port map( A1 => B(35), A2 => n224, ZN => n225);
   U32 : NOR2_X1 port map( A1 => B(55), A2 => n202, ZN => n203);
   U33 : NOR2_X1 port map( A1 => B(51), A2 => n206, ZN => n207);
   U34 : NOR2_X1 port map( A1 => B(47), A2 => n212, ZN => n213);
   U35 : OR3_X1 port map( A1 => B(57), A2 => B(58), A3 => n200, ZN => n198);
   U36 : OR3_X1 port map( A1 => B(33), A2 => B(34), A3 => n226, ZN => n224);
   U37 : OR3_X1 port map( A1 => B(37), A2 => B(38), A3 => n222, ZN => n220);
   U38 : OR3_X1 port map( A1 => B(49), A2 => B(50), A3 => n208, ZN => n206);
   U39 : OR3_X1 port map( A1 => B(41), A2 => B(42), A3 => n218, ZN => n216);
   U40 : OR3_X1 port map( A1 => B(53), A2 => B(54), A3 => n204, ZN => n202);
   U41 : OR3_X1 port map( A1 => B(21), A2 => B(22), A3 => n239, ZN => n237);
   U42 : OR3_X1 port map( A1 => B(25), A2 => B(26), A3 => n235, ZN => n233);
   U43 : OR3_X1 port map( A1 => B(17), A2 => B(18), A3 => n243, ZN => n241);
   U44 : OR3_X1 port map( A1 => B(13), A2 => B(14), A3 => n247, ZN => n245);
   U45 : OR3_X1 port map( A1 => B(29), A2 => B(30), A3 => n230, ZN => n228);
   U46 : OR3_X1 port map( A1 => B(10), A2 => B(9), A3 => n190, ZN => n249);
   U47 : OR3_X1 port map( A1 => B(45), A2 => B(46), A3 => n214, ZN => n212);
   U48 : OR3_X1 port map( A1 => B(43), A2 => B(44), A3 => n216, ZN => n214);
   U49 : OR3_X1 port map( A1 => B(47), A2 => B(48), A3 => n212, ZN => n208);
   U50 : OR3_X1 port map( A1 => B(51), A2 => B(52), A3 => n206, ZN => n204);
   U51 : XNOR2_X1 port map( A => B(16), B => n246, ZN => DIFF_16_port);
   U52 : XNOR2_X1 port map( A => B(20), B => n242, ZN => DIFF_20_port);
   U53 : XNOR2_X1 port map( A => B(24), B => n238, ZN => DIFF_24_port);
   U54 : XNOR2_X1 port map( A => B(28), B => n234, ZN => DIFF_28_port);
   U55 : XNOR2_X1 port map( A => B(40), B => n221, ZN => DIFF_40_port);
   U56 : XNOR2_X1 port map( A => B(32), B => n229, ZN => DIFF_32_port);
   U57 : XNOR2_X1 port map( A => B(36), B => n225, ZN => DIFF_36_port);
   U58 : XNOR2_X1 port map( A => B(56), B => n203, ZN => DIFF_56_port);
   U59 : XNOR2_X1 port map( A => B(52), B => n207, ZN => DIFF_52_port);
   U60 : XNOR2_X1 port map( A => B(44), B => n217, ZN => DIFF_44_port);
   U61 : OR3_X1 port map( A1 => B(39), A2 => B(40), A3 => n220, ZN => n218);
   U62 : OR3_X1 port map( A1 => B(23), A2 => B(24), A3 => n237, ZN => n235);
   U63 : OR3_X1 port map( A1 => B(19), A2 => B(20), A3 => n241, ZN => n239);
   U64 : OR3_X1 port map( A1 => B(27), A2 => B(28), A3 => n233, ZN => n230);
   U65 : OR3_X1 port map( A1 => B(15), A2 => B(16), A3 => n245, ZN => n243);
   U66 : OR3_X1 port map( A1 => B(11), A2 => B(12), A3 => n249, ZN => n247);
   U67 : OR3_X1 port map( A1 => B(35), A2 => B(36), A3 => n224, ZN => n222);
   U68 : OR3_X1 port map( A1 => B(55), A2 => B(56), A3 => n202, ZN => n200);
   U69 : OR2_X1 port map( A1 => n190, A2 => B(9), ZN => n251);
   U70 : OR2_X1 port map( A1 => n247, A2 => B(13), ZN => n248);
   U71 : OR2_X1 port map( A1 => n230, A2 => B(29), ZN => n231);
   U72 : OR2_X1 port map( A1 => n243, A2 => B(17), ZN => n244);
   U73 : OR2_X1 port map( A1 => n239, A2 => B(21), ZN => n240);
   U74 : OR2_X1 port map( A1 => n235, A2 => B(25), ZN => n236);
   U75 : OR2_X1 port map( A1 => n222, A2 => B(37), ZN => n223);
   U76 : OR2_X1 port map( A1 => n200, A2 => B(57), ZN => n201);
   U77 : OR2_X1 port map( A1 => n214, A2 => B(45), ZN => n215);
   U78 : OR2_X1 port map( A1 => n218, A2 => B(41), ZN => n219);
   U79 : OR2_X1 port map( A1 => n196, A2 => B(62), ZN => n195);
   U80 : INV_X1 port map( A => B(61), ZN => n189);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_0_DW01_sub_0 is

   port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (63 downto 0);  CO : out std_logic);

end complementer_N64_0_DW01_sub_0;

architecture SYN_rpl of complementer_N64_0_DW01_sub_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal DIFF_62_port, DIFF_61_port, DIFF_60_port, DIFF_59_port, DIFF_58_port,
      DIFF_57_port, DIFF_56_port, DIFF_55_port, DIFF_54_port, DIFF_53_port, 
      DIFF_52_port, DIFF_51_port, DIFF_50_port, DIFF_49_port, DIFF_48_port, 
      DIFF_47_port, DIFF_46_port, DIFF_45_port, DIFF_44_port, DIFF_43_port, 
      DIFF_42_port, DIFF_41_port, DIFF_40_port, DIFF_39_port, DIFF_38_port, 
      DIFF_37_port, DIFF_36_port, DIFF_35_port, DIFF_34_port, DIFF_33_port, 
      DIFF_32_port, DIFF_31_port, DIFF_30_port, DIFF_29_port, DIFF_28_port, 
      DIFF_27_port, DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, 
      DIFF_22_port, DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, 
      DIFF_17_port, DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, 
      DIFF_12_port, DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, 
      DIFF_7_port, DIFF_6_port, DIFF_5_port, DIFF_4_port, DIFF_3_port, 
      DIFF_2_port, DIFF_1_port, DIFF_63_port, n190, n191, n192, n194, n196, 
      n197, n198, n199, n200, n202, n203, n204, n206, n207, n208, n210, n211, 
      n212, n213, n214, n216, n217, n218, n220, n221, n222, n224, n225, n226, 
      n228, n229, n230, n232, n233, n234, n235, n237, n238, n239, n241, n242, 
      n243, n245, n246, n247, n249, n250, n189, n193, n195, n201, n205, n209, 
      n215, n219, n223, n227, n231, n236, n240, n244, n248, n251 : std_logic;

begin
   DIFF <= ( DIFF_63_port, DIFF_62_port, DIFF_61_port, DIFF_60_port, 
      DIFF_59_port, DIFF_58_port, DIFF_57_port, DIFF_56_port, DIFF_55_port, 
      DIFF_54_port, DIFF_53_port, DIFF_52_port, DIFF_51_port, DIFF_50_port, 
      DIFF_49_port, DIFF_48_port, DIFF_47_port, DIFF_46_port, DIFF_45_port, 
      DIFF_44_port, DIFF_43_port, DIFF_42_port, DIFF_41_port, DIFF_40_port, 
      DIFF_39_port, DIFF_38_port, DIFF_37_port, DIFF_36_port, DIFF_35_port, 
      DIFF_34_port, DIFF_33_port, DIFF_32_port, DIFF_31_port, DIFF_30_port, 
      DIFF_29_port, DIFF_28_port, DIFF_27_port, DIFF_26_port, DIFF_25_port, 
      DIFF_24_port, DIFF_23_port, DIFF_22_port, DIFF_21_port, DIFF_20_port, 
      DIFF_19_port, DIFF_18_port, DIFF_17_port, DIFF_16_port, DIFF_15_port, 
      DIFF_14_port, DIFF_13_port, DIFF_12_port, DIFF_11_port, DIFF_10_port, 
      DIFF_9_port, DIFF_8_port, DIFF_7_port, DIFF_6_port, DIFF_5_port, 
      DIFF_4_port, DIFF_3_port, DIFF_2_port, DIFF_1_port, B(0) );
   
   U81 : XOR2_X1 port map( A => n190, B => B(9), Z => DIFF_9_port);
   U82 : XOR2_X1 port map( A => n192, B => B(7), Z => DIFF_7_port);
   U85 : XOR2_X1 port map( A => n196, B => B(62), Z => DIFF_62_port);
   U86 : XOR2_X1 port map( A => n194, B => B(5), Z => DIFF_5_port);
   U87 : XOR2_X1 port map( A => n198, B => B(59), Z => DIFF_59_port);
   U89 : XOR2_X1 port map( A => n200, B => B(57), Z => DIFF_57_port);
   U90 : XOR2_X1 port map( A => n202, B => B(55), Z => DIFF_55_port);
   U92 : XOR2_X1 port map( A => n204, B => B(53), Z => DIFF_53_port);
   U93 : XOR2_X1 port map( A => n206, B => B(51), Z => DIFF_51_port);
   U95 : XOR2_X1 port map( A => n208, B => B(49), Z => DIFF_49_port);
   U96 : XOR2_X1 port map( A => n212, B => B(47), Z => DIFF_47_port);
   U98 : XOR2_X1 port map( A => n214, B => B(45), Z => DIFF_45_port);
   U99 : XOR2_X1 port map( A => n216, B => B(43), Z => DIFF_43_port);
   U101 : XOR2_X1 port map( A => n218, B => B(41), Z => DIFF_41_port);
   U102 : XOR2_X1 port map( A => n211, B => B(3), Z => DIFF_3_port);
   U103 : XOR2_X1 port map( A => n220, B => B(39), Z => DIFF_39_port);
   U105 : XOR2_X1 port map( A => n222, B => B(37), Z => DIFF_37_port);
   U106 : XOR2_X1 port map( A => n224, B => B(35), Z => DIFF_35_port);
   U108 : XOR2_X1 port map( A => n226, B => B(33), Z => DIFF_33_port);
   U109 : XOR2_X1 port map( A => n228, B => B(31), Z => DIFF_31_port);
   U111 : XOR2_X1 port map( A => n230, B => B(29), Z => DIFF_29_port);
   U112 : XOR2_X1 port map( A => n233, B => B(27), Z => DIFF_27_port);
   U114 : XOR2_X1 port map( A => n235, B => B(25), Z => DIFF_25_port);
   U115 : XOR2_X1 port map( A => n237, B => B(23), Z => DIFF_23_port);
   U117 : XOR2_X1 port map( A => n239, B => B(21), Z => DIFF_21_port);
   U119 : XOR2_X1 port map( A => n241, B => B(19), Z => DIFF_19_port);
   U121 : XOR2_X1 port map( A => n243, B => B(17), Z => DIFF_17_port);
   U122 : XOR2_X1 port map( A => n245, B => B(15), Z => DIFF_15_port);
   U124 : XOR2_X1 port map( A => n247, B => B(13), Z => DIFF_13_port);
   U125 : XOR2_X1 port map( A => n249, B => B(11), Z => DIFF_11_port);
   U1 : XOR2_X1 port map( A => B(1), B => B(0), Z => DIFF_1_port);
   U2 : XNOR2_X1 port map( A => B(48), B => n213, ZN => DIFF_48_port);
   U3 : NOR2_X1 port map( A1 => B(47), A2 => n212, ZN => n213);
   U4 : XOR2_X1 port map( A => n197, B => n251, Z => DIFF_61_port);
   U5 : NAND2_X1 port map( A1 => n197, A2 => n251, ZN => n196);
   U6 : OR3_X1 port map( A1 => B(37), A2 => B(38), A3 => n222, ZN => n220);
   U7 : OR3_X1 port map( A1 => B(47), A2 => B(48), A3 => n212, ZN => n208);
   U8 : XNOR2_X1 port map( A => n189, B => B(38), ZN => DIFF_38_port);
   U9 : NOR2_X1 port map( A1 => n222, A2 => B(37), ZN => n189);
   U10 : XNOR2_X1 port map( A => n193, B => B(6), ZN => DIFF_6_port);
   U11 : NOR2_X1 port map( A1 => n194, A2 => B(5), ZN => n193);
   U12 : XNOR2_X1 port map( A => B(4), B => n210, ZN => DIFF_4_port);
   U13 : NOR2_X1 port map( A1 => B(3), A2 => n211, ZN => n210);
   U14 : XNOR2_X1 port map( A => B(8), B => n191, ZN => DIFF_8_port);
   U15 : NOR2_X1 port map( A1 => B(7), A2 => n192, ZN => n191);
   U16 : XNOR2_X1 port map( A => B(2), B => n232, ZN => DIFF_2_port);
   U17 : NOR2_X1 port map( A1 => B(0), A2 => B(1), ZN => n232);
   U18 : OR3_X1 port map( A1 => B(5), A2 => B(6), A3 => n194, ZN => n192);
   U19 : OR3_X1 port map( A1 => B(1), A2 => B(2), A3 => B(0), ZN => n211);
   U20 : OR3_X1 port map( A1 => B(7), A2 => B(8), A3 => n192, ZN => n190);
   U21 : OR3_X1 port map( A1 => B(3), A2 => B(4), A3 => n211, ZN => n194);
   U22 : NOR3_X1 port map( A1 => B(59), A2 => B(60), A3 => n198, ZN => n197);
   U23 : XNOR2_X1 port map( A => n195, B => B(14), ZN => DIFF_14_port);
   U24 : NOR2_X1 port map( A1 => n247, A2 => B(13), ZN => n195);
   U25 : XNOR2_X1 port map( A => n201, B => B(34), ZN => DIFF_34_port);
   U26 : NOR2_X1 port map( A1 => n226, A2 => B(33), ZN => n201);
   U27 : XNOR2_X1 port map( A => n205, B => B(63), ZN => DIFF_63_port);
   U28 : NOR2_X1 port map( A1 => n196, A2 => B(62), ZN => n205);
   U29 : XNOR2_X1 port map( A => n209, B => B(58), ZN => DIFF_58_port);
   U30 : NOR2_X1 port map( A1 => n200, A2 => B(57), ZN => n209);
   U31 : XNOR2_X1 port map( A => n215, B => B(54), ZN => DIFF_54_port);
   U32 : NOR2_X1 port map( A1 => n204, A2 => B(53), ZN => n215);
   U33 : XNOR2_X1 port map( A => n219, B => B(50), ZN => DIFF_50_port);
   U34 : NOR2_X1 port map( A1 => n208, A2 => B(49), ZN => n219);
   U35 : XNOR2_X1 port map( A => n223, B => B(46), ZN => DIFF_46_port);
   U36 : NOR2_X1 port map( A1 => n214, A2 => B(45), ZN => n223);
   U37 : XNOR2_X1 port map( A => n227, B => B(42), ZN => DIFF_42_port);
   U38 : NOR2_X1 port map( A1 => n218, A2 => B(41), ZN => n227);
   U39 : XNOR2_X1 port map( A => n231, B => B(10), ZN => DIFF_10_port);
   U40 : NOR2_X1 port map( A1 => n190, A2 => B(9), ZN => n231);
   U41 : XNOR2_X1 port map( A => B(20), B => n242, ZN => DIFF_20_port);
   U42 : NOR2_X1 port map( A1 => B(19), A2 => n241, ZN => n242);
   U43 : XNOR2_X1 port map( A => B(12), B => n250, ZN => DIFF_12_port);
   U44 : NOR2_X1 port map( A1 => B(11), A2 => n249, ZN => n250);
   U45 : XNOR2_X1 port map( A => B(16), B => n246, ZN => DIFF_16_port);
   U46 : NOR2_X1 port map( A1 => B(15), A2 => n245, ZN => n246);
   U47 : XNOR2_X1 port map( A => B(24), B => n238, ZN => DIFF_24_port);
   U48 : NOR2_X1 port map( A1 => B(23), A2 => n237, ZN => n238);
   U49 : XNOR2_X1 port map( A => B(28), B => n234, ZN => DIFF_28_port);
   U50 : NOR2_X1 port map( A1 => B(27), A2 => n233, ZN => n234);
   U51 : XNOR2_X1 port map( A => B(40), B => n221, ZN => DIFF_40_port);
   U52 : NOR2_X1 port map( A1 => B(39), A2 => n220, ZN => n221);
   U53 : XNOR2_X1 port map( A => B(32), B => n229, ZN => DIFF_32_port);
   U54 : NOR2_X1 port map( A1 => B(31), A2 => n228, ZN => n229);
   U55 : XNOR2_X1 port map( A => B(36), B => n225, ZN => DIFF_36_port);
   U56 : NOR2_X1 port map( A1 => B(35), A2 => n224, ZN => n225);
   U57 : XNOR2_X1 port map( A => B(60), B => n199, ZN => DIFF_60_port);
   U58 : NOR2_X1 port map( A1 => B(59), A2 => n198, ZN => n199);
   U59 : XNOR2_X1 port map( A => B(56), B => n203, ZN => DIFF_56_port);
   U60 : NOR2_X1 port map( A1 => B(55), A2 => n202, ZN => n203);
   U61 : XNOR2_X1 port map( A => B(52), B => n207, ZN => DIFF_52_port);
   U62 : NOR2_X1 port map( A1 => B(51), A2 => n206, ZN => n207);
   U63 : XNOR2_X1 port map( A => B(44), B => n217, ZN => DIFF_44_port);
   U64 : NOR2_X1 port map( A1 => B(43), A2 => n216, ZN => n217);
   U65 : OR3_X1 port map( A1 => B(57), A2 => B(58), A3 => n200, ZN => n198);
   U66 : OR3_X1 port map( A1 => B(21), A2 => B(22), A3 => n239, ZN => n237);
   U67 : OR3_X1 port map( A1 => B(17), A2 => B(18), A3 => n243, ZN => n241);
   U68 : OR3_X1 port map( A1 => B(25), A2 => B(26), A3 => n235, ZN => n233);
   U69 : OR3_X1 port map( A1 => B(13), A2 => B(14), A3 => n247, ZN => n245);
   U70 : OR3_X1 port map( A1 => B(29), A2 => B(30), A3 => n230, ZN => n228);
   U71 : OR3_X1 port map( A1 => B(10), A2 => B(9), A3 => n190, ZN => n249);
   U72 : OR3_X1 port map( A1 => B(33), A2 => B(34), A3 => n226, ZN => n224);
   U73 : OR3_X1 port map( A1 => B(41), A2 => B(42), A3 => n218, ZN => n216);
   U74 : OR3_X1 port map( A1 => B(45), A2 => B(46), A3 => n214, ZN => n212);
   U75 : OR3_X1 port map( A1 => B(49), A2 => B(50), A3 => n208, ZN => n206);
   U76 : OR3_X1 port map( A1 => B(53), A2 => B(54), A3 => n204, ZN => n202);
   U77 : OR3_X1 port map( A1 => B(19), A2 => B(20), A3 => n241, ZN => n239);
   U78 : OR3_X1 port map( A1 => B(23), A2 => B(24), A3 => n237, ZN => n235);
   U79 : OR3_X1 port map( A1 => B(27), A2 => B(28), A3 => n233, ZN => n230);
   U80 : OR3_X1 port map( A1 => B(15), A2 => B(16), A3 => n245, ZN => n243);
   U83 : OR3_X1 port map( A1 => B(11), A2 => B(12), A3 => n249, ZN => n247);
   U84 : OR3_X1 port map( A1 => B(31), A2 => B(32), A3 => n228, ZN => n226);
   U88 : OR3_X1 port map( A1 => B(35), A2 => B(36), A3 => n224, ZN => n222);
   U91 : OR3_X1 port map( A1 => B(39), A2 => B(40), A3 => n220, ZN => n218);
   U94 : OR3_X1 port map( A1 => B(43), A2 => B(44), A3 => n216, ZN => n214);
   U97 : OR3_X1 port map( A1 => B(51), A2 => B(52), A3 => n206, ZN => n204);
   U100 : OR3_X1 port map( A1 => B(55), A2 => B(56), A3 => n202, ZN => n200);
   U104 : XNOR2_X1 port map( A => n236, B => B(30), ZN => DIFF_30_port);
   U107 : NOR2_X1 port map( A1 => n230, A2 => B(29), ZN => n236);
   U110 : XNOR2_X1 port map( A => n240, B => B(18), ZN => DIFF_18_port);
   U113 : NOR2_X1 port map( A1 => n243, A2 => B(17), ZN => n240);
   U116 : XNOR2_X1 port map( A => n244, B => B(22), ZN => DIFF_22_port);
   U118 : NOR2_X1 port map( A1 => n239, A2 => B(21), ZN => n244);
   U120 : XNOR2_X1 port map( A => n248, B => B(26), ZN => DIFF_26_port);
   U123 : NOR2_X1 port map( A1 => n235, A2 => B(25), ZN => n248);
   U126 : INV_X1 port map( A => B(61), ZN => n251);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_1 is

   port( input : in std_logic_vector (63 downto 0);  complement2 : out 
         std_logic_vector (63 downto 0));

end complementer_N64_1;

architecture SYN_beh of complementer_N64_1 is

   component complementer_N64_1_DW01_sub_0
      port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (63 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n2, n_3112 : std_logic;

begin
   
   n1 <= '0';
   n2 <= '0';
   sub_add_29_b0 : complementer_N64_1_DW01_sub_0 port map( A(63) => n1, A(62) 
                           => n1, A(61) => n1, A(60) => n1, A(59) => n1, A(58) 
                           => n1, A(57) => n1, A(56) => n1, A(55) => n1, A(54) 
                           => n1, A(53) => n1, A(52) => n1, A(51) => n1, A(50) 
                           => n1, A(49) => n1, A(48) => n1, A(47) => n1, A(46) 
                           => n1, A(45) => n1, A(44) => n1, A(43) => n1, A(42) 
                           => n1, A(41) => n1, A(40) => n1, A(39) => n1, A(38) 
                           => n1, A(37) => n1, A(36) => n1, A(35) => n1, A(34) 
                           => n1, A(33) => n1, A(32) => n1, A(31) => n1, A(30) 
                           => n1, A(29) => n1, A(28) => n1, A(27) => n1, A(26) 
                           => n1, A(25) => n1, A(24) => n1, A(23) => n1, A(22) 
                           => n1, A(21) => n1, A(20) => n1, A(19) => n1, A(18) 
                           => n1, A(17) => n1, A(16) => n1, A(15) => n1, A(14) 
                           => n1, A(13) => n1, A(12) => n1, A(11) => n1, A(10) 
                           => n1, A(9) => n1, A(8) => n1, A(7) => n1, A(6) => 
                           n1, A(5) => n1, A(4) => n1, A(3) => n1, A(2) => n1, 
                           A(1) => n1, A(0) => n2, B(63) => input(63), B(62) =>
                           input(62), B(61) => input(61), B(60) => input(60), 
                           B(59) => input(59), B(58) => input(58), B(57) => 
                           input(57), B(56) => input(56), B(55) => input(55), 
                           B(54) => input(54), B(53) => input(53), B(52) => 
                           input(52), B(51) => input(51), B(50) => input(50), 
                           B(49) => input(49), B(48) => input(48), B(47) => 
                           input(47), B(46) => input(46), B(45) => input(45), 
                           B(44) => input(44), B(43) => input(43), B(42) => 
                           input(42), B(41) => input(41), B(40) => input(40), 
                           B(39) => input(39), B(38) => input(38), B(37) => 
                           input(37), B(36) => input(36), B(35) => input(35), 
                           B(34) => input(34), B(33) => input(33), B(32) => 
                           input(32), B(31) => input(31), B(30) => input(30), 
                           B(29) => input(29), B(28) => input(28), B(27) => 
                           input(27), B(26) => input(26), B(25) => input(25), 
                           B(24) => input(24), B(23) => input(23), B(22) => 
                           input(22), B(21) => input(21), B(20) => input(20), 
                           B(19) => input(19), B(18) => input(18), B(17) => 
                           input(17), B(16) => input(16), B(15) => input(15), 
                           B(14) => input(14), B(13) => input(13), B(12) => 
                           input(12), B(11) => input(11), B(10) => input(10), 
                           B(9) => input(9), B(8) => input(8), B(7) => input(7)
                           , B(6) => input(6), B(5) => input(5), B(4) => 
                           input(4), B(3) => input(3), B(2) => input(2), B(1) 
                           => input(1), B(0) => input(0), CI => n1, DIFF(63) =>
                           complement2(63), DIFF(62) => complement2(62), 
                           DIFF(61) => complement2(61), DIFF(60) => 
                           complement2(60), DIFF(59) => complement2(59), 
                           DIFF(58) => complement2(58), DIFF(57) => 
                           complement2(57), DIFF(56) => complement2(56), 
                           DIFF(55) => complement2(55), DIFF(54) => 
                           complement2(54), DIFF(53) => complement2(53), 
                           DIFF(52) => complement2(52), DIFF(51) => 
                           complement2(51), DIFF(50) => complement2(50), 
                           DIFF(49) => complement2(49), DIFF(48) => 
                           complement2(48), DIFF(47) => complement2(47), 
                           DIFF(46) => complement2(46), DIFF(45) => 
                           complement2(45), DIFF(44) => complement2(44), 
                           DIFF(43) => complement2(43), DIFF(42) => 
                           complement2(42), DIFF(41) => complement2(41), 
                           DIFF(40) => complement2(40), DIFF(39) => 
                           complement2(39), DIFF(38) => complement2(38), 
                           DIFF(37) => complement2(37), DIFF(36) => 
                           complement2(36), DIFF(35) => complement2(35), 
                           DIFF(34) => complement2(34), DIFF(33) => 
                           complement2(33), DIFF(32) => complement2(32), 
                           DIFF(31) => complement2(31), DIFF(30) => 
                           complement2(30), DIFF(29) => complement2(29), 
                           DIFF(28) => complement2(28), DIFF(27) => 
                           complement2(27), DIFF(26) => complement2(26), 
                           DIFF(25) => complement2(25), DIFF(24) => 
                           complement2(24), DIFF(23) => complement2(23), 
                           DIFF(22) => complement2(22), DIFF(21) => 
                           complement2(21), DIFF(20) => complement2(20), 
                           DIFF(19) => complement2(19), DIFF(18) => 
                           complement2(18), DIFF(17) => complement2(17), 
                           DIFF(16) => complement2(16), DIFF(15) => 
                           complement2(15), DIFF(14) => complement2(14), 
                           DIFF(13) => complement2(13), DIFF(12) => 
                           complement2(12), DIFF(11) => complement2(11), 
                           DIFF(10) => complement2(10), DIFF(9) => 
                           complement2(9), DIFF(8) => complement2(8), DIFF(7) 
                           => complement2(7), DIFF(6) => complement2(6), 
                           DIFF(5) => complement2(5), DIFF(4) => complement2(4)
                           , DIFF(3) => complement2(3), DIFF(2) => 
                           complement2(2), DIFF(1) => complement2(1), DIFF(0) 
                           => complement2(0), CO => n_3112);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_2 is

   port( input : in std_logic_vector (63 downto 0);  complement2 : out 
         std_logic_vector (63 downto 0));

end complementer_N64_2;

architecture SYN_beh of complementer_N64_2 is

   component complementer_N64_2_DW01_sub_0
      port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (63 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n2, n_3113 : std_logic;

begin
   
   n1 <= '0';
   n2 <= '0';
   sub_add_29_b0 : complementer_N64_2_DW01_sub_0 port map( A(63) => n1, A(62) 
                           => n1, A(61) => n1, A(60) => n1, A(59) => n1, A(58) 
                           => n1, A(57) => n1, A(56) => n1, A(55) => n1, A(54) 
                           => n1, A(53) => n1, A(52) => n1, A(51) => n1, A(50) 
                           => n1, A(49) => n1, A(48) => n1, A(47) => n1, A(46) 
                           => n1, A(45) => n1, A(44) => n1, A(43) => n1, A(42) 
                           => n1, A(41) => n1, A(40) => n1, A(39) => n1, A(38) 
                           => n1, A(37) => n1, A(36) => n1, A(35) => n1, A(34) 
                           => n1, A(33) => n1, A(32) => n1, A(31) => n1, A(30) 
                           => n1, A(29) => n1, A(28) => n1, A(27) => n1, A(26) 
                           => n1, A(25) => n1, A(24) => n1, A(23) => n1, A(22) 
                           => n1, A(21) => n1, A(20) => n1, A(19) => n1, A(18) 
                           => n1, A(17) => n1, A(16) => n1, A(15) => n1, A(14) 
                           => n1, A(13) => n1, A(12) => n1, A(11) => n1, A(10) 
                           => n1, A(9) => n1, A(8) => n1, A(7) => n1, A(6) => 
                           n1, A(5) => n1, A(4) => n1, A(3) => n1, A(2) => n1, 
                           A(1) => n1, A(0) => n2, B(63) => input(63), B(62) =>
                           input(62), B(61) => input(61), B(60) => input(60), 
                           B(59) => input(59), B(58) => input(58), B(57) => 
                           input(57), B(56) => input(56), B(55) => input(55), 
                           B(54) => input(54), B(53) => input(53), B(52) => 
                           input(52), B(51) => input(51), B(50) => input(50), 
                           B(49) => input(49), B(48) => input(48), B(47) => 
                           input(47), B(46) => input(46), B(45) => input(45), 
                           B(44) => input(44), B(43) => input(43), B(42) => 
                           input(42), B(41) => input(41), B(40) => input(40), 
                           B(39) => input(39), B(38) => input(38), B(37) => 
                           input(37), B(36) => input(36), B(35) => input(35), 
                           B(34) => input(34), B(33) => input(33), B(32) => 
                           input(32), B(31) => input(31), B(30) => input(30), 
                           B(29) => input(29), B(28) => input(28), B(27) => 
                           input(27), B(26) => input(26), B(25) => input(25), 
                           B(24) => input(24), B(23) => input(23), B(22) => 
                           input(22), B(21) => input(21), B(20) => input(20), 
                           B(19) => input(19), B(18) => input(18), B(17) => 
                           input(17), B(16) => input(16), B(15) => input(15), 
                           B(14) => input(14), B(13) => input(13), B(12) => 
                           input(12), B(11) => input(11), B(10) => input(10), 
                           B(9) => input(9), B(8) => input(8), B(7) => input(7)
                           , B(6) => input(6), B(5) => input(5), B(4) => 
                           input(4), B(3) => input(3), B(2) => input(2), B(1) 
                           => input(1), B(0) => input(0), CI => n1, DIFF(63) =>
                           complement2(63), DIFF(62) => complement2(62), 
                           DIFF(61) => complement2(61), DIFF(60) => 
                           complement2(60), DIFF(59) => complement2(59), 
                           DIFF(58) => complement2(58), DIFF(57) => 
                           complement2(57), DIFF(56) => complement2(56), 
                           DIFF(55) => complement2(55), DIFF(54) => 
                           complement2(54), DIFF(53) => complement2(53), 
                           DIFF(52) => complement2(52), DIFF(51) => 
                           complement2(51), DIFF(50) => complement2(50), 
                           DIFF(49) => complement2(49), DIFF(48) => 
                           complement2(48), DIFF(47) => complement2(47), 
                           DIFF(46) => complement2(46), DIFF(45) => 
                           complement2(45), DIFF(44) => complement2(44), 
                           DIFF(43) => complement2(43), DIFF(42) => 
                           complement2(42), DIFF(41) => complement2(41), 
                           DIFF(40) => complement2(40), DIFF(39) => 
                           complement2(39), DIFF(38) => complement2(38), 
                           DIFF(37) => complement2(37), DIFF(36) => 
                           complement2(36), DIFF(35) => complement2(35), 
                           DIFF(34) => complement2(34), DIFF(33) => 
                           complement2(33), DIFF(32) => complement2(32), 
                           DIFF(31) => complement2(31), DIFF(30) => 
                           complement2(30), DIFF(29) => complement2(29), 
                           DIFF(28) => complement2(28), DIFF(27) => 
                           complement2(27), DIFF(26) => complement2(26), 
                           DIFF(25) => complement2(25), DIFF(24) => 
                           complement2(24), DIFF(23) => complement2(23), 
                           DIFF(22) => complement2(22), DIFF(21) => 
                           complement2(21), DIFF(20) => complement2(20), 
                           DIFF(19) => complement2(19), DIFF(18) => 
                           complement2(18), DIFF(17) => complement2(17), 
                           DIFF(16) => complement2(16), DIFF(15) => 
                           complement2(15), DIFF(14) => complement2(14), 
                           DIFF(13) => complement2(13), DIFF(12) => 
                           complement2(12), DIFF(11) => complement2(11), 
                           DIFF(10) => complement2(10), DIFF(9) => 
                           complement2(9), DIFF(8) => complement2(8), DIFF(7) 
                           => complement2(7), DIFF(6) => complement2(6), 
                           DIFF(5) => complement2(5), DIFF(4) => complement2(4)
                           , DIFF(3) => complement2(3), DIFF(2) => 
                           complement2(2), DIFF(1) => complement2(1), DIFF(0) 
                           => complement2(0), CO => n_3113);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_3 is

   port( input : in std_logic_vector (63 downto 0);  complement2 : out 
         std_logic_vector (63 downto 0));

end complementer_N64_3;

architecture SYN_beh of complementer_N64_3 is

   component complementer_N64_3_DW01_sub_0
      port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (63 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n2, n_3114 : std_logic;

begin
   
   n1 <= '0';
   n2 <= '0';
   sub_add_29_b0 : complementer_N64_3_DW01_sub_0 port map( A(63) => n1, A(62) 
                           => n1, A(61) => n1, A(60) => n1, A(59) => n1, A(58) 
                           => n1, A(57) => n1, A(56) => n1, A(55) => n1, A(54) 
                           => n1, A(53) => n1, A(52) => n1, A(51) => n1, A(50) 
                           => n1, A(49) => n1, A(48) => n1, A(47) => n1, A(46) 
                           => n1, A(45) => n1, A(44) => n1, A(43) => n1, A(42) 
                           => n1, A(41) => n1, A(40) => n1, A(39) => n1, A(38) 
                           => n1, A(37) => n1, A(36) => n1, A(35) => n1, A(34) 
                           => n1, A(33) => n1, A(32) => n1, A(31) => n1, A(30) 
                           => n1, A(29) => n1, A(28) => n1, A(27) => n1, A(26) 
                           => n1, A(25) => n1, A(24) => n1, A(23) => n1, A(22) 
                           => n1, A(21) => n1, A(20) => n1, A(19) => n1, A(18) 
                           => n1, A(17) => n1, A(16) => n1, A(15) => n1, A(14) 
                           => n1, A(13) => n1, A(12) => n1, A(11) => n1, A(10) 
                           => n1, A(9) => n1, A(8) => n1, A(7) => n1, A(6) => 
                           n1, A(5) => n1, A(4) => n1, A(3) => n1, A(2) => n1, 
                           A(1) => n1, A(0) => n2, B(63) => input(63), B(62) =>
                           input(62), B(61) => input(61), B(60) => input(60), 
                           B(59) => input(59), B(58) => input(58), B(57) => 
                           input(57), B(56) => input(56), B(55) => input(55), 
                           B(54) => input(54), B(53) => input(53), B(52) => 
                           input(52), B(51) => input(51), B(50) => input(50), 
                           B(49) => input(49), B(48) => input(48), B(47) => 
                           input(47), B(46) => input(46), B(45) => input(45), 
                           B(44) => input(44), B(43) => input(43), B(42) => 
                           input(42), B(41) => input(41), B(40) => input(40), 
                           B(39) => input(39), B(38) => input(38), B(37) => 
                           input(37), B(36) => input(36), B(35) => input(35), 
                           B(34) => input(34), B(33) => input(33), B(32) => 
                           input(32), B(31) => input(31), B(30) => input(30), 
                           B(29) => input(29), B(28) => input(28), B(27) => 
                           input(27), B(26) => input(26), B(25) => input(25), 
                           B(24) => input(24), B(23) => input(23), B(22) => 
                           input(22), B(21) => input(21), B(20) => input(20), 
                           B(19) => input(19), B(18) => input(18), B(17) => 
                           input(17), B(16) => input(16), B(15) => input(15), 
                           B(14) => input(14), B(13) => input(13), B(12) => 
                           input(12), B(11) => input(11), B(10) => input(10), 
                           B(9) => input(9), B(8) => input(8), B(7) => input(7)
                           , B(6) => input(6), B(5) => input(5), B(4) => 
                           input(4), B(3) => input(3), B(2) => input(2), B(1) 
                           => input(1), B(0) => input(0), CI => n1, DIFF(63) =>
                           complement2(63), DIFF(62) => complement2(62), 
                           DIFF(61) => complement2(61), DIFF(60) => 
                           complement2(60), DIFF(59) => complement2(59), 
                           DIFF(58) => complement2(58), DIFF(57) => 
                           complement2(57), DIFF(56) => complement2(56), 
                           DIFF(55) => complement2(55), DIFF(54) => 
                           complement2(54), DIFF(53) => complement2(53), 
                           DIFF(52) => complement2(52), DIFF(51) => 
                           complement2(51), DIFF(50) => complement2(50), 
                           DIFF(49) => complement2(49), DIFF(48) => 
                           complement2(48), DIFF(47) => complement2(47), 
                           DIFF(46) => complement2(46), DIFF(45) => 
                           complement2(45), DIFF(44) => complement2(44), 
                           DIFF(43) => complement2(43), DIFF(42) => 
                           complement2(42), DIFF(41) => complement2(41), 
                           DIFF(40) => complement2(40), DIFF(39) => 
                           complement2(39), DIFF(38) => complement2(38), 
                           DIFF(37) => complement2(37), DIFF(36) => 
                           complement2(36), DIFF(35) => complement2(35), 
                           DIFF(34) => complement2(34), DIFF(33) => 
                           complement2(33), DIFF(32) => complement2(32), 
                           DIFF(31) => complement2(31), DIFF(30) => 
                           complement2(30), DIFF(29) => complement2(29), 
                           DIFF(28) => complement2(28), DIFF(27) => 
                           complement2(27), DIFF(26) => complement2(26), 
                           DIFF(25) => complement2(25), DIFF(24) => 
                           complement2(24), DIFF(23) => complement2(23), 
                           DIFF(22) => complement2(22), DIFF(21) => 
                           complement2(21), DIFF(20) => complement2(20), 
                           DIFF(19) => complement2(19), DIFF(18) => 
                           complement2(18), DIFF(17) => complement2(17), 
                           DIFF(16) => complement2(16), DIFF(15) => 
                           complement2(15), DIFF(14) => complement2(14), 
                           DIFF(13) => complement2(13), DIFF(12) => 
                           complement2(12), DIFF(11) => complement2(11), 
                           DIFF(10) => complement2(10), DIFF(9) => 
                           complement2(9), DIFF(8) => complement2(8), DIFF(7) 
                           => complement2(7), DIFF(6) => complement2(6), 
                           DIFF(5) => complement2(5), DIFF(4) => complement2(4)
                           , DIFF(3) => complement2(3), DIFF(2) => 
                           complement2(2), DIFF(1) => complement2(1), DIFF(0) 
                           => complement2(0), CO => n_3114);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_4 is

   port( input : in std_logic_vector (63 downto 0);  complement2 : out 
         std_logic_vector (63 downto 0));

end complementer_N64_4;

architecture SYN_beh of complementer_N64_4 is

   component complementer_N64_4_DW01_sub_0
      port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (63 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n2, n_3115 : std_logic;

begin
   
   n1 <= '0';
   n2 <= '0';
   sub_add_29_b0 : complementer_N64_4_DW01_sub_0 port map( A(63) => n1, A(62) 
                           => n1, A(61) => n1, A(60) => n1, A(59) => n1, A(58) 
                           => n1, A(57) => n1, A(56) => n1, A(55) => n1, A(54) 
                           => n1, A(53) => n1, A(52) => n1, A(51) => n1, A(50) 
                           => n1, A(49) => n1, A(48) => n1, A(47) => n1, A(46) 
                           => n1, A(45) => n1, A(44) => n1, A(43) => n1, A(42) 
                           => n1, A(41) => n1, A(40) => n1, A(39) => n1, A(38) 
                           => n1, A(37) => n1, A(36) => n1, A(35) => n1, A(34) 
                           => n1, A(33) => n1, A(32) => n1, A(31) => n1, A(30) 
                           => n1, A(29) => n1, A(28) => n1, A(27) => n1, A(26) 
                           => n1, A(25) => n1, A(24) => n1, A(23) => n1, A(22) 
                           => n1, A(21) => n1, A(20) => n1, A(19) => n1, A(18) 
                           => n1, A(17) => n1, A(16) => n1, A(15) => n1, A(14) 
                           => n1, A(13) => n1, A(12) => n1, A(11) => n1, A(10) 
                           => n1, A(9) => n1, A(8) => n1, A(7) => n1, A(6) => 
                           n1, A(5) => n1, A(4) => n1, A(3) => n1, A(2) => n1, 
                           A(1) => n1, A(0) => n2, B(63) => input(63), B(62) =>
                           input(62), B(61) => input(61), B(60) => input(60), 
                           B(59) => input(59), B(58) => input(58), B(57) => 
                           input(57), B(56) => input(56), B(55) => input(55), 
                           B(54) => input(54), B(53) => input(53), B(52) => 
                           input(52), B(51) => input(51), B(50) => input(50), 
                           B(49) => input(49), B(48) => input(48), B(47) => 
                           input(47), B(46) => input(46), B(45) => input(45), 
                           B(44) => input(44), B(43) => input(43), B(42) => 
                           input(42), B(41) => input(41), B(40) => input(40), 
                           B(39) => input(39), B(38) => input(38), B(37) => 
                           input(37), B(36) => input(36), B(35) => input(35), 
                           B(34) => input(34), B(33) => input(33), B(32) => 
                           input(32), B(31) => input(31), B(30) => input(30), 
                           B(29) => input(29), B(28) => input(28), B(27) => 
                           input(27), B(26) => input(26), B(25) => input(25), 
                           B(24) => input(24), B(23) => input(23), B(22) => 
                           input(22), B(21) => input(21), B(20) => input(20), 
                           B(19) => input(19), B(18) => input(18), B(17) => 
                           input(17), B(16) => input(16), B(15) => input(15), 
                           B(14) => input(14), B(13) => input(13), B(12) => 
                           input(12), B(11) => input(11), B(10) => input(10), 
                           B(9) => input(9), B(8) => input(8), B(7) => input(7)
                           , B(6) => input(6), B(5) => input(5), B(4) => 
                           input(4), B(3) => input(3), B(2) => input(2), B(1) 
                           => input(1), B(0) => input(0), CI => n1, DIFF(63) =>
                           complement2(63), DIFF(62) => complement2(62), 
                           DIFF(61) => complement2(61), DIFF(60) => 
                           complement2(60), DIFF(59) => complement2(59), 
                           DIFF(58) => complement2(58), DIFF(57) => 
                           complement2(57), DIFF(56) => complement2(56), 
                           DIFF(55) => complement2(55), DIFF(54) => 
                           complement2(54), DIFF(53) => complement2(53), 
                           DIFF(52) => complement2(52), DIFF(51) => 
                           complement2(51), DIFF(50) => complement2(50), 
                           DIFF(49) => complement2(49), DIFF(48) => 
                           complement2(48), DIFF(47) => complement2(47), 
                           DIFF(46) => complement2(46), DIFF(45) => 
                           complement2(45), DIFF(44) => complement2(44), 
                           DIFF(43) => complement2(43), DIFF(42) => 
                           complement2(42), DIFF(41) => complement2(41), 
                           DIFF(40) => complement2(40), DIFF(39) => 
                           complement2(39), DIFF(38) => complement2(38), 
                           DIFF(37) => complement2(37), DIFF(36) => 
                           complement2(36), DIFF(35) => complement2(35), 
                           DIFF(34) => complement2(34), DIFF(33) => 
                           complement2(33), DIFF(32) => complement2(32), 
                           DIFF(31) => complement2(31), DIFF(30) => 
                           complement2(30), DIFF(29) => complement2(29), 
                           DIFF(28) => complement2(28), DIFF(27) => 
                           complement2(27), DIFF(26) => complement2(26), 
                           DIFF(25) => complement2(25), DIFF(24) => 
                           complement2(24), DIFF(23) => complement2(23), 
                           DIFF(22) => complement2(22), DIFF(21) => 
                           complement2(21), DIFF(20) => complement2(20), 
                           DIFF(19) => complement2(19), DIFF(18) => 
                           complement2(18), DIFF(17) => complement2(17), 
                           DIFF(16) => complement2(16), DIFF(15) => 
                           complement2(15), DIFF(14) => complement2(14), 
                           DIFF(13) => complement2(13), DIFF(12) => 
                           complement2(12), DIFF(11) => complement2(11), 
                           DIFF(10) => complement2(10), DIFF(9) => 
                           complement2(9), DIFF(8) => complement2(8), DIFF(7) 
                           => complement2(7), DIFF(6) => complement2(6), 
                           DIFF(5) => complement2(5), DIFF(4) => complement2(4)
                           , DIFF(3) => complement2(3), DIFF(2) => 
                           complement2(2), DIFF(1) => complement2(1), DIFF(0) 
                           => complement2(0), CO => n_3115);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_5 is

   port( input : in std_logic_vector (63 downto 0);  complement2 : out 
         std_logic_vector (63 downto 0));

end complementer_N64_5;

architecture SYN_beh of complementer_N64_5 is

   component complementer_N64_5_DW01_sub_0
      port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (63 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n2, n_3116 : std_logic;

begin
   
   n1 <= '0';
   n2 <= '0';
   sub_add_29_b0 : complementer_N64_5_DW01_sub_0 port map( A(63) => n1, A(62) 
                           => n1, A(61) => n1, A(60) => n1, A(59) => n1, A(58) 
                           => n1, A(57) => n1, A(56) => n1, A(55) => n1, A(54) 
                           => n1, A(53) => n1, A(52) => n1, A(51) => n1, A(50) 
                           => n1, A(49) => n1, A(48) => n1, A(47) => n1, A(46) 
                           => n1, A(45) => n1, A(44) => n1, A(43) => n1, A(42) 
                           => n1, A(41) => n1, A(40) => n1, A(39) => n1, A(38) 
                           => n1, A(37) => n1, A(36) => n1, A(35) => n1, A(34) 
                           => n1, A(33) => n1, A(32) => n1, A(31) => n1, A(30) 
                           => n1, A(29) => n1, A(28) => n1, A(27) => n1, A(26) 
                           => n1, A(25) => n1, A(24) => n1, A(23) => n1, A(22) 
                           => n1, A(21) => n1, A(20) => n1, A(19) => n1, A(18) 
                           => n1, A(17) => n1, A(16) => n1, A(15) => n1, A(14) 
                           => n1, A(13) => n1, A(12) => n1, A(11) => n1, A(10) 
                           => n1, A(9) => n1, A(8) => n1, A(7) => n1, A(6) => 
                           n1, A(5) => n1, A(4) => n1, A(3) => n1, A(2) => n1, 
                           A(1) => n1, A(0) => n2, B(63) => input(63), B(62) =>
                           input(62), B(61) => input(61), B(60) => input(60), 
                           B(59) => input(59), B(58) => input(58), B(57) => 
                           input(57), B(56) => input(56), B(55) => input(55), 
                           B(54) => input(54), B(53) => input(53), B(52) => 
                           input(52), B(51) => input(51), B(50) => input(50), 
                           B(49) => input(49), B(48) => input(48), B(47) => 
                           input(47), B(46) => input(46), B(45) => input(45), 
                           B(44) => input(44), B(43) => input(43), B(42) => 
                           input(42), B(41) => input(41), B(40) => input(40), 
                           B(39) => input(39), B(38) => input(38), B(37) => 
                           input(37), B(36) => input(36), B(35) => input(35), 
                           B(34) => input(34), B(33) => input(33), B(32) => 
                           input(32), B(31) => input(31), B(30) => input(30), 
                           B(29) => input(29), B(28) => input(28), B(27) => 
                           input(27), B(26) => input(26), B(25) => input(25), 
                           B(24) => input(24), B(23) => input(23), B(22) => 
                           input(22), B(21) => input(21), B(20) => input(20), 
                           B(19) => input(19), B(18) => input(18), B(17) => 
                           input(17), B(16) => input(16), B(15) => input(15), 
                           B(14) => input(14), B(13) => input(13), B(12) => 
                           input(12), B(11) => input(11), B(10) => input(10), 
                           B(9) => input(9), B(8) => input(8), B(7) => input(7)
                           , B(6) => input(6), B(5) => input(5), B(4) => 
                           input(4), B(3) => input(3), B(2) => input(2), B(1) 
                           => input(1), B(0) => input(0), CI => n1, DIFF(63) =>
                           complement2(63), DIFF(62) => complement2(62), 
                           DIFF(61) => complement2(61), DIFF(60) => 
                           complement2(60), DIFF(59) => complement2(59), 
                           DIFF(58) => complement2(58), DIFF(57) => 
                           complement2(57), DIFF(56) => complement2(56), 
                           DIFF(55) => complement2(55), DIFF(54) => 
                           complement2(54), DIFF(53) => complement2(53), 
                           DIFF(52) => complement2(52), DIFF(51) => 
                           complement2(51), DIFF(50) => complement2(50), 
                           DIFF(49) => complement2(49), DIFF(48) => 
                           complement2(48), DIFF(47) => complement2(47), 
                           DIFF(46) => complement2(46), DIFF(45) => 
                           complement2(45), DIFF(44) => complement2(44), 
                           DIFF(43) => complement2(43), DIFF(42) => 
                           complement2(42), DIFF(41) => complement2(41), 
                           DIFF(40) => complement2(40), DIFF(39) => 
                           complement2(39), DIFF(38) => complement2(38), 
                           DIFF(37) => complement2(37), DIFF(36) => 
                           complement2(36), DIFF(35) => complement2(35), 
                           DIFF(34) => complement2(34), DIFF(33) => 
                           complement2(33), DIFF(32) => complement2(32), 
                           DIFF(31) => complement2(31), DIFF(30) => 
                           complement2(30), DIFF(29) => complement2(29), 
                           DIFF(28) => complement2(28), DIFF(27) => 
                           complement2(27), DIFF(26) => complement2(26), 
                           DIFF(25) => complement2(25), DIFF(24) => 
                           complement2(24), DIFF(23) => complement2(23), 
                           DIFF(22) => complement2(22), DIFF(21) => 
                           complement2(21), DIFF(20) => complement2(20), 
                           DIFF(19) => complement2(19), DIFF(18) => 
                           complement2(18), DIFF(17) => complement2(17), 
                           DIFF(16) => complement2(16), DIFF(15) => 
                           complement2(15), DIFF(14) => complement2(14), 
                           DIFF(13) => complement2(13), DIFF(12) => 
                           complement2(12), DIFF(11) => complement2(11), 
                           DIFF(10) => complement2(10), DIFF(9) => 
                           complement2(9), DIFF(8) => complement2(8), DIFF(7) 
                           => complement2(7), DIFF(6) => complement2(6), 
                           DIFF(5) => complement2(5), DIFF(4) => complement2(4)
                           , DIFF(3) => complement2(3), DIFF(2) => 
                           complement2(2), DIFF(1) => complement2(1), DIFF(0) 
                           => complement2(0), CO => n_3116);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_6 is

   port( input : in std_logic_vector (63 downto 0);  complement2 : out 
         std_logic_vector (63 downto 0));

end complementer_N64_6;

architecture SYN_beh of complementer_N64_6 is

   component complementer_N64_6_DW01_sub_0
      port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (63 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n2, n_3117 : std_logic;

begin
   
   n1 <= '0';
   n2 <= '0';
   sub_add_29_b0 : complementer_N64_6_DW01_sub_0 port map( A(63) => n1, A(62) 
                           => n1, A(61) => n1, A(60) => n1, A(59) => n1, A(58) 
                           => n1, A(57) => n1, A(56) => n1, A(55) => n1, A(54) 
                           => n1, A(53) => n1, A(52) => n1, A(51) => n1, A(50) 
                           => n1, A(49) => n1, A(48) => n1, A(47) => n1, A(46) 
                           => n1, A(45) => n1, A(44) => n1, A(43) => n1, A(42) 
                           => n1, A(41) => n1, A(40) => n1, A(39) => n1, A(38) 
                           => n1, A(37) => n1, A(36) => n1, A(35) => n1, A(34) 
                           => n1, A(33) => n1, A(32) => n1, A(31) => n1, A(30) 
                           => n1, A(29) => n1, A(28) => n1, A(27) => n1, A(26) 
                           => n1, A(25) => n1, A(24) => n1, A(23) => n1, A(22) 
                           => n1, A(21) => n1, A(20) => n1, A(19) => n1, A(18) 
                           => n1, A(17) => n1, A(16) => n1, A(15) => n1, A(14) 
                           => n1, A(13) => n1, A(12) => n1, A(11) => n1, A(10) 
                           => n1, A(9) => n1, A(8) => n1, A(7) => n1, A(6) => 
                           n1, A(5) => n1, A(4) => n1, A(3) => n1, A(2) => n1, 
                           A(1) => n1, A(0) => n2, B(63) => input(63), B(62) =>
                           input(62), B(61) => input(61), B(60) => input(60), 
                           B(59) => input(59), B(58) => input(58), B(57) => 
                           input(57), B(56) => input(56), B(55) => input(55), 
                           B(54) => input(54), B(53) => input(53), B(52) => 
                           input(52), B(51) => input(51), B(50) => input(50), 
                           B(49) => input(49), B(48) => input(48), B(47) => 
                           input(47), B(46) => input(46), B(45) => input(45), 
                           B(44) => input(44), B(43) => input(43), B(42) => 
                           input(42), B(41) => input(41), B(40) => input(40), 
                           B(39) => input(39), B(38) => input(38), B(37) => 
                           input(37), B(36) => input(36), B(35) => input(35), 
                           B(34) => input(34), B(33) => input(33), B(32) => 
                           input(32), B(31) => input(31), B(30) => input(30), 
                           B(29) => input(29), B(28) => input(28), B(27) => 
                           input(27), B(26) => input(26), B(25) => input(25), 
                           B(24) => input(24), B(23) => input(23), B(22) => 
                           input(22), B(21) => input(21), B(20) => input(20), 
                           B(19) => input(19), B(18) => input(18), B(17) => 
                           input(17), B(16) => input(16), B(15) => input(15), 
                           B(14) => input(14), B(13) => input(13), B(12) => 
                           input(12), B(11) => input(11), B(10) => input(10), 
                           B(9) => input(9), B(8) => input(8), B(7) => input(7)
                           , B(6) => input(6), B(5) => input(5), B(4) => 
                           input(4), B(3) => input(3), B(2) => input(2), B(1) 
                           => input(1), B(0) => input(0), CI => n1, DIFF(63) =>
                           complement2(63), DIFF(62) => complement2(62), 
                           DIFF(61) => complement2(61), DIFF(60) => 
                           complement2(60), DIFF(59) => complement2(59), 
                           DIFF(58) => complement2(58), DIFF(57) => 
                           complement2(57), DIFF(56) => complement2(56), 
                           DIFF(55) => complement2(55), DIFF(54) => 
                           complement2(54), DIFF(53) => complement2(53), 
                           DIFF(52) => complement2(52), DIFF(51) => 
                           complement2(51), DIFF(50) => complement2(50), 
                           DIFF(49) => complement2(49), DIFF(48) => 
                           complement2(48), DIFF(47) => complement2(47), 
                           DIFF(46) => complement2(46), DIFF(45) => 
                           complement2(45), DIFF(44) => complement2(44), 
                           DIFF(43) => complement2(43), DIFF(42) => 
                           complement2(42), DIFF(41) => complement2(41), 
                           DIFF(40) => complement2(40), DIFF(39) => 
                           complement2(39), DIFF(38) => complement2(38), 
                           DIFF(37) => complement2(37), DIFF(36) => 
                           complement2(36), DIFF(35) => complement2(35), 
                           DIFF(34) => complement2(34), DIFF(33) => 
                           complement2(33), DIFF(32) => complement2(32), 
                           DIFF(31) => complement2(31), DIFF(30) => 
                           complement2(30), DIFF(29) => complement2(29), 
                           DIFF(28) => complement2(28), DIFF(27) => 
                           complement2(27), DIFF(26) => complement2(26), 
                           DIFF(25) => complement2(25), DIFF(24) => 
                           complement2(24), DIFF(23) => complement2(23), 
                           DIFF(22) => complement2(22), DIFF(21) => 
                           complement2(21), DIFF(20) => complement2(20), 
                           DIFF(19) => complement2(19), DIFF(18) => 
                           complement2(18), DIFF(17) => complement2(17), 
                           DIFF(16) => complement2(16), DIFF(15) => 
                           complement2(15), DIFF(14) => complement2(14), 
                           DIFF(13) => complement2(13), DIFF(12) => 
                           complement2(12), DIFF(11) => complement2(11), 
                           DIFF(10) => complement2(10), DIFF(9) => 
                           complement2(9), DIFF(8) => complement2(8), DIFF(7) 
                           => complement2(7), DIFF(6) => complement2(6), 
                           DIFF(5) => complement2(5), DIFF(4) => complement2(4)
                           , DIFF(3) => complement2(3), DIFF(2) => 
                           complement2(2), DIFF(1) => complement2(1), DIFF(0) 
                           => complement2(0), CO => n_3117);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_7 is

   port( input : in std_logic_vector (63 downto 0);  complement2 : out 
         std_logic_vector (63 downto 0));

end complementer_N64_7;

architecture SYN_beh of complementer_N64_7 is

   component complementer_N64_7_DW01_sub_0
      port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (63 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n2, n_3118 : std_logic;

begin
   
   n1 <= '0';
   n2 <= '0';
   sub_add_29_b0 : complementer_N64_7_DW01_sub_0 port map( A(63) => n1, A(62) 
                           => n1, A(61) => n1, A(60) => n1, A(59) => n1, A(58) 
                           => n1, A(57) => n1, A(56) => n1, A(55) => n1, A(54) 
                           => n1, A(53) => n1, A(52) => n1, A(51) => n1, A(50) 
                           => n1, A(49) => n1, A(48) => n1, A(47) => n1, A(46) 
                           => n1, A(45) => n1, A(44) => n1, A(43) => n1, A(42) 
                           => n1, A(41) => n1, A(40) => n1, A(39) => n1, A(38) 
                           => n1, A(37) => n1, A(36) => n1, A(35) => n1, A(34) 
                           => n1, A(33) => n1, A(32) => n1, A(31) => n1, A(30) 
                           => n1, A(29) => n1, A(28) => n1, A(27) => n1, A(26) 
                           => n1, A(25) => n1, A(24) => n1, A(23) => n1, A(22) 
                           => n1, A(21) => n1, A(20) => n1, A(19) => n1, A(18) 
                           => n1, A(17) => n1, A(16) => n1, A(15) => n1, A(14) 
                           => n1, A(13) => n1, A(12) => n1, A(11) => n1, A(10) 
                           => n1, A(9) => n1, A(8) => n1, A(7) => n1, A(6) => 
                           n1, A(5) => n1, A(4) => n1, A(3) => n1, A(2) => n1, 
                           A(1) => n1, A(0) => n2, B(63) => input(63), B(62) =>
                           input(62), B(61) => input(61), B(60) => input(60), 
                           B(59) => input(59), B(58) => input(58), B(57) => 
                           input(57), B(56) => input(56), B(55) => input(55), 
                           B(54) => input(54), B(53) => input(53), B(52) => 
                           input(52), B(51) => input(51), B(50) => input(50), 
                           B(49) => input(49), B(48) => input(48), B(47) => 
                           input(47), B(46) => input(46), B(45) => input(45), 
                           B(44) => input(44), B(43) => input(43), B(42) => 
                           input(42), B(41) => input(41), B(40) => input(40), 
                           B(39) => input(39), B(38) => input(38), B(37) => 
                           input(37), B(36) => input(36), B(35) => input(35), 
                           B(34) => input(34), B(33) => input(33), B(32) => 
                           input(32), B(31) => input(31), B(30) => input(30), 
                           B(29) => input(29), B(28) => input(28), B(27) => 
                           input(27), B(26) => input(26), B(25) => input(25), 
                           B(24) => input(24), B(23) => input(23), B(22) => 
                           input(22), B(21) => input(21), B(20) => input(20), 
                           B(19) => input(19), B(18) => input(18), B(17) => 
                           input(17), B(16) => input(16), B(15) => input(15), 
                           B(14) => input(14), B(13) => input(13), B(12) => 
                           input(12), B(11) => input(11), B(10) => input(10), 
                           B(9) => input(9), B(8) => input(8), B(7) => input(7)
                           , B(6) => input(6), B(5) => input(5), B(4) => 
                           input(4), B(3) => input(3), B(2) => input(2), B(1) 
                           => input(1), B(0) => input(0), CI => n1, DIFF(63) =>
                           complement2(63), DIFF(62) => complement2(62), 
                           DIFF(61) => complement2(61), DIFF(60) => 
                           complement2(60), DIFF(59) => complement2(59), 
                           DIFF(58) => complement2(58), DIFF(57) => 
                           complement2(57), DIFF(56) => complement2(56), 
                           DIFF(55) => complement2(55), DIFF(54) => 
                           complement2(54), DIFF(53) => complement2(53), 
                           DIFF(52) => complement2(52), DIFF(51) => 
                           complement2(51), DIFF(50) => complement2(50), 
                           DIFF(49) => complement2(49), DIFF(48) => 
                           complement2(48), DIFF(47) => complement2(47), 
                           DIFF(46) => complement2(46), DIFF(45) => 
                           complement2(45), DIFF(44) => complement2(44), 
                           DIFF(43) => complement2(43), DIFF(42) => 
                           complement2(42), DIFF(41) => complement2(41), 
                           DIFF(40) => complement2(40), DIFF(39) => 
                           complement2(39), DIFF(38) => complement2(38), 
                           DIFF(37) => complement2(37), DIFF(36) => 
                           complement2(36), DIFF(35) => complement2(35), 
                           DIFF(34) => complement2(34), DIFF(33) => 
                           complement2(33), DIFF(32) => complement2(32), 
                           DIFF(31) => complement2(31), DIFF(30) => 
                           complement2(30), DIFF(29) => complement2(29), 
                           DIFF(28) => complement2(28), DIFF(27) => 
                           complement2(27), DIFF(26) => complement2(26), 
                           DIFF(25) => complement2(25), DIFF(24) => 
                           complement2(24), DIFF(23) => complement2(23), 
                           DIFF(22) => complement2(22), DIFF(21) => 
                           complement2(21), DIFF(20) => complement2(20), 
                           DIFF(19) => complement2(19), DIFF(18) => 
                           complement2(18), DIFF(17) => complement2(17), 
                           DIFF(16) => complement2(16), DIFF(15) => 
                           complement2(15), DIFF(14) => complement2(14), 
                           DIFF(13) => complement2(13), DIFF(12) => 
                           complement2(12), DIFF(11) => complement2(11), 
                           DIFF(10) => complement2(10), DIFF(9) => 
                           complement2(9), DIFF(8) => complement2(8), DIFF(7) 
                           => complement2(7), DIFF(6) => complement2(6), 
                           DIFF(5) => complement2(5), DIFF(4) => complement2(4)
                           , DIFF(3) => complement2(3), DIFF(2) => 
                           complement2(2), DIFF(1) => complement2(1), DIFF(0) 
                           => complement2(0), CO => n_3118);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_8 is

   port( input : in std_logic_vector (63 downto 0);  complement2 : out 
         std_logic_vector (63 downto 0));

end complementer_N64_8;

architecture SYN_beh of complementer_N64_8 is

   component complementer_N64_8_DW01_sub_0
      port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (63 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n2, n_3119 : std_logic;

begin
   
   n1 <= '0';
   n2 <= '0';
   sub_add_29_b0 : complementer_N64_8_DW01_sub_0 port map( A(63) => n1, A(62) 
                           => n1, A(61) => n1, A(60) => n1, A(59) => n1, A(58) 
                           => n1, A(57) => n1, A(56) => n1, A(55) => n1, A(54) 
                           => n1, A(53) => n1, A(52) => n1, A(51) => n1, A(50) 
                           => n1, A(49) => n1, A(48) => n1, A(47) => n1, A(46) 
                           => n1, A(45) => n1, A(44) => n1, A(43) => n1, A(42) 
                           => n1, A(41) => n1, A(40) => n1, A(39) => n1, A(38) 
                           => n1, A(37) => n1, A(36) => n1, A(35) => n1, A(34) 
                           => n1, A(33) => n1, A(32) => n1, A(31) => n1, A(30) 
                           => n1, A(29) => n1, A(28) => n1, A(27) => n1, A(26) 
                           => n1, A(25) => n1, A(24) => n1, A(23) => n1, A(22) 
                           => n1, A(21) => n1, A(20) => n1, A(19) => n1, A(18) 
                           => n1, A(17) => n1, A(16) => n1, A(15) => n1, A(14) 
                           => n1, A(13) => n1, A(12) => n1, A(11) => n1, A(10) 
                           => n1, A(9) => n1, A(8) => n1, A(7) => n1, A(6) => 
                           n1, A(5) => n1, A(4) => n1, A(3) => n1, A(2) => n1, 
                           A(1) => n1, A(0) => n2, B(63) => input(63), B(62) =>
                           input(62), B(61) => input(61), B(60) => input(60), 
                           B(59) => input(59), B(58) => input(58), B(57) => 
                           input(57), B(56) => input(56), B(55) => input(55), 
                           B(54) => input(54), B(53) => input(53), B(52) => 
                           input(52), B(51) => input(51), B(50) => input(50), 
                           B(49) => input(49), B(48) => input(48), B(47) => 
                           input(47), B(46) => input(46), B(45) => input(45), 
                           B(44) => input(44), B(43) => input(43), B(42) => 
                           input(42), B(41) => input(41), B(40) => input(40), 
                           B(39) => input(39), B(38) => input(38), B(37) => 
                           input(37), B(36) => input(36), B(35) => input(35), 
                           B(34) => input(34), B(33) => input(33), B(32) => 
                           input(32), B(31) => input(31), B(30) => input(30), 
                           B(29) => input(29), B(28) => input(28), B(27) => 
                           input(27), B(26) => input(26), B(25) => input(25), 
                           B(24) => input(24), B(23) => input(23), B(22) => 
                           input(22), B(21) => input(21), B(20) => input(20), 
                           B(19) => input(19), B(18) => input(18), B(17) => 
                           input(17), B(16) => input(16), B(15) => input(15), 
                           B(14) => input(14), B(13) => input(13), B(12) => 
                           input(12), B(11) => input(11), B(10) => input(10), 
                           B(9) => input(9), B(8) => input(8), B(7) => input(7)
                           , B(6) => input(6), B(5) => input(5), B(4) => 
                           input(4), B(3) => input(3), B(2) => input(2), B(1) 
                           => input(1), B(0) => input(0), CI => n1, DIFF(63) =>
                           complement2(63), DIFF(62) => complement2(62), 
                           DIFF(61) => complement2(61), DIFF(60) => 
                           complement2(60), DIFF(59) => complement2(59), 
                           DIFF(58) => complement2(58), DIFF(57) => 
                           complement2(57), DIFF(56) => complement2(56), 
                           DIFF(55) => complement2(55), DIFF(54) => 
                           complement2(54), DIFF(53) => complement2(53), 
                           DIFF(52) => complement2(52), DIFF(51) => 
                           complement2(51), DIFF(50) => complement2(50), 
                           DIFF(49) => complement2(49), DIFF(48) => 
                           complement2(48), DIFF(47) => complement2(47), 
                           DIFF(46) => complement2(46), DIFF(45) => 
                           complement2(45), DIFF(44) => complement2(44), 
                           DIFF(43) => complement2(43), DIFF(42) => 
                           complement2(42), DIFF(41) => complement2(41), 
                           DIFF(40) => complement2(40), DIFF(39) => 
                           complement2(39), DIFF(38) => complement2(38), 
                           DIFF(37) => complement2(37), DIFF(36) => 
                           complement2(36), DIFF(35) => complement2(35), 
                           DIFF(34) => complement2(34), DIFF(33) => 
                           complement2(33), DIFF(32) => complement2(32), 
                           DIFF(31) => complement2(31), DIFF(30) => 
                           complement2(30), DIFF(29) => complement2(29), 
                           DIFF(28) => complement2(28), DIFF(27) => 
                           complement2(27), DIFF(26) => complement2(26), 
                           DIFF(25) => complement2(25), DIFF(24) => 
                           complement2(24), DIFF(23) => complement2(23), 
                           DIFF(22) => complement2(22), DIFF(21) => 
                           complement2(21), DIFF(20) => complement2(20), 
                           DIFF(19) => complement2(19), DIFF(18) => 
                           complement2(18), DIFF(17) => complement2(17), 
                           DIFF(16) => complement2(16), DIFF(15) => 
                           complement2(15), DIFF(14) => complement2(14), 
                           DIFF(13) => complement2(13), DIFF(12) => 
                           complement2(12), DIFF(11) => complement2(11), 
                           DIFF(10) => complement2(10), DIFF(9) => 
                           complement2(9), DIFF(8) => complement2(8), DIFF(7) 
                           => complement2(7), DIFF(6) => complement2(6), 
                           DIFF(5) => complement2(5), DIFF(4) => complement2(4)
                           , DIFF(3) => complement2(3), DIFF(2) => 
                           complement2(2), DIFF(1) => complement2(1), DIFF(0) 
                           => complement2(0), CO => n_3119);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_9 is

   port( input : in std_logic_vector (63 downto 0);  complement2 : out 
         std_logic_vector (63 downto 0));

end complementer_N64_9;

architecture SYN_beh of complementer_N64_9 is

   component complementer_N64_9_DW01_sub_0
      port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (63 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n2, n_3120 : std_logic;

begin
   
   n1 <= '0';
   n2 <= '0';
   sub_add_29_b0 : complementer_N64_9_DW01_sub_0 port map( A(63) => n1, A(62) 
                           => n1, A(61) => n1, A(60) => n1, A(59) => n1, A(58) 
                           => n1, A(57) => n1, A(56) => n1, A(55) => n1, A(54) 
                           => n1, A(53) => n1, A(52) => n1, A(51) => n1, A(50) 
                           => n1, A(49) => n1, A(48) => n1, A(47) => n1, A(46) 
                           => n1, A(45) => n1, A(44) => n1, A(43) => n1, A(42) 
                           => n1, A(41) => n1, A(40) => n1, A(39) => n1, A(38) 
                           => n1, A(37) => n1, A(36) => n1, A(35) => n1, A(34) 
                           => n1, A(33) => n1, A(32) => n1, A(31) => n1, A(30) 
                           => n1, A(29) => n1, A(28) => n1, A(27) => n1, A(26) 
                           => n1, A(25) => n1, A(24) => n1, A(23) => n1, A(22) 
                           => n1, A(21) => n1, A(20) => n1, A(19) => n1, A(18) 
                           => n1, A(17) => n1, A(16) => n1, A(15) => n1, A(14) 
                           => n1, A(13) => n1, A(12) => n1, A(11) => n1, A(10) 
                           => n1, A(9) => n1, A(8) => n1, A(7) => n1, A(6) => 
                           n1, A(5) => n1, A(4) => n1, A(3) => n1, A(2) => n1, 
                           A(1) => n1, A(0) => n2, B(63) => input(63), B(62) =>
                           input(62), B(61) => input(61), B(60) => input(60), 
                           B(59) => input(59), B(58) => input(58), B(57) => 
                           input(57), B(56) => input(56), B(55) => input(55), 
                           B(54) => input(54), B(53) => input(53), B(52) => 
                           input(52), B(51) => input(51), B(50) => input(50), 
                           B(49) => input(49), B(48) => input(48), B(47) => 
                           input(47), B(46) => input(46), B(45) => input(45), 
                           B(44) => input(44), B(43) => input(43), B(42) => 
                           input(42), B(41) => input(41), B(40) => input(40), 
                           B(39) => input(39), B(38) => input(38), B(37) => 
                           input(37), B(36) => input(36), B(35) => input(35), 
                           B(34) => input(34), B(33) => input(33), B(32) => 
                           input(32), B(31) => input(31), B(30) => input(30), 
                           B(29) => input(29), B(28) => input(28), B(27) => 
                           input(27), B(26) => input(26), B(25) => input(25), 
                           B(24) => input(24), B(23) => input(23), B(22) => 
                           input(22), B(21) => input(21), B(20) => input(20), 
                           B(19) => input(19), B(18) => input(18), B(17) => 
                           input(17), B(16) => input(16), B(15) => input(15), 
                           B(14) => input(14), B(13) => input(13), B(12) => 
                           input(12), B(11) => input(11), B(10) => input(10), 
                           B(9) => input(9), B(8) => input(8), B(7) => input(7)
                           , B(6) => input(6), B(5) => input(5), B(4) => 
                           input(4), B(3) => input(3), B(2) => input(2), B(1) 
                           => input(1), B(0) => input(0), CI => n1, DIFF(63) =>
                           complement2(63), DIFF(62) => complement2(62), 
                           DIFF(61) => complement2(61), DIFF(60) => 
                           complement2(60), DIFF(59) => complement2(59), 
                           DIFF(58) => complement2(58), DIFF(57) => 
                           complement2(57), DIFF(56) => complement2(56), 
                           DIFF(55) => complement2(55), DIFF(54) => 
                           complement2(54), DIFF(53) => complement2(53), 
                           DIFF(52) => complement2(52), DIFF(51) => 
                           complement2(51), DIFF(50) => complement2(50), 
                           DIFF(49) => complement2(49), DIFF(48) => 
                           complement2(48), DIFF(47) => complement2(47), 
                           DIFF(46) => complement2(46), DIFF(45) => 
                           complement2(45), DIFF(44) => complement2(44), 
                           DIFF(43) => complement2(43), DIFF(42) => 
                           complement2(42), DIFF(41) => complement2(41), 
                           DIFF(40) => complement2(40), DIFF(39) => 
                           complement2(39), DIFF(38) => complement2(38), 
                           DIFF(37) => complement2(37), DIFF(36) => 
                           complement2(36), DIFF(35) => complement2(35), 
                           DIFF(34) => complement2(34), DIFF(33) => 
                           complement2(33), DIFF(32) => complement2(32), 
                           DIFF(31) => complement2(31), DIFF(30) => 
                           complement2(30), DIFF(29) => complement2(29), 
                           DIFF(28) => complement2(28), DIFF(27) => 
                           complement2(27), DIFF(26) => complement2(26), 
                           DIFF(25) => complement2(25), DIFF(24) => 
                           complement2(24), DIFF(23) => complement2(23), 
                           DIFF(22) => complement2(22), DIFF(21) => 
                           complement2(21), DIFF(20) => complement2(20), 
                           DIFF(19) => complement2(19), DIFF(18) => 
                           complement2(18), DIFF(17) => complement2(17), 
                           DIFF(16) => complement2(16), DIFF(15) => 
                           complement2(15), DIFF(14) => complement2(14), 
                           DIFF(13) => complement2(13), DIFF(12) => 
                           complement2(12), DIFF(11) => complement2(11), 
                           DIFF(10) => complement2(10), DIFF(9) => 
                           complement2(9), DIFF(8) => complement2(8), DIFF(7) 
                           => complement2(7), DIFF(6) => complement2(6), 
                           DIFF(5) => complement2(5), DIFF(4) => complement2(4)
                           , DIFF(3) => complement2(3), DIFF(2) => 
                           complement2(2), DIFF(1) => complement2(1), DIFF(0) 
                           => complement2(0), CO => n_3120);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_10 is

   port( input : in std_logic_vector (63 downto 0);  complement2 : out 
         std_logic_vector (63 downto 0));

end complementer_N64_10;

architecture SYN_beh of complementer_N64_10 is

   component complementer_N64_10_DW01_sub_0
      port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (63 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n2, n_3121 : std_logic;

begin
   
   n1 <= '0';
   n2 <= '0';
   sub_add_29_b0 : complementer_N64_10_DW01_sub_0 port map( A(63) => n1, A(62) 
                           => n1, A(61) => n1, A(60) => n1, A(59) => n1, A(58) 
                           => n1, A(57) => n1, A(56) => n1, A(55) => n1, A(54) 
                           => n1, A(53) => n1, A(52) => n1, A(51) => n1, A(50) 
                           => n1, A(49) => n1, A(48) => n1, A(47) => n1, A(46) 
                           => n1, A(45) => n1, A(44) => n1, A(43) => n1, A(42) 
                           => n1, A(41) => n1, A(40) => n1, A(39) => n1, A(38) 
                           => n1, A(37) => n1, A(36) => n1, A(35) => n1, A(34) 
                           => n1, A(33) => n1, A(32) => n1, A(31) => n1, A(30) 
                           => n1, A(29) => n1, A(28) => n1, A(27) => n1, A(26) 
                           => n1, A(25) => n1, A(24) => n1, A(23) => n1, A(22) 
                           => n1, A(21) => n1, A(20) => n1, A(19) => n1, A(18) 
                           => n1, A(17) => n1, A(16) => n1, A(15) => n1, A(14) 
                           => n1, A(13) => n1, A(12) => n1, A(11) => n1, A(10) 
                           => n1, A(9) => n1, A(8) => n1, A(7) => n1, A(6) => 
                           n1, A(5) => n1, A(4) => n1, A(3) => n1, A(2) => n1, 
                           A(1) => n1, A(0) => n2, B(63) => input(63), B(62) =>
                           input(62), B(61) => input(61), B(60) => input(60), 
                           B(59) => input(59), B(58) => input(58), B(57) => 
                           input(57), B(56) => input(56), B(55) => input(55), 
                           B(54) => input(54), B(53) => input(53), B(52) => 
                           input(52), B(51) => input(51), B(50) => input(50), 
                           B(49) => input(49), B(48) => input(48), B(47) => 
                           input(47), B(46) => input(46), B(45) => input(45), 
                           B(44) => input(44), B(43) => input(43), B(42) => 
                           input(42), B(41) => input(41), B(40) => input(40), 
                           B(39) => input(39), B(38) => input(38), B(37) => 
                           input(37), B(36) => input(36), B(35) => input(35), 
                           B(34) => input(34), B(33) => input(33), B(32) => 
                           input(32), B(31) => input(31), B(30) => input(30), 
                           B(29) => input(29), B(28) => input(28), B(27) => 
                           input(27), B(26) => input(26), B(25) => input(25), 
                           B(24) => input(24), B(23) => input(23), B(22) => 
                           input(22), B(21) => input(21), B(20) => input(20), 
                           B(19) => input(19), B(18) => input(18), B(17) => 
                           input(17), B(16) => input(16), B(15) => input(15), 
                           B(14) => input(14), B(13) => input(13), B(12) => 
                           input(12), B(11) => input(11), B(10) => input(10), 
                           B(9) => input(9), B(8) => input(8), B(7) => input(7)
                           , B(6) => input(6), B(5) => input(5), B(4) => 
                           input(4), B(3) => input(3), B(2) => input(2), B(1) 
                           => input(1), B(0) => input(0), CI => n1, DIFF(63) =>
                           complement2(63), DIFF(62) => complement2(62), 
                           DIFF(61) => complement2(61), DIFF(60) => 
                           complement2(60), DIFF(59) => complement2(59), 
                           DIFF(58) => complement2(58), DIFF(57) => 
                           complement2(57), DIFF(56) => complement2(56), 
                           DIFF(55) => complement2(55), DIFF(54) => 
                           complement2(54), DIFF(53) => complement2(53), 
                           DIFF(52) => complement2(52), DIFF(51) => 
                           complement2(51), DIFF(50) => complement2(50), 
                           DIFF(49) => complement2(49), DIFF(48) => 
                           complement2(48), DIFF(47) => complement2(47), 
                           DIFF(46) => complement2(46), DIFF(45) => 
                           complement2(45), DIFF(44) => complement2(44), 
                           DIFF(43) => complement2(43), DIFF(42) => 
                           complement2(42), DIFF(41) => complement2(41), 
                           DIFF(40) => complement2(40), DIFF(39) => 
                           complement2(39), DIFF(38) => complement2(38), 
                           DIFF(37) => complement2(37), DIFF(36) => 
                           complement2(36), DIFF(35) => complement2(35), 
                           DIFF(34) => complement2(34), DIFF(33) => 
                           complement2(33), DIFF(32) => complement2(32), 
                           DIFF(31) => complement2(31), DIFF(30) => 
                           complement2(30), DIFF(29) => complement2(29), 
                           DIFF(28) => complement2(28), DIFF(27) => 
                           complement2(27), DIFF(26) => complement2(26), 
                           DIFF(25) => complement2(25), DIFF(24) => 
                           complement2(24), DIFF(23) => complement2(23), 
                           DIFF(22) => complement2(22), DIFF(21) => 
                           complement2(21), DIFF(20) => complement2(20), 
                           DIFF(19) => complement2(19), DIFF(18) => 
                           complement2(18), DIFF(17) => complement2(17), 
                           DIFF(16) => complement2(16), DIFF(15) => 
                           complement2(15), DIFF(14) => complement2(14), 
                           DIFF(13) => complement2(13), DIFF(12) => 
                           complement2(12), DIFF(11) => complement2(11), 
                           DIFF(10) => complement2(10), DIFF(9) => 
                           complement2(9), DIFF(8) => complement2(8), DIFF(7) 
                           => complement2(7), DIFF(6) => complement2(6), 
                           DIFF(5) => complement2(5), DIFF(4) => complement2(4)
                           , DIFF(3) => complement2(3), DIFF(2) => 
                           complement2(2), DIFF(1) => complement2(1), DIFF(0) 
                           => complement2(0), CO => n_3121);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_11 is

   port( input : in std_logic_vector (63 downto 0);  complement2 : out 
         std_logic_vector (63 downto 0));

end complementer_N64_11;

architecture SYN_beh of complementer_N64_11 is

   component complementer_N64_11_DW01_sub_0
      port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (63 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n2, n_3122 : std_logic;

begin
   
   n1 <= '0';
   n2 <= '0';
   sub_add_29_b0 : complementer_N64_11_DW01_sub_0 port map( A(63) => n1, A(62) 
                           => n1, A(61) => n1, A(60) => n1, A(59) => n1, A(58) 
                           => n1, A(57) => n1, A(56) => n1, A(55) => n1, A(54) 
                           => n1, A(53) => n1, A(52) => n1, A(51) => n1, A(50) 
                           => n1, A(49) => n1, A(48) => n1, A(47) => n1, A(46) 
                           => n1, A(45) => n1, A(44) => n1, A(43) => n1, A(42) 
                           => n1, A(41) => n1, A(40) => n1, A(39) => n1, A(38) 
                           => n1, A(37) => n1, A(36) => n1, A(35) => n1, A(34) 
                           => n1, A(33) => n1, A(32) => n1, A(31) => n1, A(30) 
                           => n1, A(29) => n1, A(28) => n1, A(27) => n1, A(26) 
                           => n1, A(25) => n1, A(24) => n1, A(23) => n1, A(22) 
                           => n1, A(21) => n1, A(20) => n1, A(19) => n1, A(18) 
                           => n1, A(17) => n1, A(16) => n1, A(15) => n1, A(14) 
                           => n1, A(13) => n1, A(12) => n1, A(11) => n1, A(10) 
                           => n1, A(9) => n1, A(8) => n1, A(7) => n1, A(6) => 
                           n1, A(5) => n1, A(4) => n1, A(3) => n1, A(2) => n1, 
                           A(1) => n1, A(0) => n2, B(63) => input(63), B(62) =>
                           input(62), B(61) => input(61), B(60) => input(60), 
                           B(59) => input(59), B(58) => input(58), B(57) => 
                           input(57), B(56) => input(56), B(55) => input(55), 
                           B(54) => input(54), B(53) => input(53), B(52) => 
                           input(52), B(51) => input(51), B(50) => input(50), 
                           B(49) => input(49), B(48) => input(48), B(47) => 
                           input(47), B(46) => input(46), B(45) => input(45), 
                           B(44) => input(44), B(43) => input(43), B(42) => 
                           input(42), B(41) => input(41), B(40) => input(40), 
                           B(39) => input(39), B(38) => input(38), B(37) => 
                           input(37), B(36) => input(36), B(35) => input(35), 
                           B(34) => input(34), B(33) => input(33), B(32) => 
                           input(32), B(31) => input(31), B(30) => input(30), 
                           B(29) => input(29), B(28) => input(28), B(27) => 
                           input(27), B(26) => input(26), B(25) => input(25), 
                           B(24) => input(24), B(23) => input(23), B(22) => 
                           input(22), B(21) => input(21), B(20) => input(20), 
                           B(19) => input(19), B(18) => input(18), B(17) => 
                           input(17), B(16) => input(16), B(15) => input(15), 
                           B(14) => input(14), B(13) => input(13), B(12) => 
                           input(12), B(11) => input(11), B(10) => input(10), 
                           B(9) => input(9), B(8) => input(8), B(7) => input(7)
                           , B(6) => input(6), B(5) => input(5), B(4) => 
                           input(4), B(3) => input(3), B(2) => input(2), B(1) 
                           => input(1), B(0) => input(0), CI => n1, DIFF(63) =>
                           complement2(63), DIFF(62) => complement2(62), 
                           DIFF(61) => complement2(61), DIFF(60) => 
                           complement2(60), DIFF(59) => complement2(59), 
                           DIFF(58) => complement2(58), DIFF(57) => 
                           complement2(57), DIFF(56) => complement2(56), 
                           DIFF(55) => complement2(55), DIFF(54) => 
                           complement2(54), DIFF(53) => complement2(53), 
                           DIFF(52) => complement2(52), DIFF(51) => 
                           complement2(51), DIFF(50) => complement2(50), 
                           DIFF(49) => complement2(49), DIFF(48) => 
                           complement2(48), DIFF(47) => complement2(47), 
                           DIFF(46) => complement2(46), DIFF(45) => 
                           complement2(45), DIFF(44) => complement2(44), 
                           DIFF(43) => complement2(43), DIFF(42) => 
                           complement2(42), DIFF(41) => complement2(41), 
                           DIFF(40) => complement2(40), DIFF(39) => 
                           complement2(39), DIFF(38) => complement2(38), 
                           DIFF(37) => complement2(37), DIFF(36) => 
                           complement2(36), DIFF(35) => complement2(35), 
                           DIFF(34) => complement2(34), DIFF(33) => 
                           complement2(33), DIFF(32) => complement2(32), 
                           DIFF(31) => complement2(31), DIFF(30) => 
                           complement2(30), DIFF(29) => complement2(29), 
                           DIFF(28) => complement2(28), DIFF(27) => 
                           complement2(27), DIFF(26) => complement2(26), 
                           DIFF(25) => complement2(25), DIFF(24) => 
                           complement2(24), DIFF(23) => complement2(23), 
                           DIFF(22) => complement2(22), DIFF(21) => 
                           complement2(21), DIFF(20) => complement2(20), 
                           DIFF(19) => complement2(19), DIFF(18) => 
                           complement2(18), DIFF(17) => complement2(17), 
                           DIFF(16) => complement2(16), DIFF(15) => 
                           complement2(15), DIFF(14) => complement2(14), 
                           DIFF(13) => complement2(13), DIFF(12) => 
                           complement2(12), DIFF(11) => complement2(11), 
                           DIFF(10) => complement2(10), DIFF(9) => 
                           complement2(9), DIFF(8) => complement2(8), DIFF(7) 
                           => complement2(7), DIFF(6) => complement2(6), 
                           DIFF(5) => complement2(5), DIFF(4) => complement2(4)
                           , DIFF(3) => complement2(3), DIFF(2) => 
                           complement2(2), DIFF(1) => complement2(1), DIFF(0) 
                           => complement2(0), CO => n_3122);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_12 is

   port( input : in std_logic_vector (63 downto 0);  complement2 : out 
         std_logic_vector (63 downto 0));

end complementer_N64_12;

architecture SYN_beh of complementer_N64_12 is

   component complementer_N64_12_DW01_sub_0
      port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (63 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n2, n_3123 : std_logic;

begin
   
   n1 <= '0';
   n2 <= '0';
   sub_add_29_b0 : complementer_N64_12_DW01_sub_0 port map( A(63) => n1, A(62) 
                           => n1, A(61) => n1, A(60) => n1, A(59) => n1, A(58) 
                           => n1, A(57) => n1, A(56) => n1, A(55) => n1, A(54) 
                           => n1, A(53) => n1, A(52) => n1, A(51) => n1, A(50) 
                           => n1, A(49) => n1, A(48) => n1, A(47) => n1, A(46) 
                           => n1, A(45) => n1, A(44) => n1, A(43) => n1, A(42) 
                           => n1, A(41) => n1, A(40) => n1, A(39) => n1, A(38) 
                           => n1, A(37) => n1, A(36) => n1, A(35) => n1, A(34) 
                           => n1, A(33) => n1, A(32) => n1, A(31) => n1, A(30) 
                           => n1, A(29) => n1, A(28) => n1, A(27) => n1, A(26) 
                           => n1, A(25) => n1, A(24) => n1, A(23) => n1, A(22) 
                           => n1, A(21) => n1, A(20) => n1, A(19) => n1, A(18) 
                           => n1, A(17) => n1, A(16) => n1, A(15) => n1, A(14) 
                           => n1, A(13) => n1, A(12) => n1, A(11) => n1, A(10) 
                           => n1, A(9) => n1, A(8) => n1, A(7) => n1, A(6) => 
                           n1, A(5) => n1, A(4) => n1, A(3) => n1, A(2) => n1, 
                           A(1) => n1, A(0) => n2, B(63) => input(63), B(62) =>
                           input(62), B(61) => input(61), B(60) => input(60), 
                           B(59) => input(59), B(58) => input(58), B(57) => 
                           input(57), B(56) => input(56), B(55) => input(55), 
                           B(54) => input(54), B(53) => input(53), B(52) => 
                           input(52), B(51) => input(51), B(50) => input(50), 
                           B(49) => input(49), B(48) => input(48), B(47) => 
                           input(47), B(46) => input(46), B(45) => input(45), 
                           B(44) => input(44), B(43) => input(43), B(42) => 
                           input(42), B(41) => input(41), B(40) => input(40), 
                           B(39) => input(39), B(38) => input(38), B(37) => 
                           input(37), B(36) => input(36), B(35) => input(35), 
                           B(34) => input(34), B(33) => input(33), B(32) => 
                           input(32), B(31) => input(31), B(30) => input(30), 
                           B(29) => input(29), B(28) => input(28), B(27) => 
                           input(27), B(26) => input(26), B(25) => input(25), 
                           B(24) => input(24), B(23) => input(23), B(22) => 
                           input(22), B(21) => input(21), B(20) => input(20), 
                           B(19) => input(19), B(18) => input(18), B(17) => 
                           input(17), B(16) => input(16), B(15) => input(15), 
                           B(14) => input(14), B(13) => input(13), B(12) => 
                           input(12), B(11) => input(11), B(10) => input(10), 
                           B(9) => input(9), B(8) => input(8), B(7) => input(7)
                           , B(6) => input(6), B(5) => input(5), B(4) => 
                           input(4), B(3) => input(3), B(2) => input(2), B(1) 
                           => input(1), B(0) => input(0), CI => n1, DIFF(63) =>
                           complement2(63), DIFF(62) => complement2(62), 
                           DIFF(61) => complement2(61), DIFF(60) => 
                           complement2(60), DIFF(59) => complement2(59), 
                           DIFF(58) => complement2(58), DIFF(57) => 
                           complement2(57), DIFF(56) => complement2(56), 
                           DIFF(55) => complement2(55), DIFF(54) => 
                           complement2(54), DIFF(53) => complement2(53), 
                           DIFF(52) => complement2(52), DIFF(51) => 
                           complement2(51), DIFF(50) => complement2(50), 
                           DIFF(49) => complement2(49), DIFF(48) => 
                           complement2(48), DIFF(47) => complement2(47), 
                           DIFF(46) => complement2(46), DIFF(45) => 
                           complement2(45), DIFF(44) => complement2(44), 
                           DIFF(43) => complement2(43), DIFF(42) => 
                           complement2(42), DIFF(41) => complement2(41), 
                           DIFF(40) => complement2(40), DIFF(39) => 
                           complement2(39), DIFF(38) => complement2(38), 
                           DIFF(37) => complement2(37), DIFF(36) => 
                           complement2(36), DIFF(35) => complement2(35), 
                           DIFF(34) => complement2(34), DIFF(33) => 
                           complement2(33), DIFF(32) => complement2(32), 
                           DIFF(31) => complement2(31), DIFF(30) => 
                           complement2(30), DIFF(29) => complement2(29), 
                           DIFF(28) => complement2(28), DIFF(27) => 
                           complement2(27), DIFF(26) => complement2(26), 
                           DIFF(25) => complement2(25), DIFF(24) => 
                           complement2(24), DIFF(23) => complement2(23), 
                           DIFF(22) => complement2(22), DIFF(21) => 
                           complement2(21), DIFF(20) => complement2(20), 
                           DIFF(19) => complement2(19), DIFF(18) => 
                           complement2(18), DIFF(17) => complement2(17), 
                           DIFF(16) => complement2(16), DIFF(15) => 
                           complement2(15), DIFF(14) => complement2(14), 
                           DIFF(13) => complement2(13), DIFF(12) => 
                           complement2(12), DIFF(11) => complement2(11), 
                           DIFF(10) => complement2(10), DIFF(9) => 
                           complement2(9), DIFF(8) => complement2(8), DIFF(7) 
                           => complement2(7), DIFF(6) => complement2(6), 
                           DIFF(5) => complement2(5), DIFF(4) => complement2(4)
                           , DIFF(3) => complement2(3), DIFF(2) => 
                           complement2(2), DIFF(1) => complement2(1), DIFF(0) 
                           => complement2(0), CO => n_3123);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_13 is

   port( input : in std_logic_vector (63 downto 0);  complement2 : out 
         std_logic_vector (63 downto 0));

end complementer_N64_13;

architecture SYN_beh of complementer_N64_13 is

   component complementer_N64_13_DW01_sub_0
      port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (63 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n2, n_3124 : std_logic;

begin
   
   n1 <= '0';
   n2 <= '0';
   sub_add_29_b0 : complementer_N64_13_DW01_sub_0 port map( A(63) => n1, A(62) 
                           => n1, A(61) => n1, A(60) => n1, A(59) => n1, A(58) 
                           => n1, A(57) => n1, A(56) => n1, A(55) => n1, A(54) 
                           => n1, A(53) => n1, A(52) => n1, A(51) => n1, A(50) 
                           => n1, A(49) => n1, A(48) => n1, A(47) => n1, A(46) 
                           => n1, A(45) => n1, A(44) => n1, A(43) => n1, A(42) 
                           => n1, A(41) => n1, A(40) => n1, A(39) => n1, A(38) 
                           => n1, A(37) => n1, A(36) => n1, A(35) => n1, A(34) 
                           => n1, A(33) => n1, A(32) => n1, A(31) => n1, A(30) 
                           => n1, A(29) => n1, A(28) => n1, A(27) => n1, A(26) 
                           => n1, A(25) => n1, A(24) => n1, A(23) => n1, A(22) 
                           => n1, A(21) => n1, A(20) => n1, A(19) => n1, A(18) 
                           => n1, A(17) => n1, A(16) => n1, A(15) => n1, A(14) 
                           => n1, A(13) => n1, A(12) => n1, A(11) => n1, A(10) 
                           => n1, A(9) => n1, A(8) => n1, A(7) => n1, A(6) => 
                           n1, A(5) => n1, A(4) => n1, A(3) => n1, A(2) => n1, 
                           A(1) => n1, A(0) => n2, B(63) => input(63), B(62) =>
                           input(62), B(61) => input(61), B(60) => input(60), 
                           B(59) => input(59), B(58) => input(58), B(57) => 
                           input(57), B(56) => input(56), B(55) => input(55), 
                           B(54) => input(54), B(53) => input(53), B(52) => 
                           input(52), B(51) => input(51), B(50) => input(50), 
                           B(49) => input(49), B(48) => input(48), B(47) => 
                           input(47), B(46) => input(46), B(45) => input(45), 
                           B(44) => input(44), B(43) => input(43), B(42) => 
                           input(42), B(41) => input(41), B(40) => input(40), 
                           B(39) => input(39), B(38) => input(38), B(37) => 
                           input(37), B(36) => input(36), B(35) => input(35), 
                           B(34) => input(34), B(33) => input(33), B(32) => 
                           input(32), B(31) => input(31), B(30) => input(30), 
                           B(29) => input(29), B(28) => input(28), B(27) => 
                           input(27), B(26) => input(26), B(25) => input(25), 
                           B(24) => input(24), B(23) => input(23), B(22) => 
                           input(22), B(21) => input(21), B(20) => input(20), 
                           B(19) => input(19), B(18) => input(18), B(17) => 
                           input(17), B(16) => input(16), B(15) => input(15), 
                           B(14) => input(14), B(13) => input(13), B(12) => 
                           input(12), B(11) => input(11), B(10) => input(10), 
                           B(9) => input(9), B(8) => input(8), B(7) => input(7)
                           , B(6) => input(6), B(5) => input(5), B(4) => 
                           input(4), B(3) => input(3), B(2) => input(2), B(1) 
                           => input(1), B(0) => input(0), CI => n1, DIFF(63) =>
                           complement2(63), DIFF(62) => complement2(62), 
                           DIFF(61) => complement2(61), DIFF(60) => 
                           complement2(60), DIFF(59) => complement2(59), 
                           DIFF(58) => complement2(58), DIFF(57) => 
                           complement2(57), DIFF(56) => complement2(56), 
                           DIFF(55) => complement2(55), DIFF(54) => 
                           complement2(54), DIFF(53) => complement2(53), 
                           DIFF(52) => complement2(52), DIFF(51) => 
                           complement2(51), DIFF(50) => complement2(50), 
                           DIFF(49) => complement2(49), DIFF(48) => 
                           complement2(48), DIFF(47) => complement2(47), 
                           DIFF(46) => complement2(46), DIFF(45) => 
                           complement2(45), DIFF(44) => complement2(44), 
                           DIFF(43) => complement2(43), DIFF(42) => 
                           complement2(42), DIFF(41) => complement2(41), 
                           DIFF(40) => complement2(40), DIFF(39) => 
                           complement2(39), DIFF(38) => complement2(38), 
                           DIFF(37) => complement2(37), DIFF(36) => 
                           complement2(36), DIFF(35) => complement2(35), 
                           DIFF(34) => complement2(34), DIFF(33) => 
                           complement2(33), DIFF(32) => complement2(32), 
                           DIFF(31) => complement2(31), DIFF(30) => 
                           complement2(30), DIFF(29) => complement2(29), 
                           DIFF(28) => complement2(28), DIFF(27) => 
                           complement2(27), DIFF(26) => complement2(26), 
                           DIFF(25) => complement2(25), DIFF(24) => 
                           complement2(24), DIFF(23) => complement2(23), 
                           DIFF(22) => complement2(22), DIFF(21) => 
                           complement2(21), DIFF(20) => complement2(20), 
                           DIFF(19) => complement2(19), DIFF(18) => 
                           complement2(18), DIFF(17) => complement2(17), 
                           DIFF(16) => complement2(16), DIFF(15) => 
                           complement2(15), DIFF(14) => complement2(14), 
                           DIFF(13) => complement2(13), DIFF(12) => 
                           complement2(12), DIFF(11) => complement2(11), 
                           DIFF(10) => complement2(10), DIFF(9) => 
                           complement2(9), DIFF(8) => complement2(8), DIFF(7) 
                           => complement2(7), DIFF(6) => complement2(6), 
                           DIFF(5) => complement2(5), DIFF(4) => complement2(4)
                           , DIFF(3) => complement2(3), DIFF(2) => 
                           complement2(2), DIFF(1) => complement2(1), DIFF(0) 
                           => complement2(0), CO => n_3124);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_14 is

   port( input : in std_logic_vector (63 downto 0);  complement2 : out 
         std_logic_vector (63 downto 0));

end complementer_N64_14;

architecture SYN_beh of complementer_N64_14 is

   component complementer_N64_14_DW01_sub_0
      port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (63 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n2, n_3125 : std_logic;

begin
   
   n1 <= '0';
   n2 <= '0';
   sub_add_29_b0 : complementer_N64_14_DW01_sub_0 port map( A(63) => n1, A(62) 
                           => n1, A(61) => n1, A(60) => n1, A(59) => n1, A(58) 
                           => n1, A(57) => n1, A(56) => n1, A(55) => n1, A(54) 
                           => n1, A(53) => n1, A(52) => n1, A(51) => n1, A(50) 
                           => n1, A(49) => n1, A(48) => n1, A(47) => n1, A(46) 
                           => n1, A(45) => n1, A(44) => n1, A(43) => n1, A(42) 
                           => n1, A(41) => n1, A(40) => n1, A(39) => n1, A(38) 
                           => n1, A(37) => n1, A(36) => n1, A(35) => n1, A(34) 
                           => n1, A(33) => n1, A(32) => n1, A(31) => n1, A(30) 
                           => n1, A(29) => n1, A(28) => n1, A(27) => n1, A(26) 
                           => n1, A(25) => n1, A(24) => n1, A(23) => n1, A(22) 
                           => n1, A(21) => n1, A(20) => n1, A(19) => n1, A(18) 
                           => n1, A(17) => n1, A(16) => n1, A(15) => n1, A(14) 
                           => n1, A(13) => n1, A(12) => n1, A(11) => n1, A(10) 
                           => n1, A(9) => n1, A(8) => n1, A(7) => n1, A(6) => 
                           n1, A(5) => n1, A(4) => n1, A(3) => n1, A(2) => n1, 
                           A(1) => n1, A(0) => n2, B(63) => input(63), B(62) =>
                           input(62), B(61) => input(61), B(60) => input(60), 
                           B(59) => input(59), B(58) => input(58), B(57) => 
                           input(57), B(56) => input(56), B(55) => input(55), 
                           B(54) => input(54), B(53) => input(53), B(52) => 
                           input(52), B(51) => input(51), B(50) => input(50), 
                           B(49) => input(49), B(48) => input(48), B(47) => 
                           input(47), B(46) => input(46), B(45) => input(45), 
                           B(44) => input(44), B(43) => input(43), B(42) => 
                           input(42), B(41) => input(41), B(40) => input(40), 
                           B(39) => input(39), B(38) => input(38), B(37) => 
                           input(37), B(36) => input(36), B(35) => input(35), 
                           B(34) => input(34), B(33) => input(33), B(32) => 
                           input(32), B(31) => input(31), B(30) => input(30), 
                           B(29) => input(29), B(28) => input(28), B(27) => 
                           input(27), B(26) => input(26), B(25) => input(25), 
                           B(24) => input(24), B(23) => input(23), B(22) => 
                           input(22), B(21) => input(21), B(20) => input(20), 
                           B(19) => input(19), B(18) => input(18), B(17) => 
                           input(17), B(16) => input(16), B(15) => input(15), 
                           B(14) => input(14), B(13) => input(13), B(12) => 
                           input(12), B(11) => input(11), B(10) => input(10), 
                           B(9) => input(9), B(8) => input(8), B(7) => input(7)
                           , B(6) => input(6), B(5) => input(5), B(4) => 
                           input(4), B(3) => input(3), B(2) => input(2), B(1) 
                           => input(1), B(0) => input(0), CI => n1, DIFF(63) =>
                           complement2(63), DIFF(62) => complement2(62), 
                           DIFF(61) => complement2(61), DIFF(60) => 
                           complement2(60), DIFF(59) => complement2(59), 
                           DIFF(58) => complement2(58), DIFF(57) => 
                           complement2(57), DIFF(56) => complement2(56), 
                           DIFF(55) => complement2(55), DIFF(54) => 
                           complement2(54), DIFF(53) => complement2(53), 
                           DIFF(52) => complement2(52), DIFF(51) => 
                           complement2(51), DIFF(50) => complement2(50), 
                           DIFF(49) => complement2(49), DIFF(48) => 
                           complement2(48), DIFF(47) => complement2(47), 
                           DIFF(46) => complement2(46), DIFF(45) => 
                           complement2(45), DIFF(44) => complement2(44), 
                           DIFF(43) => complement2(43), DIFF(42) => 
                           complement2(42), DIFF(41) => complement2(41), 
                           DIFF(40) => complement2(40), DIFF(39) => 
                           complement2(39), DIFF(38) => complement2(38), 
                           DIFF(37) => complement2(37), DIFF(36) => 
                           complement2(36), DIFF(35) => complement2(35), 
                           DIFF(34) => complement2(34), DIFF(33) => 
                           complement2(33), DIFF(32) => complement2(32), 
                           DIFF(31) => complement2(31), DIFF(30) => 
                           complement2(30), DIFF(29) => complement2(29), 
                           DIFF(28) => complement2(28), DIFF(27) => 
                           complement2(27), DIFF(26) => complement2(26), 
                           DIFF(25) => complement2(25), DIFF(24) => 
                           complement2(24), DIFF(23) => complement2(23), 
                           DIFF(22) => complement2(22), DIFF(21) => 
                           complement2(21), DIFF(20) => complement2(20), 
                           DIFF(19) => complement2(19), DIFF(18) => 
                           complement2(18), DIFF(17) => complement2(17), 
                           DIFF(16) => complement2(16), DIFF(15) => 
                           complement2(15), DIFF(14) => complement2(14), 
                           DIFF(13) => complement2(13), DIFF(12) => 
                           complement2(12), DIFF(11) => complement2(11), 
                           DIFF(10) => complement2(10), DIFF(9) => 
                           complement2(9), DIFF(8) => complement2(8), DIFF(7) 
                           => complement2(7), DIFF(6) => complement2(6), 
                           DIFF(5) => complement2(5), DIFF(4) => complement2(4)
                           , DIFF(3) => complement2(3), DIFF(2) => 
                           complement2(2), DIFF(1) => complement2(1), DIFF(0) 
                           => complement2(0), CO => n_3125);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_15 is

   port( input : in std_logic_vector (63 downto 0);  complement2 : out 
         std_logic_vector (63 downto 0));

end complementer_N64_15;

architecture SYN_beh of complementer_N64_15 is

   component complementer_N64_15_DW01_sub_0
      port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (63 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n2, n_3126 : std_logic;

begin
   
   n1 <= '0';
   n2 <= '0';
   sub_add_29_b0 : complementer_N64_15_DW01_sub_0 port map( A(63) => n1, A(62) 
                           => n1, A(61) => n1, A(60) => n1, A(59) => n1, A(58) 
                           => n1, A(57) => n1, A(56) => n1, A(55) => n1, A(54) 
                           => n1, A(53) => n1, A(52) => n1, A(51) => n1, A(50) 
                           => n1, A(49) => n1, A(48) => n1, A(47) => n1, A(46) 
                           => n1, A(45) => n1, A(44) => n1, A(43) => n1, A(42) 
                           => n1, A(41) => n1, A(40) => n1, A(39) => n1, A(38) 
                           => n1, A(37) => n1, A(36) => n1, A(35) => n1, A(34) 
                           => n1, A(33) => n1, A(32) => n1, A(31) => n1, A(30) 
                           => n1, A(29) => n1, A(28) => n1, A(27) => n1, A(26) 
                           => n1, A(25) => n1, A(24) => n1, A(23) => n1, A(22) 
                           => n1, A(21) => n1, A(20) => n1, A(19) => n1, A(18) 
                           => n1, A(17) => n1, A(16) => n1, A(15) => n1, A(14) 
                           => n1, A(13) => n1, A(12) => n1, A(11) => n1, A(10) 
                           => n1, A(9) => n1, A(8) => n1, A(7) => n1, A(6) => 
                           n1, A(5) => n1, A(4) => n1, A(3) => n1, A(2) => n1, 
                           A(1) => n1, A(0) => n2, B(63) => input(63), B(62) =>
                           input(62), B(61) => input(61), B(60) => input(60), 
                           B(59) => input(59), B(58) => input(58), B(57) => 
                           input(57), B(56) => input(56), B(55) => input(55), 
                           B(54) => input(54), B(53) => input(53), B(52) => 
                           input(52), B(51) => input(51), B(50) => input(50), 
                           B(49) => input(49), B(48) => input(48), B(47) => 
                           input(47), B(46) => input(46), B(45) => input(45), 
                           B(44) => input(44), B(43) => input(43), B(42) => 
                           input(42), B(41) => input(41), B(40) => input(40), 
                           B(39) => input(39), B(38) => input(38), B(37) => 
                           input(37), B(36) => input(36), B(35) => input(35), 
                           B(34) => input(34), B(33) => input(33), B(32) => 
                           input(32), B(31) => input(31), B(30) => input(30), 
                           B(29) => input(29), B(28) => input(28), B(27) => 
                           input(27), B(26) => input(26), B(25) => input(25), 
                           B(24) => input(24), B(23) => input(23), B(22) => 
                           input(22), B(21) => input(21), B(20) => input(20), 
                           B(19) => input(19), B(18) => input(18), B(17) => 
                           input(17), B(16) => input(16), B(15) => input(15), 
                           B(14) => input(14), B(13) => input(13), B(12) => 
                           input(12), B(11) => input(11), B(10) => input(10), 
                           B(9) => input(9), B(8) => input(8), B(7) => input(7)
                           , B(6) => input(6), B(5) => input(5), B(4) => 
                           input(4), B(3) => input(3), B(2) => input(2), B(1) 
                           => input(1), B(0) => input(0), CI => n1, DIFF(63) =>
                           complement2(63), DIFF(62) => complement2(62), 
                           DIFF(61) => complement2(61), DIFF(60) => 
                           complement2(60), DIFF(59) => complement2(59), 
                           DIFF(58) => complement2(58), DIFF(57) => 
                           complement2(57), DIFF(56) => complement2(56), 
                           DIFF(55) => complement2(55), DIFF(54) => 
                           complement2(54), DIFF(53) => complement2(53), 
                           DIFF(52) => complement2(52), DIFF(51) => 
                           complement2(51), DIFF(50) => complement2(50), 
                           DIFF(49) => complement2(49), DIFF(48) => 
                           complement2(48), DIFF(47) => complement2(47), 
                           DIFF(46) => complement2(46), DIFF(45) => 
                           complement2(45), DIFF(44) => complement2(44), 
                           DIFF(43) => complement2(43), DIFF(42) => 
                           complement2(42), DIFF(41) => complement2(41), 
                           DIFF(40) => complement2(40), DIFF(39) => 
                           complement2(39), DIFF(38) => complement2(38), 
                           DIFF(37) => complement2(37), DIFF(36) => 
                           complement2(36), DIFF(35) => complement2(35), 
                           DIFF(34) => complement2(34), DIFF(33) => 
                           complement2(33), DIFF(32) => complement2(32), 
                           DIFF(31) => complement2(31), DIFF(30) => 
                           complement2(30), DIFF(29) => complement2(29), 
                           DIFF(28) => complement2(28), DIFF(27) => 
                           complement2(27), DIFF(26) => complement2(26), 
                           DIFF(25) => complement2(25), DIFF(24) => 
                           complement2(24), DIFF(23) => complement2(23), 
                           DIFF(22) => complement2(22), DIFF(21) => 
                           complement2(21), DIFF(20) => complement2(20), 
                           DIFF(19) => complement2(19), DIFF(18) => 
                           complement2(18), DIFF(17) => complement2(17), 
                           DIFF(16) => complement2(16), DIFF(15) => 
                           complement2(15), DIFF(14) => complement2(14), 
                           DIFF(13) => complement2(13), DIFF(12) => 
                           complement2(12), DIFF(11) => complement2(11), 
                           DIFF(10) => complement2(10), DIFF(9) => 
                           complement2(9), DIFF(8) => complement2(8), DIFF(7) 
                           => complement2(7), DIFF(6) => complement2(6), 
                           DIFF(5) => complement2(5), DIFF(4) => complement2(4)
                           , DIFF(3) => complement2(3), DIFF(2) => 
                           complement2(2), DIFF(1) => complement2(1), DIFF(0) 
                           => complement2(0), CO => n_3126);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_16 is

   port( input : in std_logic_vector (63 downto 0);  complement2 : out 
         std_logic_vector (63 downto 0));

end complementer_N64_16;

architecture SYN_beh of complementer_N64_16 is

   component complementer_N64_16_DW01_sub_0
      port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (63 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n2, n_3127 : std_logic;

begin
   
   n1 <= '0';
   n2 <= '0';
   sub_add_29_b0 : complementer_N64_16_DW01_sub_0 port map( A(63) => n1, A(62) 
                           => n1, A(61) => n1, A(60) => n1, A(59) => n1, A(58) 
                           => n1, A(57) => n1, A(56) => n1, A(55) => n1, A(54) 
                           => n1, A(53) => n1, A(52) => n1, A(51) => n1, A(50) 
                           => n1, A(49) => n1, A(48) => n1, A(47) => n1, A(46) 
                           => n1, A(45) => n1, A(44) => n1, A(43) => n1, A(42) 
                           => n1, A(41) => n1, A(40) => n1, A(39) => n1, A(38) 
                           => n1, A(37) => n1, A(36) => n1, A(35) => n1, A(34) 
                           => n1, A(33) => n1, A(32) => n1, A(31) => n1, A(30) 
                           => n1, A(29) => n1, A(28) => n1, A(27) => n1, A(26) 
                           => n1, A(25) => n1, A(24) => n1, A(23) => n1, A(22) 
                           => n1, A(21) => n1, A(20) => n1, A(19) => n1, A(18) 
                           => n1, A(17) => n1, A(16) => n1, A(15) => n1, A(14) 
                           => n1, A(13) => n1, A(12) => n1, A(11) => n1, A(10) 
                           => n1, A(9) => n1, A(8) => n1, A(7) => n1, A(6) => 
                           n1, A(5) => n1, A(4) => n1, A(3) => n1, A(2) => n1, 
                           A(1) => n1, A(0) => n2, B(63) => input(63), B(62) =>
                           input(62), B(61) => input(61), B(60) => input(60), 
                           B(59) => input(59), B(58) => input(58), B(57) => 
                           input(57), B(56) => input(56), B(55) => input(55), 
                           B(54) => input(54), B(53) => input(53), B(52) => 
                           input(52), B(51) => input(51), B(50) => input(50), 
                           B(49) => input(49), B(48) => input(48), B(47) => 
                           input(47), B(46) => input(46), B(45) => input(45), 
                           B(44) => input(44), B(43) => input(43), B(42) => 
                           input(42), B(41) => input(41), B(40) => input(40), 
                           B(39) => input(39), B(38) => input(38), B(37) => 
                           input(37), B(36) => input(36), B(35) => input(35), 
                           B(34) => input(34), B(33) => input(33), B(32) => 
                           input(32), B(31) => input(31), B(30) => input(30), 
                           B(29) => input(29), B(28) => input(28), B(27) => 
                           input(27), B(26) => input(26), B(25) => input(25), 
                           B(24) => input(24), B(23) => input(23), B(22) => 
                           input(22), B(21) => input(21), B(20) => input(20), 
                           B(19) => input(19), B(18) => input(18), B(17) => 
                           input(17), B(16) => input(16), B(15) => input(15), 
                           B(14) => input(14), B(13) => input(13), B(12) => 
                           input(12), B(11) => input(11), B(10) => input(10), 
                           B(9) => input(9), B(8) => input(8), B(7) => input(7)
                           , B(6) => input(6), B(5) => input(5), B(4) => 
                           input(4), B(3) => input(3), B(2) => input(2), B(1) 
                           => input(1), B(0) => input(0), CI => n1, DIFF(63) =>
                           complement2(63), DIFF(62) => complement2(62), 
                           DIFF(61) => complement2(61), DIFF(60) => 
                           complement2(60), DIFF(59) => complement2(59), 
                           DIFF(58) => complement2(58), DIFF(57) => 
                           complement2(57), DIFF(56) => complement2(56), 
                           DIFF(55) => complement2(55), DIFF(54) => 
                           complement2(54), DIFF(53) => complement2(53), 
                           DIFF(52) => complement2(52), DIFF(51) => 
                           complement2(51), DIFF(50) => complement2(50), 
                           DIFF(49) => complement2(49), DIFF(48) => 
                           complement2(48), DIFF(47) => complement2(47), 
                           DIFF(46) => complement2(46), DIFF(45) => 
                           complement2(45), DIFF(44) => complement2(44), 
                           DIFF(43) => complement2(43), DIFF(42) => 
                           complement2(42), DIFF(41) => complement2(41), 
                           DIFF(40) => complement2(40), DIFF(39) => 
                           complement2(39), DIFF(38) => complement2(38), 
                           DIFF(37) => complement2(37), DIFF(36) => 
                           complement2(36), DIFF(35) => complement2(35), 
                           DIFF(34) => complement2(34), DIFF(33) => 
                           complement2(33), DIFF(32) => complement2(32), 
                           DIFF(31) => complement2(31), DIFF(30) => 
                           complement2(30), DIFF(29) => complement2(29), 
                           DIFF(28) => complement2(28), DIFF(27) => 
                           complement2(27), DIFF(26) => complement2(26), 
                           DIFF(25) => complement2(25), DIFF(24) => 
                           complement2(24), DIFF(23) => complement2(23), 
                           DIFF(22) => complement2(22), DIFF(21) => 
                           complement2(21), DIFF(20) => complement2(20), 
                           DIFF(19) => complement2(19), DIFF(18) => 
                           complement2(18), DIFF(17) => complement2(17), 
                           DIFF(16) => complement2(16), DIFF(15) => 
                           complement2(15), DIFF(14) => complement2(14), 
                           DIFF(13) => complement2(13), DIFF(12) => 
                           complement2(12), DIFF(11) => complement2(11), 
                           DIFF(10) => complement2(10), DIFF(9) => 
                           complement2(9), DIFF(8) => complement2(8), DIFF(7) 
                           => complement2(7), DIFF(6) => complement2(6), 
                           DIFF(5) => complement2(5), DIFF(4) => complement2(4)
                           , DIFF(3) => complement2(3), DIFF(2) => 
                           complement2(2), DIFF(1) => complement2(1), DIFF(0) 
                           => complement2(0), CO => n_3127);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_17 is

   port( input : in std_logic_vector (63 downto 0);  complement2 : out 
         std_logic_vector (63 downto 0));

end complementer_N64_17;

architecture SYN_beh of complementer_N64_17 is

   component complementer_N64_17_DW01_sub_0
      port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (63 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n2, n_3128 : std_logic;

begin
   
   n1 <= '0';
   n2 <= '0';
   sub_add_29_b0 : complementer_N64_17_DW01_sub_0 port map( A(63) => n1, A(62) 
                           => n1, A(61) => n1, A(60) => n1, A(59) => n1, A(58) 
                           => n1, A(57) => n1, A(56) => n1, A(55) => n1, A(54) 
                           => n1, A(53) => n1, A(52) => n1, A(51) => n1, A(50) 
                           => n1, A(49) => n1, A(48) => n1, A(47) => n1, A(46) 
                           => n1, A(45) => n1, A(44) => n1, A(43) => n1, A(42) 
                           => n1, A(41) => n1, A(40) => n1, A(39) => n1, A(38) 
                           => n1, A(37) => n1, A(36) => n1, A(35) => n1, A(34) 
                           => n1, A(33) => n1, A(32) => n1, A(31) => n1, A(30) 
                           => n1, A(29) => n1, A(28) => n1, A(27) => n1, A(26) 
                           => n1, A(25) => n1, A(24) => n1, A(23) => n1, A(22) 
                           => n1, A(21) => n1, A(20) => n1, A(19) => n1, A(18) 
                           => n1, A(17) => n1, A(16) => n1, A(15) => n1, A(14) 
                           => n1, A(13) => n1, A(12) => n1, A(11) => n1, A(10) 
                           => n1, A(9) => n1, A(8) => n1, A(7) => n1, A(6) => 
                           n1, A(5) => n1, A(4) => n1, A(3) => n1, A(2) => n1, 
                           A(1) => n1, A(0) => n2, B(63) => input(63), B(62) =>
                           input(62), B(61) => input(61), B(60) => input(60), 
                           B(59) => input(59), B(58) => input(58), B(57) => 
                           input(57), B(56) => input(56), B(55) => input(55), 
                           B(54) => input(54), B(53) => input(53), B(52) => 
                           input(52), B(51) => input(51), B(50) => input(50), 
                           B(49) => input(49), B(48) => input(48), B(47) => 
                           input(47), B(46) => input(46), B(45) => input(45), 
                           B(44) => input(44), B(43) => input(43), B(42) => 
                           input(42), B(41) => input(41), B(40) => input(40), 
                           B(39) => input(39), B(38) => input(38), B(37) => 
                           input(37), B(36) => input(36), B(35) => input(35), 
                           B(34) => input(34), B(33) => input(33), B(32) => 
                           input(32), B(31) => input(31), B(30) => input(30), 
                           B(29) => input(29), B(28) => input(28), B(27) => 
                           input(27), B(26) => input(26), B(25) => input(25), 
                           B(24) => input(24), B(23) => input(23), B(22) => 
                           input(22), B(21) => input(21), B(20) => input(20), 
                           B(19) => input(19), B(18) => input(18), B(17) => 
                           input(17), B(16) => input(16), B(15) => input(15), 
                           B(14) => input(14), B(13) => input(13), B(12) => 
                           input(12), B(11) => input(11), B(10) => input(10), 
                           B(9) => input(9), B(8) => input(8), B(7) => input(7)
                           , B(6) => input(6), B(5) => input(5), B(4) => 
                           input(4), B(3) => input(3), B(2) => input(2), B(1) 
                           => input(1), B(0) => input(0), CI => n1, DIFF(63) =>
                           complement2(63), DIFF(62) => complement2(62), 
                           DIFF(61) => complement2(61), DIFF(60) => 
                           complement2(60), DIFF(59) => complement2(59), 
                           DIFF(58) => complement2(58), DIFF(57) => 
                           complement2(57), DIFF(56) => complement2(56), 
                           DIFF(55) => complement2(55), DIFF(54) => 
                           complement2(54), DIFF(53) => complement2(53), 
                           DIFF(52) => complement2(52), DIFF(51) => 
                           complement2(51), DIFF(50) => complement2(50), 
                           DIFF(49) => complement2(49), DIFF(48) => 
                           complement2(48), DIFF(47) => complement2(47), 
                           DIFF(46) => complement2(46), DIFF(45) => 
                           complement2(45), DIFF(44) => complement2(44), 
                           DIFF(43) => complement2(43), DIFF(42) => 
                           complement2(42), DIFF(41) => complement2(41), 
                           DIFF(40) => complement2(40), DIFF(39) => 
                           complement2(39), DIFF(38) => complement2(38), 
                           DIFF(37) => complement2(37), DIFF(36) => 
                           complement2(36), DIFF(35) => complement2(35), 
                           DIFF(34) => complement2(34), DIFF(33) => 
                           complement2(33), DIFF(32) => complement2(32), 
                           DIFF(31) => complement2(31), DIFF(30) => 
                           complement2(30), DIFF(29) => complement2(29), 
                           DIFF(28) => complement2(28), DIFF(27) => 
                           complement2(27), DIFF(26) => complement2(26), 
                           DIFF(25) => complement2(25), DIFF(24) => 
                           complement2(24), DIFF(23) => complement2(23), 
                           DIFF(22) => complement2(22), DIFF(21) => 
                           complement2(21), DIFF(20) => complement2(20), 
                           DIFF(19) => complement2(19), DIFF(18) => 
                           complement2(18), DIFF(17) => complement2(17), 
                           DIFF(16) => complement2(16), DIFF(15) => 
                           complement2(15), DIFF(14) => complement2(14), 
                           DIFF(13) => complement2(13), DIFF(12) => 
                           complement2(12), DIFF(11) => complement2(11), 
                           DIFF(10) => complement2(10), DIFF(9) => 
                           complement2(9), DIFF(8) => complement2(8), DIFF(7) 
                           => complement2(7), DIFF(6) => complement2(6), 
                           DIFF(5) => complement2(5), DIFF(4) => complement2(4)
                           , DIFF(3) => complement2(3), DIFF(2) => 
                           complement2(2), DIFF(1) => complement2(1), DIFF(0) 
                           => complement2(0), CO => n_3128);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_18 is

   port( input : in std_logic_vector (63 downto 0);  complement2 : out 
         std_logic_vector (63 downto 0));

end complementer_N64_18;

architecture SYN_beh of complementer_N64_18 is

   component complementer_N64_18_DW01_sub_0
      port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (63 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n2, n_3129 : std_logic;

begin
   
   n1 <= '0';
   n2 <= '0';
   sub_add_29_b0 : complementer_N64_18_DW01_sub_0 port map( A(63) => n1, A(62) 
                           => n1, A(61) => n1, A(60) => n1, A(59) => n1, A(58) 
                           => n1, A(57) => n1, A(56) => n1, A(55) => n1, A(54) 
                           => n1, A(53) => n1, A(52) => n1, A(51) => n1, A(50) 
                           => n1, A(49) => n1, A(48) => n1, A(47) => n1, A(46) 
                           => n1, A(45) => n1, A(44) => n1, A(43) => n1, A(42) 
                           => n1, A(41) => n1, A(40) => n1, A(39) => n1, A(38) 
                           => n1, A(37) => n1, A(36) => n1, A(35) => n1, A(34) 
                           => n1, A(33) => n1, A(32) => n1, A(31) => n1, A(30) 
                           => n1, A(29) => n1, A(28) => n1, A(27) => n1, A(26) 
                           => n1, A(25) => n1, A(24) => n1, A(23) => n1, A(22) 
                           => n1, A(21) => n1, A(20) => n1, A(19) => n1, A(18) 
                           => n1, A(17) => n1, A(16) => n1, A(15) => n1, A(14) 
                           => n1, A(13) => n1, A(12) => n1, A(11) => n1, A(10) 
                           => n1, A(9) => n1, A(8) => n1, A(7) => n1, A(6) => 
                           n1, A(5) => n1, A(4) => n1, A(3) => n1, A(2) => n1, 
                           A(1) => n1, A(0) => n2, B(63) => input(63), B(62) =>
                           input(62), B(61) => input(61), B(60) => input(60), 
                           B(59) => input(59), B(58) => input(58), B(57) => 
                           input(57), B(56) => input(56), B(55) => input(55), 
                           B(54) => input(54), B(53) => input(53), B(52) => 
                           input(52), B(51) => input(51), B(50) => input(50), 
                           B(49) => input(49), B(48) => input(48), B(47) => 
                           input(47), B(46) => input(46), B(45) => input(45), 
                           B(44) => input(44), B(43) => input(43), B(42) => 
                           input(42), B(41) => input(41), B(40) => input(40), 
                           B(39) => input(39), B(38) => input(38), B(37) => 
                           input(37), B(36) => input(36), B(35) => input(35), 
                           B(34) => input(34), B(33) => input(33), B(32) => 
                           input(32), B(31) => input(31), B(30) => input(30), 
                           B(29) => input(29), B(28) => input(28), B(27) => 
                           input(27), B(26) => input(26), B(25) => input(25), 
                           B(24) => input(24), B(23) => input(23), B(22) => 
                           input(22), B(21) => input(21), B(20) => input(20), 
                           B(19) => input(19), B(18) => input(18), B(17) => 
                           input(17), B(16) => input(16), B(15) => input(15), 
                           B(14) => input(14), B(13) => input(13), B(12) => 
                           input(12), B(11) => input(11), B(10) => input(10), 
                           B(9) => input(9), B(8) => input(8), B(7) => input(7)
                           , B(6) => input(6), B(5) => input(5), B(4) => 
                           input(4), B(3) => input(3), B(2) => input(2), B(1) 
                           => input(1), B(0) => input(0), CI => n1, DIFF(63) =>
                           complement2(63), DIFF(62) => complement2(62), 
                           DIFF(61) => complement2(61), DIFF(60) => 
                           complement2(60), DIFF(59) => complement2(59), 
                           DIFF(58) => complement2(58), DIFF(57) => 
                           complement2(57), DIFF(56) => complement2(56), 
                           DIFF(55) => complement2(55), DIFF(54) => 
                           complement2(54), DIFF(53) => complement2(53), 
                           DIFF(52) => complement2(52), DIFF(51) => 
                           complement2(51), DIFF(50) => complement2(50), 
                           DIFF(49) => complement2(49), DIFF(48) => 
                           complement2(48), DIFF(47) => complement2(47), 
                           DIFF(46) => complement2(46), DIFF(45) => 
                           complement2(45), DIFF(44) => complement2(44), 
                           DIFF(43) => complement2(43), DIFF(42) => 
                           complement2(42), DIFF(41) => complement2(41), 
                           DIFF(40) => complement2(40), DIFF(39) => 
                           complement2(39), DIFF(38) => complement2(38), 
                           DIFF(37) => complement2(37), DIFF(36) => 
                           complement2(36), DIFF(35) => complement2(35), 
                           DIFF(34) => complement2(34), DIFF(33) => 
                           complement2(33), DIFF(32) => complement2(32), 
                           DIFF(31) => complement2(31), DIFF(30) => 
                           complement2(30), DIFF(29) => complement2(29), 
                           DIFF(28) => complement2(28), DIFF(27) => 
                           complement2(27), DIFF(26) => complement2(26), 
                           DIFF(25) => complement2(25), DIFF(24) => 
                           complement2(24), DIFF(23) => complement2(23), 
                           DIFF(22) => complement2(22), DIFF(21) => 
                           complement2(21), DIFF(20) => complement2(20), 
                           DIFF(19) => complement2(19), DIFF(18) => 
                           complement2(18), DIFF(17) => complement2(17), 
                           DIFF(16) => complement2(16), DIFF(15) => 
                           complement2(15), DIFF(14) => complement2(14), 
                           DIFF(13) => complement2(13), DIFF(12) => 
                           complement2(12), DIFF(11) => complement2(11), 
                           DIFF(10) => complement2(10), DIFF(9) => 
                           complement2(9), DIFF(8) => complement2(8), DIFF(7) 
                           => complement2(7), DIFF(6) => complement2(6), 
                           DIFF(5) => complement2(5), DIFF(4) => complement2(4)
                           , DIFF(3) => complement2(3), DIFF(2) => 
                           complement2(2), DIFF(1) => complement2(1), DIFF(0) 
                           => complement2(0), CO => n_3129);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_19 is

   port( input : in std_logic_vector (63 downto 0);  complement2 : out 
         std_logic_vector (63 downto 0));

end complementer_N64_19;

architecture SYN_beh of complementer_N64_19 is

   component complementer_N64_19_DW01_sub_0
      port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (63 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n2, n_3130 : std_logic;

begin
   
   n1 <= '0';
   n2 <= '0';
   sub_add_29_b0 : complementer_N64_19_DW01_sub_0 port map( A(63) => n1, A(62) 
                           => n1, A(61) => n1, A(60) => n1, A(59) => n1, A(58) 
                           => n1, A(57) => n1, A(56) => n1, A(55) => n1, A(54) 
                           => n1, A(53) => n1, A(52) => n1, A(51) => n1, A(50) 
                           => n1, A(49) => n1, A(48) => n1, A(47) => n1, A(46) 
                           => n1, A(45) => n1, A(44) => n1, A(43) => n1, A(42) 
                           => n1, A(41) => n1, A(40) => n1, A(39) => n1, A(38) 
                           => n1, A(37) => n1, A(36) => n1, A(35) => n1, A(34) 
                           => n1, A(33) => n1, A(32) => n1, A(31) => n1, A(30) 
                           => n1, A(29) => n1, A(28) => n1, A(27) => n1, A(26) 
                           => n1, A(25) => n1, A(24) => n1, A(23) => n1, A(22) 
                           => n1, A(21) => n1, A(20) => n1, A(19) => n1, A(18) 
                           => n1, A(17) => n1, A(16) => n1, A(15) => n1, A(14) 
                           => n1, A(13) => n1, A(12) => n1, A(11) => n1, A(10) 
                           => n1, A(9) => n1, A(8) => n1, A(7) => n1, A(6) => 
                           n1, A(5) => n1, A(4) => n1, A(3) => n1, A(2) => n1, 
                           A(1) => n1, A(0) => n2, B(63) => input(63), B(62) =>
                           input(62), B(61) => input(61), B(60) => input(60), 
                           B(59) => input(59), B(58) => input(58), B(57) => 
                           input(57), B(56) => input(56), B(55) => input(55), 
                           B(54) => input(54), B(53) => input(53), B(52) => 
                           input(52), B(51) => input(51), B(50) => input(50), 
                           B(49) => input(49), B(48) => input(48), B(47) => 
                           input(47), B(46) => input(46), B(45) => input(45), 
                           B(44) => input(44), B(43) => input(43), B(42) => 
                           input(42), B(41) => input(41), B(40) => input(40), 
                           B(39) => input(39), B(38) => input(38), B(37) => 
                           input(37), B(36) => input(36), B(35) => input(35), 
                           B(34) => input(34), B(33) => input(33), B(32) => 
                           input(32), B(31) => input(31), B(30) => input(30), 
                           B(29) => input(29), B(28) => input(28), B(27) => 
                           input(27), B(26) => input(26), B(25) => input(25), 
                           B(24) => input(24), B(23) => input(23), B(22) => 
                           input(22), B(21) => input(21), B(20) => input(20), 
                           B(19) => input(19), B(18) => input(18), B(17) => 
                           input(17), B(16) => input(16), B(15) => input(15), 
                           B(14) => input(14), B(13) => input(13), B(12) => 
                           input(12), B(11) => input(11), B(10) => input(10), 
                           B(9) => input(9), B(8) => input(8), B(7) => input(7)
                           , B(6) => input(6), B(5) => input(5), B(4) => 
                           input(4), B(3) => input(3), B(2) => input(2), B(1) 
                           => input(1), B(0) => input(0), CI => n1, DIFF(63) =>
                           complement2(63), DIFF(62) => complement2(62), 
                           DIFF(61) => complement2(61), DIFF(60) => 
                           complement2(60), DIFF(59) => complement2(59), 
                           DIFF(58) => complement2(58), DIFF(57) => 
                           complement2(57), DIFF(56) => complement2(56), 
                           DIFF(55) => complement2(55), DIFF(54) => 
                           complement2(54), DIFF(53) => complement2(53), 
                           DIFF(52) => complement2(52), DIFF(51) => 
                           complement2(51), DIFF(50) => complement2(50), 
                           DIFF(49) => complement2(49), DIFF(48) => 
                           complement2(48), DIFF(47) => complement2(47), 
                           DIFF(46) => complement2(46), DIFF(45) => 
                           complement2(45), DIFF(44) => complement2(44), 
                           DIFF(43) => complement2(43), DIFF(42) => 
                           complement2(42), DIFF(41) => complement2(41), 
                           DIFF(40) => complement2(40), DIFF(39) => 
                           complement2(39), DIFF(38) => complement2(38), 
                           DIFF(37) => complement2(37), DIFF(36) => 
                           complement2(36), DIFF(35) => complement2(35), 
                           DIFF(34) => complement2(34), DIFF(33) => 
                           complement2(33), DIFF(32) => complement2(32), 
                           DIFF(31) => complement2(31), DIFF(30) => 
                           complement2(30), DIFF(29) => complement2(29), 
                           DIFF(28) => complement2(28), DIFF(27) => 
                           complement2(27), DIFF(26) => complement2(26), 
                           DIFF(25) => complement2(25), DIFF(24) => 
                           complement2(24), DIFF(23) => complement2(23), 
                           DIFF(22) => complement2(22), DIFF(21) => 
                           complement2(21), DIFF(20) => complement2(20), 
                           DIFF(19) => complement2(19), DIFF(18) => 
                           complement2(18), DIFF(17) => complement2(17), 
                           DIFF(16) => complement2(16), DIFF(15) => 
                           complement2(15), DIFF(14) => complement2(14), 
                           DIFF(13) => complement2(13), DIFF(12) => 
                           complement2(12), DIFF(11) => complement2(11), 
                           DIFF(10) => complement2(10), DIFF(9) => 
                           complement2(9), DIFF(8) => complement2(8), DIFF(7) 
                           => complement2(7), DIFF(6) => complement2(6), 
                           DIFF(5) => complement2(5), DIFF(4) => complement2(4)
                           , DIFF(3) => complement2(3), DIFF(2) => 
                           complement2(2), DIFF(1) => complement2(1), DIFF(0) 
                           => complement2(0), CO => n_3130);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_20 is

   port( input : in std_logic_vector (63 downto 0);  complement2 : out 
         std_logic_vector (63 downto 0));

end complementer_N64_20;

architecture SYN_beh of complementer_N64_20 is

   component complementer_N64_20_DW01_sub_0
      port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (63 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n2, n_3131 : std_logic;

begin
   
   n1 <= '0';
   n2 <= '0';
   sub_add_29_b0 : complementer_N64_20_DW01_sub_0 port map( A(63) => n1, A(62) 
                           => n1, A(61) => n1, A(60) => n1, A(59) => n1, A(58) 
                           => n1, A(57) => n1, A(56) => n1, A(55) => n1, A(54) 
                           => n1, A(53) => n1, A(52) => n1, A(51) => n1, A(50) 
                           => n1, A(49) => n1, A(48) => n1, A(47) => n1, A(46) 
                           => n1, A(45) => n1, A(44) => n1, A(43) => n1, A(42) 
                           => n1, A(41) => n1, A(40) => n1, A(39) => n1, A(38) 
                           => n1, A(37) => n1, A(36) => n1, A(35) => n1, A(34) 
                           => n1, A(33) => n1, A(32) => n1, A(31) => n1, A(30) 
                           => n1, A(29) => n1, A(28) => n1, A(27) => n1, A(26) 
                           => n1, A(25) => n1, A(24) => n1, A(23) => n1, A(22) 
                           => n1, A(21) => n1, A(20) => n1, A(19) => n1, A(18) 
                           => n1, A(17) => n1, A(16) => n1, A(15) => n1, A(14) 
                           => n1, A(13) => n1, A(12) => n1, A(11) => n1, A(10) 
                           => n1, A(9) => n1, A(8) => n1, A(7) => n1, A(6) => 
                           n1, A(5) => n1, A(4) => n1, A(3) => n1, A(2) => n1, 
                           A(1) => n1, A(0) => n2, B(63) => input(63), B(62) =>
                           input(62), B(61) => input(61), B(60) => input(60), 
                           B(59) => input(59), B(58) => input(58), B(57) => 
                           input(57), B(56) => input(56), B(55) => input(55), 
                           B(54) => input(54), B(53) => input(53), B(52) => 
                           input(52), B(51) => input(51), B(50) => input(50), 
                           B(49) => input(49), B(48) => input(48), B(47) => 
                           input(47), B(46) => input(46), B(45) => input(45), 
                           B(44) => input(44), B(43) => input(43), B(42) => 
                           input(42), B(41) => input(41), B(40) => input(40), 
                           B(39) => input(39), B(38) => input(38), B(37) => 
                           input(37), B(36) => input(36), B(35) => input(35), 
                           B(34) => input(34), B(33) => input(33), B(32) => 
                           input(32), B(31) => input(31), B(30) => input(30), 
                           B(29) => input(29), B(28) => input(28), B(27) => 
                           input(27), B(26) => input(26), B(25) => input(25), 
                           B(24) => input(24), B(23) => input(23), B(22) => 
                           input(22), B(21) => input(21), B(20) => input(20), 
                           B(19) => input(19), B(18) => input(18), B(17) => 
                           input(17), B(16) => input(16), B(15) => input(15), 
                           B(14) => input(14), B(13) => input(13), B(12) => 
                           input(12), B(11) => input(11), B(10) => input(10), 
                           B(9) => input(9), B(8) => input(8), B(7) => input(7)
                           , B(6) => input(6), B(5) => input(5), B(4) => 
                           input(4), B(3) => input(3), B(2) => input(2), B(1) 
                           => input(1), B(0) => input(0), CI => n1, DIFF(63) =>
                           complement2(63), DIFF(62) => complement2(62), 
                           DIFF(61) => complement2(61), DIFF(60) => 
                           complement2(60), DIFF(59) => complement2(59), 
                           DIFF(58) => complement2(58), DIFF(57) => 
                           complement2(57), DIFF(56) => complement2(56), 
                           DIFF(55) => complement2(55), DIFF(54) => 
                           complement2(54), DIFF(53) => complement2(53), 
                           DIFF(52) => complement2(52), DIFF(51) => 
                           complement2(51), DIFF(50) => complement2(50), 
                           DIFF(49) => complement2(49), DIFF(48) => 
                           complement2(48), DIFF(47) => complement2(47), 
                           DIFF(46) => complement2(46), DIFF(45) => 
                           complement2(45), DIFF(44) => complement2(44), 
                           DIFF(43) => complement2(43), DIFF(42) => 
                           complement2(42), DIFF(41) => complement2(41), 
                           DIFF(40) => complement2(40), DIFF(39) => 
                           complement2(39), DIFF(38) => complement2(38), 
                           DIFF(37) => complement2(37), DIFF(36) => 
                           complement2(36), DIFF(35) => complement2(35), 
                           DIFF(34) => complement2(34), DIFF(33) => 
                           complement2(33), DIFF(32) => complement2(32), 
                           DIFF(31) => complement2(31), DIFF(30) => 
                           complement2(30), DIFF(29) => complement2(29), 
                           DIFF(28) => complement2(28), DIFF(27) => 
                           complement2(27), DIFF(26) => complement2(26), 
                           DIFF(25) => complement2(25), DIFF(24) => 
                           complement2(24), DIFF(23) => complement2(23), 
                           DIFF(22) => complement2(22), DIFF(21) => 
                           complement2(21), DIFF(20) => complement2(20), 
                           DIFF(19) => complement2(19), DIFF(18) => 
                           complement2(18), DIFF(17) => complement2(17), 
                           DIFF(16) => complement2(16), DIFF(15) => 
                           complement2(15), DIFF(14) => complement2(14), 
                           DIFF(13) => complement2(13), DIFF(12) => 
                           complement2(12), DIFF(11) => complement2(11), 
                           DIFF(10) => complement2(10), DIFF(9) => 
                           complement2(9), DIFF(8) => complement2(8), DIFF(7) 
                           => complement2(7), DIFF(6) => complement2(6), 
                           DIFF(5) => complement2(5), DIFF(4) => complement2(4)
                           , DIFF(3) => complement2(3), DIFF(2) => 
                           complement2(2), DIFF(1) => complement2(1), DIFF(0) 
                           => complement2(0), CO => n_3131);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_21 is

   port( input : in std_logic_vector (63 downto 0);  complement2 : out 
         std_logic_vector (63 downto 0));

end complementer_N64_21;

architecture SYN_beh of complementer_N64_21 is

   component complementer_N64_21_DW01_sub_0
      port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (63 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n2, n_3132 : std_logic;

begin
   
   n1 <= '0';
   n2 <= '0';
   sub_add_29_b0 : complementer_N64_21_DW01_sub_0 port map( A(63) => n1, A(62) 
                           => n1, A(61) => n1, A(60) => n1, A(59) => n1, A(58) 
                           => n1, A(57) => n1, A(56) => n1, A(55) => n1, A(54) 
                           => n1, A(53) => n1, A(52) => n1, A(51) => n1, A(50) 
                           => n1, A(49) => n1, A(48) => n1, A(47) => n1, A(46) 
                           => n1, A(45) => n1, A(44) => n1, A(43) => n1, A(42) 
                           => n1, A(41) => n1, A(40) => n1, A(39) => n1, A(38) 
                           => n1, A(37) => n1, A(36) => n1, A(35) => n1, A(34) 
                           => n1, A(33) => n1, A(32) => n1, A(31) => n1, A(30) 
                           => n1, A(29) => n1, A(28) => n1, A(27) => n1, A(26) 
                           => n1, A(25) => n1, A(24) => n1, A(23) => n1, A(22) 
                           => n1, A(21) => n1, A(20) => n1, A(19) => n1, A(18) 
                           => n1, A(17) => n1, A(16) => n1, A(15) => n1, A(14) 
                           => n1, A(13) => n1, A(12) => n1, A(11) => n1, A(10) 
                           => n1, A(9) => n1, A(8) => n1, A(7) => n1, A(6) => 
                           n1, A(5) => n1, A(4) => n1, A(3) => n1, A(2) => n1, 
                           A(1) => n1, A(0) => n2, B(63) => input(63), B(62) =>
                           input(62), B(61) => input(61), B(60) => input(60), 
                           B(59) => input(59), B(58) => input(58), B(57) => 
                           input(57), B(56) => input(56), B(55) => input(55), 
                           B(54) => input(54), B(53) => input(53), B(52) => 
                           input(52), B(51) => input(51), B(50) => input(50), 
                           B(49) => input(49), B(48) => input(48), B(47) => 
                           input(47), B(46) => input(46), B(45) => input(45), 
                           B(44) => input(44), B(43) => input(43), B(42) => 
                           input(42), B(41) => input(41), B(40) => input(40), 
                           B(39) => input(39), B(38) => input(38), B(37) => 
                           input(37), B(36) => input(36), B(35) => input(35), 
                           B(34) => input(34), B(33) => input(33), B(32) => 
                           input(32), B(31) => input(31), B(30) => input(30), 
                           B(29) => input(29), B(28) => input(28), B(27) => 
                           input(27), B(26) => input(26), B(25) => input(25), 
                           B(24) => input(24), B(23) => input(23), B(22) => 
                           input(22), B(21) => input(21), B(20) => input(20), 
                           B(19) => input(19), B(18) => input(18), B(17) => 
                           input(17), B(16) => input(16), B(15) => input(15), 
                           B(14) => input(14), B(13) => input(13), B(12) => 
                           input(12), B(11) => input(11), B(10) => input(10), 
                           B(9) => input(9), B(8) => input(8), B(7) => input(7)
                           , B(6) => input(6), B(5) => input(5), B(4) => 
                           input(4), B(3) => input(3), B(2) => input(2), B(1) 
                           => input(1), B(0) => input(0), CI => n1, DIFF(63) =>
                           complement2(63), DIFF(62) => complement2(62), 
                           DIFF(61) => complement2(61), DIFF(60) => 
                           complement2(60), DIFF(59) => complement2(59), 
                           DIFF(58) => complement2(58), DIFF(57) => 
                           complement2(57), DIFF(56) => complement2(56), 
                           DIFF(55) => complement2(55), DIFF(54) => 
                           complement2(54), DIFF(53) => complement2(53), 
                           DIFF(52) => complement2(52), DIFF(51) => 
                           complement2(51), DIFF(50) => complement2(50), 
                           DIFF(49) => complement2(49), DIFF(48) => 
                           complement2(48), DIFF(47) => complement2(47), 
                           DIFF(46) => complement2(46), DIFF(45) => 
                           complement2(45), DIFF(44) => complement2(44), 
                           DIFF(43) => complement2(43), DIFF(42) => 
                           complement2(42), DIFF(41) => complement2(41), 
                           DIFF(40) => complement2(40), DIFF(39) => 
                           complement2(39), DIFF(38) => complement2(38), 
                           DIFF(37) => complement2(37), DIFF(36) => 
                           complement2(36), DIFF(35) => complement2(35), 
                           DIFF(34) => complement2(34), DIFF(33) => 
                           complement2(33), DIFF(32) => complement2(32), 
                           DIFF(31) => complement2(31), DIFF(30) => 
                           complement2(30), DIFF(29) => complement2(29), 
                           DIFF(28) => complement2(28), DIFF(27) => 
                           complement2(27), DIFF(26) => complement2(26), 
                           DIFF(25) => complement2(25), DIFF(24) => 
                           complement2(24), DIFF(23) => complement2(23), 
                           DIFF(22) => complement2(22), DIFF(21) => 
                           complement2(21), DIFF(20) => complement2(20), 
                           DIFF(19) => complement2(19), DIFF(18) => 
                           complement2(18), DIFF(17) => complement2(17), 
                           DIFF(16) => complement2(16), DIFF(15) => 
                           complement2(15), DIFF(14) => complement2(14), 
                           DIFF(13) => complement2(13), DIFF(12) => 
                           complement2(12), DIFF(11) => complement2(11), 
                           DIFF(10) => complement2(10), DIFF(9) => 
                           complement2(9), DIFF(8) => complement2(8), DIFF(7) 
                           => complement2(7), DIFF(6) => complement2(6), 
                           DIFF(5) => complement2(5), DIFF(4) => complement2(4)
                           , DIFF(3) => complement2(3), DIFF(2) => 
                           complement2(2), DIFF(1) => complement2(1), DIFF(0) 
                           => complement2(0), CO => n_3132);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_22 is

   port( input : in std_logic_vector (63 downto 0);  complement2 : out 
         std_logic_vector (63 downto 0));

end complementer_N64_22;

architecture SYN_beh of complementer_N64_22 is

   component complementer_N64_22_DW01_sub_0
      port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (63 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n2, n_3133 : std_logic;

begin
   
   n1 <= '0';
   n2 <= '0';
   sub_add_29_b0 : complementer_N64_22_DW01_sub_0 port map( A(63) => n1, A(62) 
                           => n1, A(61) => n1, A(60) => n1, A(59) => n1, A(58) 
                           => n1, A(57) => n1, A(56) => n1, A(55) => n1, A(54) 
                           => n1, A(53) => n1, A(52) => n1, A(51) => n1, A(50) 
                           => n1, A(49) => n1, A(48) => n1, A(47) => n1, A(46) 
                           => n1, A(45) => n1, A(44) => n1, A(43) => n1, A(42) 
                           => n1, A(41) => n1, A(40) => n1, A(39) => n1, A(38) 
                           => n1, A(37) => n1, A(36) => n1, A(35) => n1, A(34) 
                           => n1, A(33) => n1, A(32) => n1, A(31) => n1, A(30) 
                           => n1, A(29) => n1, A(28) => n1, A(27) => n1, A(26) 
                           => n1, A(25) => n1, A(24) => n1, A(23) => n1, A(22) 
                           => n1, A(21) => n1, A(20) => n1, A(19) => n1, A(18) 
                           => n1, A(17) => n1, A(16) => n1, A(15) => n1, A(14) 
                           => n1, A(13) => n1, A(12) => n1, A(11) => n1, A(10) 
                           => n1, A(9) => n1, A(8) => n1, A(7) => n1, A(6) => 
                           n1, A(5) => n1, A(4) => n1, A(3) => n1, A(2) => n1, 
                           A(1) => n1, A(0) => n2, B(63) => input(63), B(62) =>
                           input(62), B(61) => input(61), B(60) => input(60), 
                           B(59) => input(59), B(58) => input(58), B(57) => 
                           input(57), B(56) => input(56), B(55) => input(55), 
                           B(54) => input(54), B(53) => input(53), B(52) => 
                           input(52), B(51) => input(51), B(50) => input(50), 
                           B(49) => input(49), B(48) => input(48), B(47) => 
                           input(47), B(46) => input(46), B(45) => input(45), 
                           B(44) => input(44), B(43) => input(43), B(42) => 
                           input(42), B(41) => input(41), B(40) => input(40), 
                           B(39) => input(39), B(38) => input(38), B(37) => 
                           input(37), B(36) => input(36), B(35) => input(35), 
                           B(34) => input(34), B(33) => input(33), B(32) => 
                           input(32), B(31) => input(31), B(30) => input(30), 
                           B(29) => input(29), B(28) => input(28), B(27) => 
                           input(27), B(26) => input(26), B(25) => input(25), 
                           B(24) => input(24), B(23) => input(23), B(22) => 
                           input(22), B(21) => input(21), B(20) => input(20), 
                           B(19) => input(19), B(18) => input(18), B(17) => 
                           input(17), B(16) => input(16), B(15) => input(15), 
                           B(14) => input(14), B(13) => input(13), B(12) => 
                           input(12), B(11) => input(11), B(10) => input(10), 
                           B(9) => input(9), B(8) => input(8), B(7) => input(7)
                           , B(6) => input(6), B(5) => input(5), B(4) => 
                           input(4), B(3) => input(3), B(2) => input(2), B(1) 
                           => input(1), B(0) => input(0), CI => n1, DIFF(63) =>
                           complement2(63), DIFF(62) => complement2(62), 
                           DIFF(61) => complement2(61), DIFF(60) => 
                           complement2(60), DIFF(59) => complement2(59), 
                           DIFF(58) => complement2(58), DIFF(57) => 
                           complement2(57), DIFF(56) => complement2(56), 
                           DIFF(55) => complement2(55), DIFF(54) => 
                           complement2(54), DIFF(53) => complement2(53), 
                           DIFF(52) => complement2(52), DIFF(51) => 
                           complement2(51), DIFF(50) => complement2(50), 
                           DIFF(49) => complement2(49), DIFF(48) => 
                           complement2(48), DIFF(47) => complement2(47), 
                           DIFF(46) => complement2(46), DIFF(45) => 
                           complement2(45), DIFF(44) => complement2(44), 
                           DIFF(43) => complement2(43), DIFF(42) => 
                           complement2(42), DIFF(41) => complement2(41), 
                           DIFF(40) => complement2(40), DIFF(39) => 
                           complement2(39), DIFF(38) => complement2(38), 
                           DIFF(37) => complement2(37), DIFF(36) => 
                           complement2(36), DIFF(35) => complement2(35), 
                           DIFF(34) => complement2(34), DIFF(33) => 
                           complement2(33), DIFF(32) => complement2(32), 
                           DIFF(31) => complement2(31), DIFF(30) => 
                           complement2(30), DIFF(29) => complement2(29), 
                           DIFF(28) => complement2(28), DIFF(27) => 
                           complement2(27), DIFF(26) => complement2(26), 
                           DIFF(25) => complement2(25), DIFF(24) => 
                           complement2(24), DIFF(23) => complement2(23), 
                           DIFF(22) => complement2(22), DIFF(21) => 
                           complement2(21), DIFF(20) => complement2(20), 
                           DIFF(19) => complement2(19), DIFF(18) => 
                           complement2(18), DIFF(17) => complement2(17), 
                           DIFF(16) => complement2(16), DIFF(15) => 
                           complement2(15), DIFF(14) => complement2(14), 
                           DIFF(13) => complement2(13), DIFF(12) => 
                           complement2(12), DIFF(11) => complement2(11), 
                           DIFF(10) => complement2(10), DIFF(9) => 
                           complement2(9), DIFF(8) => complement2(8), DIFF(7) 
                           => complement2(7), DIFF(6) => complement2(6), 
                           DIFF(5) => complement2(5), DIFF(4) => complement2(4)
                           , DIFF(3) => complement2(3), DIFF(2) => 
                           complement2(2), DIFF(1) => complement2(1), DIFF(0) 
                           => complement2(0), CO => n_3133);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_23 is

   port( input : in std_logic_vector (63 downto 0);  complement2 : out 
         std_logic_vector (63 downto 0));

end complementer_N64_23;

architecture SYN_beh of complementer_N64_23 is

   component complementer_N64_23_DW01_sub_0
      port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (63 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n2, n_3134 : std_logic;

begin
   
   n1 <= '0';
   n2 <= '0';
   sub_add_29_b0 : complementer_N64_23_DW01_sub_0 port map( A(63) => n1, A(62) 
                           => n1, A(61) => n1, A(60) => n1, A(59) => n1, A(58) 
                           => n1, A(57) => n1, A(56) => n1, A(55) => n1, A(54) 
                           => n1, A(53) => n1, A(52) => n1, A(51) => n1, A(50) 
                           => n1, A(49) => n1, A(48) => n1, A(47) => n1, A(46) 
                           => n1, A(45) => n1, A(44) => n1, A(43) => n1, A(42) 
                           => n1, A(41) => n1, A(40) => n1, A(39) => n1, A(38) 
                           => n1, A(37) => n1, A(36) => n1, A(35) => n1, A(34) 
                           => n1, A(33) => n1, A(32) => n1, A(31) => n1, A(30) 
                           => n1, A(29) => n1, A(28) => n1, A(27) => n1, A(26) 
                           => n1, A(25) => n1, A(24) => n1, A(23) => n1, A(22) 
                           => n1, A(21) => n1, A(20) => n1, A(19) => n1, A(18) 
                           => n1, A(17) => n1, A(16) => n1, A(15) => n1, A(14) 
                           => n1, A(13) => n1, A(12) => n1, A(11) => n1, A(10) 
                           => n1, A(9) => n1, A(8) => n1, A(7) => n1, A(6) => 
                           n1, A(5) => n1, A(4) => n1, A(3) => n1, A(2) => n1, 
                           A(1) => n1, A(0) => n2, B(63) => input(63), B(62) =>
                           input(62), B(61) => input(61), B(60) => input(60), 
                           B(59) => input(59), B(58) => input(58), B(57) => 
                           input(57), B(56) => input(56), B(55) => input(55), 
                           B(54) => input(54), B(53) => input(53), B(52) => 
                           input(52), B(51) => input(51), B(50) => input(50), 
                           B(49) => input(49), B(48) => input(48), B(47) => 
                           input(47), B(46) => input(46), B(45) => input(45), 
                           B(44) => input(44), B(43) => input(43), B(42) => 
                           input(42), B(41) => input(41), B(40) => input(40), 
                           B(39) => input(39), B(38) => input(38), B(37) => 
                           input(37), B(36) => input(36), B(35) => input(35), 
                           B(34) => input(34), B(33) => input(33), B(32) => 
                           input(32), B(31) => input(31), B(30) => input(30), 
                           B(29) => input(29), B(28) => input(28), B(27) => 
                           input(27), B(26) => input(26), B(25) => input(25), 
                           B(24) => input(24), B(23) => input(23), B(22) => 
                           input(22), B(21) => input(21), B(20) => input(20), 
                           B(19) => input(19), B(18) => input(18), B(17) => 
                           input(17), B(16) => input(16), B(15) => input(15), 
                           B(14) => input(14), B(13) => input(13), B(12) => 
                           input(12), B(11) => input(11), B(10) => input(10), 
                           B(9) => input(9), B(8) => input(8), B(7) => input(7)
                           , B(6) => input(6), B(5) => input(5), B(4) => 
                           input(4), B(3) => input(3), B(2) => input(2), B(1) 
                           => input(1), B(0) => input(0), CI => n1, DIFF(63) =>
                           complement2(63), DIFF(62) => complement2(62), 
                           DIFF(61) => complement2(61), DIFF(60) => 
                           complement2(60), DIFF(59) => complement2(59), 
                           DIFF(58) => complement2(58), DIFF(57) => 
                           complement2(57), DIFF(56) => complement2(56), 
                           DIFF(55) => complement2(55), DIFF(54) => 
                           complement2(54), DIFF(53) => complement2(53), 
                           DIFF(52) => complement2(52), DIFF(51) => 
                           complement2(51), DIFF(50) => complement2(50), 
                           DIFF(49) => complement2(49), DIFF(48) => 
                           complement2(48), DIFF(47) => complement2(47), 
                           DIFF(46) => complement2(46), DIFF(45) => 
                           complement2(45), DIFF(44) => complement2(44), 
                           DIFF(43) => complement2(43), DIFF(42) => 
                           complement2(42), DIFF(41) => complement2(41), 
                           DIFF(40) => complement2(40), DIFF(39) => 
                           complement2(39), DIFF(38) => complement2(38), 
                           DIFF(37) => complement2(37), DIFF(36) => 
                           complement2(36), DIFF(35) => complement2(35), 
                           DIFF(34) => complement2(34), DIFF(33) => 
                           complement2(33), DIFF(32) => complement2(32), 
                           DIFF(31) => complement2(31), DIFF(30) => 
                           complement2(30), DIFF(29) => complement2(29), 
                           DIFF(28) => complement2(28), DIFF(27) => 
                           complement2(27), DIFF(26) => complement2(26), 
                           DIFF(25) => complement2(25), DIFF(24) => 
                           complement2(24), DIFF(23) => complement2(23), 
                           DIFF(22) => complement2(22), DIFF(21) => 
                           complement2(21), DIFF(20) => complement2(20), 
                           DIFF(19) => complement2(19), DIFF(18) => 
                           complement2(18), DIFF(17) => complement2(17), 
                           DIFF(16) => complement2(16), DIFF(15) => 
                           complement2(15), DIFF(14) => complement2(14), 
                           DIFF(13) => complement2(13), DIFF(12) => 
                           complement2(12), DIFF(11) => complement2(11), 
                           DIFF(10) => complement2(10), DIFF(9) => 
                           complement2(9), DIFF(8) => complement2(8), DIFF(7) 
                           => complement2(7), DIFF(6) => complement2(6), 
                           DIFF(5) => complement2(5), DIFF(4) => complement2(4)
                           , DIFF(3) => complement2(3), DIFF(2) => 
                           complement2(2), DIFF(1) => complement2(1), DIFF(0) 
                           => complement2(0), CO => n_3134);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_24 is

   port( input : in std_logic_vector (63 downto 0);  complement2 : out 
         std_logic_vector (63 downto 0));

end complementer_N64_24;

architecture SYN_beh of complementer_N64_24 is

   component complementer_N64_24_DW01_sub_0
      port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (63 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n2, n_3135 : std_logic;

begin
   
   n1 <= '0';
   n2 <= '0';
   sub_add_29_b0 : complementer_N64_24_DW01_sub_0 port map( A(63) => n1, A(62) 
                           => n1, A(61) => n1, A(60) => n1, A(59) => n1, A(58) 
                           => n1, A(57) => n1, A(56) => n1, A(55) => n1, A(54) 
                           => n1, A(53) => n1, A(52) => n1, A(51) => n1, A(50) 
                           => n1, A(49) => n1, A(48) => n1, A(47) => n1, A(46) 
                           => n1, A(45) => n1, A(44) => n1, A(43) => n1, A(42) 
                           => n1, A(41) => n1, A(40) => n1, A(39) => n1, A(38) 
                           => n1, A(37) => n1, A(36) => n1, A(35) => n1, A(34) 
                           => n1, A(33) => n1, A(32) => n1, A(31) => n1, A(30) 
                           => n1, A(29) => n1, A(28) => n1, A(27) => n1, A(26) 
                           => n1, A(25) => n1, A(24) => n1, A(23) => n1, A(22) 
                           => n1, A(21) => n1, A(20) => n1, A(19) => n1, A(18) 
                           => n1, A(17) => n1, A(16) => n1, A(15) => n1, A(14) 
                           => n1, A(13) => n1, A(12) => n1, A(11) => n1, A(10) 
                           => n1, A(9) => n1, A(8) => n1, A(7) => n1, A(6) => 
                           n1, A(5) => n1, A(4) => n1, A(3) => n1, A(2) => n1, 
                           A(1) => n1, A(0) => n2, B(63) => input(63), B(62) =>
                           input(62), B(61) => input(61), B(60) => input(60), 
                           B(59) => input(59), B(58) => input(58), B(57) => 
                           input(57), B(56) => input(56), B(55) => input(55), 
                           B(54) => input(54), B(53) => input(53), B(52) => 
                           input(52), B(51) => input(51), B(50) => input(50), 
                           B(49) => input(49), B(48) => input(48), B(47) => 
                           input(47), B(46) => input(46), B(45) => input(45), 
                           B(44) => input(44), B(43) => input(43), B(42) => 
                           input(42), B(41) => input(41), B(40) => input(40), 
                           B(39) => input(39), B(38) => input(38), B(37) => 
                           input(37), B(36) => input(36), B(35) => input(35), 
                           B(34) => input(34), B(33) => input(33), B(32) => 
                           input(32), B(31) => input(31), B(30) => input(30), 
                           B(29) => input(29), B(28) => input(28), B(27) => 
                           input(27), B(26) => input(26), B(25) => input(25), 
                           B(24) => input(24), B(23) => input(23), B(22) => 
                           input(22), B(21) => input(21), B(20) => input(20), 
                           B(19) => input(19), B(18) => input(18), B(17) => 
                           input(17), B(16) => input(16), B(15) => input(15), 
                           B(14) => input(14), B(13) => input(13), B(12) => 
                           input(12), B(11) => input(11), B(10) => input(10), 
                           B(9) => input(9), B(8) => input(8), B(7) => input(7)
                           , B(6) => input(6), B(5) => input(5), B(4) => 
                           input(4), B(3) => input(3), B(2) => input(2), B(1) 
                           => input(1), B(0) => input(0), CI => n1, DIFF(63) =>
                           complement2(63), DIFF(62) => complement2(62), 
                           DIFF(61) => complement2(61), DIFF(60) => 
                           complement2(60), DIFF(59) => complement2(59), 
                           DIFF(58) => complement2(58), DIFF(57) => 
                           complement2(57), DIFF(56) => complement2(56), 
                           DIFF(55) => complement2(55), DIFF(54) => 
                           complement2(54), DIFF(53) => complement2(53), 
                           DIFF(52) => complement2(52), DIFF(51) => 
                           complement2(51), DIFF(50) => complement2(50), 
                           DIFF(49) => complement2(49), DIFF(48) => 
                           complement2(48), DIFF(47) => complement2(47), 
                           DIFF(46) => complement2(46), DIFF(45) => 
                           complement2(45), DIFF(44) => complement2(44), 
                           DIFF(43) => complement2(43), DIFF(42) => 
                           complement2(42), DIFF(41) => complement2(41), 
                           DIFF(40) => complement2(40), DIFF(39) => 
                           complement2(39), DIFF(38) => complement2(38), 
                           DIFF(37) => complement2(37), DIFF(36) => 
                           complement2(36), DIFF(35) => complement2(35), 
                           DIFF(34) => complement2(34), DIFF(33) => 
                           complement2(33), DIFF(32) => complement2(32), 
                           DIFF(31) => complement2(31), DIFF(30) => 
                           complement2(30), DIFF(29) => complement2(29), 
                           DIFF(28) => complement2(28), DIFF(27) => 
                           complement2(27), DIFF(26) => complement2(26), 
                           DIFF(25) => complement2(25), DIFF(24) => 
                           complement2(24), DIFF(23) => complement2(23), 
                           DIFF(22) => complement2(22), DIFF(21) => 
                           complement2(21), DIFF(20) => complement2(20), 
                           DIFF(19) => complement2(19), DIFF(18) => 
                           complement2(18), DIFF(17) => complement2(17), 
                           DIFF(16) => complement2(16), DIFF(15) => 
                           complement2(15), DIFF(14) => complement2(14), 
                           DIFF(13) => complement2(13), DIFF(12) => 
                           complement2(12), DIFF(11) => complement2(11), 
                           DIFF(10) => complement2(10), DIFF(9) => 
                           complement2(9), DIFF(8) => complement2(8), DIFF(7) 
                           => complement2(7), DIFF(6) => complement2(6), 
                           DIFF(5) => complement2(5), DIFF(4) => complement2(4)
                           , DIFF(3) => complement2(3), DIFF(2) => 
                           complement2(2), DIFF(1) => complement2(1), DIFF(0) 
                           => complement2(0), CO => n_3135);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_25 is

   port( input : in std_logic_vector (63 downto 0);  complement2 : out 
         std_logic_vector (63 downto 0));

end complementer_N64_25;

architecture SYN_beh of complementer_N64_25 is

   component complementer_N64_25_DW01_sub_0
      port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (63 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n2, n_3136 : std_logic;

begin
   
   n1 <= '0';
   n2 <= '0';
   sub_add_29_b0 : complementer_N64_25_DW01_sub_0 port map( A(63) => n1, A(62) 
                           => n1, A(61) => n1, A(60) => n1, A(59) => n1, A(58) 
                           => n1, A(57) => n1, A(56) => n1, A(55) => n1, A(54) 
                           => n1, A(53) => n1, A(52) => n1, A(51) => n1, A(50) 
                           => n1, A(49) => n1, A(48) => n1, A(47) => n1, A(46) 
                           => n1, A(45) => n1, A(44) => n1, A(43) => n1, A(42) 
                           => n1, A(41) => n1, A(40) => n1, A(39) => n1, A(38) 
                           => n1, A(37) => n1, A(36) => n1, A(35) => n1, A(34) 
                           => n1, A(33) => n1, A(32) => n1, A(31) => n1, A(30) 
                           => n1, A(29) => n1, A(28) => n1, A(27) => n1, A(26) 
                           => n1, A(25) => n1, A(24) => n1, A(23) => n1, A(22) 
                           => n1, A(21) => n1, A(20) => n1, A(19) => n1, A(18) 
                           => n1, A(17) => n1, A(16) => n1, A(15) => n1, A(14) 
                           => n1, A(13) => n1, A(12) => n1, A(11) => n1, A(10) 
                           => n1, A(9) => n1, A(8) => n1, A(7) => n1, A(6) => 
                           n1, A(5) => n1, A(4) => n1, A(3) => n1, A(2) => n1, 
                           A(1) => n1, A(0) => n2, B(63) => input(63), B(62) =>
                           input(62), B(61) => input(61), B(60) => input(60), 
                           B(59) => input(59), B(58) => input(58), B(57) => 
                           input(57), B(56) => input(56), B(55) => input(55), 
                           B(54) => input(54), B(53) => input(53), B(52) => 
                           input(52), B(51) => input(51), B(50) => input(50), 
                           B(49) => input(49), B(48) => input(48), B(47) => 
                           input(47), B(46) => input(46), B(45) => input(45), 
                           B(44) => input(44), B(43) => input(43), B(42) => 
                           input(42), B(41) => input(41), B(40) => input(40), 
                           B(39) => input(39), B(38) => input(38), B(37) => 
                           input(37), B(36) => input(36), B(35) => input(35), 
                           B(34) => input(34), B(33) => input(33), B(32) => 
                           input(32), B(31) => input(31), B(30) => input(30), 
                           B(29) => input(29), B(28) => input(28), B(27) => 
                           input(27), B(26) => input(26), B(25) => input(25), 
                           B(24) => input(24), B(23) => input(23), B(22) => 
                           input(22), B(21) => input(21), B(20) => input(20), 
                           B(19) => input(19), B(18) => input(18), B(17) => 
                           input(17), B(16) => input(16), B(15) => input(15), 
                           B(14) => input(14), B(13) => input(13), B(12) => 
                           input(12), B(11) => input(11), B(10) => input(10), 
                           B(9) => input(9), B(8) => input(8), B(7) => input(7)
                           , B(6) => input(6), B(5) => input(5), B(4) => 
                           input(4), B(3) => input(3), B(2) => input(2), B(1) 
                           => input(1), B(0) => input(0), CI => n1, DIFF(63) =>
                           complement2(63), DIFF(62) => complement2(62), 
                           DIFF(61) => complement2(61), DIFF(60) => 
                           complement2(60), DIFF(59) => complement2(59), 
                           DIFF(58) => complement2(58), DIFF(57) => 
                           complement2(57), DIFF(56) => complement2(56), 
                           DIFF(55) => complement2(55), DIFF(54) => 
                           complement2(54), DIFF(53) => complement2(53), 
                           DIFF(52) => complement2(52), DIFF(51) => 
                           complement2(51), DIFF(50) => complement2(50), 
                           DIFF(49) => complement2(49), DIFF(48) => 
                           complement2(48), DIFF(47) => complement2(47), 
                           DIFF(46) => complement2(46), DIFF(45) => 
                           complement2(45), DIFF(44) => complement2(44), 
                           DIFF(43) => complement2(43), DIFF(42) => 
                           complement2(42), DIFF(41) => complement2(41), 
                           DIFF(40) => complement2(40), DIFF(39) => 
                           complement2(39), DIFF(38) => complement2(38), 
                           DIFF(37) => complement2(37), DIFF(36) => 
                           complement2(36), DIFF(35) => complement2(35), 
                           DIFF(34) => complement2(34), DIFF(33) => 
                           complement2(33), DIFF(32) => complement2(32), 
                           DIFF(31) => complement2(31), DIFF(30) => 
                           complement2(30), DIFF(29) => complement2(29), 
                           DIFF(28) => complement2(28), DIFF(27) => 
                           complement2(27), DIFF(26) => complement2(26), 
                           DIFF(25) => complement2(25), DIFF(24) => 
                           complement2(24), DIFF(23) => complement2(23), 
                           DIFF(22) => complement2(22), DIFF(21) => 
                           complement2(21), DIFF(20) => complement2(20), 
                           DIFF(19) => complement2(19), DIFF(18) => 
                           complement2(18), DIFF(17) => complement2(17), 
                           DIFF(16) => complement2(16), DIFF(15) => 
                           complement2(15), DIFF(14) => complement2(14), 
                           DIFF(13) => complement2(13), DIFF(12) => 
                           complement2(12), DIFF(11) => complement2(11), 
                           DIFF(10) => complement2(10), DIFF(9) => 
                           complement2(9), DIFF(8) => complement2(8), DIFF(7) 
                           => complement2(7), DIFF(6) => complement2(6), 
                           DIFF(5) => complement2(5), DIFF(4) => complement2(4)
                           , DIFF(3) => complement2(3), DIFF(2) => 
                           complement2(2), DIFF(1) => complement2(1), DIFF(0) 
                           => complement2(0), CO => n_3136);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_26 is

   port( input : in std_logic_vector (63 downto 0);  complement2 : out 
         std_logic_vector (63 downto 0));

end complementer_N64_26;

architecture SYN_beh of complementer_N64_26 is

   component complementer_N64_26_DW01_sub_0
      port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (63 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n2, n_3137 : std_logic;

begin
   
   n1 <= '0';
   n2 <= '0';
   sub_add_29_b0 : complementer_N64_26_DW01_sub_0 port map( A(63) => n1, A(62) 
                           => n1, A(61) => n1, A(60) => n1, A(59) => n1, A(58) 
                           => n1, A(57) => n1, A(56) => n1, A(55) => n1, A(54) 
                           => n1, A(53) => n1, A(52) => n1, A(51) => n1, A(50) 
                           => n1, A(49) => n1, A(48) => n1, A(47) => n1, A(46) 
                           => n1, A(45) => n1, A(44) => n1, A(43) => n1, A(42) 
                           => n1, A(41) => n1, A(40) => n1, A(39) => n1, A(38) 
                           => n1, A(37) => n1, A(36) => n1, A(35) => n1, A(34) 
                           => n1, A(33) => n1, A(32) => n1, A(31) => n1, A(30) 
                           => n1, A(29) => n1, A(28) => n1, A(27) => n1, A(26) 
                           => n1, A(25) => n1, A(24) => n1, A(23) => n1, A(22) 
                           => n1, A(21) => n1, A(20) => n1, A(19) => n1, A(18) 
                           => n1, A(17) => n1, A(16) => n1, A(15) => n1, A(14) 
                           => n1, A(13) => n1, A(12) => n1, A(11) => n1, A(10) 
                           => n1, A(9) => n1, A(8) => n1, A(7) => n1, A(6) => 
                           n1, A(5) => n1, A(4) => n1, A(3) => n1, A(2) => n1, 
                           A(1) => n1, A(0) => n2, B(63) => input(63), B(62) =>
                           input(62), B(61) => input(61), B(60) => input(60), 
                           B(59) => input(59), B(58) => input(58), B(57) => 
                           input(57), B(56) => input(56), B(55) => input(55), 
                           B(54) => input(54), B(53) => input(53), B(52) => 
                           input(52), B(51) => input(51), B(50) => input(50), 
                           B(49) => input(49), B(48) => input(48), B(47) => 
                           input(47), B(46) => input(46), B(45) => input(45), 
                           B(44) => input(44), B(43) => input(43), B(42) => 
                           input(42), B(41) => input(41), B(40) => input(40), 
                           B(39) => input(39), B(38) => input(38), B(37) => 
                           input(37), B(36) => input(36), B(35) => input(35), 
                           B(34) => input(34), B(33) => input(33), B(32) => 
                           input(32), B(31) => input(31), B(30) => input(30), 
                           B(29) => input(29), B(28) => input(28), B(27) => 
                           input(27), B(26) => input(26), B(25) => input(25), 
                           B(24) => input(24), B(23) => input(23), B(22) => 
                           input(22), B(21) => input(21), B(20) => input(20), 
                           B(19) => input(19), B(18) => input(18), B(17) => 
                           input(17), B(16) => input(16), B(15) => input(15), 
                           B(14) => input(14), B(13) => input(13), B(12) => 
                           input(12), B(11) => input(11), B(10) => input(10), 
                           B(9) => input(9), B(8) => input(8), B(7) => input(7)
                           , B(6) => input(6), B(5) => input(5), B(4) => 
                           input(4), B(3) => input(3), B(2) => input(2), B(1) 
                           => input(1), B(0) => input(0), CI => n1, DIFF(63) =>
                           complement2(63), DIFF(62) => complement2(62), 
                           DIFF(61) => complement2(61), DIFF(60) => 
                           complement2(60), DIFF(59) => complement2(59), 
                           DIFF(58) => complement2(58), DIFF(57) => 
                           complement2(57), DIFF(56) => complement2(56), 
                           DIFF(55) => complement2(55), DIFF(54) => 
                           complement2(54), DIFF(53) => complement2(53), 
                           DIFF(52) => complement2(52), DIFF(51) => 
                           complement2(51), DIFF(50) => complement2(50), 
                           DIFF(49) => complement2(49), DIFF(48) => 
                           complement2(48), DIFF(47) => complement2(47), 
                           DIFF(46) => complement2(46), DIFF(45) => 
                           complement2(45), DIFF(44) => complement2(44), 
                           DIFF(43) => complement2(43), DIFF(42) => 
                           complement2(42), DIFF(41) => complement2(41), 
                           DIFF(40) => complement2(40), DIFF(39) => 
                           complement2(39), DIFF(38) => complement2(38), 
                           DIFF(37) => complement2(37), DIFF(36) => 
                           complement2(36), DIFF(35) => complement2(35), 
                           DIFF(34) => complement2(34), DIFF(33) => 
                           complement2(33), DIFF(32) => complement2(32), 
                           DIFF(31) => complement2(31), DIFF(30) => 
                           complement2(30), DIFF(29) => complement2(29), 
                           DIFF(28) => complement2(28), DIFF(27) => 
                           complement2(27), DIFF(26) => complement2(26), 
                           DIFF(25) => complement2(25), DIFF(24) => 
                           complement2(24), DIFF(23) => complement2(23), 
                           DIFF(22) => complement2(22), DIFF(21) => 
                           complement2(21), DIFF(20) => complement2(20), 
                           DIFF(19) => complement2(19), DIFF(18) => 
                           complement2(18), DIFF(17) => complement2(17), 
                           DIFF(16) => complement2(16), DIFF(15) => 
                           complement2(15), DIFF(14) => complement2(14), 
                           DIFF(13) => complement2(13), DIFF(12) => 
                           complement2(12), DIFF(11) => complement2(11), 
                           DIFF(10) => complement2(10), DIFF(9) => 
                           complement2(9), DIFF(8) => complement2(8), DIFF(7) 
                           => complement2(7), DIFF(6) => complement2(6), 
                           DIFF(5) => complement2(5), DIFF(4) => complement2(4)
                           , DIFF(3) => complement2(3), DIFF(2) => 
                           complement2(2), DIFF(1) => complement2(1), DIFF(0) 
                           => complement2(0), CO => n_3137);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_27 is

   port( input : in std_logic_vector (63 downto 0);  complement2 : out 
         std_logic_vector (63 downto 0));

end complementer_N64_27;

architecture SYN_beh of complementer_N64_27 is

   component complementer_N64_27_DW01_sub_0
      port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (63 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n2, n_3138 : std_logic;

begin
   
   n1 <= '0';
   n2 <= '0';
   sub_add_29_b0 : complementer_N64_27_DW01_sub_0 port map( A(63) => n1, A(62) 
                           => n1, A(61) => n1, A(60) => n1, A(59) => n1, A(58) 
                           => n1, A(57) => n1, A(56) => n1, A(55) => n1, A(54) 
                           => n1, A(53) => n1, A(52) => n1, A(51) => n1, A(50) 
                           => n1, A(49) => n1, A(48) => n1, A(47) => n1, A(46) 
                           => n1, A(45) => n1, A(44) => n1, A(43) => n1, A(42) 
                           => n1, A(41) => n1, A(40) => n1, A(39) => n1, A(38) 
                           => n1, A(37) => n1, A(36) => n1, A(35) => n1, A(34) 
                           => n1, A(33) => n1, A(32) => n1, A(31) => n1, A(30) 
                           => n1, A(29) => n1, A(28) => n1, A(27) => n1, A(26) 
                           => n1, A(25) => n1, A(24) => n1, A(23) => n1, A(22) 
                           => n1, A(21) => n1, A(20) => n1, A(19) => n1, A(18) 
                           => n1, A(17) => n1, A(16) => n1, A(15) => n1, A(14) 
                           => n1, A(13) => n1, A(12) => n1, A(11) => n1, A(10) 
                           => n1, A(9) => n1, A(8) => n1, A(7) => n1, A(6) => 
                           n1, A(5) => n1, A(4) => n1, A(3) => n1, A(2) => n1, 
                           A(1) => n1, A(0) => n2, B(63) => input(63), B(62) =>
                           input(62), B(61) => input(61), B(60) => input(60), 
                           B(59) => input(59), B(58) => input(58), B(57) => 
                           input(57), B(56) => input(56), B(55) => input(55), 
                           B(54) => input(54), B(53) => input(53), B(52) => 
                           input(52), B(51) => input(51), B(50) => input(50), 
                           B(49) => input(49), B(48) => input(48), B(47) => 
                           input(47), B(46) => input(46), B(45) => input(45), 
                           B(44) => input(44), B(43) => input(43), B(42) => 
                           input(42), B(41) => input(41), B(40) => input(40), 
                           B(39) => input(39), B(38) => input(38), B(37) => 
                           input(37), B(36) => input(36), B(35) => input(35), 
                           B(34) => input(34), B(33) => input(33), B(32) => 
                           input(32), B(31) => input(31), B(30) => input(30), 
                           B(29) => input(29), B(28) => input(28), B(27) => 
                           input(27), B(26) => input(26), B(25) => input(25), 
                           B(24) => input(24), B(23) => input(23), B(22) => 
                           input(22), B(21) => input(21), B(20) => input(20), 
                           B(19) => input(19), B(18) => input(18), B(17) => 
                           input(17), B(16) => input(16), B(15) => input(15), 
                           B(14) => input(14), B(13) => input(13), B(12) => 
                           input(12), B(11) => input(11), B(10) => input(10), 
                           B(9) => input(9), B(8) => input(8), B(7) => input(7)
                           , B(6) => input(6), B(5) => input(5), B(4) => 
                           input(4), B(3) => input(3), B(2) => input(2), B(1) 
                           => input(1), B(0) => input(0), CI => n1, DIFF(63) =>
                           complement2(63), DIFF(62) => complement2(62), 
                           DIFF(61) => complement2(61), DIFF(60) => 
                           complement2(60), DIFF(59) => complement2(59), 
                           DIFF(58) => complement2(58), DIFF(57) => 
                           complement2(57), DIFF(56) => complement2(56), 
                           DIFF(55) => complement2(55), DIFF(54) => 
                           complement2(54), DIFF(53) => complement2(53), 
                           DIFF(52) => complement2(52), DIFF(51) => 
                           complement2(51), DIFF(50) => complement2(50), 
                           DIFF(49) => complement2(49), DIFF(48) => 
                           complement2(48), DIFF(47) => complement2(47), 
                           DIFF(46) => complement2(46), DIFF(45) => 
                           complement2(45), DIFF(44) => complement2(44), 
                           DIFF(43) => complement2(43), DIFF(42) => 
                           complement2(42), DIFF(41) => complement2(41), 
                           DIFF(40) => complement2(40), DIFF(39) => 
                           complement2(39), DIFF(38) => complement2(38), 
                           DIFF(37) => complement2(37), DIFF(36) => 
                           complement2(36), DIFF(35) => complement2(35), 
                           DIFF(34) => complement2(34), DIFF(33) => 
                           complement2(33), DIFF(32) => complement2(32), 
                           DIFF(31) => complement2(31), DIFF(30) => 
                           complement2(30), DIFF(29) => complement2(29), 
                           DIFF(28) => complement2(28), DIFF(27) => 
                           complement2(27), DIFF(26) => complement2(26), 
                           DIFF(25) => complement2(25), DIFF(24) => 
                           complement2(24), DIFF(23) => complement2(23), 
                           DIFF(22) => complement2(22), DIFF(21) => 
                           complement2(21), DIFF(20) => complement2(20), 
                           DIFF(19) => complement2(19), DIFF(18) => 
                           complement2(18), DIFF(17) => complement2(17), 
                           DIFF(16) => complement2(16), DIFF(15) => 
                           complement2(15), DIFF(14) => complement2(14), 
                           DIFF(13) => complement2(13), DIFF(12) => 
                           complement2(12), DIFF(11) => complement2(11), 
                           DIFF(10) => complement2(10), DIFF(9) => 
                           complement2(9), DIFF(8) => complement2(8), DIFF(7) 
                           => complement2(7), DIFF(6) => complement2(6), 
                           DIFF(5) => complement2(5), DIFF(4) => complement2(4)
                           , DIFF(3) => complement2(3), DIFF(2) => 
                           complement2(2), DIFF(1) => complement2(1), DIFF(0) 
                           => complement2(0), CO => n_3138);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_28 is

   port( input : in std_logic_vector (63 downto 0);  complement2 : out 
         std_logic_vector (63 downto 0));

end complementer_N64_28;

architecture SYN_beh of complementer_N64_28 is

   component complementer_N64_28_DW01_sub_0
      port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (63 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n2, n_3139 : std_logic;

begin
   
   n1 <= '0';
   n2 <= '0';
   sub_add_29_b0 : complementer_N64_28_DW01_sub_0 port map( A(63) => n1, A(62) 
                           => n1, A(61) => n1, A(60) => n1, A(59) => n1, A(58) 
                           => n1, A(57) => n1, A(56) => n1, A(55) => n1, A(54) 
                           => n1, A(53) => n1, A(52) => n1, A(51) => n1, A(50) 
                           => n1, A(49) => n1, A(48) => n1, A(47) => n1, A(46) 
                           => n1, A(45) => n1, A(44) => n1, A(43) => n1, A(42) 
                           => n1, A(41) => n1, A(40) => n1, A(39) => n1, A(38) 
                           => n1, A(37) => n1, A(36) => n1, A(35) => n1, A(34) 
                           => n1, A(33) => n1, A(32) => n1, A(31) => n1, A(30) 
                           => n1, A(29) => n1, A(28) => n1, A(27) => n1, A(26) 
                           => n1, A(25) => n1, A(24) => n1, A(23) => n1, A(22) 
                           => n1, A(21) => n1, A(20) => n1, A(19) => n1, A(18) 
                           => n1, A(17) => n1, A(16) => n1, A(15) => n1, A(14) 
                           => n1, A(13) => n1, A(12) => n1, A(11) => n1, A(10) 
                           => n1, A(9) => n1, A(8) => n1, A(7) => n1, A(6) => 
                           n1, A(5) => n1, A(4) => n1, A(3) => n1, A(2) => n1, 
                           A(1) => n1, A(0) => n2, B(63) => input(63), B(62) =>
                           input(62), B(61) => input(61), B(60) => input(60), 
                           B(59) => input(59), B(58) => input(58), B(57) => 
                           input(57), B(56) => input(56), B(55) => input(55), 
                           B(54) => input(54), B(53) => input(53), B(52) => 
                           input(52), B(51) => input(51), B(50) => input(50), 
                           B(49) => input(49), B(48) => input(48), B(47) => 
                           input(47), B(46) => input(46), B(45) => input(45), 
                           B(44) => input(44), B(43) => input(43), B(42) => 
                           input(42), B(41) => input(41), B(40) => input(40), 
                           B(39) => input(39), B(38) => input(38), B(37) => 
                           input(37), B(36) => input(36), B(35) => input(35), 
                           B(34) => input(34), B(33) => input(33), B(32) => 
                           input(32), B(31) => input(31), B(30) => input(30), 
                           B(29) => input(29), B(28) => input(28), B(27) => 
                           input(27), B(26) => input(26), B(25) => input(25), 
                           B(24) => input(24), B(23) => input(23), B(22) => 
                           input(22), B(21) => input(21), B(20) => input(20), 
                           B(19) => input(19), B(18) => input(18), B(17) => 
                           input(17), B(16) => input(16), B(15) => input(15), 
                           B(14) => input(14), B(13) => input(13), B(12) => 
                           input(12), B(11) => input(11), B(10) => input(10), 
                           B(9) => input(9), B(8) => input(8), B(7) => input(7)
                           , B(6) => input(6), B(5) => input(5), B(4) => 
                           input(4), B(3) => input(3), B(2) => input(2), B(1) 
                           => input(1), B(0) => input(0), CI => n1, DIFF(63) =>
                           complement2(63), DIFF(62) => complement2(62), 
                           DIFF(61) => complement2(61), DIFF(60) => 
                           complement2(60), DIFF(59) => complement2(59), 
                           DIFF(58) => complement2(58), DIFF(57) => 
                           complement2(57), DIFF(56) => complement2(56), 
                           DIFF(55) => complement2(55), DIFF(54) => 
                           complement2(54), DIFF(53) => complement2(53), 
                           DIFF(52) => complement2(52), DIFF(51) => 
                           complement2(51), DIFF(50) => complement2(50), 
                           DIFF(49) => complement2(49), DIFF(48) => 
                           complement2(48), DIFF(47) => complement2(47), 
                           DIFF(46) => complement2(46), DIFF(45) => 
                           complement2(45), DIFF(44) => complement2(44), 
                           DIFF(43) => complement2(43), DIFF(42) => 
                           complement2(42), DIFF(41) => complement2(41), 
                           DIFF(40) => complement2(40), DIFF(39) => 
                           complement2(39), DIFF(38) => complement2(38), 
                           DIFF(37) => complement2(37), DIFF(36) => 
                           complement2(36), DIFF(35) => complement2(35), 
                           DIFF(34) => complement2(34), DIFF(33) => 
                           complement2(33), DIFF(32) => complement2(32), 
                           DIFF(31) => complement2(31), DIFF(30) => 
                           complement2(30), DIFF(29) => complement2(29), 
                           DIFF(28) => complement2(28), DIFF(27) => 
                           complement2(27), DIFF(26) => complement2(26), 
                           DIFF(25) => complement2(25), DIFF(24) => 
                           complement2(24), DIFF(23) => complement2(23), 
                           DIFF(22) => complement2(22), DIFF(21) => 
                           complement2(21), DIFF(20) => complement2(20), 
                           DIFF(19) => complement2(19), DIFF(18) => 
                           complement2(18), DIFF(17) => complement2(17), 
                           DIFF(16) => complement2(16), DIFF(15) => 
                           complement2(15), DIFF(14) => complement2(14), 
                           DIFF(13) => complement2(13), DIFF(12) => 
                           complement2(12), DIFF(11) => complement2(11), 
                           DIFF(10) => complement2(10), DIFF(9) => 
                           complement2(9), DIFF(8) => complement2(8), DIFF(7) 
                           => complement2(7), DIFF(6) => complement2(6), 
                           DIFF(5) => complement2(5), DIFF(4) => complement2(4)
                           , DIFF(3) => complement2(3), DIFF(2) => 
                           complement2(2), DIFF(1) => complement2(1), DIFF(0) 
                           => complement2(0), CO => n_3139);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity FA_0 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_0;

architecture SYN_BEHAVIORAL of FA_0 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n2, n4 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n3, B2 => Ci, ZN => n2);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U5 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_29 is

   port( input : in std_logic_vector (63 downto 0);  complement2 : out 
         std_logic_vector (63 downto 0));

end complementer_N64_29;

architecture SYN_beh of complementer_N64_29 is

   component complementer_N64_29_DW01_sub_0
      port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (63 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n2, n_3140 : std_logic;

begin
   
   n1 <= '0';
   n2 <= '0';
   sub_add_29_b0 : complementer_N64_29_DW01_sub_0 port map( A(63) => n1, A(62) 
                           => n1, A(61) => n1, A(60) => n1, A(59) => n1, A(58) 
                           => n1, A(57) => n1, A(56) => n1, A(55) => n1, A(54) 
                           => n1, A(53) => n1, A(52) => n1, A(51) => n1, A(50) 
                           => n1, A(49) => n1, A(48) => n1, A(47) => n1, A(46) 
                           => n1, A(45) => n1, A(44) => n1, A(43) => n1, A(42) 
                           => n1, A(41) => n1, A(40) => n1, A(39) => n1, A(38) 
                           => n1, A(37) => n1, A(36) => n1, A(35) => n1, A(34) 
                           => n1, A(33) => n1, A(32) => n1, A(31) => n1, A(30) 
                           => n1, A(29) => n1, A(28) => n1, A(27) => n1, A(26) 
                           => n1, A(25) => n1, A(24) => n1, A(23) => n1, A(22) 
                           => n1, A(21) => n1, A(20) => n1, A(19) => n1, A(18) 
                           => n1, A(17) => n1, A(16) => n1, A(15) => n1, A(14) 
                           => n1, A(13) => n1, A(12) => n1, A(11) => n1, A(10) 
                           => n1, A(9) => n1, A(8) => n1, A(7) => n1, A(6) => 
                           n1, A(5) => n1, A(4) => n1, A(3) => n1, A(2) => n1, 
                           A(1) => n1, A(0) => n2, B(63) => input(63), B(62) =>
                           input(62), B(61) => input(61), B(60) => input(60), 
                           B(59) => input(59), B(58) => input(58), B(57) => 
                           input(57), B(56) => input(56), B(55) => input(55), 
                           B(54) => input(54), B(53) => input(53), B(52) => 
                           input(52), B(51) => input(51), B(50) => input(50), 
                           B(49) => input(49), B(48) => input(48), B(47) => 
                           input(47), B(46) => input(46), B(45) => input(45), 
                           B(44) => input(44), B(43) => input(43), B(42) => 
                           input(42), B(41) => input(41), B(40) => input(40), 
                           B(39) => input(39), B(38) => input(38), B(37) => 
                           input(37), B(36) => input(36), B(35) => input(35), 
                           B(34) => input(34), B(33) => input(33), B(32) => 
                           input(32), B(31) => input(31), B(30) => input(30), 
                           B(29) => input(29), B(28) => input(28), B(27) => 
                           input(27), B(26) => input(26), B(25) => input(25), 
                           B(24) => input(24), B(23) => input(23), B(22) => 
                           input(22), B(21) => input(21), B(20) => input(20), 
                           B(19) => input(19), B(18) => input(18), B(17) => 
                           input(17), B(16) => input(16), B(15) => input(15), 
                           B(14) => input(14), B(13) => input(13), B(12) => 
                           input(12), B(11) => input(11), B(10) => input(10), 
                           B(9) => input(9), B(8) => input(8), B(7) => input(7)
                           , B(6) => input(6), B(5) => input(5), B(4) => 
                           input(4), B(3) => input(3), B(2) => input(2), B(1) 
                           => input(1), B(0) => input(0), CI => n1, DIFF(63) =>
                           complement2(63), DIFF(62) => complement2(62), 
                           DIFF(61) => complement2(61), DIFF(60) => 
                           complement2(60), DIFF(59) => complement2(59), 
                           DIFF(58) => complement2(58), DIFF(57) => 
                           complement2(57), DIFF(56) => complement2(56), 
                           DIFF(55) => complement2(55), DIFF(54) => 
                           complement2(54), DIFF(53) => complement2(53), 
                           DIFF(52) => complement2(52), DIFF(51) => 
                           complement2(51), DIFF(50) => complement2(50), 
                           DIFF(49) => complement2(49), DIFF(48) => 
                           complement2(48), DIFF(47) => complement2(47), 
                           DIFF(46) => complement2(46), DIFF(45) => 
                           complement2(45), DIFF(44) => complement2(44), 
                           DIFF(43) => complement2(43), DIFF(42) => 
                           complement2(42), DIFF(41) => complement2(41), 
                           DIFF(40) => complement2(40), DIFF(39) => 
                           complement2(39), DIFF(38) => complement2(38), 
                           DIFF(37) => complement2(37), DIFF(36) => 
                           complement2(36), DIFF(35) => complement2(35), 
                           DIFF(34) => complement2(34), DIFF(33) => 
                           complement2(33), DIFF(32) => complement2(32), 
                           DIFF(31) => complement2(31), DIFF(30) => 
                           complement2(30), DIFF(29) => complement2(29), 
                           DIFF(28) => complement2(28), DIFF(27) => 
                           complement2(27), DIFF(26) => complement2(26), 
                           DIFF(25) => complement2(25), DIFF(24) => 
                           complement2(24), DIFF(23) => complement2(23), 
                           DIFF(22) => complement2(22), DIFF(21) => 
                           complement2(21), DIFF(20) => complement2(20), 
                           DIFF(19) => complement2(19), DIFF(18) => 
                           complement2(18), DIFF(17) => complement2(17), 
                           DIFF(16) => complement2(16), DIFF(15) => 
                           complement2(15), DIFF(14) => complement2(14), 
                           DIFF(13) => complement2(13), DIFF(12) => 
                           complement2(12), DIFF(11) => complement2(11), 
                           DIFF(10) => complement2(10), DIFF(9) => 
                           complement2(9), DIFF(8) => complement2(8), DIFF(7) 
                           => complement2(7), DIFF(6) => complement2(6), 
                           DIFF(5) => complement2(5), DIFF(4) => complement2(4)
                           , DIFF(3) => complement2(3), DIFF(2) => 
                           complement2(2), DIFF(1) => complement2(1), DIFF(0) 
                           => complement2(0), CO => n_3140);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_30 is

   port( input : in std_logic_vector (63 downto 0);  complement2 : out 
         std_logic_vector (63 downto 0));

end complementer_N64_30;

architecture SYN_beh of complementer_N64_30 is

   component complementer_N64_30_DW01_sub_0
      port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (63 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n2, n_3141 : std_logic;

begin
   
   n1 <= '0';
   n2 <= '0';
   sub_add_29_b0 : complementer_N64_30_DW01_sub_0 port map( A(63) => n1, A(62) 
                           => n1, A(61) => n1, A(60) => n1, A(59) => n1, A(58) 
                           => n1, A(57) => n1, A(56) => n1, A(55) => n1, A(54) 
                           => n1, A(53) => n1, A(52) => n1, A(51) => n1, A(50) 
                           => n1, A(49) => n1, A(48) => n1, A(47) => n1, A(46) 
                           => n1, A(45) => n1, A(44) => n1, A(43) => n1, A(42) 
                           => n1, A(41) => n1, A(40) => n1, A(39) => n1, A(38) 
                           => n1, A(37) => n1, A(36) => n1, A(35) => n1, A(34) 
                           => n1, A(33) => n1, A(32) => n1, A(31) => n1, A(30) 
                           => n1, A(29) => n1, A(28) => n1, A(27) => n1, A(26) 
                           => n1, A(25) => n1, A(24) => n1, A(23) => n1, A(22) 
                           => n1, A(21) => n1, A(20) => n1, A(19) => n1, A(18) 
                           => n1, A(17) => n1, A(16) => n1, A(15) => n1, A(14) 
                           => n1, A(13) => n1, A(12) => n1, A(11) => n1, A(10) 
                           => n1, A(9) => n1, A(8) => n1, A(7) => n1, A(6) => 
                           n1, A(5) => n1, A(4) => n1, A(3) => n1, A(2) => n1, 
                           A(1) => n1, A(0) => n2, B(63) => input(63), B(62) =>
                           input(62), B(61) => input(61), B(60) => input(60), 
                           B(59) => input(59), B(58) => input(58), B(57) => 
                           input(57), B(56) => input(56), B(55) => input(55), 
                           B(54) => input(54), B(53) => input(53), B(52) => 
                           input(52), B(51) => input(51), B(50) => input(50), 
                           B(49) => input(49), B(48) => input(48), B(47) => 
                           input(47), B(46) => input(46), B(45) => input(45), 
                           B(44) => input(44), B(43) => input(43), B(42) => 
                           input(42), B(41) => input(41), B(40) => input(40), 
                           B(39) => input(39), B(38) => input(38), B(37) => 
                           input(37), B(36) => input(36), B(35) => input(35), 
                           B(34) => input(34), B(33) => input(33), B(32) => 
                           input(32), B(31) => input(31), B(30) => input(30), 
                           B(29) => input(29), B(28) => input(28), B(27) => 
                           input(27), B(26) => input(26), B(25) => input(25), 
                           B(24) => input(24), B(23) => input(23), B(22) => 
                           input(22), B(21) => input(21), B(20) => input(20), 
                           B(19) => input(19), B(18) => input(18), B(17) => 
                           input(17), B(16) => input(16), B(15) => input(15), 
                           B(14) => input(14), B(13) => input(13), B(12) => 
                           input(12), B(11) => input(11), B(10) => input(10), 
                           B(9) => input(9), B(8) => input(8), B(7) => input(7)
                           , B(6) => input(6), B(5) => input(5), B(4) => 
                           input(4), B(3) => input(3), B(2) => input(2), B(1) 
                           => input(1), B(0) => input(0), CI => n1, DIFF(63) =>
                           complement2(63), DIFF(62) => complement2(62), 
                           DIFF(61) => complement2(61), DIFF(60) => 
                           complement2(60), DIFF(59) => complement2(59), 
                           DIFF(58) => complement2(58), DIFF(57) => 
                           complement2(57), DIFF(56) => complement2(56), 
                           DIFF(55) => complement2(55), DIFF(54) => 
                           complement2(54), DIFF(53) => complement2(53), 
                           DIFF(52) => complement2(52), DIFF(51) => 
                           complement2(51), DIFF(50) => complement2(50), 
                           DIFF(49) => complement2(49), DIFF(48) => 
                           complement2(48), DIFF(47) => complement2(47), 
                           DIFF(46) => complement2(46), DIFF(45) => 
                           complement2(45), DIFF(44) => complement2(44), 
                           DIFF(43) => complement2(43), DIFF(42) => 
                           complement2(42), DIFF(41) => complement2(41), 
                           DIFF(40) => complement2(40), DIFF(39) => 
                           complement2(39), DIFF(38) => complement2(38), 
                           DIFF(37) => complement2(37), DIFF(36) => 
                           complement2(36), DIFF(35) => complement2(35), 
                           DIFF(34) => complement2(34), DIFF(33) => 
                           complement2(33), DIFF(32) => complement2(32), 
                           DIFF(31) => complement2(31), DIFF(30) => 
                           complement2(30), DIFF(29) => complement2(29), 
                           DIFF(28) => complement2(28), DIFF(27) => 
                           complement2(27), DIFF(26) => complement2(26), 
                           DIFF(25) => complement2(25), DIFF(24) => 
                           complement2(24), DIFF(23) => complement2(23), 
                           DIFF(22) => complement2(22), DIFF(21) => 
                           complement2(21), DIFF(20) => complement2(20), 
                           DIFF(19) => complement2(19), DIFF(18) => 
                           complement2(18), DIFF(17) => complement2(17), 
                           DIFF(16) => complement2(16), DIFF(15) => 
                           complement2(15), DIFF(14) => complement2(14), 
                           DIFF(13) => complement2(13), DIFF(12) => 
                           complement2(12), DIFF(11) => complement2(11), 
                           DIFF(10) => complement2(10), DIFF(9) => 
                           complement2(9), DIFF(8) => complement2(8), DIFF(7) 
                           => complement2(7), DIFF(6) => complement2(6), 
                           DIFF(5) => complement2(5), DIFF(4) => complement2(4)
                           , DIFF(3) => complement2(3), DIFF(2) => 
                           complement2(2), DIFF(1) => complement2(1), DIFF(0) 
                           => complement2(0), CO => n_3141);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_31 is

   port( input : in std_logic_vector (63 downto 0);  complement2 : out 
         std_logic_vector (63 downto 0));

end complementer_N64_31;

architecture SYN_beh of complementer_N64_31 is

   component complementer_N64_31_DW01_sub_0
      port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (63 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n2, n_3142 : std_logic;

begin
   
   n1 <= '0';
   n2 <= '0';
   sub_add_29_b0 : complementer_N64_31_DW01_sub_0 port map( A(63) => n1, A(62) 
                           => n1, A(61) => n1, A(60) => n1, A(59) => n1, A(58) 
                           => n1, A(57) => n1, A(56) => n1, A(55) => n1, A(54) 
                           => n1, A(53) => n1, A(52) => n1, A(51) => n1, A(50) 
                           => n1, A(49) => n1, A(48) => n1, A(47) => n1, A(46) 
                           => n1, A(45) => n1, A(44) => n1, A(43) => n1, A(42) 
                           => n1, A(41) => n1, A(40) => n1, A(39) => n1, A(38) 
                           => n1, A(37) => n1, A(36) => n1, A(35) => n1, A(34) 
                           => n1, A(33) => n1, A(32) => n1, A(31) => n1, A(30) 
                           => n1, A(29) => n1, A(28) => n1, A(27) => n1, A(26) 
                           => n1, A(25) => n1, A(24) => n1, A(23) => n1, A(22) 
                           => n1, A(21) => n1, A(20) => n1, A(19) => n1, A(18) 
                           => n1, A(17) => n1, A(16) => n1, A(15) => n1, A(14) 
                           => n1, A(13) => n1, A(12) => n1, A(11) => n1, A(10) 
                           => n1, A(9) => n1, A(8) => n1, A(7) => n1, A(6) => 
                           n1, A(5) => n1, A(4) => n1, A(3) => n1, A(2) => n1, 
                           A(1) => n1, A(0) => n2, B(63) => input(63), B(62) =>
                           input(62), B(61) => input(61), B(60) => input(60), 
                           B(59) => input(59), B(58) => input(58), B(57) => 
                           input(57), B(56) => input(56), B(55) => input(55), 
                           B(54) => input(54), B(53) => input(53), B(52) => 
                           input(52), B(51) => input(51), B(50) => input(50), 
                           B(49) => input(49), B(48) => input(48), B(47) => 
                           input(47), B(46) => input(46), B(45) => input(45), 
                           B(44) => input(44), B(43) => input(43), B(42) => 
                           input(42), B(41) => input(41), B(40) => input(40), 
                           B(39) => input(39), B(38) => input(38), B(37) => 
                           input(37), B(36) => input(36), B(35) => input(35), 
                           B(34) => input(34), B(33) => input(33), B(32) => 
                           input(32), B(31) => input(31), B(30) => input(30), 
                           B(29) => input(29), B(28) => input(28), B(27) => 
                           input(27), B(26) => input(26), B(25) => input(25), 
                           B(24) => input(24), B(23) => input(23), B(22) => 
                           input(22), B(21) => input(21), B(20) => input(20), 
                           B(19) => input(19), B(18) => input(18), B(17) => 
                           input(17), B(16) => input(16), B(15) => input(15), 
                           B(14) => input(14), B(13) => input(13), B(12) => 
                           input(12), B(11) => input(11), B(10) => input(10), 
                           B(9) => input(9), B(8) => input(8), B(7) => input(7)
                           , B(6) => input(6), B(5) => input(5), B(4) => 
                           input(4), B(3) => input(3), B(2) => input(2), B(1) 
                           => input(1), B(0) => input(0), CI => n1, DIFF(63) =>
                           complement2(63), DIFF(62) => complement2(62), 
                           DIFF(61) => complement2(61), DIFF(60) => 
                           complement2(60), DIFF(59) => complement2(59), 
                           DIFF(58) => complement2(58), DIFF(57) => 
                           complement2(57), DIFF(56) => complement2(56), 
                           DIFF(55) => complement2(55), DIFF(54) => 
                           complement2(54), DIFF(53) => complement2(53), 
                           DIFF(52) => complement2(52), DIFF(51) => 
                           complement2(51), DIFF(50) => complement2(50), 
                           DIFF(49) => complement2(49), DIFF(48) => 
                           complement2(48), DIFF(47) => complement2(47), 
                           DIFF(46) => complement2(46), DIFF(45) => 
                           complement2(45), DIFF(44) => complement2(44), 
                           DIFF(43) => complement2(43), DIFF(42) => 
                           complement2(42), DIFF(41) => complement2(41), 
                           DIFF(40) => complement2(40), DIFF(39) => 
                           complement2(39), DIFF(38) => complement2(38), 
                           DIFF(37) => complement2(37), DIFF(36) => 
                           complement2(36), DIFF(35) => complement2(35), 
                           DIFF(34) => complement2(34), DIFF(33) => 
                           complement2(33), DIFF(32) => complement2(32), 
                           DIFF(31) => complement2(31), DIFF(30) => 
                           complement2(30), DIFF(29) => complement2(29), 
                           DIFF(28) => complement2(28), DIFF(27) => 
                           complement2(27), DIFF(26) => complement2(26), 
                           DIFF(25) => complement2(25), DIFF(24) => 
                           complement2(24), DIFF(23) => complement2(23), 
                           DIFF(22) => complement2(22), DIFF(21) => 
                           complement2(21), DIFF(20) => complement2(20), 
                           DIFF(19) => complement2(19), DIFF(18) => 
                           complement2(18), DIFF(17) => complement2(17), 
                           DIFF(16) => complement2(16), DIFF(15) => 
                           complement2(15), DIFF(14) => complement2(14), 
                           DIFF(13) => complement2(13), DIFF(12) => 
                           complement2(12), DIFF(11) => complement2(11), 
                           DIFF(10) => complement2(10), DIFF(9) => 
                           complement2(9), DIFF(8) => complement2(8), DIFF(7) 
                           => complement2(7), DIFF(6) => complement2(6), 
                           DIFF(5) => complement2(5), DIFF(4) => complement2(4)
                           , DIFF(3) => complement2(3), DIFF(2) => 
                           complement2(2), DIFF(1) => complement2(1), DIFF(0) 
                           => complement2(0), CO => n_3142);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity complementer_N64_0 is

   port( input : in std_logic_vector (63 downto 0);  complement2 : out 
         std_logic_vector (63 downto 0));

end complementer_N64_0;

architecture SYN_beh of complementer_N64_0 is

   component complementer_N64_0_DW01_sub_0
      port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (63 downto 0);  CO : out std_logic);
   end component;
   
   signal n3, n4, n_3143 : std_logic;

begin
   
   n3 <= '0';
   n4 <= '0';
   sub_add_29_b0 : complementer_N64_0_DW01_sub_0 port map( A(63) => n4, A(62) 
                           => n4, A(61) => n4, A(60) => n4, A(59) => n4, A(58) 
                           => n4, A(57) => n4, A(56) => n4, A(55) => n4, A(54) 
                           => n4, A(53) => n4, A(52) => n4, A(51) => n4, A(50) 
                           => n4, A(49) => n4, A(48) => n4, A(47) => n4, A(46) 
                           => n4, A(45) => n4, A(44) => n4, A(43) => n4, A(42) 
                           => n4, A(41) => n4, A(40) => n4, A(39) => n4, A(38) 
                           => n4, A(37) => n4, A(36) => n4, A(35) => n4, A(34) 
                           => n4, A(33) => n4, A(32) => n4, A(31) => n4, A(30) 
                           => n4, A(29) => n4, A(28) => n4, A(27) => n4, A(26) 
                           => n4, A(25) => n4, A(24) => n4, A(23) => n4, A(22) 
                           => n4, A(21) => n4, A(20) => n4, A(19) => n4, A(18) 
                           => n4, A(17) => n4, A(16) => n4, A(15) => n4, A(14) 
                           => n4, A(13) => n4, A(12) => n4, A(11) => n4, A(10) 
                           => n4, A(9) => n4, A(8) => n4, A(7) => n4, A(6) => 
                           n4, A(5) => n4, A(4) => n4, A(3) => n4, A(2) => n4, 
                           A(1) => n4, A(0) => n3, B(63) => input(63), B(62) =>
                           input(62), B(61) => input(61), B(60) => input(60), 
                           B(59) => input(59), B(58) => input(58), B(57) => 
                           input(57), B(56) => input(56), B(55) => input(55), 
                           B(54) => input(54), B(53) => input(53), B(52) => 
                           input(52), B(51) => input(51), B(50) => input(50), 
                           B(49) => input(49), B(48) => input(48), B(47) => 
                           input(47), B(46) => input(46), B(45) => input(45), 
                           B(44) => input(44), B(43) => input(43), B(42) => 
                           input(42), B(41) => input(41), B(40) => input(40), 
                           B(39) => input(39), B(38) => input(38), B(37) => 
                           input(37), B(36) => input(36), B(35) => input(35), 
                           B(34) => input(34), B(33) => input(33), B(32) => 
                           input(32), B(31) => input(31), B(30) => input(30), 
                           B(29) => input(29), B(28) => input(28), B(27) => 
                           input(27), B(26) => input(26), B(25) => input(25), 
                           B(24) => input(24), B(23) => input(23), B(22) => 
                           input(22), B(21) => input(21), B(20) => input(20), 
                           B(19) => input(19), B(18) => input(18), B(17) => 
                           input(17), B(16) => input(16), B(15) => input(15), 
                           B(14) => input(14), B(13) => input(13), B(12) => 
                           input(12), B(11) => input(11), B(10) => input(10), 
                           B(9) => input(9), B(8) => input(8), B(7) => input(7)
                           , B(6) => input(6), B(5) => input(5), B(4) => 
                           input(4), B(3) => input(3), B(2) => input(2), B(1) 
                           => input(1), B(0) => input(0), CI => n4, DIFF(63) =>
                           complement2(63), DIFF(62) => complement2(62), 
                           DIFF(61) => complement2(61), DIFF(60) => 
                           complement2(60), DIFF(59) => complement2(59), 
                           DIFF(58) => complement2(58), DIFF(57) => 
                           complement2(57), DIFF(56) => complement2(56), 
                           DIFF(55) => complement2(55), DIFF(54) => 
                           complement2(54), DIFF(53) => complement2(53), 
                           DIFF(52) => complement2(52), DIFF(51) => 
                           complement2(51), DIFF(50) => complement2(50), 
                           DIFF(49) => complement2(49), DIFF(48) => 
                           complement2(48), DIFF(47) => complement2(47), 
                           DIFF(46) => complement2(46), DIFF(45) => 
                           complement2(45), DIFF(44) => complement2(44), 
                           DIFF(43) => complement2(43), DIFF(42) => 
                           complement2(42), DIFF(41) => complement2(41), 
                           DIFF(40) => complement2(40), DIFF(39) => 
                           complement2(39), DIFF(38) => complement2(38), 
                           DIFF(37) => complement2(37), DIFF(36) => 
                           complement2(36), DIFF(35) => complement2(35), 
                           DIFF(34) => complement2(34), DIFF(33) => 
                           complement2(33), DIFF(32) => complement2(32), 
                           DIFF(31) => complement2(31), DIFF(30) => 
                           complement2(30), DIFF(29) => complement2(29), 
                           DIFF(28) => complement2(28), DIFF(27) => 
                           complement2(27), DIFF(26) => complement2(26), 
                           DIFF(25) => complement2(25), DIFF(24) => 
                           complement2(24), DIFF(23) => complement2(23), 
                           DIFF(22) => complement2(22), DIFF(21) => 
                           complement2(21), DIFF(20) => complement2(20), 
                           DIFF(19) => complement2(19), DIFF(18) => 
                           complement2(18), DIFF(17) => complement2(17), 
                           DIFF(16) => complement2(16), DIFF(15) => 
                           complement2(15), DIFF(14) => complement2(14), 
                           DIFF(13) => complement2(13), DIFF(12) => 
                           complement2(12), DIFF(11) => complement2(11), 
                           DIFF(10) => complement2(10), DIFF(9) => 
                           complement2(9), DIFF(8) => complement2(8), DIFF(7) 
                           => complement2(7), DIFF(6) => complement2(6), 
                           DIFF(5) => complement2(5), DIFF(4) => complement2(4)
                           , DIFF(3) => complement2(3), DIFF(2) => 
                           complement2(2), DIFF(1) => complement2(1), DIFF(0) 
                           => complement2(0), CO => n_3143);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity shifter_N64_0 is

   port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
         std_logic_vector (63 downto 0));

end shifter_N64_0;

architecture SYN_beh of shifter_N64_0 is

signal X_Logic0_port : std_logic;

begin
   shiftLeftOnePos <= ( input(62), input(61), input(60), input(59), input(58), 
      input(57), input(56), input(55), input(54), input(53), input(52), 
      input(51), input(50), input(49), input(48), input(47), input(46), 
      input(45), input(44), input(43), input(42), input(41), input(40), 
      input(39), input(38), input(37), input(36), input(35), input(34), 
      input(33), input(32), input(31), input(30), input(29), input(28), 
      input(27), input(26), input(25), input(24), input(23), input(22), 
      input(21), input(20), input(19), input(18), input(17), input(16), 
      input(15), input(14), input(13), input(12), input(11), input(10), 
      input(9), input(8), input(7), input(6), input(5), input(4), input(3), 
      input(2), input(1), input(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity ShiftnCompl_N64_1 is

   port( plusA : in std_logic_vector (63 downto 0);  plus2A_out, minus2A_out, 
         plus4A_out, minus4A_out : out std_logic_vector (63 downto 0));

end ShiftnCompl_N64_1;

architecture SYN_struct of ShiftnCompl_N64_1 is

   component complementer_N64_1
      port( input : in std_logic_vector (63 downto 0);  complement2 : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component complementer_N64_2
      port( input : in std_logic_vector (63 downto 0);  complement2 : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component shifter_N64_1
      port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component shifter_N64_2
      port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
            std_logic_vector (63 downto 0));
   end component;
   
   signal plus2A_out_63_port, plus2A_out_62_port, plus2A_out_61_port, 
      plus2A_out_60_port, plus2A_out_59_port, plus2A_out_58_port, 
      plus2A_out_57_port, plus2A_out_56_port, plus2A_out_55_port, 
      plus2A_out_54_port, plus2A_out_53_port, plus2A_out_52_port, 
      plus2A_out_51_port, plus2A_out_50_port, plus2A_out_49_port, 
      plus2A_out_48_port, plus2A_out_47_port, plus2A_out_46_port, 
      plus2A_out_45_port, plus2A_out_44_port, plus2A_out_43_port, 
      plus2A_out_42_port, plus2A_out_41_port, plus2A_out_40_port, 
      plus2A_out_39_port, plus2A_out_38_port, plus2A_out_37_port, 
      plus2A_out_36_port, plus2A_out_35_port, plus2A_out_34_port, 
      plus2A_out_33_port, plus2A_out_32_port, plus2A_out_31_port, 
      plus2A_out_30_port, plus2A_out_29_port, plus2A_out_28_port, 
      plus2A_out_27_port, plus2A_out_26_port, plus2A_out_25_port, 
      plus2A_out_24_port, plus2A_out_23_port, plus2A_out_22_port, 
      plus2A_out_21_port, plus2A_out_20_port, plus2A_out_19_port, 
      plus2A_out_18_port, plus2A_out_17_port, plus2A_out_16_port, 
      plus2A_out_15_port, plus2A_out_14_port, plus2A_out_13_port, 
      plus2A_out_12_port, plus2A_out_11_port, plus2A_out_10_port, 
      plus2A_out_9_port, plus2A_out_8_port, plus2A_out_7_port, 
      plus2A_out_6_port, plus2A_out_5_port, plus2A_out_4_port, 
      plus2A_out_3_port, plus2A_out_2_port, plus2A_out_1_port, 
      plus2A_out_0_port, plus4A_out_63_port, plus4A_out_62_port, 
      plus4A_out_61_port, plus4A_out_60_port, plus4A_out_59_port, 
      plus4A_out_58_port, plus4A_out_57_port, plus4A_out_56_port, 
      plus4A_out_55_port, plus4A_out_54_port, plus4A_out_53_port, 
      plus4A_out_52_port, plus4A_out_51_port, plus4A_out_50_port, 
      plus4A_out_49_port, plus4A_out_48_port, plus4A_out_47_port, 
      plus4A_out_46_port, plus4A_out_45_port, plus4A_out_44_port, 
      plus4A_out_43_port, plus4A_out_42_port, plus4A_out_41_port, 
      plus4A_out_40_port, plus4A_out_39_port, plus4A_out_38_port, 
      plus4A_out_37_port, plus4A_out_36_port, plus4A_out_35_port, 
      plus4A_out_34_port, plus4A_out_33_port, plus4A_out_32_port, 
      plus4A_out_31_port, plus4A_out_30_port, plus4A_out_29_port, 
      plus4A_out_28_port, plus4A_out_27_port, plus4A_out_26_port, 
      plus4A_out_25_port, plus4A_out_24_port, plus4A_out_23_port, 
      plus4A_out_22_port, plus4A_out_21_port, plus4A_out_20_port, 
      plus4A_out_19_port, plus4A_out_18_port, plus4A_out_17_port, 
      plus4A_out_16_port, plus4A_out_15_port, plus4A_out_14_port, 
      plus4A_out_13_port, plus4A_out_12_port, plus4A_out_11_port, 
      plus4A_out_10_port, plus4A_out_9_port, plus4A_out_8_port, 
      plus4A_out_7_port, plus4A_out_6_port, plus4A_out_5_port, 
      plus4A_out_4_port, plus4A_out_3_port, plus4A_out_2_port, 
      plus4A_out_1_port, plus4A_out_0_port, n_3144, n_3145 : std_logic;

begin
   plus2A_out <= ( plus2A_out_63_port, plus2A_out_62_port, plus2A_out_61_port, 
      plus2A_out_60_port, plus2A_out_59_port, plus2A_out_58_port, 
      plus2A_out_57_port, plus2A_out_56_port, plus2A_out_55_port, 
      plus2A_out_54_port, plus2A_out_53_port, plus2A_out_52_port, 
      plus2A_out_51_port, plus2A_out_50_port, plus2A_out_49_port, 
      plus2A_out_48_port, plus2A_out_47_port, plus2A_out_46_port, 
      plus2A_out_45_port, plus2A_out_44_port, plus2A_out_43_port, 
      plus2A_out_42_port, plus2A_out_41_port, plus2A_out_40_port, 
      plus2A_out_39_port, plus2A_out_38_port, plus2A_out_37_port, 
      plus2A_out_36_port, plus2A_out_35_port, plus2A_out_34_port, 
      plus2A_out_33_port, plus2A_out_32_port, plus2A_out_31_port, 
      plus2A_out_30_port, plus2A_out_29_port, plus2A_out_28_port, 
      plus2A_out_27_port, plus2A_out_26_port, plus2A_out_25_port, 
      plus2A_out_24_port, plus2A_out_23_port, plus2A_out_22_port, 
      plus2A_out_21_port, plus2A_out_20_port, plus2A_out_19_port, 
      plus2A_out_18_port, plus2A_out_17_port, plus2A_out_16_port, 
      plus2A_out_15_port, plus2A_out_14_port, plus2A_out_13_port, 
      plus2A_out_12_port, plus2A_out_11_port, plus2A_out_10_port, 
      plus2A_out_9_port, plus2A_out_8_port, plus2A_out_7_port, 
      plus2A_out_6_port, plus2A_out_5_port, plus2A_out_4_port, 
      plus2A_out_3_port, plus2A_out_2_port, plus2A_out_1_port, 
      plus2A_out_0_port );
   plus4A_out <= ( plus4A_out_63_port, plus4A_out_62_port, plus4A_out_61_port, 
      plus4A_out_60_port, plus4A_out_59_port, plus4A_out_58_port, 
      plus4A_out_57_port, plus4A_out_56_port, plus4A_out_55_port, 
      plus4A_out_54_port, plus4A_out_53_port, plus4A_out_52_port, 
      plus4A_out_51_port, plus4A_out_50_port, plus4A_out_49_port, 
      plus4A_out_48_port, plus4A_out_47_port, plus4A_out_46_port, 
      plus4A_out_45_port, plus4A_out_44_port, plus4A_out_43_port, 
      plus4A_out_42_port, plus4A_out_41_port, plus4A_out_40_port, 
      plus4A_out_39_port, plus4A_out_38_port, plus4A_out_37_port, 
      plus4A_out_36_port, plus4A_out_35_port, plus4A_out_34_port, 
      plus4A_out_33_port, plus4A_out_32_port, plus4A_out_31_port, 
      plus4A_out_30_port, plus4A_out_29_port, plus4A_out_28_port, 
      plus4A_out_27_port, plus4A_out_26_port, plus4A_out_25_port, 
      plus4A_out_24_port, plus4A_out_23_port, plus4A_out_22_port, 
      plus4A_out_21_port, plus4A_out_20_port, plus4A_out_19_port, 
      plus4A_out_18_port, plus4A_out_17_port, plus4A_out_16_port, 
      plus4A_out_15_port, plus4A_out_14_port, plus4A_out_13_port, 
      plus4A_out_12_port, plus4A_out_11_port, plus4A_out_10_port, 
      plus4A_out_9_port, plus4A_out_8_port, plus4A_out_7_port, 
      plus4A_out_6_port, plus4A_out_5_port, plus4A_out_4_port, 
      plus4A_out_3_port, plus4A_out_2_port, plus4A_out_1_port, 
      plus4A_out_0_port );
   
   plus2A_out_0_port <= '0';
   plus4A_out_0_port <= '0';
   shifter_1 : shifter_N64_2 port map( input(63) => plusA(63), input(62) => 
                           plusA(62), input(61) => plusA(61), input(60) => 
                           plusA(60), input(59) => plusA(59), input(58) => 
                           plusA(58), input(57) => plusA(57), input(56) => 
                           plusA(56), input(55) => plusA(55), input(54) => 
                           plusA(54), input(53) => plusA(53), input(52) => 
                           plusA(52), input(51) => plusA(51), input(50) => 
                           plusA(50), input(49) => plusA(49), input(48) => 
                           plusA(48), input(47) => plusA(47), input(46) => 
                           plusA(46), input(45) => plusA(45), input(44) => 
                           plusA(44), input(43) => plusA(43), input(42) => 
                           plusA(42), input(41) => plusA(41), input(40) => 
                           plusA(40), input(39) => plusA(39), input(38) => 
                           plusA(38), input(37) => plusA(37), input(36) => 
                           plusA(36), input(35) => plusA(35), input(34) => 
                           plusA(34), input(33) => plusA(33), input(32) => 
                           plusA(32), input(31) => plusA(31), input(30) => 
                           plusA(30), input(29) => plusA(29), input(28) => 
                           plusA(28), input(27) => plusA(27), input(26) => 
                           plusA(26), input(25) => plusA(25), input(24) => 
                           plusA(24), input(23) => plusA(23), input(22) => 
                           plusA(22), input(21) => plusA(21), input(20) => 
                           plusA(20), input(19) => plusA(19), input(18) => 
                           plusA(18), input(17) => plusA(17), input(16) => 
                           plusA(16), input(15) => plusA(15), input(14) => 
                           plusA(14), input(13) => plusA(13), input(12) => 
                           plusA(12), input(11) => plusA(11), input(10) => 
                           plusA(10), input(9) => plusA(9), input(8) => 
                           plusA(8), input(7) => plusA(7), input(6) => plusA(6)
                           , input(5) => plusA(5), input(4) => plusA(4), 
                           input(3) => plusA(3), input(2) => plusA(2), input(1)
                           => plusA(1), input(0) => plusA(0), 
                           shiftLeftOnePos(63) => plus2A_out_63_port, 
                           shiftLeftOnePos(62) => plus2A_out_62_port, 
                           shiftLeftOnePos(61) => plus2A_out_61_port, 
                           shiftLeftOnePos(60) => plus2A_out_60_port, 
                           shiftLeftOnePos(59) => plus2A_out_59_port, 
                           shiftLeftOnePos(58) => plus2A_out_58_port, 
                           shiftLeftOnePos(57) => plus2A_out_57_port, 
                           shiftLeftOnePos(56) => plus2A_out_56_port, 
                           shiftLeftOnePos(55) => plus2A_out_55_port, 
                           shiftLeftOnePos(54) => plus2A_out_54_port, 
                           shiftLeftOnePos(53) => plus2A_out_53_port, 
                           shiftLeftOnePos(52) => plus2A_out_52_port, 
                           shiftLeftOnePos(51) => plus2A_out_51_port, 
                           shiftLeftOnePos(50) => plus2A_out_50_port, 
                           shiftLeftOnePos(49) => plus2A_out_49_port, 
                           shiftLeftOnePos(48) => plus2A_out_48_port, 
                           shiftLeftOnePos(47) => plus2A_out_47_port, 
                           shiftLeftOnePos(46) => plus2A_out_46_port, 
                           shiftLeftOnePos(45) => plus2A_out_45_port, 
                           shiftLeftOnePos(44) => plus2A_out_44_port, 
                           shiftLeftOnePos(43) => plus2A_out_43_port, 
                           shiftLeftOnePos(42) => plus2A_out_42_port, 
                           shiftLeftOnePos(41) => plus2A_out_41_port, 
                           shiftLeftOnePos(40) => plus2A_out_40_port, 
                           shiftLeftOnePos(39) => plus2A_out_39_port, 
                           shiftLeftOnePos(38) => plus2A_out_38_port, 
                           shiftLeftOnePos(37) => plus2A_out_37_port, 
                           shiftLeftOnePos(36) => plus2A_out_36_port, 
                           shiftLeftOnePos(35) => plus2A_out_35_port, 
                           shiftLeftOnePos(34) => plus2A_out_34_port, 
                           shiftLeftOnePos(33) => plus2A_out_33_port, 
                           shiftLeftOnePos(32) => plus2A_out_32_port, 
                           shiftLeftOnePos(31) => plus2A_out_31_port, 
                           shiftLeftOnePos(30) => plus2A_out_30_port, 
                           shiftLeftOnePos(29) => plus2A_out_29_port, 
                           shiftLeftOnePos(28) => plus2A_out_28_port, 
                           shiftLeftOnePos(27) => plus2A_out_27_port, 
                           shiftLeftOnePos(26) => plus2A_out_26_port, 
                           shiftLeftOnePos(25) => plus2A_out_25_port, 
                           shiftLeftOnePos(24) => plus2A_out_24_port, 
                           shiftLeftOnePos(23) => plus2A_out_23_port, 
                           shiftLeftOnePos(22) => plus2A_out_22_port, 
                           shiftLeftOnePos(21) => plus2A_out_21_port, 
                           shiftLeftOnePos(20) => plus2A_out_20_port, 
                           shiftLeftOnePos(19) => plus2A_out_19_port, 
                           shiftLeftOnePos(18) => plus2A_out_18_port, 
                           shiftLeftOnePos(17) => plus2A_out_17_port, 
                           shiftLeftOnePos(16) => plus2A_out_16_port, 
                           shiftLeftOnePos(15) => plus2A_out_15_port, 
                           shiftLeftOnePos(14) => plus2A_out_14_port, 
                           shiftLeftOnePos(13) => plus2A_out_13_port, 
                           shiftLeftOnePos(12) => plus2A_out_12_port, 
                           shiftLeftOnePos(11) => plus2A_out_11_port, 
                           shiftLeftOnePos(10) => plus2A_out_10_port, 
                           shiftLeftOnePos(9) => plus2A_out_9_port, 
                           shiftLeftOnePos(8) => plus2A_out_8_port, 
                           shiftLeftOnePos(7) => plus2A_out_7_port, 
                           shiftLeftOnePos(6) => plus2A_out_6_port, 
                           shiftLeftOnePos(5) => plus2A_out_5_port, 
                           shiftLeftOnePos(4) => plus2A_out_4_port, 
                           shiftLeftOnePos(3) => plus2A_out_3_port, 
                           shiftLeftOnePos(2) => plus2A_out_2_port, 
                           shiftLeftOnePos(1) => plus2A_out_1_port, 
                           shiftLeftOnePos(0) => n_3144);
   shifter_2 : shifter_N64_1 port map( input(63) => plus2A_out_63_port, 
                           input(62) => plus2A_out_62_port, input(61) => 
                           plus2A_out_61_port, input(60) => plus2A_out_60_port,
                           input(59) => plus2A_out_59_port, input(58) => 
                           plus2A_out_58_port, input(57) => plus2A_out_57_port,
                           input(56) => plus2A_out_56_port, input(55) => 
                           plus2A_out_55_port, input(54) => plus2A_out_54_port,
                           input(53) => plus2A_out_53_port, input(52) => 
                           plus2A_out_52_port, input(51) => plus2A_out_51_port,
                           input(50) => plus2A_out_50_port, input(49) => 
                           plus2A_out_49_port, input(48) => plus2A_out_48_port,
                           input(47) => plus2A_out_47_port, input(46) => 
                           plus2A_out_46_port, input(45) => plus2A_out_45_port,
                           input(44) => plus2A_out_44_port, input(43) => 
                           plus2A_out_43_port, input(42) => plus2A_out_42_port,
                           input(41) => plus2A_out_41_port, input(40) => 
                           plus2A_out_40_port, input(39) => plus2A_out_39_port,
                           input(38) => plus2A_out_38_port, input(37) => 
                           plus2A_out_37_port, input(36) => plus2A_out_36_port,
                           input(35) => plus2A_out_35_port, input(34) => 
                           plus2A_out_34_port, input(33) => plus2A_out_33_port,
                           input(32) => plus2A_out_32_port, input(31) => 
                           plus2A_out_31_port, input(30) => plus2A_out_30_port,
                           input(29) => plus2A_out_29_port, input(28) => 
                           plus2A_out_28_port, input(27) => plus2A_out_27_port,
                           input(26) => plus2A_out_26_port, input(25) => 
                           plus2A_out_25_port, input(24) => plus2A_out_24_port,
                           input(23) => plus2A_out_23_port, input(22) => 
                           plus2A_out_22_port, input(21) => plus2A_out_21_port,
                           input(20) => plus2A_out_20_port, input(19) => 
                           plus2A_out_19_port, input(18) => plus2A_out_18_port,
                           input(17) => plus2A_out_17_port, input(16) => 
                           plus2A_out_16_port, input(15) => plus2A_out_15_port,
                           input(14) => plus2A_out_14_port, input(13) => 
                           plus2A_out_13_port, input(12) => plus2A_out_12_port,
                           input(11) => plus2A_out_11_port, input(10) => 
                           plus2A_out_10_port, input(9) => plus2A_out_9_port, 
                           input(8) => plus2A_out_8_port, input(7) => 
                           plus2A_out_7_port, input(6) => plus2A_out_6_port, 
                           input(5) => plus2A_out_5_port, input(4) => 
                           plus2A_out_4_port, input(3) => plus2A_out_3_port, 
                           input(2) => plus2A_out_2_port, input(1) => 
                           plus2A_out_1_port, input(0) => plus2A_out_0_port, 
                           shiftLeftOnePos(63) => plus4A_out_63_port, 
                           shiftLeftOnePos(62) => plus4A_out_62_port, 
                           shiftLeftOnePos(61) => plus4A_out_61_port, 
                           shiftLeftOnePos(60) => plus4A_out_60_port, 
                           shiftLeftOnePos(59) => plus4A_out_59_port, 
                           shiftLeftOnePos(58) => plus4A_out_58_port, 
                           shiftLeftOnePos(57) => plus4A_out_57_port, 
                           shiftLeftOnePos(56) => plus4A_out_56_port, 
                           shiftLeftOnePos(55) => plus4A_out_55_port, 
                           shiftLeftOnePos(54) => plus4A_out_54_port, 
                           shiftLeftOnePos(53) => plus4A_out_53_port, 
                           shiftLeftOnePos(52) => plus4A_out_52_port, 
                           shiftLeftOnePos(51) => plus4A_out_51_port, 
                           shiftLeftOnePos(50) => plus4A_out_50_port, 
                           shiftLeftOnePos(49) => plus4A_out_49_port, 
                           shiftLeftOnePos(48) => plus4A_out_48_port, 
                           shiftLeftOnePos(47) => plus4A_out_47_port, 
                           shiftLeftOnePos(46) => plus4A_out_46_port, 
                           shiftLeftOnePos(45) => plus4A_out_45_port, 
                           shiftLeftOnePos(44) => plus4A_out_44_port, 
                           shiftLeftOnePos(43) => plus4A_out_43_port, 
                           shiftLeftOnePos(42) => plus4A_out_42_port, 
                           shiftLeftOnePos(41) => plus4A_out_41_port, 
                           shiftLeftOnePos(40) => plus4A_out_40_port, 
                           shiftLeftOnePos(39) => plus4A_out_39_port, 
                           shiftLeftOnePos(38) => plus4A_out_38_port, 
                           shiftLeftOnePos(37) => plus4A_out_37_port, 
                           shiftLeftOnePos(36) => plus4A_out_36_port, 
                           shiftLeftOnePos(35) => plus4A_out_35_port, 
                           shiftLeftOnePos(34) => plus4A_out_34_port, 
                           shiftLeftOnePos(33) => plus4A_out_33_port, 
                           shiftLeftOnePos(32) => plus4A_out_32_port, 
                           shiftLeftOnePos(31) => plus4A_out_31_port, 
                           shiftLeftOnePos(30) => plus4A_out_30_port, 
                           shiftLeftOnePos(29) => plus4A_out_29_port, 
                           shiftLeftOnePos(28) => plus4A_out_28_port, 
                           shiftLeftOnePos(27) => plus4A_out_27_port, 
                           shiftLeftOnePos(26) => plus4A_out_26_port, 
                           shiftLeftOnePos(25) => plus4A_out_25_port, 
                           shiftLeftOnePos(24) => plus4A_out_24_port, 
                           shiftLeftOnePos(23) => plus4A_out_23_port, 
                           shiftLeftOnePos(22) => plus4A_out_22_port, 
                           shiftLeftOnePos(21) => plus4A_out_21_port, 
                           shiftLeftOnePos(20) => plus4A_out_20_port, 
                           shiftLeftOnePos(19) => plus4A_out_19_port, 
                           shiftLeftOnePos(18) => plus4A_out_18_port, 
                           shiftLeftOnePos(17) => plus4A_out_17_port, 
                           shiftLeftOnePos(16) => plus4A_out_16_port, 
                           shiftLeftOnePos(15) => plus4A_out_15_port, 
                           shiftLeftOnePos(14) => plus4A_out_14_port, 
                           shiftLeftOnePos(13) => plus4A_out_13_port, 
                           shiftLeftOnePos(12) => plus4A_out_12_port, 
                           shiftLeftOnePos(11) => plus4A_out_11_port, 
                           shiftLeftOnePos(10) => plus4A_out_10_port, 
                           shiftLeftOnePos(9) => plus4A_out_9_port, 
                           shiftLeftOnePos(8) => plus4A_out_8_port, 
                           shiftLeftOnePos(7) => plus4A_out_7_port, 
                           shiftLeftOnePos(6) => plus4A_out_6_port, 
                           shiftLeftOnePos(5) => plus4A_out_5_port, 
                           shiftLeftOnePos(4) => plus4A_out_4_port, 
                           shiftLeftOnePos(3) => plus4A_out_3_port, 
                           shiftLeftOnePos(2) => plus4A_out_2_port, 
                           shiftLeftOnePos(1) => plus4A_out_1_port, 
                           shiftLeftOnePos(0) => n_3145);
   complementer_1 : complementer_N64_2 port map( input(63) => 
                           plus2A_out_63_port, input(62) => plus2A_out_62_port,
                           input(61) => plus2A_out_61_port, input(60) => 
                           plus2A_out_60_port, input(59) => plus2A_out_59_port,
                           input(58) => plus2A_out_58_port, input(57) => 
                           plus2A_out_57_port, input(56) => plus2A_out_56_port,
                           input(55) => plus2A_out_55_port, input(54) => 
                           plus2A_out_54_port, input(53) => plus2A_out_53_port,
                           input(52) => plus2A_out_52_port, input(51) => 
                           plus2A_out_51_port, input(50) => plus2A_out_50_port,
                           input(49) => plus2A_out_49_port, input(48) => 
                           plus2A_out_48_port, input(47) => plus2A_out_47_port,
                           input(46) => plus2A_out_46_port, input(45) => 
                           plus2A_out_45_port, input(44) => plus2A_out_44_port,
                           input(43) => plus2A_out_43_port, input(42) => 
                           plus2A_out_42_port, input(41) => plus2A_out_41_port,
                           input(40) => plus2A_out_40_port, input(39) => 
                           plus2A_out_39_port, input(38) => plus2A_out_38_port,
                           input(37) => plus2A_out_37_port, input(36) => 
                           plus2A_out_36_port, input(35) => plus2A_out_35_port,
                           input(34) => plus2A_out_34_port, input(33) => 
                           plus2A_out_33_port, input(32) => plus2A_out_32_port,
                           input(31) => plus2A_out_31_port, input(30) => 
                           plus2A_out_30_port, input(29) => plus2A_out_29_port,
                           input(28) => plus2A_out_28_port, input(27) => 
                           plus2A_out_27_port, input(26) => plus2A_out_26_port,
                           input(25) => plus2A_out_25_port, input(24) => 
                           plus2A_out_24_port, input(23) => plus2A_out_23_port,
                           input(22) => plus2A_out_22_port, input(21) => 
                           plus2A_out_21_port, input(20) => plus2A_out_20_port,
                           input(19) => plus2A_out_19_port, input(18) => 
                           plus2A_out_18_port, input(17) => plus2A_out_17_port,
                           input(16) => plus2A_out_16_port, input(15) => 
                           plus2A_out_15_port, input(14) => plus2A_out_14_port,
                           input(13) => plus2A_out_13_port, input(12) => 
                           plus2A_out_12_port, input(11) => plus2A_out_11_port,
                           input(10) => plus2A_out_10_port, input(9) => 
                           plus2A_out_9_port, input(8) => plus2A_out_8_port, 
                           input(7) => plus2A_out_7_port, input(6) => 
                           plus2A_out_6_port, input(5) => plus2A_out_5_port, 
                           input(4) => plus2A_out_4_port, input(3) => 
                           plus2A_out_3_port, input(2) => plus2A_out_2_port, 
                           input(1) => plus2A_out_1_port, input(0) => 
                           plus2A_out_0_port, complement2(63) => 
                           minus2A_out(63), complement2(62) => minus2A_out(62),
                           complement2(61) => minus2A_out(61), complement2(60) 
                           => minus2A_out(60), complement2(59) => 
                           minus2A_out(59), complement2(58) => minus2A_out(58),
                           complement2(57) => minus2A_out(57), complement2(56) 
                           => minus2A_out(56), complement2(55) => 
                           minus2A_out(55), complement2(54) => minus2A_out(54),
                           complement2(53) => minus2A_out(53), complement2(52) 
                           => minus2A_out(52), complement2(51) => 
                           minus2A_out(51), complement2(50) => minus2A_out(50),
                           complement2(49) => minus2A_out(49), complement2(48) 
                           => minus2A_out(48), complement2(47) => 
                           minus2A_out(47), complement2(46) => minus2A_out(46),
                           complement2(45) => minus2A_out(45), complement2(44) 
                           => minus2A_out(44), complement2(43) => 
                           minus2A_out(43), complement2(42) => minus2A_out(42),
                           complement2(41) => minus2A_out(41), complement2(40) 
                           => minus2A_out(40), complement2(39) => 
                           minus2A_out(39), complement2(38) => minus2A_out(38),
                           complement2(37) => minus2A_out(37), complement2(36) 
                           => minus2A_out(36), complement2(35) => 
                           minus2A_out(35), complement2(34) => minus2A_out(34),
                           complement2(33) => minus2A_out(33), complement2(32) 
                           => minus2A_out(32), complement2(31) => 
                           minus2A_out(31), complement2(30) => minus2A_out(30),
                           complement2(29) => minus2A_out(29), complement2(28) 
                           => minus2A_out(28), complement2(27) => 
                           minus2A_out(27), complement2(26) => minus2A_out(26),
                           complement2(25) => minus2A_out(25), complement2(24) 
                           => minus2A_out(24), complement2(23) => 
                           minus2A_out(23), complement2(22) => minus2A_out(22),
                           complement2(21) => minus2A_out(21), complement2(20) 
                           => minus2A_out(20), complement2(19) => 
                           minus2A_out(19), complement2(18) => minus2A_out(18),
                           complement2(17) => minus2A_out(17), complement2(16) 
                           => minus2A_out(16), complement2(15) => 
                           minus2A_out(15), complement2(14) => minus2A_out(14),
                           complement2(13) => minus2A_out(13), complement2(12) 
                           => minus2A_out(12), complement2(11) => 
                           minus2A_out(11), complement2(10) => minus2A_out(10),
                           complement2(9) => minus2A_out(9), complement2(8) => 
                           minus2A_out(8), complement2(7) => minus2A_out(7), 
                           complement2(6) => minus2A_out(6), complement2(5) => 
                           minus2A_out(5), complement2(4) => minus2A_out(4), 
                           complement2(3) => minus2A_out(3), complement2(2) => 
                           minus2A_out(2), complement2(1) => minus2A_out(1), 
                           complement2(0) => minus2A_out(0));
   complementer_2 : complementer_N64_1 port map( input(63) => 
                           plus4A_out_63_port, input(62) => plus4A_out_62_port,
                           input(61) => plus4A_out_61_port, input(60) => 
                           plus4A_out_60_port, input(59) => plus4A_out_59_port,
                           input(58) => plus4A_out_58_port, input(57) => 
                           plus4A_out_57_port, input(56) => plus4A_out_56_port,
                           input(55) => plus4A_out_55_port, input(54) => 
                           plus4A_out_54_port, input(53) => plus4A_out_53_port,
                           input(52) => plus4A_out_52_port, input(51) => 
                           plus4A_out_51_port, input(50) => plus4A_out_50_port,
                           input(49) => plus4A_out_49_port, input(48) => 
                           plus4A_out_48_port, input(47) => plus4A_out_47_port,
                           input(46) => plus4A_out_46_port, input(45) => 
                           plus4A_out_45_port, input(44) => plus4A_out_44_port,
                           input(43) => plus4A_out_43_port, input(42) => 
                           plus4A_out_42_port, input(41) => plus4A_out_41_port,
                           input(40) => plus4A_out_40_port, input(39) => 
                           plus4A_out_39_port, input(38) => plus4A_out_38_port,
                           input(37) => plus4A_out_37_port, input(36) => 
                           plus4A_out_36_port, input(35) => plus4A_out_35_port,
                           input(34) => plus4A_out_34_port, input(33) => 
                           plus4A_out_33_port, input(32) => plus4A_out_32_port,
                           input(31) => plus4A_out_31_port, input(30) => 
                           plus4A_out_30_port, input(29) => plus4A_out_29_port,
                           input(28) => plus4A_out_28_port, input(27) => 
                           plus4A_out_27_port, input(26) => plus4A_out_26_port,
                           input(25) => plus4A_out_25_port, input(24) => 
                           plus4A_out_24_port, input(23) => plus4A_out_23_port,
                           input(22) => plus4A_out_22_port, input(21) => 
                           plus4A_out_21_port, input(20) => plus4A_out_20_port,
                           input(19) => plus4A_out_19_port, input(18) => 
                           plus4A_out_18_port, input(17) => plus4A_out_17_port,
                           input(16) => plus4A_out_16_port, input(15) => 
                           plus4A_out_15_port, input(14) => plus4A_out_14_port,
                           input(13) => plus4A_out_13_port, input(12) => 
                           plus4A_out_12_port, input(11) => plus4A_out_11_port,
                           input(10) => plus4A_out_10_port, input(9) => 
                           plus4A_out_9_port, input(8) => plus4A_out_8_port, 
                           input(7) => plus4A_out_7_port, input(6) => 
                           plus4A_out_6_port, input(5) => plus4A_out_5_port, 
                           input(4) => plus4A_out_4_port, input(3) => 
                           plus4A_out_3_port, input(2) => plus4A_out_2_port, 
                           input(1) => plus4A_out_1_port, input(0) => 
                           plus4A_out_0_port, complement2(63) => 
                           minus4A_out(63), complement2(62) => minus4A_out(62),
                           complement2(61) => minus4A_out(61), complement2(60) 
                           => minus4A_out(60), complement2(59) => 
                           minus4A_out(59), complement2(58) => minus4A_out(58),
                           complement2(57) => minus4A_out(57), complement2(56) 
                           => minus4A_out(56), complement2(55) => 
                           minus4A_out(55), complement2(54) => minus4A_out(54),
                           complement2(53) => minus4A_out(53), complement2(52) 
                           => minus4A_out(52), complement2(51) => 
                           minus4A_out(51), complement2(50) => minus4A_out(50),
                           complement2(49) => minus4A_out(49), complement2(48) 
                           => minus4A_out(48), complement2(47) => 
                           minus4A_out(47), complement2(46) => minus4A_out(46),
                           complement2(45) => minus4A_out(45), complement2(44) 
                           => minus4A_out(44), complement2(43) => 
                           minus4A_out(43), complement2(42) => minus4A_out(42),
                           complement2(41) => minus4A_out(41), complement2(40) 
                           => minus4A_out(40), complement2(39) => 
                           minus4A_out(39), complement2(38) => minus4A_out(38),
                           complement2(37) => minus4A_out(37), complement2(36) 
                           => minus4A_out(36), complement2(35) => 
                           minus4A_out(35), complement2(34) => minus4A_out(34),
                           complement2(33) => minus4A_out(33), complement2(32) 
                           => minus4A_out(32), complement2(31) => 
                           minus4A_out(31), complement2(30) => minus4A_out(30),
                           complement2(29) => minus4A_out(29), complement2(28) 
                           => minus4A_out(28), complement2(27) => 
                           minus4A_out(27), complement2(26) => minus4A_out(26),
                           complement2(25) => minus4A_out(25), complement2(24) 
                           => minus4A_out(24), complement2(23) => 
                           minus4A_out(23), complement2(22) => minus4A_out(22),
                           complement2(21) => minus4A_out(21), complement2(20) 
                           => minus4A_out(20), complement2(19) => 
                           minus4A_out(19), complement2(18) => minus4A_out(18),
                           complement2(17) => minus4A_out(17), complement2(16) 
                           => minus4A_out(16), complement2(15) => 
                           minus4A_out(15), complement2(14) => minus4A_out(14),
                           complement2(13) => minus4A_out(13), complement2(12) 
                           => minus4A_out(12), complement2(11) => 
                           minus4A_out(11), complement2(10) => minus4A_out(10),
                           complement2(9) => minus4A_out(9), complement2(8) => 
                           minus4A_out(8), complement2(7) => minus4A_out(7), 
                           complement2(6) => minus4A_out(6), complement2(5) => 
                           minus4A_out(5), complement2(4) => minus4A_out(4), 
                           complement2(3) => minus4A_out(3), complement2(2) => 
                           minus4A_out(2), complement2(1) => minus4A_out(1), 
                           complement2(0) => minus4A_out(0));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity ShiftnCompl_N64_2 is

   port( plusA : in std_logic_vector (63 downto 0);  plus2A_out, minus2A_out, 
         plus4A_out, minus4A_out : out std_logic_vector (63 downto 0));

end ShiftnCompl_N64_2;

architecture SYN_struct of ShiftnCompl_N64_2 is

   component complementer_N64_3
      port( input : in std_logic_vector (63 downto 0);  complement2 : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component complementer_N64_4
      port( input : in std_logic_vector (63 downto 0);  complement2 : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component shifter_N64_3
      port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component shifter_N64_4
      port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
            std_logic_vector (63 downto 0));
   end component;
   
   signal plus2A_out_63_port, plus2A_out_62_port, plus2A_out_61_port, 
      plus2A_out_60_port, plus2A_out_59_port, plus2A_out_58_port, 
      plus2A_out_57_port, plus2A_out_56_port, plus2A_out_55_port, 
      plus2A_out_54_port, plus2A_out_53_port, plus2A_out_52_port, 
      plus2A_out_51_port, plus2A_out_50_port, plus2A_out_49_port, 
      plus2A_out_48_port, plus2A_out_47_port, plus2A_out_46_port, 
      plus2A_out_45_port, plus2A_out_44_port, plus2A_out_43_port, 
      plus2A_out_42_port, plus2A_out_41_port, plus2A_out_40_port, 
      plus2A_out_39_port, plus2A_out_38_port, plus2A_out_37_port, 
      plus2A_out_36_port, plus2A_out_35_port, plus2A_out_34_port, 
      plus2A_out_33_port, plus2A_out_32_port, plus2A_out_31_port, 
      plus2A_out_30_port, plus2A_out_29_port, plus2A_out_28_port, 
      plus2A_out_27_port, plus2A_out_26_port, plus2A_out_25_port, 
      plus2A_out_24_port, plus2A_out_23_port, plus2A_out_22_port, 
      plus2A_out_21_port, plus2A_out_20_port, plus2A_out_19_port, 
      plus2A_out_18_port, plus2A_out_17_port, plus2A_out_16_port, 
      plus2A_out_15_port, plus2A_out_14_port, plus2A_out_13_port, 
      plus2A_out_12_port, plus2A_out_11_port, plus2A_out_10_port, 
      plus2A_out_9_port, plus2A_out_8_port, plus2A_out_7_port, 
      plus2A_out_6_port, plus2A_out_5_port, plus2A_out_4_port, 
      plus2A_out_3_port, plus2A_out_2_port, plus2A_out_1_port, 
      plus2A_out_0_port, plus4A_out_63_port, plus4A_out_62_port, 
      plus4A_out_61_port, plus4A_out_60_port, plus4A_out_59_port, 
      plus4A_out_58_port, plus4A_out_57_port, plus4A_out_56_port, 
      plus4A_out_55_port, plus4A_out_54_port, plus4A_out_53_port, 
      plus4A_out_52_port, plus4A_out_51_port, plus4A_out_50_port, 
      plus4A_out_49_port, plus4A_out_48_port, plus4A_out_47_port, 
      plus4A_out_46_port, plus4A_out_45_port, plus4A_out_44_port, 
      plus4A_out_43_port, plus4A_out_42_port, plus4A_out_41_port, 
      plus4A_out_40_port, plus4A_out_39_port, plus4A_out_38_port, 
      plus4A_out_37_port, plus4A_out_36_port, plus4A_out_35_port, 
      plus4A_out_34_port, plus4A_out_33_port, plus4A_out_32_port, 
      plus4A_out_31_port, plus4A_out_30_port, plus4A_out_29_port, 
      plus4A_out_28_port, plus4A_out_27_port, plus4A_out_26_port, 
      plus4A_out_25_port, plus4A_out_24_port, plus4A_out_23_port, 
      plus4A_out_22_port, plus4A_out_21_port, plus4A_out_20_port, 
      plus4A_out_19_port, plus4A_out_18_port, plus4A_out_17_port, 
      plus4A_out_16_port, plus4A_out_15_port, plus4A_out_14_port, 
      plus4A_out_13_port, plus4A_out_12_port, plus4A_out_11_port, 
      plus4A_out_10_port, plus4A_out_9_port, plus4A_out_8_port, 
      plus4A_out_7_port, plus4A_out_6_port, plus4A_out_5_port, 
      plus4A_out_4_port, plus4A_out_3_port, plus4A_out_2_port, 
      plus4A_out_1_port, plus4A_out_0_port, n_3146, n_3147 : std_logic;

begin
   plus2A_out <= ( plus2A_out_63_port, plus2A_out_62_port, plus2A_out_61_port, 
      plus2A_out_60_port, plus2A_out_59_port, plus2A_out_58_port, 
      plus2A_out_57_port, plus2A_out_56_port, plus2A_out_55_port, 
      plus2A_out_54_port, plus2A_out_53_port, plus2A_out_52_port, 
      plus2A_out_51_port, plus2A_out_50_port, plus2A_out_49_port, 
      plus2A_out_48_port, plus2A_out_47_port, plus2A_out_46_port, 
      plus2A_out_45_port, plus2A_out_44_port, plus2A_out_43_port, 
      plus2A_out_42_port, plus2A_out_41_port, plus2A_out_40_port, 
      plus2A_out_39_port, plus2A_out_38_port, plus2A_out_37_port, 
      plus2A_out_36_port, plus2A_out_35_port, plus2A_out_34_port, 
      plus2A_out_33_port, plus2A_out_32_port, plus2A_out_31_port, 
      plus2A_out_30_port, plus2A_out_29_port, plus2A_out_28_port, 
      plus2A_out_27_port, plus2A_out_26_port, plus2A_out_25_port, 
      plus2A_out_24_port, plus2A_out_23_port, plus2A_out_22_port, 
      plus2A_out_21_port, plus2A_out_20_port, plus2A_out_19_port, 
      plus2A_out_18_port, plus2A_out_17_port, plus2A_out_16_port, 
      plus2A_out_15_port, plus2A_out_14_port, plus2A_out_13_port, 
      plus2A_out_12_port, plus2A_out_11_port, plus2A_out_10_port, 
      plus2A_out_9_port, plus2A_out_8_port, plus2A_out_7_port, 
      plus2A_out_6_port, plus2A_out_5_port, plus2A_out_4_port, 
      plus2A_out_3_port, plus2A_out_2_port, plus2A_out_1_port, 
      plus2A_out_0_port );
   plus4A_out <= ( plus4A_out_63_port, plus4A_out_62_port, plus4A_out_61_port, 
      plus4A_out_60_port, plus4A_out_59_port, plus4A_out_58_port, 
      plus4A_out_57_port, plus4A_out_56_port, plus4A_out_55_port, 
      plus4A_out_54_port, plus4A_out_53_port, plus4A_out_52_port, 
      plus4A_out_51_port, plus4A_out_50_port, plus4A_out_49_port, 
      plus4A_out_48_port, plus4A_out_47_port, plus4A_out_46_port, 
      plus4A_out_45_port, plus4A_out_44_port, plus4A_out_43_port, 
      plus4A_out_42_port, plus4A_out_41_port, plus4A_out_40_port, 
      plus4A_out_39_port, plus4A_out_38_port, plus4A_out_37_port, 
      plus4A_out_36_port, plus4A_out_35_port, plus4A_out_34_port, 
      plus4A_out_33_port, plus4A_out_32_port, plus4A_out_31_port, 
      plus4A_out_30_port, plus4A_out_29_port, plus4A_out_28_port, 
      plus4A_out_27_port, plus4A_out_26_port, plus4A_out_25_port, 
      plus4A_out_24_port, plus4A_out_23_port, plus4A_out_22_port, 
      plus4A_out_21_port, plus4A_out_20_port, plus4A_out_19_port, 
      plus4A_out_18_port, plus4A_out_17_port, plus4A_out_16_port, 
      plus4A_out_15_port, plus4A_out_14_port, plus4A_out_13_port, 
      plus4A_out_12_port, plus4A_out_11_port, plus4A_out_10_port, 
      plus4A_out_9_port, plus4A_out_8_port, plus4A_out_7_port, 
      plus4A_out_6_port, plus4A_out_5_port, plus4A_out_4_port, 
      plus4A_out_3_port, plus4A_out_2_port, plus4A_out_1_port, 
      plus4A_out_0_port );
   
   plus2A_out_0_port <= '0';
   plus4A_out_0_port <= '0';
   shifter_1 : shifter_N64_4 port map( input(63) => plusA(63), input(62) => 
                           plusA(62), input(61) => plusA(61), input(60) => 
                           plusA(60), input(59) => plusA(59), input(58) => 
                           plusA(58), input(57) => plusA(57), input(56) => 
                           plusA(56), input(55) => plusA(55), input(54) => 
                           plusA(54), input(53) => plusA(53), input(52) => 
                           plusA(52), input(51) => plusA(51), input(50) => 
                           plusA(50), input(49) => plusA(49), input(48) => 
                           plusA(48), input(47) => plusA(47), input(46) => 
                           plusA(46), input(45) => plusA(45), input(44) => 
                           plusA(44), input(43) => plusA(43), input(42) => 
                           plusA(42), input(41) => plusA(41), input(40) => 
                           plusA(40), input(39) => plusA(39), input(38) => 
                           plusA(38), input(37) => plusA(37), input(36) => 
                           plusA(36), input(35) => plusA(35), input(34) => 
                           plusA(34), input(33) => plusA(33), input(32) => 
                           plusA(32), input(31) => plusA(31), input(30) => 
                           plusA(30), input(29) => plusA(29), input(28) => 
                           plusA(28), input(27) => plusA(27), input(26) => 
                           plusA(26), input(25) => plusA(25), input(24) => 
                           plusA(24), input(23) => plusA(23), input(22) => 
                           plusA(22), input(21) => plusA(21), input(20) => 
                           plusA(20), input(19) => plusA(19), input(18) => 
                           plusA(18), input(17) => plusA(17), input(16) => 
                           plusA(16), input(15) => plusA(15), input(14) => 
                           plusA(14), input(13) => plusA(13), input(12) => 
                           plusA(12), input(11) => plusA(11), input(10) => 
                           plusA(10), input(9) => plusA(9), input(8) => 
                           plusA(8), input(7) => plusA(7), input(6) => plusA(6)
                           , input(5) => plusA(5), input(4) => plusA(4), 
                           input(3) => plusA(3), input(2) => plusA(2), input(1)
                           => plusA(1), input(0) => plusA(0), 
                           shiftLeftOnePos(63) => plus2A_out_63_port, 
                           shiftLeftOnePos(62) => plus2A_out_62_port, 
                           shiftLeftOnePos(61) => plus2A_out_61_port, 
                           shiftLeftOnePos(60) => plus2A_out_60_port, 
                           shiftLeftOnePos(59) => plus2A_out_59_port, 
                           shiftLeftOnePos(58) => plus2A_out_58_port, 
                           shiftLeftOnePos(57) => plus2A_out_57_port, 
                           shiftLeftOnePos(56) => plus2A_out_56_port, 
                           shiftLeftOnePos(55) => plus2A_out_55_port, 
                           shiftLeftOnePos(54) => plus2A_out_54_port, 
                           shiftLeftOnePos(53) => plus2A_out_53_port, 
                           shiftLeftOnePos(52) => plus2A_out_52_port, 
                           shiftLeftOnePos(51) => plus2A_out_51_port, 
                           shiftLeftOnePos(50) => plus2A_out_50_port, 
                           shiftLeftOnePos(49) => plus2A_out_49_port, 
                           shiftLeftOnePos(48) => plus2A_out_48_port, 
                           shiftLeftOnePos(47) => plus2A_out_47_port, 
                           shiftLeftOnePos(46) => plus2A_out_46_port, 
                           shiftLeftOnePos(45) => plus2A_out_45_port, 
                           shiftLeftOnePos(44) => plus2A_out_44_port, 
                           shiftLeftOnePos(43) => plus2A_out_43_port, 
                           shiftLeftOnePos(42) => plus2A_out_42_port, 
                           shiftLeftOnePos(41) => plus2A_out_41_port, 
                           shiftLeftOnePos(40) => plus2A_out_40_port, 
                           shiftLeftOnePos(39) => plus2A_out_39_port, 
                           shiftLeftOnePos(38) => plus2A_out_38_port, 
                           shiftLeftOnePos(37) => plus2A_out_37_port, 
                           shiftLeftOnePos(36) => plus2A_out_36_port, 
                           shiftLeftOnePos(35) => plus2A_out_35_port, 
                           shiftLeftOnePos(34) => plus2A_out_34_port, 
                           shiftLeftOnePos(33) => plus2A_out_33_port, 
                           shiftLeftOnePos(32) => plus2A_out_32_port, 
                           shiftLeftOnePos(31) => plus2A_out_31_port, 
                           shiftLeftOnePos(30) => plus2A_out_30_port, 
                           shiftLeftOnePos(29) => plus2A_out_29_port, 
                           shiftLeftOnePos(28) => plus2A_out_28_port, 
                           shiftLeftOnePos(27) => plus2A_out_27_port, 
                           shiftLeftOnePos(26) => plus2A_out_26_port, 
                           shiftLeftOnePos(25) => plus2A_out_25_port, 
                           shiftLeftOnePos(24) => plus2A_out_24_port, 
                           shiftLeftOnePos(23) => plus2A_out_23_port, 
                           shiftLeftOnePos(22) => plus2A_out_22_port, 
                           shiftLeftOnePos(21) => plus2A_out_21_port, 
                           shiftLeftOnePos(20) => plus2A_out_20_port, 
                           shiftLeftOnePos(19) => plus2A_out_19_port, 
                           shiftLeftOnePos(18) => plus2A_out_18_port, 
                           shiftLeftOnePos(17) => plus2A_out_17_port, 
                           shiftLeftOnePos(16) => plus2A_out_16_port, 
                           shiftLeftOnePos(15) => plus2A_out_15_port, 
                           shiftLeftOnePos(14) => plus2A_out_14_port, 
                           shiftLeftOnePos(13) => plus2A_out_13_port, 
                           shiftLeftOnePos(12) => plus2A_out_12_port, 
                           shiftLeftOnePos(11) => plus2A_out_11_port, 
                           shiftLeftOnePos(10) => plus2A_out_10_port, 
                           shiftLeftOnePos(9) => plus2A_out_9_port, 
                           shiftLeftOnePos(8) => plus2A_out_8_port, 
                           shiftLeftOnePos(7) => plus2A_out_7_port, 
                           shiftLeftOnePos(6) => plus2A_out_6_port, 
                           shiftLeftOnePos(5) => plus2A_out_5_port, 
                           shiftLeftOnePos(4) => plus2A_out_4_port, 
                           shiftLeftOnePos(3) => plus2A_out_3_port, 
                           shiftLeftOnePos(2) => plus2A_out_2_port, 
                           shiftLeftOnePos(1) => plus2A_out_1_port, 
                           shiftLeftOnePos(0) => n_3146);
   shifter_2 : shifter_N64_3 port map( input(63) => plus2A_out_63_port, 
                           input(62) => plus2A_out_62_port, input(61) => 
                           plus2A_out_61_port, input(60) => plus2A_out_60_port,
                           input(59) => plus2A_out_59_port, input(58) => 
                           plus2A_out_58_port, input(57) => plus2A_out_57_port,
                           input(56) => plus2A_out_56_port, input(55) => 
                           plus2A_out_55_port, input(54) => plus2A_out_54_port,
                           input(53) => plus2A_out_53_port, input(52) => 
                           plus2A_out_52_port, input(51) => plus2A_out_51_port,
                           input(50) => plus2A_out_50_port, input(49) => 
                           plus2A_out_49_port, input(48) => plus2A_out_48_port,
                           input(47) => plus2A_out_47_port, input(46) => 
                           plus2A_out_46_port, input(45) => plus2A_out_45_port,
                           input(44) => plus2A_out_44_port, input(43) => 
                           plus2A_out_43_port, input(42) => plus2A_out_42_port,
                           input(41) => plus2A_out_41_port, input(40) => 
                           plus2A_out_40_port, input(39) => plus2A_out_39_port,
                           input(38) => plus2A_out_38_port, input(37) => 
                           plus2A_out_37_port, input(36) => plus2A_out_36_port,
                           input(35) => plus2A_out_35_port, input(34) => 
                           plus2A_out_34_port, input(33) => plus2A_out_33_port,
                           input(32) => plus2A_out_32_port, input(31) => 
                           plus2A_out_31_port, input(30) => plus2A_out_30_port,
                           input(29) => plus2A_out_29_port, input(28) => 
                           plus2A_out_28_port, input(27) => plus2A_out_27_port,
                           input(26) => plus2A_out_26_port, input(25) => 
                           plus2A_out_25_port, input(24) => plus2A_out_24_port,
                           input(23) => plus2A_out_23_port, input(22) => 
                           plus2A_out_22_port, input(21) => plus2A_out_21_port,
                           input(20) => plus2A_out_20_port, input(19) => 
                           plus2A_out_19_port, input(18) => plus2A_out_18_port,
                           input(17) => plus2A_out_17_port, input(16) => 
                           plus2A_out_16_port, input(15) => plus2A_out_15_port,
                           input(14) => plus2A_out_14_port, input(13) => 
                           plus2A_out_13_port, input(12) => plus2A_out_12_port,
                           input(11) => plus2A_out_11_port, input(10) => 
                           plus2A_out_10_port, input(9) => plus2A_out_9_port, 
                           input(8) => plus2A_out_8_port, input(7) => 
                           plus2A_out_7_port, input(6) => plus2A_out_6_port, 
                           input(5) => plus2A_out_5_port, input(4) => 
                           plus2A_out_4_port, input(3) => plus2A_out_3_port, 
                           input(2) => plus2A_out_2_port, input(1) => 
                           plus2A_out_1_port, input(0) => plus2A_out_0_port, 
                           shiftLeftOnePos(63) => plus4A_out_63_port, 
                           shiftLeftOnePos(62) => plus4A_out_62_port, 
                           shiftLeftOnePos(61) => plus4A_out_61_port, 
                           shiftLeftOnePos(60) => plus4A_out_60_port, 
                           shiftLeftOnePos(59) => plus4A_out_59_port, 
                           shiftLeftOnePos(58) => plus4A_out_58_port, 
                           shiftLeftOnePos(57) => plus4A_out_57_port, 
                           shiftLeftOnePos(56) => plus4A_out_56_port, 
                           shiftLeftOnePos(55) => plus4A_out_55_port, 
                           shiftLeftOnePos(54) => plus4A_out_54_port, 
                           shiftLeftOnePos(53) => plus4A_out_53_port, 
                           shiftLeftOnePos(52) => plus4A_out_52_port, 
                           shiftLeftOnePos(51) => plus4A_out_51_port, 
                           shiftLeftOnePos(50) => plus4A_out_50_port, 
                           shiftLeftOnePos(49) => plus4A_out_49_port, 
                           shiftLeftOnePos(48) => plus4A_out_48_port, 
                           shiftLeftOnePos(47) => plus4A_out_47_port, 
                           shiftLeftOnePos(46) => plus4A_out_46_port, 
                           shiftLeftOnePos(45) => plus4A_out_45_port, 
                           shiftLeftOnePos(44) => plus4A_out_44_port, 
                           shiftLeftOnePos(43) => plus4A_out_43_port, 
                           shiftLeftOnePos(42) => plus4A_out_42_port, 
                           shiftLeftOnePos(41) => plus4A_out_41_port, 
                           shiftLeftOnePos(40) => plus4A_out_40_port, 
                           shiftLeftOnePos(39) => plus4A_out_39_port, 
                           shiftLeftOnePos(38) => plus4A_out_38_port, 
                           shiftLeftOnePos(37) => plus4A_out_37_port, 
                           shiftLeftOnePos(36) => plus4A_out_36_port, 
                           shiftLeftOnePos(35) => plus4A_out_35_port, 
                           shiftLeftOnePos(34) => plus4A_out_34_port, 
                           shiftLeftOnePos(33) => plus4A_out_33_port, 
                           shiftLeftOnePos(32) => plus4A_out_32_port, 
                           shiftLeftOnePos(31) => plus4A_out_31_port, 
                           shiftLeftOnePos(30) => plus4A_out_30_port, 
                           shiftLeftOnePos(29) => plus4A_out_29_port, 
                           shiftLeftOnePos(28) => plus4A_out_28_port, 
                           shiftLeftOnePos(27) => plus4A_out_27_port, 
                           shiftLeftOnePos(26) => plus4A_out_26_port, 
                           shiftLeftOnePos(25) => plus4A_out_25_port, 
                           shiftLeftOnePos(24) => plus4A_out_24_port, 
                           shiftLeftOnePos(23) => plus4A_out_23_port, 
                           shiftLeftOnePos(22) => plus4A_out_22_port, 
                           shiftLeftOnePos(21) => plus4A_out_21_port, 
                           shiftLeftOnePos(20) => plus4A_out_20_port, 
                           shiftLeftOnePos(19) => plus4A_out_19_port, 
                           shiftLeftOnePos(18) => plus4A_out_18_port, 
                           shiftLeftOnePos(17) => plus4A_out_17_port, 
                           shiftLeftOnePos(16) => plus4A_out_16_port, 
                           shiftLeftOnePos(15) => plus4A_out_15_port, 
                           shiftLeftOnePos(14) => plus4A_out_14_port, 
                           shiftLeftOnePos(13) => plus4A_out_13_port, 
                           shiftLeftOnePos(12) => plus4A_out_12_port, 
                           shiftLeftOnePos(11) => plus4A_out_11_port, 
                           shiftLeftOnePos(10) => plus4A_out_10_port, 
                           shiftLeftOnePos(9) => plus4A_out_9_port, 
                           shiftLeftOnePos(8) => plus4A_out_8_port, 
                           shiftLeftOnePos(7) => plus4A_out_7_port, 
                           shiftLeftOnePos(6) => plus4A_out_6_port, 
                           shiftLeftOnePos(5) => plus4A_out_5_port, 
                           shiftLeftOnePos(4) => plus4A_out_4_port, 
                           shiftLeftOnePos(3) => plus4A_out_3_port, 
                           shiftLeftOnePos(2) => plus4A_out_2_port, 
                           shiftLeftOnePos(1) => plus4A_out_1_port, 
                           shiftLeftOnePos(0) => n_3147);
   complementer_1 : complementer_N64_4 port map( input(63) => 
                           plus2A_out_63_port, input(62) => plus2A_out_62_port,
                           input(61) => plus2A_out_61_port, input(60) => 
                           plus2A_out_60_port, input(59) => plus2A_out_59_port,
                           input(58) => plus2A_out_58_port, input(57) => 
                           plus2A_out_57_port, input(56) => plus2A_out_56_port,
                           input(55) => plus2A_out_55_port, input(54) => 
                           plus2A_out_54_port, input(53) => plus2A_out_53_port,
                           input(52) => plus2A_out_52_port, input(51) => 
                           plus2A_out_51_port, input(50) => plus2A_out_50_port,
                           input(49) => plus2A_out_49_port, input(48) => 
                           plus2A_out_48_port, input(47) => plus2A_out_47_port,
                           input(46) => plus2A_out_46_port, input(45) => 
                           plus2A_out_45_port, input(44) => plus2A_out_44_port,
                           input(43) => plus2A_out_43_port, input(42) => 
                           plus2A_out_42_port, input(41) => plus2A_out_41_port,
                           input(40) => plus2A_out_40_port, input(39) => 
                           plus2A_out_39_port, input(38) => plus2A_out_38_port,
                           input(37) => plus2A_out_37_port, input(36) => 
                           plus2A_out_36_port, input(35) => plus2A_out_35_port,
                           input(34) => plus2A_out_34_port, input(33) => 
                           plus2A_out_33_port, input(32) => plus2A_out_32_port,
                           input(31) => plus2A_out_31_port, input(30) => 
                           plus2A_out_30_port, input(29) => plus2A_out_29_port,
                           input(28) => plus2A_out_28_port, input(27) => 
                           plus2A_out_27_port, input(26) => plus2A_out_26_port,
                           input(25) => plus2A_out_25_port, input(24) => 
                           plus2A_out_24_port, input(23) => plus2A_out_23_port,
                           input(22) => plus2A_out_22_port, input(21) => 
                           plus2A_out_21_port, input(20) => plus2A_out_20_port,
                           input(19) => plus2A_out_19_port, input(18) => 
                           plus2A_out_18_port, input(17) => plus2A_out_17_port,
                           input(16) => plus2A_out_16_port, input(15) => 
                           plus2A_out_15_port, input(14) => plus2A_out_14_port,
                           input(13) => plus2A_out_13_port, input(12) => 
                           plus2A_out_12_port, input(11) => plus2A_out_11_port,
                           input(10) => plus2A_out_10_port, input(9) => 
                           plus2A_out_9_port, input(8) => plus2A_out_8_port, 
                           input(7) => plus2A_out_7_port, input(6) => 
                           plus2A_out_6_port, input(5) => plus2A_out_5_port, 
                           input(4) => plus2A_out_4_port, input(3) => 
                           plus2A_out_3_port, input(2) => plus2A_out_2_port, 
                           input(1) => plus2A_out_1_port, input(0) => 
                           plus2A_out_0_port, complement2(63) => 
                           minus2A_out(63), complement2(62) => minus2A_out(62),
                           complement2(61) => minus2A_out(61), complement2(60) 
                           => minus2A_out(60), complement2(59) => 
                           minus2A_out(59), complement2(58) => minus2A_out(58),
                           complement2(57) => minus2A_out(57), complement2(56) 
                           => minus2A_out(56), complement2(55) => 
                           minus2A_out(55), complement2(54) => minus2A_out(54),
                           complement2(53) => minus2A_out(53), complement2(52) 
                           => minus2A_out(52), complement2(51) => 
                           minus2A_out(51), complement2(50) => minus2A_out(50),
                           complement2(49) => minus2A_out(49), complement2(48) 
                           => minus2A_out(48), complement2(47) => 
                           minus2A_out(47), complement2(46) => minus2A_out(46),
                           complement2(45) => minus2A_out(45), complement2(44) 
                           => minus2A_out(44), complement2(43) => 
                           minus2A_out(43), complement2(42) => minus2A_out(42),
                           complement2(41) => minus2A_out(41), complement2(40) 
                           => minus2A_out(40), complement2(39) => 
                           minus2A_out(39), complement2(38) => minus2A_out(38),
                           complement2(37) => minus2A_out(37), complement2(36) 
                           => minus2A_out(36), complement2(35) => 
                           minus2A_out(35), complement2(34) => minus2A_out(34),
                           complement2(33) => minus2A_out(33), complement2(32) 
                           => minus2A_out(32), complement2(31) => 
                           minus2A_out(31), complement2(30) => minus2A_out(30),
                           complement2(29) => minus2A_out(29), complement2(28) 
                           => minus2A_out(28), complement2(27) => 
                           minus2A_out(27), complement2(26) => minus2A_out(26),
                           complement2(25) => minus2A_out(25), complement2(24) 
                           => minus2A_out(24), complement2(23) => 
                           minus2A_out(23), complement2(22) => minus2A_out(22),
                           complement2(21) => minus2A_out(21), complement2(20) 
                           => minus2A_out(20), complement2(19) => 
                           minus2A_out(19), complement2(18) => minus2A_out(18),
                           complement2(17) => minus2A_out(17), complement2(16) 
                           => minus2A_out(16), complement2(15) => 
                           minus2A_out(15), complement2(14) => minus2A_out(14),
                           complement2(13) => minus2A_out(13), complement2(12) 
                           => minus2A_out(12), complement2(11) => 
                           minus2A_out(11), complement2(10) => minus2A_out(10),
                           complement2(9) => minus2A_out(9), complement2(8) => 
                           minus2A_out(8), complement2(7) => minus2A_out(7), 
                           complement2(6) => minus2A_out(6), complement2(5) => 
                           minus2A_out(5), complement2(4) => minus2A_out(4), 
                           complement2(3) => minus2A_out(3), complement2(2) => 
                           minus2A_out(2), complement2(1) => minus2A_out(1), 
                           complement2(0) => minus2A_out(0));
   complementer_2 : complementer_N64_3 port map( input(63) => 
                           plus4A_out_63_port, input(62) => plus4A_out_62_port,
                           input(61) => plus4A_out_61_port, input(60) => 
                           plus4A_out_60_port, input(59) => plus4A_out_59_port,
                           input(58) => plus4A_out_58_port, input(57) => 
                           plus4A_out_57_port, input(56) => plus4A_out_56_port,
                           input(55) => plus4A_out_55_port, input(54) => 
                           plus4A_out_54_port, input(53) => plus4A_out_53_port,
                           input(52) => plus4A_out_52_port, input(51) => 
                           plus4A_out_51_port, input(50) => plus4A_out_50_port,
                           input(49) => plus4A_out_49_port, input(48) => 
                           plus4A_out_48_port, input(47) => plus4A_out_47_port,
                           input(46) => plus4A_out_46_port, input(45) => 
                           plus4A_out_45_port, input(44) => plus4A_out_44_port,
                           input(43) => plus4A_out_43_port, input(42) => 
                           plus4A_out_42_port, input(41) => plus4A_out_41_port,
                           input(40) => plus4A_out_40_port, input(39) => 
                           plus4A_out_39_port, input(38) => plus4A_out_38_port,
                           input(37) => plus4A_out_37_port, input(36) => 
                           plus4A_out_36_port, input(35) => plus4A_out_35_port,
                           input(34) => plus4A_out_34_port, input(33) => 
                           plus4A_out_33_port, input(32) => plus4A_out_32_port,
                           input(31) => plus4A_out_31_port, input(30) => 
                           plus4A_out_30_port, input(29) => plus4A_out_29_port,
                           input(28) => plus4A_out_28_port, input(27) => 
                           plus4A_out_27_port, input(26) => plus4A_out_26_port,
                           input(25) => plus4A_out_25_port, input(24) => 
                           plus4A_out_24_port, input(23) => plus4A_out_23_port,
                           input(22) => plus4A_out_22_port, input(21) => 
                           plus4A_out_21_port, input(20) => plus4A_out_20_port,
                           input(19) => plus4A_out_19_port, input(18) => 
                           plus4A_out_18_port, input(17) => plus4A_out_17_port,
                           input(16) => plus4A_out_16_port, input(15) => 
                           plus4A_out_15_port, input(14) => plus4A_out_14_port,
                           input(13) => plus4A_out_13_port, input(12) => 
                           plus4A_out_12_port, input(11) => plus4A_out_11_port,
                           input(10) => plus4A_out_10_port, input(9) => 
                           plus4A_out_9_port, input(8) => plus4A_out_8_port, 
                           input(7) => plus4A_out_7_port, input(6) => 
                           plus4A_out_6_port, input(5) => plus4A_out_5_port, 
                           input(4) => plus4A_out_4_port, input(3) => 
                           plus4A_out_3_port, input(2) => plus4A_out_2_port, 
                           input(1) => plus4A_out_1_port, input(0) => 
                           plus4A_out_0_port, complement2(63) => 
                           minus4A_out(63), complement2(62) => minus4A_out(62),
                           complement2(61) => minus4A_out(61), complement2(60) 
                           => minus4A_out(60), complement2(59) => 
                           minus4A_out(59), complement2(58) => minus4A_out(58),
                           complement2(57) => minus4A_out(57), complement2(56) 
                           => minus4A_out(56), complement2(55) => 
                           minus4A_out(55), complement2(54) => minus4A_out(54),
                           complement2(53) => minus4A_out(53), complement2(52) 
                           => minus4A_out(52), complement2(51) => 
                           minus4A_out(51), complement2(50) => minus4A_out(50),
                           complement2(49) => minus4A_out(49), complement2(48) 
                           => minus4A_out(48), complement2(47) => 
                           minus4A_out(47), complement2(46) => minus4A_out(46),
                           complement2(45) => minus4A_out(45), complement2(44) 
                           => minus4A_out(44), complement2(43) => 
                           minus4A_out(43), complement2(42) => minus4A_out(42),
                           complement2(41) => minus4A_out(41), complement2(40) 
                           => minus4A_out(40), complement2(39) => 
                           minus4A_out(39), complement2(38) => minus4A_out(38),
                           complement2(37) => minus4A_out(37), complement2(36) 
                           => minus4A_out(36), complement2(35) => 
                           minus4A_out(35), complement2(34) => minus4A_out(34),
                           complement2(33) => minus4A_out(33), complement2(32) 
                           => minus4A_out(32), complement2(31) => 
                           minus4A_out(31), complement2(30) => minus4A_out(30),
                           complement2(29) => minus4A_out(29), complement2(28) 
                           => minus4A_out(28), complement2(27) => 
                           minus4A_out(27), complement2(26) => minus4A_out(26),
                           complement2(25) => minus4A_out(25), complement2(24) 
                           => minus4A_out(24), complement2(23) => 
                           minus4A_out(23), complement2(22) => minus4A_out(22),
                           complement2(21) => minus4A_out(21), complement2(20) 
                           => minus4A_out(20), complement2(19) => 
                           minus4A_out(19), complement2(18) => minus4A_out(18),
                           complement2(17) => minus4A_out(17), complement2(16) 
                           => minus4A_out(16), complement2(15) => 
                           minus4A_out(15), complement2(14) => minus4A_out(14),
                           complement2(13) => minus4A_out(13), complement2(12) 
                           => minus4A_out(12), complement2(11) => 
                           minus4A_out(11), complement2(10) => minus4A_out(10),
                           complement2(9) => minus4A_out(9), complement2(8) => 
                           minus4A_out(8), complement2(7) => minus4A_out(7), 
                           complement2(6) => minus4A_out(6), complement2(5) => 
                           minus4A_out(5), complement2(4) => minus4A_out(4), 
                           complement2(3) => minus4A_out(3), complement2(2) => 
                           minus4A_out(2), complement2(1) => minus4A_out(1), 
                           complement2(0) => minus4A_out(0));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity ShiftnCompl_N64_3 is

   port( plusA : in std_logic_vector (63 downto 0);  plus2A_out, minus2A_out, 
         plus4A_out, minus4A_out : out std_logic_vector (63 downto 0));

end ShiftnCompl_N64_3;

architecture SYN_struct of ShiftnCompl_N64_3 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component complementer_N64_5
      port( input : in std_logic_vector (63 downto 0);  complement2 : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component complementer_N64_6
      port( input : in std_logic_vector (63 downto 0);  complement2 : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component shifter_N64_5
      port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component shifter_N64_6
      port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
            std_logic_vector (63 downto 0));
   end component;
   
   signal plus2A_out_63_port, plus2A_out_62_port, plus2A_out_61_port, 
      plus2A_out_60_port, plus2A_out_59_port, plus2A_out_58_port, n26, n27, 
      plus2A_out_55_port, plus2A_out_54_port, plus2A_out_53_port, 
      plus2A_out_52_port, plus2A_out_51_port, plus2A_out_50_port, 
      plus2A_out_49_port, plus2A_out_48_port, plus2A_out_47_port, 
      plus2A_out_46_port, plus2A_out_45_port, plus2A_out_44_port, 
      plus2A_out_43_port, plus2A_out_42_port, plus2A_out_41_port, 
      plus2A_out_40_port, plus2A_out_39_port, plus2A_out_38_port, 
      plus2A_out_37_port, plus2A_out_36_port, plus2A_out_35_port, 
      plus2A_out_34_port, plus2A_out_33_port, plus2A_out_32_port, 
      plus2A_out_31_port, plus2A_out_30_port, plus2A_out_29_port, 
      plus2A_out_28_port, plus2A_out_27_port, plus2A_out_26_port, 
      plus2A_out_25_port, plus2A_out_24_port, plus2A_out_23_port, 
      plus2A_out_22_port, plus2A_out_21_port, plus2A_out_20_port, 
      plus2A_out_19_port, plus2A_out_18_port, plus2A_out_17_port, 
      plus2A_out_16_port, plus2A_out_15_port, plus2A_out_14_port, 
      plus2A_out_13_port, plus2A_out_12_port, plus2A_out_11_port, 
      plus2A_out_10_port, plus2A_out_9_port, plus2A_out_8_port, 
      plus2A_out_7_port, plus2A_out_6_port, plus2A_out_5_port, 
      plus2A_out_4_port, plus2A_out_3_port, plus2A_out_2_port, 
      plus2A_out_1_port, plus2A_out_0_port, plus4A_out_63_port, 
      plus4A_out_62_port, plus4A_out_61_port, plus4A_out_60_port, 
      plus4A_out_59_port, plus4A_out_58_port, plus4A_out_57_port, n28, n29, 
      plus4A_out_54_port, n30, n31, n32, plus4A_out_50_port, n33, n34, n35, 
      plus4A_out_46_port, n36, n37, n38, plus4A_out_42_port, n39, n40, n41, 
      plus4A_out_38_port, n42, n43, n44, plus4A_out_34_port, n45, n46, n47, 
      plus4A_out_30_port, n48, n49, n50, plus4A_out_26_port, plus4A_out_25_port
      , plus4A_out_24_port, plus4A_out_23_port, plus4A_out_22_port, 
      plus4A_out_21_port, plus4A_out_20_port, plus4A_out_19_port, 
      plus4A_out_18_port, plus4A_out_17_port, plus4A_out_16_port, 
      plus4A_out_15_port, plus4A_out_14_port, plus4A_out_13_port, 
      plus4A_out_12_port, plus4A_out_11_port, plus4A_out_10_port, 
      plus4A_out_9_port, plus4A_out_8_port, plus4A_out_7_port, 
      plus4A_out_6_port, plus4A_out_5_port, plus4A_out_4_port, 
      plus4A_out_3_port, plus4A_out_2_port, plus4A_out_1_port, 
      plus4A_out_0_port, plus4A_out_27_port, plus4A_out_28_port, 
      plus4A_out_29_port, plus4A_out_31_port, plus4A_out_32_port, 
      plus4A_out_33_port, plus4A_out_35_port, plus4A_out_36_port, 
      plus4A_out_37_port, plus4A_out_39_port, plus4A_out_40_port, 
      plus4A_out_41_port, plus4A_out_43_port, plus4A_out_44_port, 
      plus4A_out_45_port, plus4A_out_47_port, plus4A_out_48_port, 
      plus4A_out_49_port, plus4A_out_51_port, plus4A_out_52_port, 
      plus4A_out_53_port, plus4A_out_55_port, plus4A_out_56_port, 
      plus2A_out_56_port, plus2A_out_57_port, n_3148, n_3149 : std_logic;

begin
   plus2A_out <= ( plus2A_out_63_port, plus2A_out_62_port, plus2A_out_61_port, 
      plus2A_out_60_port, plus2A_out_59_port, plus2A_out_58_port, 
      plus2A_out_57_port, plus2A_out_56_port, plus2A_out_55_port, 
      plus2A_out_54_port, plus2A_out_53_port, plus2A_out_52_port, 
      plus2A_out_51_port, plus2A_out_50_port, plus2A_out_49_port, 
      plus2A_out_48_port, plus2A_out_47_port, plus2A_out_46_port, 
      plus2A_out_45_port, plus2A_out_44_port, plus2A_out_43_port, 
      plus2A_out_42_port, plus2A_out_41_port, plus2A_out_40_port, 
      plus2A_out_39_port, plus2A_out_38_port, plus2A_out_37_port, 
      plus2A_out_36_port, plus2A_out_35_port, plus2A_out_34_port, 
      plus2A_out_33_port, plus2A_out_32_port, plus2A_out_31_port, 
      plus2A_out_30_port, plus2A_out_29_port, plus2A_out_28_port, 
      plus2A_out_27_port, plus2A_out_26_port, plus2A_out_25_port, 
      plus2A_out_24_port, plus2A_out_23_port, plus2A_out_22_port, 
      plus2A_out_21_port, plus2A_out_20_port, plus2A_out_19_port, 
      plus2A_out_18_port, plus2A_out_17_port, plus2A_out_16_port, 
      plus2A_out_15_port, plus2A_out_14_port, plus2A_out_13_port, 
      plus2A_out_12_port, plus2A_out_11_port, plus2A_out_10_port, 
      plus2A_out_9_port, plus2A_out_8_port, plus2A_out_7_port, 
      plus2A_out_6_port, plus2A_out_5_port, plus2A_out_4_port, 
      plus2A_out_3_port, plus2A_out_2_port, plus2A_out_1_port, 
      plus2A_out_0_port );
   plus4A_out <= ( plus4A_out_63_port, plus4A_out_62_port, plus4A_out_61_port, 
      plus4A_out_60_port, plus4A_out_59_port, plus4A_out_58_port, 
      plus4A_out_57_port, plus4A_out_56_port, plus4A_out_55_port, 
      plus4A_out_54_port, plus4A_out_53_port, plus4A_out_52_port, 
      plus4A_out_51_port, plus4A_out_50_port, plus4A_out_49_port, 
      plus4A_out_48_port, plus4A_out_47_port, plus4A_out_46_port, 
      plus4A_out_45_port, plus4A_out_44_port, plus4A_out_43_port, 
      plus4A_out_42_port, plus4A_out_41_port, plus4A_out_40_port, 
      plus4A_out_39_port, plus4A_out_38_port, plus4A_out_37_port, 
      plus4A_out_36_port, plus4A_out_35_port, plus4A_out_34_port, 
      plus4A_out_33_port, plus4A_out_32_port, plus4A_out_31_port, 
      plus4A_out_30_port, plus4A_out_29_port, plus4A_out_28_port, 
      plus4A_out_27_port, plus4A_out_26_port, plus4A_out_25_port, 
      plus4A_out_24_port, plus4A_out_23_port, plus4A_out_22_port, 
      plus4A_out_21_port, plus4A_out_20_port, plus4A_out_19_port, 
      plus4A_out_18_port, plus4A_out_17_port, plus4A_out_16_port, 
      plus4A_out_15_port, plus4A_out_14_port, plus4A_out_13_port, 
      plus4A_out_12_port, plus4A_out_11_port, plus4A_out_10_port, 
      plus4A_out_9_port, plus4A_out_8_port, plus4A_out_7_port, 
      plus4A_out_6_port, plus4A_out_5_port, plus4A_out_4_port, 
      plus4A_out_3_port, plus4A_out_2_port, plus4A_out_1_port, 
      plus4A_out_0_port );
   
   plus2A_out_0_port <= '0';
   plus4A_out_0_port <= '0';
   shifter_1 : shifter_N64_6 port map( input(63) => plusA(63), input(62) => 
                           plusA(62), input(61) => plusA(61), input(60) => 
                           plusA(60), input(59) => plusA(59), input(58) => 
                           plusA(58), input(57) => plusA(57), input(56) => 
                           plusA(56), input(55) => plusA(55), input(54) => 
                           plusA(54), input(53) => plusA(53), input(52) => 
                           plusA(52), input(51) => plusA(51), input(50) => 
                           plusA(50), input(49) => plusA(49), input(48) => 
                           plusA(48), input(47) => plusA(47), input(46) => 
                           plusA(46), input(45) => plusA(45), input(44) => 
                           plusA(44), input(43) => plusA(43), input(42) => 
                           plusA(42), input(41) => plusA(41), input(40) => 
                           plusA(40), input(39) => plusA(39), input(38) => 
                           plusA(38), input(37) => plusA(37), input(36) => 
                           plusA(36), input(35) => plusA(35), input(34) => 
                           plusA(34), input(33) => plusA(33), input(32) => 
                           plusA(32), input(31) => plusA(31), input(30) => 
                           plusA(30), input(29) => plusA(29), input(28) => 
                           plusA(28), input(27) => plusA(27), input(26) => 
                           plusA(26), input(25) => plusA(25), input(24) => 
                           plusA(24), input(23) => plusA(23), input(22) => 
                           plusA(22), input(21) => plusA(21), input(20) => 
                           plusA(20), input(19) => plusA(19), input(18) => 
                           plusA(18), input(17) => plusA(17), input(16) => 
                           plusA(16), input(15) => plusA(15), input(14) => 
                           plusA(14), input(13) => plusA(13), input(12) => 
                           plusA(12), input(11) => plusA(11), input(10) => 
                           plusA(10), input(9) => plusA(9), input(8) => 
                           plusA(8), input(7) => plusA(7), input(6) => plusA(6)
                           , input(5) => plusA(5), input(4) => plusA(4), 
                           input(3) => plusA(3), input(2) => plusA(2), input(1)
                           => plusA(1), input(0) => plusA(0), 
                           shiftLeftOnePos(63) => plus2A_out_63_port, 
                           shiftLeftOnePos(62) => plus2A_out_62_port, 
                           shiftLeftOnePos(61) => plus2A_out_61_port, 
                           shiftLeftOnePos(60) => plus2A_out_60_port, 
                           shiftLeftOnePos(59) => plus2A_out_59_port, 
                           shiftLeftOnePos(58) => plus2A_out_58_port, 
                           shiftLeftOnePos(57) => n26, shiftLeftOnePos(56) => 
                           n27, shiftLeftOnePos(55) => plus2A_out_55_port, 
                           shiftLeftOnePos(54) => plus2A_out_54_port, 
                           shiftLeftOnePos(53) => plus2A_out_53_port, 
                           shiftLeftOnePos(52) => plus2A_out_52_port, 
                           shiftLeftOnePos(51) => plus2A_out_51_port, 
                           shiftLeftOnePos(50) => plus2A_out_50_port, 
                           shiftLeftOnePos(49) => plus2A_out_49_port, 
                           shiftLeftOnePos(48) => plus2A_out_48_port, 
                           shiftLeftOnePos(47) => plus2A_out_47_port, 
                           shiftLeftOnePos(46) => plus2A_out_46_port, 
                           shiftLeftOnePos(45) => plus2A_out_45_port, 
                           shiftLeftOnePos(44) => plus2A_out_44_port, 
                           shiftLeftOnePos(43) => plus2A_out_43_port, 
                           shiftLeftOnePos(42) => plus2A_out_42_port, 
                           shiftLeftOnePos(41) => plus2A_out_41_port, 
                           shiftLeftOnePos(40) => plus2A_out_40_port, 
                           shiftLeftOnePos(39) => plus2A_out_39_port, 
                           shiftLeftOnePos(38) => plus2A_out_38_port, 
                           shiftLeftOnePos(37) => plus2A_out_37_port, 
                           shiftLeftOnePos(36) => plus2A_out_36_port, 
                           shiftLeftOnePos(35) => plus2A_out_35_port, 
                           shiftLeftOnePos(34) => plus2A_out_34_port, 
                           shiftLeftOnePos(33) => plus2A_out_33_port, 
                           shiftLeftOnePos(32) => plus2A_out_32_port, 
                           shiftLeftOnePos(31) => plus2A_out_31_port, 
                           shiftLeftOnePos(30) => plus2A_out_30_port, 
                           shiftLeftOnePos(29) => plus2A_out_29_port, 
                           shiftLeftOnePos(28) => plus2A_out_28_port, 
                           shiftLeftOnePos(27) => plus2A_out_27_port, 
                           shiftLeftOnePos(26) => plus2A_out_26_port, 
                           shiftLeftOnePos(25) => plus2A_out_25_port, 
                           shiftLeftOnePos(24) => plus2A_out_24_port, 
                           shiftLeftOnePos(23) => plus2A_out_23_port, 
                           shiftLeftOnePos(22) => plus2A_out_22_port, 
                           shiftLeftOnePos(21) => plus2A_out_21_port, 
                           shiftLeftOnePos(20) => plus2A_out_20_port, 
                           shiftLeftOnePos(19) => plus2A_out_19_port, 
                           shiftLeftOnePos(18) => plus2A_out_18_port, 
                           shiftLeftOnePos(17) => plus2A_out_17_port, 
                           shiftLeftOnePos(16) => plus2A_out_16_port, 
                           shiftLeftOnePos(15) => plus2A_out_15_port, 
                           shiftLeftOnePos(14) => plus2A_out_14_port, 
                           shiftLeftOnePos(13) => plus2A_out_13_port, 
                           shiftLeftOnePos(12) => plus2A_out_12_port, 
                           shiftLeftOnePos(11) => plus2A_out_11_port, 
                           shiftLeftOnePos(10) => plus2A_out_10_port, 
                           shiftLeftOnePos(9) => plus2A_out_9_port, 
                           shiftLeftOnePos(8) => plus2A_out_8_port, 
                           shiftLeftOnePos(7) => plus2A_out_7_port, 
                           shiftLeftOnePos(6) => plus2A_out_6_port, 
                           shiftLeftOnePos(5) => plus2A_out_5_port, 
                           shiftLeftOnePos(4) => plus2A_out_4_port, 
                           shiftLeftOnePos(3) => plus2A_out_3_port, 
                           shiftLeftOnePos(2) => plus2A_out_2_port, 
                           shiftLeftOnePos(1) => plus2A_out_1_port, 
                           shiftLeftOnePos(0) => n_3148);
   shifter_2 : shifter_N64_5 port map( input(63) => plus2A_out_63_port, 
                           input(62) => plus2A_out_62_port, input(61) => 
                           plus2A_out_61_port, input(60) => plus2A_out_60_port,
                           input(59) => plus2A_out_59_port, input(58) => 
                           plus2A_out_58_port, input(57) => plus2A_out_57_port,
                           input(56) => plus2A_out_56_port, input(55) => 
                           plus2A_out_55_port, input(54) => plus2A_out_54_port,
                           input(53) => plus2A_out_53_port, input(52) => 
                           plus2A_out_52_port, input(51) => plus2A_out_51_port,
                           input(50) => plus2A_out_50_port, input(49) => 
                           plus2A_out_49_port, input(48) => plus2A_out_48_port,
                           input(47) => plus2A_out_47_port, input(46) => 
                           plus2A_out_46_port, input(45) => plus2A_out_45_port,
                           input(44) => plus2A_out_44_port, input(43) => 
                           plus2A_out_43_port, input(42) => plus2A_out_42_port,
                           input(41) => plus2A_out_41_port, input(40) => 
                           plus2A_out_40_port, input(39) => plus2A_out_39_port,
                           input(38) => plus2A_out_38_port, input(37) => 
                           plus2A_out_37_port, input(36) => plus2A_out_36_port,
                           input(35) => plus2A_out_35_port, input(34) => 
                           plus2A_out_34_port, input(33) => plus2A_out_33_port,
                           input(32) => plus2A_out_32_port, input(31) => 
                           plus2A_out_31_port, input(30) => plus2A_out_30_port,
                           input(29) => plus2A_out_29_port, input(28) => 
                           plus2A_out_28_port, input(27) => plus2A_out_27_port,
                           input(26) => plus2A_out_26_port, input(25) => 
                           plus2A_out_25_port, input(24) => plus2A_out_24_port,
                           input(23) => plus2A_out_23_port, input(22) => 
                           plus2A_out_22_port, input(21) => plus2A_out_21_port,
                           input(20) => plus2A_out_20_port, input(19) => 
                           plus2A_out_19_port, input(18) => plus2A_out_18_port,
                           input(17) => plus2A_out_17_port, input(16) => 
                           plus2A_out_16_port, input(15) => plus2A_out_15_port,
                           input(14) => plus2A_out_14_port, input(13) => 
                           plus2A_out_13_port, input(12) => plus2A_out_12_port,
                           input(11) => plus2A_out_11_port, input(10) => 
                           plus2A_out_10_port, input(9) => plus2A_out_9_port, 
                           input(8) => plus2A_out_8_port, input(7) => 
                           plus2A_out_7_port, input(6) => plus2A_out_6_port, 
                           input(5) => plus2A_out_5_port, input(4) => 
                           plus2A_out_4_port, input(3) => plus2A_out_3_port, 
                           input(2) => plus2A_out_2_port, input(1) => 
                           plus2A_out_1_port, input(0) => plus2A_out_0_port, 
                           shiftLeftOnePos(63) => plus4A_out_63_port, 
                           shiftLeftOnePos(62) => plus4A_out_62_port, 
                           shiftLeftOnePos(61) => plus4A_out_61_port, 
                           shiftLeftOnePos(60) => plus4A_out_60_port, 
                           shiftLeftOnePos(59) => plus4A_out_59_port, 
                           shiftLeftOnePos(58) => plus4A_out_58_port, 
                           shiftLeftOnePos(57) => plus4A_out_57_port, 
                           shiftLeftOnePos(56) => n28, shiftLeftOnePos(55) => 
                           n29, shiftLeftOnePos(54) => plus4A_out_54_port, 
                           shiftLeftOnePos(53) => n30, shiftLeftOnePos(52) => 
                           n31, shiftLeftOnePos(51) => n32, shiftLeftOnePos(50)
                           => plus4A_out_50_port, shiftLeftOnePos(49) => n33, 
                           shiftLeftOnePos(48) => n34, shiftLeftOnePos(47) => 
                           n35, shiftLeftOnePos(46) => plus4A_out_46_port, 
                           shiftLeftOnePos(45) => n36, shiftLeftOnePos(44) => 
                           n37, shiftLeftOnePos(43) => n38, shiftLeftOnePos(42)
                           => plus4A_out_42_port, shiftLeftOnePos(41) => n39, 
                           shiftLeftOnePos(40) => n40, shiftLeftOnePos(39) => 
                           n41, shiftLeftOnePos(38) => plus4A_out_38_port, 
                           shiftLeftOnePos(37) => n42, shiftLeftOnePos(36) => 
                           n43, shiftLeftOnePos(35) => n44, shiftLeftOnePos(34)
                           => plus4A_out_34_port, shiftLeftOnePos(33) => n45, 
                           shiftLeftOnePos(32) => n46, shiftLeftOnePos(31) => 
                           n47, shiftLeftOnePos(30) => plus4A_out_30_port, 
                           shiftLeftOnePos(29) => n48, shiftLeftOnePos(28) => 
                           n49, shiftLeftOnePos(27) => n50, shiftLeftOnePos(26)
                           => plus4A_out_26_port, shiftLeftOnePos(25) => 
                           plus4A_out_25_port, shiftLeftOnePos(24) => 
                           plus4A_out_24_port, shiftLeftOnePos(23) => 
                           plus4A_out_23_port, shiftLeftOnePos(22) => 
                           plus4A_out_22_port, shiftLeftOnePos(21) => 
                           plus4A_out_21_port, shiftLeftOnePos(20) => 
                           plus4A_out_20_port, shiftLeftOnePos(19) => 
                           plus4A_out_19_port, shiftLeftOnePos(18) => 
                           plus4A_out_18_port, shiftLeftOnePos(17) => 
                           plus4A_out_17_port, shiftLeftOnePos(16) => 
                           plus4A_out_16_port, shiftLeftOnePos(15) => 
                           plus4A_out_15_port, shiftLeftOnePos(14) => 
                           plus4A_out_14_port, shiftLeftOnePos(13) => 
                           plus4A_out_13_port, shiftLeftOnePos(12) => 
                           plus4A_out_12_port, shiftLeftOnePos(11) => 
                           plus4A_out_11_port, shiftLeftOnePos(10) => 
                           plus4A_out_10_port, shiftLeftOnePos(9) => 
                           plus4A_out_9_port, shiftLeftOnePos(8) => 
                           plus4A_out_8_port, shiftLeftOnePos(7) => 
                           plus4A_out_7_port, shiftLeftOnePos(6) => 
                           plus4A_out_6_port, shiftLeftOnePos(5) => 
                           plus4A_out_5_port, shiftLeftOnePos(4) => 
                           plus4A_out_4_port, shiftLeftOnePos(3) => 
                           plus4A_out_3_port, shiftLeftOnePos(2) => 
                           plus4A_out_2_port, shiftLeftOnePos(1) => 
                           plus4A_out_1_port, shiftLeftOnePos(0) => n_3149);
   complementer_1 : complementer_N64_6 port map( input(63) => 
                           plus2A_out_63_port, input(62) => plus2A_out_62_port,
                           input(61) => plus2A_out_61_port, input(60) => 
                           plus2A_out_60_port, input(59) => plus2A_out_59_port,
                           input(58) => plus2A_out_58_port, input(57) => 
                           plus2A_out_57_port, input(56) => plus2A_out_56_port,
                           input(55) => plus2A_out_55_port, input(54) => 
                           plus2A_out_54_port, input(53) => plus2A_out_53_port,
                           input(52) => plus2A_out_52_port, input(51) => 
                           plus2A_out_51_port, input(50) => plus2A_out_50_port,
                           input(49) => plus2A_out_49_port, input(48) => 
                           plus2A_out_48_port, input(47) => plus2A_out_47_port,
                           input(46) => plus2A_out_46_port, input(45) => 
                           plus2A_out_45_port, input(44) => plus2A_out_44_port,
                           input(43) => plus2A_out_43_port, input(42) => 
                           plus2A_out_42_port, input(41) => plus2A_out_41_port,
                           input(40) => plus2A_out_40_port, input(39) => 
                           plus2A_out_39_port, input(38) => plus2A_out_38_port,
                           input(37) => plus2A_out_37_port, input(36) => 
                           plus2A_out_36_port, input(35) => plus2A_out_35_port,
                           input(34) => plus2A_out_34_port, input(33) => 
                           plus2A_out_33_port, input(32) => plus2A_out_32_port,
                           input(31) => plus2A_out_31_port, input(30) => 
                           plus2A_out_30_port, input(29) => plus2A_out_29_port,
                           input(28) => plus2A_out_28_port, input(27) => 
                           plus2A_out_27_port, input(26) => plus2A_out_26_port,
                           input(25) => plus2A_out_25_port, input(24) => 
                           plus2A_out_24_port, input(23) => plus2A_out_23_port,
                           input(22) => plus2A_out_22_port, input(21) => 
                           plus2A_out_21_port, input(20) => plus2A_out_20_port,
                           input(19) => plus2A_out_19_port, input(18) => 
                           plus2A_out_18_port, input(17) => plus2A_out_17_port,
                           input(16) => plus2A_out_16_port, input(15) => 
                           plus2A_out_15_port, input(14) => plus2A_out_14_port,
                           input(13) => plus2A_out_13_port, input(12) => 
                           plus2A_out_12_port, input(11) => plus2A_out_11_port,
                           input(10) => plus2A_out_10_port, input(9) => 
                           plus2A_out_9_port, input(8) => plus2A_out_8_port, 
                           input(7) => plus2A_out_7_port, input(6) => 
                           plus2A_out_6_port, input(5) => plus2A_out_5_port, 
                           input(4) => plus2A_out_4_port, input(3) => 
                           plus2A_out_3_port, input(2) => plus2A_out_2_port, 
                           input(1) => plus2A_out_1_port, input(0) => 
                           plus2A_out_0_port, complement2(63) => 
                           minus2A_out(63), complement2(62) => minus2A_out(62),
                           complement2(61) => minus2A_out(61), complement2(60) 
                           => minus2A_out(60), complement2(59) => 
                           minus2A_out(59), complement2(58) => minus2A_out(58),
                           complement2(57) => minus2A_out(57), complement2(56) 
                           => minus2A_out(56), complement2(55) => 
                           minus2A_out(55), complement2(54) => minus2A_out(54),
                           complement2(53) => minus2A_out(53), complement2(52) 
                           => minus2A_out(52), complement2(51) => 
                           minus2A_out(51), complement2(50) => minus2A_out(50),
                           complement2(49) => minus2A_out(49), complement2(48) 
                           => minus2A_out(48), complement2(47) => 
                           minus2A_out(47), complement2(46) => minus2A_out(46),
                           complement2(45) => minus2A_out(45), complement2(44) 
                           => minus2A_out(44), complement2(43) => 
                           minus2A_out(43), complement2(42) => minus2A_out(42),
                           complement2(41) => minus2A_out(41), complement2(40) 
                           => minus2A_out(40), complement2(39) => 
                           minus2A_out(39), complement2(38) => minus2A_out(38),
                           complement2(37) => minus2A_out(37), complement2(36) 
                           => minus2A_out(36), complement2(35) => 
                           minus2A_out(35), complement2(34) => minus2A_out(34),
                           complement2(33) => minus2A_out(33), complement2(32) 
                           => minus2A_out(32), complement2(31) => 
                           minus2A_out(31), complement2(30) => minus2A_out(30),
                           complement2(29) => minus2A_out(29), complement2(28) 
                           => minus2A_out(28), complement2(27) => 
                           minus2A_out(27), complement2(26) => minus2A_out(26),
                           complement2(25) => minus2A_out(25), complement2(24) 
                           => minus2A_out(24), complement2(23) => 
                           minus2A_out(23), complement2(22) => minus2A_out(22),
                           complement2(21) => minus2A_out(21), complement2(20) 
                           => minus2A_out(20), complement2(19) => 
                           minus2A_out(19), complement2(18) => minus2A_out(18),
                           complement2(17) => minus2A_out(17), complement2(16) 
                           => minus2A_out(16), complement2(15) => 
                           minus2A_out(15), complement2(14) => minus2A_out(14),
                           complement2(13) => minus2A_out(13), complement2(12) 
                           => minus2A_out(12), complement2(11) => 
                           minus2A_out(11), complement2(10) => minus2A_out(10),
                           complement2(9) => minus2A_out(9), complement2(8) => 
                           minus2A_out(8), complement2(7) => minus2A_out(7), 
                           complement2(6) => minus2A_out(6), complement2(5) => 
                           minus2A_out(5), complement2(4) => minus2A_out(4), 
                           complement2(3) => minus2A_out(3), complement2(2) => 
                           minus2A_out(2), complement2(1) => minus2A_out(1), 
                           complement2(0) => minus2A_out(0));
   complementer_2 : complementer_N64_5 port map( input(63) => 
                           plus4A_out_63_port, input(62) => plus4A_out_62_port,
                           input(61) => plus4A_out_61_port, input(60) => 
                           plus4A_out_60_port, input(59) => plus4A_out_59_port,
                           input(58) => plus4A_out_58_port, input(57) => 
                           plus4A_out_57_port, input(56) => plus4A_out_56_port,
                           input(55) => plus4A_out_55_port, input(54) => 
                           plus4A_out_54_port, input(53) => plus4A_out_53_port,
                           input(52) => plus4A_out_52_port, input(51) => 
                           plus4A_out_51_port, input(50) => plus4A_out_50_port,
                           input(49) => plus4A_out_49_port, input(48) => 
                           plus4A_out_48_port, input(47) => plus4A_out_47_port,
                           input(46) => plus4A_out_46_port, input(45) => 
                           plus4A_out_45_port, input(44) => plus4A_out_44_port,
                           input(43) => plus4A_out_43_port, input(42) => 
                           plus4A_out_42_port, input(41) => plus4A_out_41_port,
                           input(40) => plus4A_out_40_port, input(39) => 
                           plus4A_out_39_port, input(38) => plus4A_out_38_port,
                           input(37) => plus4A_out_37_port, input(36) => 
                           plus4A_out_36_port, input(35) => plus4A_out_35_port,
                           input(34) => plus4A_out_34_port, input(33) => 
                           plus4A_out_33_port, input(32) => plus4A_out_32_port,
                           input(31) => plus4A_out_31_port, input(30) => 
                           plus4A_out_30_port, input(29) => plus4A_out_29_port,
                           input(28) => plus4A_out_28_port, input(27) => 
                           plus4A_out_27_port, input(26) => plus4A_out_26_port,
                           input(25) => plus4A_out_25_port, input(24) => 
                           plus4A_out_24_port, input(23) => plus4A_out_23_port,
                           input(22) => plus4A_out_22_port, input(21) => 
                           plus4A_out_21_port, input(20) => plus4A_out_20_port,
                           input(19) => plus4A_out_19_port, input(18) => 
                           plus4A_out_18_port, input(17) => plus4A_out_17_port,
                           input(16) => plus4A_out_16_port, input(15) => 
                           plus4A_out_15_port, input(14) => plus4A_out_14_port,
                           input(13) => plus4A_out_13_port, input(12) => 
                           plus4A_out_12_port, input(11) => plus4A_out_11_port,
                           input(10) => plus4A_out_10_port, input(9) => 
                           plus4A_out_9_port, input(8) => plus4A_out_8_port, 
                           input(7) => plus4A_out_7_port, input(6) => 
                           plus4A_out_6_port, input(5) => plus4A_out_5_port, 
                           input(4) => plus4A_out_4_port, input(3) => 
                           plus4A_out_3_port, input(2) => plus4A_out_2_port, 
                           input(1) => plus4A_out_1_port, input(0) => 
                           plus4A_out_0_port, complement2(63) => 
                           minus4A_out(63), complement2(62) => minus4A_out(62),
                           complement2(61) => minus4A_out(61), complement2(60) 
                           => minus4A_out(60), complement2(59) => 
                           minus4A_out(59), complement2(58) => minus4A_out(58),
                           complement2(57) => minus4A_out(57), complement2(56) 
                           => minus4A_out(56), complement2(55) => 
                           minus4A_out(55), complement2(54) => minus4A_out(54),
                           complement2(53) => minus4A_out(53), complement2(52) 
                           => minus4A_out(52), complement2(51) => 
                           minus4A_out(51), complement2(50) => minus4A_out(50),
                           complement2(49) => minus4A_out(49), complement2(48) 
                           => minus4A_out(48), complement2(47) => 
                           minus4A_out(47), complement2(46) => minus4A_out(46),
                           complement2(45) => minus4A_out(45), complement2(44) 
                           => minus4A_out(44), complement2(43) => 
                           minus4A_out(43), complement2(42) => minus4A_out(42),
                           complement2(41) => minus4A_out(41), complement2(40) 
                           => minus4A_out(40), complement2(39) => 
                           minus4A_out(39), complement2(38) => minus4A_out(38),
                           complement2(37) => minus4A_out(37), complement2(36) 
                           => minus4A_out(36), complement2(35) => 
                           minus4A_out(35), complement2(34) => minus4A_out(34),
                           complement2(33) => minus4A_out(33), complement2(32) 
                           => minus4A_out(32), complement2(31) => 
                           minus4A_out(31), complement2(30) => minus4A_out(30),
                           complement2(29) => minus4A_out(29), complement2(28) 
                           => minus4A_out(28), complement2(27) => 
                           minus4A_out(27), complement2(26) => minus4A_out(26),
                           complement2(25) => minus4A_out(25), complement2(24) 
                           => minus4A_out(24), complement2(23) => 
                           minus4A_out(23), complement2(22) => minus4A_out(22),
                           complement2(21) => minus4A_out(21), complement2(20) 
                           => minus4A_out(20), complement2(19) => 
                           minus4A_out(19), complement2(18) => minus4A_out(18),
                           complement2(17) => minus4A_out(17), complement2(16) 
                           => minus4A_out(16), complement2(15) => 
                           minus4A_out(15), complement2(14) => minus4A_out(14),
                           complement2(13) => minus4A_out(13), complement2(12) 
                           => minus4A_out(12), complement2(11) => 
                           minus4A_out(11), complement2(10) => minus4A_out(10),
                           complement2(9) => minus4A_out(9), complement2(8) => 
                           minus4A_out(8), complement2(7) => minus4A_out(7), 
                           complement2(6) => minus4A_out(6), complement2(5) => 
                           minus4A_out(5), complement2(4) => minus4A_out(4), 
                           complement2(3) => minus4A_out(3), complement2(2) => 
                           minus4A_out(2), complement2(1) => minus4A_out(1), 
                           complement2(0) => minus4A_out(0));
   U3 : BUF_X1 port map( A => n47, Z => plus4A_out_31_port);
   U4 : BUF_X1 port map( A => n50, Z => plus4A_out_27_port);
   U5 : BUF_X1 port map( A => n45, Z => plus4A_out_33_port);
   U6 : BUF_X1 port map( A => n48, Z => plus4A_out_29_port);
   U7 : BUF_X1 port map( A => n46, Z => plus4A_out_32_port);
   U8 : BUF_X1 port map( A => n49, Z => plus4A_out_28_port);
   U9 : BUF_X1 port map( A => n38, Z => plus4A_out_43_port);
   U10 : BUF_X1 port map( A => n41, Z => plus4A_out_39_port);
   U11 : BUF_X1 port map( A => n44, Z => plus4A_out_35_port);
   U12 : BUF_X1 port map( A => n36, Z => plus4A_out_45_port);
   U13 : BUF_X1 port map( A => n39, Z => plus4A_out_41_port);
   U14 : BUF_X1 port map( A => n42, Z => plus4A_out_37_port);
   U15 : BUF_X1 port map( A => n37, Z => plus4A_out_44_port);
   U16 : BUF_X1 port map( A => n40, Z => plus4A_out_40_port);
   U17 : BUF_X1 port map( A => n43, Z => plus4A_out_36_port);
   U18 : BUF_X1 port map( A => n27, Z => plus2A_out_56_port);
   U19 : BUF_X1 port map( A => n26, Z => plus2A_out_57_port);
   U20 : BUF_X1 port map( A => n32, Z => plus4A_out_51_port);
   U21 : BUF_X1 port map( A => n35, Z => plus4A_out_47_port);
   U22 : BUF_X1 port map( A => n29, Z => plus4A_out_55_port);
   U23 : BUF_X1 port map( A => n30, Z => plus4A_out_53_port);
   U24 : BUF_X1 port map( A => n33, Z => plus4A_out_49_port);
   U25 : BUF_X1 port map( A => n28, Z => plus4A_out_56_port);
   U26 : BUF_X1 port map( A => n31, Z => plus4A_out_52_port);
   U27 : BUF_X1 port map( A => n34, Z => plus4A_out_48_port);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity ShiftnCompl_N64_4 is

   port( plusA : in std_logic_vector (63 downto 0);  plus2A_out, minus2A_out, 
         plus4A_out, minus4A_out : out std_logic_vector (63 downto 0));

end ShiftnCompl_N64_4;

architecture SYN_struct of ShiftnCompl_N64_4 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component complementer_N64_7
      port( input : in std_logic_vector (63 downto 0);  complement2 : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component complementer_N64_8
      port( input : in std_logic_vector (63 downto 0);  complement2 : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component shifter_N64_7
      port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component shifter_N64_8
      port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
            std_logic_vector (63 downto 0));
   end component;
   
   signal plus2A_out_63_port, plus2A_out_62_port, plus2A_out_61_port, 
      plus2A_out_60_port, plus2A_out_59_port, plus2A_out_58_port, n2, 
      plus2A_out_56_port, plus2A_out_55_port, plus2A_out_54_port, 
      plus2A_out_53_port, plus2A_out_52_port, plus2A_out_51_port, 
      plus2A_out_50_port, plus2A_out_49_port, plus2A_out_48_port, 
      plus2A_out_47_port, plus2A_out_46_port, plus2A_out_45_port, 
      plus2A_out_44_port, plus2A_out_43_port, plus2A_out_42_port, 
      plus2A_out_41_port, plus2A_out_40_port, plus2A_out_39_port, 
      plus2A_out_38_port, plus2A_out_37_port, plus2A_out_36_port, 
      plus2A_out_35_port, plus2A_out_34_port, plus2A_out_33_port, 
      plus2A_out_32_port, plus2A_out_31_port, plus2A_out_30_port, 
      plus2A_out_29_port, plus2A_out_28_port, plus2A_out_27_port, 
      plus2A_out_26_port, plus2A_out_25_port, plus2A_out_24_port, 
      plus2A_out_23_port, plus2A_out_22_port, plus2A_out_21_port, 
      plus2A_out_20_port, plus2A_out_19_port, plus2A_out_18_port, 
      plus2A_out_17_port, plus2A_out_16_port, plus2A_out_15_port, 
      plus2A_out_14_port, plus2A_out_13_port, plus2A_out_12_port, 
      plus2A_out_11_port, plus2A_out_10_port, plus2A_out_9_port, 
      plus2A_out_8_port, plus2A_out_7_port, plus2A_out_6_port, 
      plus2A_out_5_port, plus2A_out_4_port, plus2A_out_3_port, 
      plus2A_out_2_port, plus2A_out_1_port, plus2A_out_0_port, 
      plus4A_out_63_port, plus4A_out_62_port, plus4A_out_61_port, 
      plus4A_out_60_port, plus4A_out_59_port, plus4A_out_58_port, 
      plus4A_out_57_port, plus4A_out_56_port, plus4A_out_55_port, 
      plus4A_out_54_port, plus4A_out_53_port, plus4A_out_52_port, 
      plus4A_out_51_port, plus4A_out_50_port, plus4A_out_49_port, 
      plus4A_out_48_port, plus4A_out_47_port, plus4A_out_46_port, 
      plus4A_out_45_port, plus4A_out_44_port, plus4A_out_43_port, 
      plus4A_out_42_port, plus4A_out_41_port, plus4A_out_40_port, 
      plus4A_out_39_port, plus4A_out_38_port, plus4A_out_37_port, 
      plus4A_out_36_port, plus4A_out_35_port, plus4A_out_34_port, 
      plus4A_out_33_port, plus4A_out_32_port, plus4A_out_31_port, 
      plus4A_out_30_port, plus4A_out_29_port, plus4A_out_28_port, 
      plus4A_out_27_port, plus4A_out_26_port, plus4A_out_25_port, 
      plus4A_out_24_port, plus4A_out_23_port, plus4A_out_22_port, 
      plus4A_out_21_port, plus4A_out_20_port, plus4A_out_19_port, 
      plus4A_out_18_port, plus4A_out_17_port, plus4A_out_16_port, 
      plus4A_out_15_port, plus4A_out_14_port, plus4A_out_13_port, 
      plus4A_out_12_port, plus4A_out_11_port, plus4A_out_10_port, 
      plus4A_out_9_port, plus4A_out_8_port, plus4A_out_7_port, 
      plus4A_out_6_port, plus4A_out_5_port, plus4A_out_4_port, 
      plus4A_out_3_port, plus4A_out_2_port, plus4A_out_1_port, 
      plus4A_out_0_port, plus2A_out_57_port, n_3150, n_3151 : std_logic;

begin
   plus2A_out <= ( plus2A_out_63_port, plus2A_out_62_port, plus2A_out_61_port, 
      plus2A_out_60_port, plus2A_out_59_port, plus2A_out_58_port, 
      plus2A_out_57_port, plus2A_out_56_port, plus2A_out_55_port, 
      plus2A_out_54_port, plus2A_out_53_port, plus2A_out_52_port, 
      plus2A_out_51_port, plus2A_out_50_port, plus2A_out_49_port, 
      plus2A_out_48_port, plus2A_out_47_port, plus2A_out_46_port, 
      plus2A_out_45_port, plus2A_out_44_port, plus2A_out_43_port, 
      plus2A_out_42_port, plus2A_out_41_port, plus2A_out_40_port, 
      plus2A_out_39_port, plus2A_out_38_port, plus2A_out_37_port, 
      plus2A_out_36_port, plus2A_out_35_port, plus2A_out_34_port, 
      plus2A_out_33_port, plus2A_out_32_port, plus2A_out_31_port, 
      plus2A_out_30_port, plus2A_out_29_port, plus2A_out_28_port, 
      plus2A_out_27_port, plus2A_out_26_port, plus2A_out_25_port, 
      plus2A_out_24_port, plus2A_out_23_port, plus2A_out_22_port, 
      plus2A_out_21_port, plus2A_out_20_port, plus2A_out_19_port, 
      plus2A_out_18_port, plus2A_out_17_port, plus2A_out_16_port, 
      plus2A_out_15_port, plus2A_out_14_port, plus2A_out_13_port, 
      plus2A_out_12_port, plus2A_out_11_port, plus2A_out_10_port, 
      plus2A_out_9_port, plus2A_out_8_port, plus2A_out_7_port, 
      plus2A_out_6_port, plus2A_out_5_port, plus2A_out_4_port, 
      plus2A_out_3_port, plus2A_out_2_port, plus2A_out_1_port, 
      plus2A_out_0_port );
   plus4A_out <= ( plus4A_out_63_port, plus4A_out_62_port, plus4A_out_61_port, 
      plus4A_out_60_port, plus4A_out_59_port, plus4A_out_58_port, 
      plus4A_out_57_port, plus4A_out_56_port, plus4A_out_55_port, 
      plus4A_out_54_port, plus4A_out_53_port, plus4A_out_52_port, 
      plus4A_out_51_port, plus4A_out_50_port, plus4A_out_49_port, 
      plus4A_out_48_port, plus4A_out_47_port, plus4A_out_46_port, 
      plus4A_out_45_port, plus4A_out_44_port, plus4A_out_43_port, 
      plus4A_out_42_port, plus4A_out_41_port, plus4A_out_40_port, 
      plus4A_out_39_port, plus4A_out_38_port, plus4A_out_37_port, 
      plus4A_out_36_port, plus4A_out_35_port, plus4A_out_34_port, 
      plus4A_out_33_port, plus4A_out_32_port, plus4A_out_31_port, 
      plus4A_out_30_port, plus4A_out_29_port, plus4A_out_28_port, 
      plus4A_out_27_port, plus4A_out_26_port, plus4A_out_25_port, 
      plus4A_out_24_port, plus4A_out_23_port, plus4A_out_22_port, 
      plus4A_out_21_port, plus4A_out_20_port, plus4A_out_19_port, 
      plus4A_out_18_port, plus4A_out_17_port, plus4A_out_16_port, 
      plus4A_out_15_port, plus4A_out_14_port, plus4A_out_13_port, 
      plus4A_out_12_port, plus4A_out_11_port, plus4A_out_10_port, 
      plus4A_out_9_port, plus4A_out_8_port, plus4A_out_7_port, 
      plus4A_out_6_port, plus4A_out_5_port, plus4A_out_4_port, 
      plus4A_out_3_port, plus4A_out_2_port, plus4A_out_1_port, 
      plus4A_out_0_port );
   
   plus2A_out_0_port <= '0';
   plus4A_out_0_port <= '0';
   shifter_1 : shifter_N64_8 port map( input(63) => plusA(63), input(62) => 
                           plusA(62), input(61) => plusA(61), input(60) => 
                           plusA(60), input(59) => plusA(59), input(58) => 
                           plusA(58), input(57) => plusA(57), input(56) => 
                           plusA(56), input(55) => plusA(55), input(54) => 
                           plusA(54), input(53) => plusA(53), input(52) => 
                           plusA(52), input(51) => plusA(51), input(50) => 
                           plusA(50), input(49) => plusA(49), input(48) => 
                           plusA(48), input(47) => plusA(47), input(46) => 
                           plusA(46), input(45) => plusA(45), input(44) => 
                           plusA(44), input(43) => plusA(43), input(42) => 
                           plusA(42), input(41) => plusA(41), input(40) => 
                           plusA(40), input(39) => plusA(39), input(38) => 
                           plusA(38), input(37) => plusA(37), input(36) => 
                           plusA(36), input(35) => plusA(35), input(34) => 
                           plusA(34), input(33) => plusA(33), input(32) => 
                           plusA(32), input(31) => plusA(31), input(30) => 
                           plusA(30), input(29) => plusA(29), input(28) => 
                           plusA(28), input(27) => plusA(27), input(26) => 
                           plusA(26), input(25) => plusA(25), input(24) => 
                           plusA(24), input(23) => plusA(23), input(22) => 
                           plusA(22), input(21) => plusA(21), input(20) => 
                           plusA(20), input(19) => plusA(19), input(18) => 
                           plusA(18), input(17) => plusA(17), input(16) => 
                           plusA(16), input(15) => plusA(15), input(14) => 
                           plusA(14), input(13) => plusA(13), input(12) => 
                           plusA(12), input(11) => plusA(11), input(10) => 
                           plusA(10), input(9) => plusA(9), input(8) => 
                           plusA(8), input(7) => plusA(7), input(6) => plusA(6)
                           , input(5) => plusA(5), input(4) => plusA(4), 
                           input(3) => plusA(3), input(2) => plusA(2), input(1)
                           => plusA(1), input(0) => plusA(0), 
                           shiftLeftOnePos(63) => plus2A_out_63_port, 
                           shiftLeftOnePos(62) => plus2A_out_62_port, 
                           shiftLeftOnePos(61) => plus2A_out_61_port, 
                           shiftLeftOnePos(60) => plus2A_out_60_port, 
                           shiftLeftOnePos(59) => plus2A_out_59_port, 
                           shiftLeftOnePos(58) => plus2A_out_58_port, 
                           shiftLeftOnePos(57) => n2, shiftLeftOnePos(56) => 
                           plus2A_out_56_port, shiftLeftOnePos(55) => 
                           plus2A_out_55_port, shiftLeftOnePos(54) => 
                           plus2A_out_54_port, shiftLeftOnePos(53) => 
                           plus2A_out_53_port, shiftLeftOnePos(52) => 
                           plus2A_out_52_port, shiftLeftOnePos(51) => 
                           plus2A_out_51_port, shiftLeftOnePos(50) => 
                           plus2A_out_50_port, shiftLeftOnePos(49) => 
                           plus2A_out_49_port, shiftLeftOnePos(48) => 
                           plus2A_out_48_port, shiftLeftOnePos(47) => 
                           plus2A_out_47_port, shiftLeftOnePos(46) => 
                           plus2A_out_46_port, shiftLeftOnePos(45) => 
                           plus2A_out_45_port, shiftLeftOnePos(44) => 
                           plus2A_out_44_port, shiftLeftOnePos(43) => 
                           plus2A_out_43_port, shiftLeftOnePos(42) => 
                           plus2A_out_42_port, shiftLeftOnePos(41) => 
                           plus2A_out_41_port, shiftLeftOnePos(40) => 
                           plus2A_out_40_port, shiftLeftOnePos(39) => 
                           plus2A_out_39_port, shiftLeftOnePos(38) => 
                           plus2A_out_38_port, shiftLeftOnePos(37) => 
                           plus2A_out_37_port, shiftLeftOnePos(36) => 
                           plus2A_out_36_port, shiftLeftOnePos(35) => 
                           plus2A_out_35_port, shiftLeftOnePos(34) => 
                           plus2A_out_34_port, shiftLeftOnePos(33) => 
                           plus2A_out_33_port, shiftLeftOnePos(32) => 
                           plus2A_out_32_port, shiftLeftOnePos(31) => 
                           plus2A_out_31_port, shiftLeftOnePos(30) => 
                           plus2A_out_30_port, shiftLeftOnePos(29) => 
                           plus2A_out_29_port, shiftLeftOnePos(28) => 
                           plus2A_out_28_port, shiftLeftOnePos(27) => 
                           plus2A_out_27_port, shiftLeftOnePos(26) => 
                           plus2A_out_26_port, shiftLeftOnePos(25) => 
                           plus2A_out_25_port, shiftLeftOnePos(24) => 
                           plus2A_out_24_port, shiftLeftOnePos(23) => 
                           plus2A_out_23_port, shiftLeftOnePos(22) => 
                           plus2A_out_22_port, shiftLeftOnePos(21) => 
                           plus2A_out_21_port, shiftLeftOnePos(20) => 
                           plus2A_out_20_port, shiftLeftOnePos(19) => 
                           plus2A_out_19_port, shiftLeftOnePos(18) => 
                           plus2A_out_18_port, shiftLeftOnePos(17) => 
                           plus2A_out_17_port, shiftLeftOnePos(16) => 
                           plus2A_out_16_port, shiftLeftOnePos(15) => 
                           plus2A_out_15_port, shiftLeftOnePos(14) => 
                           plus2A_out_14_port, shiftLeftOnePos(13) => 
                           plus2A_out_13_port, shiftLeftOnePos(12) => 
                           plus2A_out_12_port, shiftLeftOnePos(11) => 
                           plus2A_out_11_port, shiftLeftOnePos(10) => 
                           plus2A_out_10_port, shiftLeftOnePos(9) => 
                           plus2A_out_9_port, shiftLeftOnePos(8) => 
                           plus2A_out_8_port, shiftLeftOnePos(7) => 
                           plus2A_out_7_port, shiftLeftOnePos(6) => 
                           plus2A_out_6_port, shiftLeftOnePos(5) => 
                           plus2A_out_5_port, shiftLeftOnePos(4) => 
                           plus2A_out_4_port, shiftLeftOnePos(3) => 
                           plus2A_out_3_port, shiftLeftOnePos(2) => 
                           plus2A_out_2_port, shiftLeftOnePos(1) => 
                           plus2A_out_1_port, shiftLeftOnePos(0) => n_3150);
   shifter_2 : shifter_N64_7 port map( input(63) => plus2A_out_63_port, 
                           input(62) => plus2A_out_62_port, input(61) => 
                           plus2A_out_61_port, input(60) => plus2A_out_60_port,
                           input(59) => plus2A_out_59_port, input(58) => 
                           plus2A_out_58_port, input(57) => plus2A_out_57_port,
                           input(56) => plus2A_out_56_port, input(55) => 
                           plus2A_out_55_port, input(54) => plus2A_out_54_port,
                           input(53) => plus2A_out_53_port, input(52) => 
                           plus2A_out_52_port, input(51) => plus2A_out_51_port,
                           input(50) => plus2A_out_50_port, input(49) => 
                           plus2A_out_49_port, input(48) => plus2A_out_48_port,
                           input(47) => plus2A_out_47_port, input(46) => 
                           plus2A_out_46_port, input(45) => plus2A_out_45_port,
                           input(44) => plus2A_out_44_port, input(43) => 
                           plus2A_out_43_port, input(42) => plus2A_out_42_port,
                           input(41) => plus2A_out_41_port, input(40) => 
                           plus2A_out_40_port, input(39) => plus2A_out_39_port,
                           input(38) => plus2A_out_38_port, input(37) => 
                           plus2A_out_37_port, input(36) => plus2A_out_36_port,
                           input(35) => plus2A_out_35_port, input(34) => 
                           plus2A_out_34_port, input(33) => plus2A_out_33_port,
                           input(32) => plus2A_out_32_port, input(31) => 
                           plus2A_out_31_port, input(30) => plus2A_out_30_port,
                           input(29) => plus2A_out_29_port, input(28) => 
                           plus2A_out_28_port, input(27) => plus2A_out_27_port,
                           input(26) => plus2A_out_26_port, input(25) => 
                           plus2A_out_25_port, input(24) => plus2A_out_24_port,
                           input(23) => plus2A_out_23_port, input(22) => 
                           plus2A_out_22_port, input(21) => plus2A_out_21_port,
                           input(20) => plus2A_out_20_port, input(19) => 
                           plus2A_out_19_port, input(18) => plus2A_out_18_port,
                           input(17) => plus2A_out_17_port, input(16) => 
                           plus2A_out_16_port, input(15) => plus2A_out_15_port,
                           input(14) => plus2A_out_14_port, input(13) => 
                           plus2A_out_13_port, input(12) => plus2A_out_12_port,
                           input(11) => plus2A_out_11_port, input(10) => 
                           plus2A_out_10_port, input(9) => plus2A_out_9_port, 
                           input(8) => plus2A_out_8_port, input(7) => 
                           plus2A_out_7_port, input(6) => plus2A_out_6_port, 
                           input(5) => plus2A_out_5_port, input(4) => 
                           plus2A_out_4_port, input(3) => plus2A_out_3_port, 
                           input(2) => plus2A_out_2_port, input(1) => 
                           plus2A_out_1_port, input(0) => plus2A_out_0_port, 
                           shiftLeftOnePos(63) => plus4A_out_63_port, 
                           shiftLeftOnePos(62) => plus4A_out_62_port, 
                           shiftLeftOnePos(61) => plus4A_out_61_port, 
                           shiftLeftOnePos(60) => plus4A_out_60_port, 
                           shiftLeftOnePos(59) => plus4A_out_59_port, 
                           shiftLeftOnePos(58) => plus4A_out_58_port, 
                           shiftLeftOnePos(57) => plus4A_out_57_port, 
                           shiftLeftOnePos(56) => plus4A_out_56_port, 
                           shiftLeftOnePos(55) => plus4A_out_55_port, 
                           shiftLeftOnePos(54) => plus4A_out_54_port, 
                           shiftLeftOnePos(53) => plus4A_out_53_port, 
                           shiftLeftOnePos(52) => plus4A_out_52_port, 
                           shiftLeftOnePos(51) => plus4A_out_51_port, 
                           shiftLeftOnePos(50) => plus4A_out_50_port, 
                           shiftLeftOnePos(49) => plus4A_out_49_port, 
                           shiftLeftOnePos(48) => plus4A_out_48_port, 
                           shiftLeftOnePos(47) => plus4A_out_47_port, 
                           shiftLeftOnePos(46) => plus4A_out_46_port, 
                           shiftLeftOnePos(45) => plus4A_out_45_port, 
                           shiftLeftOnePos(44) => plus4A_out_44_port, 
                           shiftLeftOnePos(43) => plus4A_out_43_port, 
                           shiftLeftOnePos(42) => plus4A_out_42_port, 
                           shiftLeftOnePos(41) => plus4A_out_41_port, 
                           shiftLeftOnePos(40) => plus4A_out_40_port, 
                           shiftLeftOnePos(39) => plus4A_out_39_port, 
                           shiftLeftOnePos(38) => plus4A_out_38_port, 
                           shiftLeftOnePos(37) => plus4A_out_37_port, 
                           shiftLeftOnePos(36) => plus4A_out_36_port, 
                           shiftLeftOnePos(35) => plus4A_out_35_port, 
                           shiftLeftOnePos(34) => plus4A_out_34_port, 
                           shiftLeftOnePos(33) => plus4A_out_33_port, 
                           shiftLeftOnePos(32) => plus4A_out_32_port, 
                           shiftLeftOnePos(31) => plus4A_out_31_port, 
                           shiftLeftOnePos(30) => plus4A_out_30_port, 
                           shiftLeftOnePos(29) => plus4A_out_29_port, 
                           shiftLeftOnePos(28) => plus4A_out_28_port, 
                           shiftLeftOnePos(27) => plus4A_out_27_port, 
                           shiftLeftOnePos(26) => plus4A_out_26_port, 
                           shiftLeftOnePos(25) => plus4A_out_25_port, 
                           shiftLeftOnePos(24) => plus4A_out_24_port, 
                           shiftLeftOnePos(23) => plus4A_out_23_port, 
                           shiftLeftOnePos(22) => plus4A_out_22_port, 
                           shiftLeftOnePos(21) => plus4A_out_21_port, 
                           shiftLeftOnePos(20) => plus4A_out_20_port, 
                           shiftLeftOnePos(19) => plus4A_out_19_port, 
                           shiftLeftOnePos(18) => plus4A_out_18_port, 
                           shiftLeftOnePos(17) => plus4A_out_17_port, 
                           shiftLeftOnePos(16) => plus4A_out_16_port, 
                           shiftLeftOnePos(15) => plus4A_out_15_port, 
                           shiftLeftOnePos(14) => plus4A_out_14_port, 
                           shiftLeftOnePos(13) => plus4A_out_13_port, 
                           shiftLeftOnePos(12) => plus4A_out_12_port, 
                           shiftLeftOnePos(11) => plus4A_out_11_port, 
                           shiftLeftOnePos(10) => plus4A_out_10_port, 
                           shiftLeftOnePos(9) => plus4A_out_9_port, 
                           shiftLeftOnePos(8) => plus4A_out_8_port, 
                           shiftLeftOnePos(7) => plus4A_out_7_port, 
                           shiftLeftOnePos(6) => plus4A_out_6_port, 
                           shiftLeftOnePos(5) => plus4A_out_5_port, 
                           shiftLeftOnePos(4) => plus4A_out_4_port, 
                           shiftLeftOnePos(3) => plus4A_out_3_port, 
                           shiftLeftOnePos(2) => plus4A_out_2_port, 
                           shiftLeftOnePos(1) => plus4A_out_1_port, 
                           shiftLeftOnePos(0) => n_3151);
   complementer_1 : complementer_N64_8 port map( input(63) => 
                           plus2A_out_63_port, input(62) => plus2A_out_62_port,
                           input(61) => plus2A_out_61_port, input(60) => 
                           plus2A_out_60_port, input(59) => plus2A_out_59_port,
                           input(58) => plus2A_out_58_port, input(57) => 
                           plus2A_out_57_port, input(56) => plus2A_out_56_port,
                           input(55) => plus2A_out_55_port, input(54) => 
                           plus2A_out_54_port, input(53) => plus2A_out_53_port,
                           input(52) => plus2A_out_52_port, input(51) => 
                           plus2A_out_51_port, input(50) => plus2A_out_50_port,
                           input(49) => plus2A_out_49_port, input(48) => 
                           plus2A_out_48_port, input(47) => plus2A_out_47_port,
                           input(46) => plus2A_out_46_port, input(45) => 
                           plus2A_out_45_port, input(44) => plus2A_out_44_port,
                           input(43) => plus2A_out_43_port, input(42) => 
                           plus2A_out_42_port, input(41) => plus2A_out_41_port,
                           input(40) => plus2A_out_40_port, input(39) => 
                           plus2A_out_39_port, input(38) => plus2A_out_38_port,
                           input(37) => plus2A_out_37_port, input(36) => 
                           plus2A_out_36_port, input(35) => plus2A_out_35_port,
                           input(34) => plus2A_out_34_port, input(33) => 
                           plus2A_out_33_port, input(32) => plus2A_out_32_port,
                           input(31) => plus2A_out_31_port, input(30) => 
                           plus2A_out_30_port, input(29) => plus2A_out_29_port,
                           input(28) => plus2A_out_28_port, input(27) => 
                           plus2A_out_27_port, input(26) => plus2A_out_26_port,
                           input(25) => plus2A_out_25_port, input(24) => 
                           plus2A_out_24_port, input(23) => plus2A_out_23_port,
                           input(22) => plus2A_out_22_port, input(21) => 
                           plus2A_out_21_port, input(20) => plus2A_out_20_port,
                           input(19) => plus2A_out_19_port, input(18) => 
                           plus2A_out_18_port, input(17) => plus2A_out_17_port,
                           input(16) => plus2A_out_16_port, input(15) => 
                           plus2A_out_15_port, input(14) => plus2A_out_14_port,
                           input(13) => plus2A_out_13_port, input(12) => 
                           plus2A_out_12_port, input(11) => plus2A_out_11_port,
                           input(10) => plus2A_out_10_port, input(9) => 
                           plus2A_out_9_port, input(8) => plus2A_out_8_port, 
                           input(7) => plus2A_out_7_port, input(6) => 
                           plus2A_out_6_port, input(5) => plus2A_out_5_port, 
                           input(4) => plus2A_out_4_port, input(3) => 
                           plus2A_out_3_port, input(2) => plus2A_out_2_port, 
                           input(1) => plus2A_out_1_port, input(0) => 
                           plus2A_out_0_port, complement2(63) => 
                           minus2A_out(63), complement2(62) => minus2A_out(62),
                           complement2(61) => minus2A_out(61), complement2(60) 
                           => minus2A_out(60), complement2(59) => 
                           minus2A_out(59), complement2(58) => minus2A_out(58),
                           complement2(57) => minus2A_out(57), complement2(56) 
                           => minus2A_out(56), complement2(55) => 
                           minus2A_out(55), complement2(54) => minus2A_out(54),
                           complement2(53) => minus2A_out(53), complement2(52) 
                           => minus2A_out(52), complement2(51) => 
                           minus2A_out(51), complement2(50) => minus2A_out(50),
                           complement2(49) => minus2A_out(49), complement2(48) 
                           => minus2A_out(48), complement2(47) => 
                           minus2A_out(47), complement2(46) => minus2A_out(46),
                           complement2(45) => minus2A_out(45), complement2(44) 
                           => minus2A_out(44), complement2(43) => 
                           minus2A_out(43), complement2(42) => minus2A_out(42),
                           complement2(41) => minus2A_out(41), complement2(40) 
                           => minus2A_out(40), complement2(39) => 
                           minus2A_out(39), complement2(38) => minus2A_out(38),
                           complement2(37) => minus2A_out(37), complement2(36) 
                           => minus2A_out(36), complement2(35) => 
                           minus2A_out(35), complement2(34) => minus2A_out(34),
                           complement2(33) => minus2A_out(33), complement2(32) 
                           => minus2A_out(32), complement2(31) => 
                           minus2A_out(31), complement2(30) => minus2A_out(30),
                           complement2(29) => minus2A_out(29), complement2(28) 
                           => minus2A_out(28), complement2(27) => 
                           minus2A_out(27), complement2(26) => minus2A_out(26),
                           complement2(25) => minus2A_out(25), complement2(24) 
                           => minus2A_out(24), complement2(23) => 
                           minus2A_out(23), complement2(22) => minus2A_out(22),
                           complement2(21) => minus2A_out(21), complement2(20) 
                           => minus2A_out(20), complement2(19) => 
                           minus2A_out(19), complement2(18) => minus2A_out(18),
                           complement2(17) => minus2A_out(17), complement2(16) 
                           => minus2A_out(16), complement2(15) => 
                           minus2A_out(15), complement2(14) => minus2A_out(14),
                           complement2(13) => minus2A_out(13), complement2(12) 
                           => minus2A_out(12), complement2(11) => 
                           minus2A_out(11), complement2(10) => minus2A_out(10),
                           complement2(9) => minus2A_out(9), complement2(8) => 
                           minus2A_out(8), complement2(7) => minus2A_out(7), 
                           complement2(6) => minus2A_out(6), complement2(5) => 
                           minus2A_out(5), complement2(4) => minus2A_out(4), 
                           complement2(3) => minus2A_out(3), complement2(2) => 
                           minus2A_out(2), complement2(1) => minus2A_out(1), 
                           complement2(0) => minus2A_out(0));
   complementer_2 : complementer_N64_7 port map( input(63) => 
                           plus4A_out_63_port, input(62) => plus4A_out_62_port,
                           input(61) => plus4A_out_61_port, input(60) => 
                           plus4A_out_60_port, input(59) => plus4A_out_59_port,
                           input(58) => plus4A_out_58_port, input(57) => 
                           plus4A_out_57_port, input(56) => plus4A_out_56_port,
                           input(55) => plus4A_out_55_port, input(54) => 
                           plus4A_out_54_port, input(53) => plus4A_out_53_port,
                           input(52) => plus4A_out_52_port, input(51) => 
                           plus4A_out_51_port, input(50) => plus4A_out_50_port,
                           input(49) => plus4A_out_49_port, input(48) => 
                           plus4A_out_48_port, input(47) => plus4A_out_47_port,
                           input(46) => plus4A_out_46_port, input(45) => 
                           plus4A_out_45_port, input(44) => plus4A_out_44_port,
                           input(43) => plus4A_out_43_port, input(42) => 
                           plus4A_out_42_port, input(41) => plus4A_out_41_port,
                           input(40) => plus4A_out_40_port, input(39) => 
                           plus4A_out_39_port, input(38) => plus4A_out_38_port,
                           input(37) => plus4A_out_37_port, input(36) => 
                           plus4A_out_36_port, input(35) => plus4A_out_35_port,
                           input(34) => plus4A_out_34_port, input(33) => 
                           plus4A_out_33_port, input(32) => plus4A_out_32_port,
                           input(31) => plus4A_out_31_port, input(30) => 
                           plus4A_out_30_port, input(29) => plus4A_out_29_port,
                           input(28) => plus4A_out_28_port, input(27) => 
                           plus4A_out_27_port, input(26) => plus4A_out_26_port,
                           input(25) => plus4A_out_25_port, input(24) => 
                           plus4A_out_24_port, input(23) => plus4A_out_23_port,
                           input(22) => plus4A_out_22_port, input(21) => 
                           plus4A_out_21_port, input(20) => plus4A_out_20_port,
                           input(19) => plus4A_out_19_port, input(18) => 
                           plus4A_out_18_port, input(17) => plus4A_out_17_port,
                           input(16) => plus4A_out_16_port, input(15) => 
                           plus4A_out_15_port, input(14) => plus4A_out_14_port,
                           input(13) => plus4A_out_13_port, input(12) => 
                           plus4A_out_12_port, input(11) => plus4A_out_11_port,
                           input(10) => plus4A_out_10_port, input(9) => 
                           plus4A_out_9_port, input(8) => plus4A_out_8_port, 
                           input(7) => plus4A_out_7_port, input(6) => 
                           plus4A_out_6_port, input(5) => plus4A_out_5_port, 
                           input(4) => plus4A_out_4_port, input(3) => 
                           plus4A_out_3_port, input(2) => plus4A_out_2_port, 
                           input(1) => plus4A_out_1_port, input(0) => 
                           plus4A_out_0_port, complement2(63) => 
                           minus4A_out(63), complement2(62) => minus4A_out(62),
                           complement2(61) => minus4A_out(61), complement2(60) 
                           => minus4A_out(60), complement2(59) => 
                           minus4A_out(59), complement2(58) => minus4A_out(58),
                           complement2(57) => minus4A_out(57), complement2(56) 
                           => minus4A_out(56), complement2(55) => 
                           minus4A_out(55), complement2(54) => minus4A_out(54),
                           complement2(53) => minus4A_out(53), complement2(52) 
                           => minus4A_out(52), complement2(51) => 
                           minus4A_out(51), complement2(50) => minus4A_out(50),
                           complement2(49) => minus4A_out(49), complement2(48) 
                           => minus4A_out(48), complement2(47) => 
                           minus4A_out(47), complement2(46) => minus4A_out(46),
                           complement2(45) => minus4A_out(45), complement2(44) 
                           => minus4A_out(44), complement2(43) => 
                           minus4A_out(43), complement2(42) => minus4A_out(42),
                           complement2(41) => minus4A_out(41), complement2(40) 
                           => minus4A_out(40), complement2(39) => 
                           minus4A_out(39), complement2(38) => minus4A_out(38),
                           complement2(37) => minus4A_out(37), complement2(36) 
                           => minus4A_out(36), complement2(35) => 
                           minus4A_out(35), complement2(34) => minus4A_out(34),
                           complement2(33) => minus4A_out(33), complement2(32) 
                           => minus4A_out(32), complement2(31) => 
                           minus4A_out(31), complement2(30) => minus4A_out(30),
                           complement2(29) => minus4A_out(29), complement2(28) 
                           => minus4A_out(28), complement2(27) => 
                           minus4A_out(27), complement2(26) => minus4A_out(26),
                           complement2(25) => minus4A_out(25), complement2(24) 
                           => minus4A_out(24), complement2(23) => 
                           minus4A_out(23), complement2(22) => minus4A_out(22),
                           complement2(21) => minus4A_out(21), complement2(20) 
                           => minus4A_out(20), complement2(19) => 
                           minus4A_out(19), complement2(18) => minus4A_out(18),
                           complement2(17) => minus4A_out(17), complement2(16) 
                           => minus4A_out(16), complement2(15) => 
                           minus4A_out(15), complement2(14) => minus4A_out(14),
                           complement2(13) => minus4A_out(13), complement2(12) 
                           => minus4A_out(12), complement2(11) => 
                           minus4A_out(11), complement2(10) => minus4A_out(10),
                           complement2(9) => minus4A_out(9), complement2(8) => 
                           minus4A_out(8), complement2(7) => minus4A_out(7), 
                           complement2(6) => minus4A_out(6), complement2(5) => 
                           minus4A_out(5), complement2(4) => minus4A_out(4), 
                           complement2(3) => minus4A_out(3), complement2(2) => 
                           minus4A_out(2), complement2(1) => minus4A_out(1), 
                           complement2(0) => minus4A_out(0));
   U3 : BUF_X1 port map( A => n2, Z => plus2A_out_57_port);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity ShiftnCompl_N64_5 is

   port( plusA : in std_logic_vector (63 downto 0);  plus2A_out, minus2A_out, 
         plus4A_out, minus4A_out : out std_logic_vector (63 downto 0));

end ShiftnCompl_N64_5;

architecture SYN_struct of ShiftnCompl_N64_5 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component complementer_N64_9
      port( input : in std_logic_vector (63 downto 0);  complement2 : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component complementer_N64_10
      port( input : in std_logic_vector (63 downto 0);  complement2 : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component shifter_N64_9
      port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component shifter_N64_10
      port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
            std_logic_vector (63 downto 0));
   end component;
   
   signal plus2A_out_63_port, plus2A_out_62_port, plus2A_out_61_port, 
      plus2A_out_60_port, plus2A_out_59_port, plus2A_out_58_port, n32, 
      plus2A_out_56_port, plus2A_out_55_port, plus2A_out_54_port, 
      plus2A_out_53_port, plus2A_out_52_port, n33, n34, n35, n36, n37, n38, n39
      , n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, 
      n54, n55, n56, n57, n58, n59, n60, n61, n62, plus2A_out_21_port, 
      plus2A_out_20_port, plus2A_out_19_port, plus2A_out_18_port, 
      plus2A_out_17_port, plus2A_out_16_port, plus2A_out_15_port, 
      plus2A_out_14_port, plus2A_out_13_port, plus2A_out_12_port, 
      plus2A_out_11_port, plus2A_out_10_port, plus2A_out_9_port, 
      plus2A_out_8_port, plus2A_out_7_port, plus2A_out_6_port, 
      plus2A_out_5_port, plus2A_out_4_port, plus2A_out_3_port, 
      plus2A_out_2_port, plus2A_out_1_port, plus2A_out_0_port, 
      plus4A_out_63_port, plus4A_out_62_port, plus4A_out_61_port, 
      plus4A_out_60_port, plus4A_out_59_port, plus4A_out_58_port, 
      plus4A_out_57_port, plus4A_out_56_port, plus4A_out_55_port, 
      plus4A_out_54_port, plus4A_out_53_port, plus4A_out_52_port, 
      plus4A_out_51_port, plus4A_out_50_port, plus4A_out_49_port, 
      plus4A_out_48_port, plus4A_out_47_port, plus4A_out_46_port, 
      plus4A_out_45_port, plus4A_out_44_port, plus4A_out_43_port, 
      plus4A_out_42_port, plus4A_out_41_port, plus4A_out_40_port, 
      plus4A_out_39_port, plus4A_out_38_port, plus4A_out_37_port, 
      plus4A_out_36_port, plus4A_out_35_port, plus4A_out_34_port, 
      plus4A_out_33_port, plus4A_out_32_port, plus4A_out_31_port, 
      plus4A_out_30_port, plus4A_out_29_port, plus4A_out_28_port, 
      plus4A_out_27_port, plus4A_out_26_port, plus4A_out_25_port, 
      plus4A_out_24_port, plus4A_out_23_port, plus4A_out_22_port, 
      plus4A_out_21_port, plus4A_out_20_port, plus4A_out_19_port, 
      plus4A_out_18_port, plus4A_out_17_port, plus4A_out_16_port, 
      plus4A_out_15_port, plus4A_out_14_port, plus4A_out_13_port, 
      plus4A_out_12_port, plus4A_out_11_port, plus4A_out_10_port, 
      plus4A_out_9_port, plus4A_out_8_port, plus4A_out_7_port, 
      plus4A_out_6_port, plus4A_out_5_port, plus4A_out_4_port, 
      plus4A_out_3_port, plus4A_out_2_port, plus4A_out_1_port, 
      plus4A_out_0_port, plus2A_out_22_port, plus2A_out_23_port, 
      plus2A_out_24_port, plus2A_out_25_port, plus2A_out_26_port, 
      plus2A_out_27_port, plus2A_out_28_port, plus2A_out_29_port, 
      plus2A_out_30_port, plus2A_out_31_port, plus2A_out_32_port, 
      plus2A_out_33_port, plus2A_out_34_port, plus2A_out_35_port, 
      plus2A_out_36_port, plus2A_out_37_port, plus2A_out_38_port, 
      plus2A_out_39_port, plus2A_out_40_port, plus2A_out_41_port, 
      plus2A_out_42_port, plus2A_out_43_port, plus2A_out_44_port, 
      plus2A_out_45_port, plus2A_out_46_port, plus2A_out_47_port, 
      plus2A_out_48_port, plus2A_out_49_port, plus2A_out_50_port, 
      plus2A_out_51_port, plus2A_out_57_port, n_3152, n_3153 : std_logic;

begin
   plus2A_out <= ( plus2A_out_63_port, plus2A_out_62_port, plus2A_out_61_port, 
      plus2A_out_60_port, plus2A_out_59_port, plus2A_out_58_port, 
      plus2A_out_57_port, plus2A_out_56_port, plus2A_out_55_port, 
      plus2A_out_54_port, plus2A_out_53_port, plus2A_out_52_port, 
      plus2A_out_51_port, plus2A_out_50_port, plus2A_out_49_port, 
      plus2A_out_48_port, plus2A_out_47_port, plus2A_out_46_port, 
      plus2A_out_45_port, plus2A_out_44_port, plus2A_out_43_port, 
      plus2A_out_42_port, plus2A_out_41_port, plus2A_out_40_port, 
      plus2A_out_39_port, plus2A_out_38_port, plus2A_out_37_port, 
      plus2A_out_36_port, plus2A_out_35_port, plus2A_out_34_port, 
      plus2A_out_33_port, plus2A_out_32_port, plus2A_out_31_port, 
      plus2A_out_30_port, plus2A_out_29_port, plus2A_out_28_port, 
      plus2A_out_27_port, plus2A_out_26_port, plus2A_out_25_port, 
      plus2A_out_24_port, plus2A_out_23_port, plus2A_out_22_port, 
      plus2A_out_21_port, plus2A_out_20_port, plus2A_out_19_port, 
      plus2A_out_18_port, plus2A_out_17_port, plus2A_out_16_port, 
      plus2A_out_15_port, plus2A_out_14_port, plus2A_out_13_port, 
      plus2A_out_12_port, plus2A_out_11_port, plus2A_out_10_port, 
      plus2A_out_9_port, plus2A_out_8_port, plus2A_out_7_port, 
      plus2A_out_6_port, plus2A_out_5_port, plus2A_out_4_port, 
      plus2A_out_3_port, plus2A_out_2_port, plus2A_out_1_port, 
      plus2A_out_0_port );
   plus4A_out <= ( plus4A_out_63_port, plus4A_out_62_port, plus4A_out_61_port, 
      plus4A_out_60_port, plus4A_out_59_port, plus4A_out_58_port, 
      plus4A_out_57_port, plus4A_out_56_port, plus4A_out_55_port, 
      plus4A_out_54_port, plus4A_out_53_port, plus4A_out_52_port, 
      plus4A_out_51_port, plus4A_out_50_port, plus4A_out_49_port, 
      plus4A_out_48_port, plus4A_out_47_port, plus4A_out_46_port, 
      plus4A_out_45_port, plus4A_out_44_port, plus4A_out_43_port, 
      plus4A_out_42_port, plus4A_out_41_port, plus4A_out_40_port, 
      plus4A_out_39_port, plus4A_out_38_port, plus4A_out_37_port, 
      plus4A_out_36_port, plus4A_out_35_port, plus4A_out_34_port, 
      plus4A_out_33_port, plus4A_out_32_port, plus4A_out_31_port, 
      plus4A_out_30_port, plus4A_out_29_port, plus4A_out_28_port, 
      plus4A_out_27_port, plus4A_out_26_port, plus4A_out_25_port, 
      plus4A_out_24_port, plus4A_out_23_port, plus4A_out_22_port, 
      plus4A_out_21_port, plus4A_out_20_port, plus4A_out_19_port, 
      plus4A_out_18_port, plus4A_out_17_port, plus4A_out_16_port, 
      plus4A_out_15_port, plus4A_out_14_port, plus4A_out_13_port, 
      plus4A_out_12_port, plus4A_out_11_port, plus4A_out_10_port, 
      plus4A_out_9_port, plus4A_out_8_port, plus4A_out_7_port, 
      plus4A_out_6_port, plus4A_out_5_port, plus4A_out_4_port, 
      plus4A_out_3_port, plus4A_out_2_port, plus4A_out_1_port, 
      plus4A_out_0_port );
   
   plus2A_out_0_port <= '0';
   plus4A_out_0_port <= '0';
   shifter_1 : shifter_N64_10 port map( input(63) => plusA(63), input(62) => 
                           plusA(62), input(61) => plusA(61), input(60) => 
                           plusA(60), input(59) => plusA(59), input(58) => 
                           plusA(58), input(57) => plusA(57), input(56) => 
                           plusA(56), input(55) => plusA(55), input(54) => 
                           plusA(54), input(53) => plusA(53), input(52) => 
                           plusA(52), input(51) => plusA(51), input(50) => 
                           plusA(50), input(49) => plusA(49), input(48) => 
                           plusA(48), input(47) => plusA(47), input(46) => 
                           plusA(46), input(45) => plusA(45), input(44) => 
                           plusA(44), input(43) => plusA(43), input(42) => 
                           plusA(42), input(41) => plusA(41), input(40) => 
                           plusA(40), input(39) => plusA(39), input(38) => 
                           plusA(38), input(37) => plusA(37), input(36) => 
                           plusA(36), input(35) => plusA(35), input(34) => 
                           plusA(34), input(33) => plusA(33), input(32) => 
                           plusA(32), input(31) => plusA(31), input(30) => 
                           plusA(30), input(29) => plusA(29), input(28) => 
                           plusA(28), input(27) => plusA(27), input(26) => 
                           plusA(26), input(25) => plusA(25), input(24) => 
                           plusA(24), input(23) => plusA(23), input(22) => 
                           plusA(22), input(21) => plusA(21), input(20) => 
                           plusA(20), input(19) => plusA(19), input(18) => 
                           plusA(18), input(17) => plusA(17), input(16) => 
                           plusA(16), input(15) => plusA(15), input(14) => 
                           plusA(14), input(13) => plusA(13), input(12) => 
                           plusA(12), input(11) => plusA(11), input(10) => 
                           plusA(10), input(9) => plusA(9), input(8) => 
                           plusA(8), input(7) => plusA(7), input(6) => plusA(6)
                           , input(5) => plusA(5), input(4) => plusA(4), 
                           input(3) => plusA(3), input(2) => plusA(2), input(1)
                           => plusA(1), input(0) => plusA(0), 
                           shiftLeftOnePos(63) => plus2A_out_63_port, 
                           shiftLeftOnePos(62) => plus2A_out_62_port, 
                           shiftLeftOnePos(61) => plus2A_out_61_port, 
                           shiftLeftOnePos(60) => plus2A_out_60_port, 
                           shiftLeftOnePos(59) => plus2A_out_59_port, 
                           shiftLeftOnePos(58) => plus2A_out_58_port, 
                           shiftLeftOnePos(57) => n32, shiftLeftOnePos(56) => 
                           plus2A_out_56_port, shiftLeftOnePos(55) => 
                           plus2A_out_55_port, shiftLeftOnePos(54) => 
                           plus2A_out_54_port, shiftLeftOnePos(53) => 
                           plus2A_out_53_port, shiftLeftOnePos(52) => 
                           plus2A_out_52_port, shiftLeftOnePos(51) => n33, 
                           shiftLeftOnePos(50) => n34, shiftLeftOnePos(49) => 
                           n35, shiftLeftOnePos(48) => n36, shiftLeftOnePos(47)
                           => n37, shiftLeftOnePos(46) => n38, 
                           shiftLeftOnePos(45) => n39, shiftLeftOnePos(44) => 
                           n40, shiftLeftOnePos(43) => n41, shiftLeftOnePos(42)
                           => n42, shiftLeftOnePos(41) => n43, 
                           shiftLeftOnePos(40) => n44, shiftLeftOnePos(39) => 
                           n45, shiftLeftOnePos(38) => n46, shiftLeftOnePos(37)
                           => n47, shiftLeftOnePos(36) => n48, 
                           shiftLeftOnePos(35) => n49, shiftLeftOnePos(34) => 
                           n50, shiftLeftOnePos(33) => n51, shiftLeftOnePos(32)
                           => n52, shiftLeftOnePos(31) => n53, 
                           shiftLeftOnePos(30) => n54, shiftLeftOnePos(29) => 
                           n55, shiftLeftOnePos(28) => n56, shiftLeftOnePos(27)
                           => n57, shiftLeftOnePos(26) => n58, 
                           shiftLeftOnePos(25) => n59, shiftLeftOnePos(24) => 
                           n60, shiftLeftOnePos(23) => n61, shiftLeftOnePos(22)
                           => n62, shiftLeftOnePos(21) => plus2A_out_21_port, 
                           shiftLeftOnePos(20) => plus2A_out_20_port, 
                           shiftLeftOnePos(19) => plus2A_out_19_port, 
                           shiftLeftOnePos(18) => plus2A_out_18_port, 
                           shiftLeftOnePos(17) => plus2A_out_17_port, 
                           shiftLeftOnePos(16) => plus2A_out_16_port, 
                           shiftLeftOnePos(15) => plus2A_out_15_port, 
                           shiftLeftOnePos(14) => plus2A_out_14_port, 
                           shiftLeftOnePos(13) => plus2A_out_13_port, 
                           shiftLeftOnePos(12) => plus2A_out_12_port, 
                           shiftLeftOnePos(11) => plus2A_out_11_port, 
                           shiftLeftOnePos(10) => plus2A_out_10_port, 
                           shiftLeftOnePos(9) => plus2A_out_9_port, 
                           shiftLeftOnePos(8) => plus2A_out_8_port, 
                           shiftLeftOnePos(7) => plus2A_out_7_port, 
                           shiftLeftOnePos(6) => plus2A_out_6_port, 
                           shiftLeftOnePos(5) => plus2A_out_5_port, 
                           shiftLeftOnePos(4) => plus2A_out_4_port, 
                           shiftLeftOnePos(3) => plus2A_out_3_port, 
                           shiftLeftOnePos(2) => plus2A_out_2_port, 
                           shiftLeftOnePos(1) => plus2A_out_1_port, 
                           shiftLeftOnePos(0) => n_3152);
   shifter_2 : shifter_N64_9 port map( input(63) => plus2A_out_63_port, 
                           input(62) => plus2A_out_62_port, input(61) => 
                           plus2A_out_61_port, input(60) => plus2A_out_60_port,
                           input(59) => plus2A_out_59_port, input(58) => 
                           plus2A_out_58_port, input(57) => plus2A_out_57_port,
                           input(56) => plus2A_out_56_port, input(55) => 
                           plus2A_out_55_port, input(54) => plus2A_out_54_port,
                           input(53) => plus2A_out_53_port, input(52) => 
                           plus2A_out_52_port, input(51) => plus2A_out_51_port,
                           input(50) => plus2A_out_50_port, input(49) => 
                           plus2A_out_49_port, input(48) => plus2A_out_48_port,
                           input(47) => plus2A_out_47_port, input(46) => 
                           plus2A_out_46_port, input(45) => plus2A_out_45_port,
                           input(44) => plus2A_out_44_port, input(43) => 
                           plus2A_out_43_port, input(42) => plus2A_out_42_port,
                           input(41) => plus2A_out_41_port, input(40) => 
                           plus2A_out_40_port, input(39) => plus2A_out_39_port,
                           input(38) => plus2A_out_38_port, input(37) => 
                           plus2A_out_37_port, input(36) => plus2A_out_36_port,
                           input(35) => plus2A_out_35_port, input(34) => 
                           plus2A_out_34_port, input(33) => plus2A_out_33_port,
                           input(32) => plus2A_out_32_port, input(31) => 
                           plus2A_out_31_port, input(30) => plus2A_out_30_port,
                           input(29) => plus2A_out_29_port, input(28) => 
                           plus2A_out_28_port, input(27) => plus2A_out_27_port,
                           input(26) => plus2A_out_26_port, input(25) => 
                           plus2A_out_25_port, input(24) => plus2A_out_24_port,
                           input(23) => plus2A_out_23_port, input(22) => 
                           plus2A_out_22_port, input(21) => plus2A_out_21_port,
                           input(20) => plus2A_out_20_port, input(19) => 
                           plus2A_out_19_port, input(18) => plus2A_out_18_port,
                           input(17) => plus2A_out_17_port, input(16) => 
                           plus2A_out_16_port, input(15) => plus2A_out_15_port,
                           input(14) => plus2A_out_14_port, input(13) => 
                           plus2A_out_13_port, input(12) => plus2A_out_12_port,
                           input(11) => plus2A_out_11_port, input(10) => 
                           plus2A_out_10_port, input(9) => plus2A_out_9_port, 
                           input(8) => plus2A_out_8_port, input(7) => 
                           plus2A_out_7_port, input(6) => plus2A_out_6_port, 
                           input(5) => plus2A_out_5_port, input(4) => 
                           plus2A_out_4_port, input(3) => plus2A_out_3_port, 
                           input(2) => plus2A_out_2_port, input(1) => 
                           plus2A_out_1_port, input(0) => plus2A_out_0_port, 
                           shiftLeftOnePos(63) => plus4A_out_63_port, 
                           shiftLeftOnePos(62) => plus4A_out_62_port, 
                           shiftLeftOnePos(61) => plus4A_out_61_port, 
                           shiftLeftOnePos(60) => plus4A_out_60_port, 
                           shiftLeftOnePos(59) => plus4A_out_59_port, 
                           shiftLeftOnePos(58) => plus4A_out_58_port, 
                           shiftLeftOnePos(57) => plus4A_out_57_port, 
                           shiftLeftOnePos(56) => plus4A_out_56_port, 
                           shiftLeftOnePos(55) => plus4A_out_55_port, 
                           shiftLeftOnePos(54) => plus4A_out_54_port, 
                           shiftLeftOnePos(53) => plus4A_out_53_port, 
                           shiftLeftOnePos(52) => plus4A_out_52_port, 
                           shiftLeftOnePos(51) => plus4A_out_51_port, 
                           shiftLeftOnePos(50) => plus4A_out_50_port, 
                           shiftLeftOnePos(49) => plus4A_out_49_port, 
                           shiftLeftOnePos(48) => plus4A_out_48_port, 
                           shiftLeftOnePos(47) => plus4A_out_47_port, 
                           shiftLeftOnePos(46) => plus4A_out_46_port, 
                           shiftLeftOnePos(45) => plus4A_out_45_port, 
                           shiftLeftOnePos(44) => plus4A_out_44_port, 
                           shiftLeftOnePos(43) => plus4A_out_43_port, 
                           shiftLeftOnePos(42) => plus4A_out_42_port, 
                           shiftLeftOnePos(41) => plus4A_out_41_port, 
                           shiftLeftOnePos(40) => plus4A_out_40_port, 
                           shiftLeftOnePos(39) => plus4A_out_39_port, 
                           shiftLeftOnePos(38) => plus4A_out_38_port, 
                           shiftLeftOnePos(37) => plus4A_out_37_port, 
                           shiftLeftOnePos(36) => plus4A_out_36_port, 
                           shiftLeftOnePos(35) => plus4A_out_35_port, 
                           shiftLeftOnePos(34) => plus4A_out_34_port, 
                           shiftLeftOnePos(33) => plus4A_out_33_port, 
                           shiftLeftOnePos(32) => plus4A_out_32_port, 
                           shiftLeftOnePos(31) => plus4A_out_31_port, 
                           shiftLeftOnePos(30) => plus4A_out_30_port, 
                           shiftLeftOnePos(29) => plus4A_out_29_port, 
                           shiftLeftOnePos(28) => plus4A_out_28_port, 
                           shiftLeftOnePos(27) => plus4A_out_27_port, 
                           shiftLeftOnePos(26) => plus4A_out_26_port, 
                           shiftLeftOnePos(25) => plus4A_out_25_port, 
                           shiftLeftOnePos(24) => plus4A_out_24_port, 
                           shiftLeftOnePos(23) => plus4A_out_23_port, 
                           shiftLeftOnePos(22) => plus4A_out_22_port, 
                           shiftLeftOnePos(21) => plus4A_out_21_port, 
                           shiftLeftOnePos(20) => plus4A_out_20_port, 
                           shiftLeftOnePos(19) => plus4A_out_19_port, 
                           shiftLeftOnePos(18) => plus4A_out_18_port, 
                           shiftLeftOnePos(17) => plus4A_out_17_port, 
                           shiftLeftOnePos(16) => plus4A_out_16_port, 
                           shiftLeftOnePos(15) => plus4A_out_15_port, 
                           shiftLeftOnePos(14) => plus4A_out_14_port, 
                           shiftLeftOnePos(13) => plus4A_out_13_port, 
                           shiftLeftOnePos(12) => plus4A_out_12_port, 
                           shiftLeftOnePos(11) => plus4A_out_11_port, 
                           shiftLeftOnePos(10) => plus4A_out_10_port, 
                           shiftLeftOnePos(9) => plus4A_out_9_port, 
                           shiftLeftOnePos(8) => plus4A_out_8_port, 
                           shiftLeftOnePos(7) => plus4A_out_7_port, 
                           shiftLeftOnePos(6) => plus4A_out_6_port, 
                           shiftLeftOnePos(5) => plus4A_out_5_port, 
                           shiftLeftOnePos(4) => plus4A_out_4_port, 
                           shiftLeftOnePos(3) => plus4A_out_3_port, 
                           shiftLeftOnePos(2) => plus4A_out_2_port, 
                           shiftLeftOnePos(1) => plus4A_out_1_port, 
                           shiftLeftOnePos(0) => n_3153);
   complementer_1 : complementer_N64_10 port map( input(63) => 
                           plus2A_out_63_port, input(62) => plus2A_out_62_port,
                           input(61) => plus2A_out_61_port, input(60) => 
                           plus2A_out_60_port, input(59) => plus2A_out_59_port,
                           input(58) => plus2A_out_58_port, input(57) => 
                           plus2A_out_57_port, input(56) => plus2A_out_56_port,
                           input(55) => plus2A_out_55_port, input(54) => 
                           plus2A_out_54_port, input(53) => plus2A_out_53_port,
                           input(52) => plus2A_out_52_port, input(51) => 
                           plus2A_out_51_port, input(50) => plus2A_out_50_port,
                           input(49) => plus2A_out_49_port, input(48) => 
                           plus2A_out_48_port, input(47) => plus2A_out_47_port,
                           input(46) => plus2A_out_46_port, input(45) => 
                           plus2A_out_45_port, input(44) => plus2A_out_44_port,
                           input(43) => plus2A_out_43_port, input(42) => 
                           plus2A_out_42_port, input(41) => plus2A_out_41_port,
                           input(40) => plus2A_out_40_port, input(39) => 
                           plus2A_out_39_port, input(38) => plus2A_out_38_port,
                           input(37) => plus2A_out_37_port, input(36) => 
                           plus2A_out_36_port, input(35) => plus2A_out_35_port,
                           input(34) => plus2A_out_34_port, input(33) => 
                           plus2A_out_33_port, input(32) => plus2A_out_32_port,
                           input(31) => plus2A_out_31_port, input(30) => 
                           plus2A_out_30_port, input(29) => plus2A_out_29_port,
                           input(28) => plus2A_out_28_port, input(27) => 
                           plus2A_out_27_port, input(26) => plus2A_out_26_port,
                           input(25) => plus2A_out_25_port, input(24) => 
                           plus2A_out_24_port, input(23) => plus2A_out_23_port,
                           input(22) => plus2A_out_22_port, input(21) => 
                           plus2A_out_21_port, input(20) => plus2A_out_20_port,
                           input(19) => plus2A_out_19_port, input(18) => 
                           plus2A_out_18_port, input(17) => plus2A_out_17_port,
                           input(16) => plus2A_out_16_port, input(15) => 
                           plus2A_out_15_port, input(14) => plus2A_out_14_port,
                           input(13) => plus2A_out_13_port, input(12) => 
                           plus2A_out_12_port, input(11) => plus2A_out_11_port,
                           input(10) => plus2A_out_10_port, input(9) => 
                           plus2A_out_9_port, input(8) => plus2A_out_8_port, 
                           input(7) => plus2A_out_7_port, input(6) => 
                           plus2A_out_6_port, input(5) => plus2A_out_5_port, 
                           input(4) => plus2A_out_4_port, input(3) => 
                           plus2A_out_3_port, input(2) => plus2A_out_2_port, 
                           input(1) => plus2A_out_1_port, input(0) => 
                           plus2A_out_0_port, complement2(63) => 
                           minus2A_out(63), complement2(62) => minus2A_out(62),
                           complement2(61) => minus2A_out(61), complement2(60) 
                           => minus2A_out(60), complement2(59) => 
                           minus2A_out(59), complement2(58) => minus2A_out(58),
                           complement2(57) => minus2A_out(57), complement2(56) 
                           => minus2A_out(56), complement2(55) => 
                           minus2A_out(55), complement2(54) => minus2A_out(54),
                           complement2(53) => minus2A_out(53), complement2(52) 
                           => minus2A_out(52), complement2(51) => 
                           minus2A_out(51), complement2(50) => minus2A_out(50),
                           complement2(49) => minus2A_out(49), complement2(48) 
                           => minus2A_out(48), complement2(47) => 
                           minus2A_out(47), complement2(46) => minus2A_out(46),
                           complement2(45) => minus2A_out(45), complement2(44) 
                           => minus2A_out(44), complement2(43) => 
                           minus2A_out(43), complement2(42) => minus2A_out(42),
                           complement2(41) => minus2A_out(41), complement2(40) 
                           => minus2A_out(40), complement2(39) => 
                           minus2A_out(39), complement2(38) => minus2A_out(38),
                           complement2(37) => minus2A_out(37), complement2(36) 
                           => minus2A_out(36), complement2(35) => 
                           minus2A_out(35), complement2(34) => minus2A_out(34),
                           complement2(33) => minus2A_out(33), complement2(32) 
                           => minus2A_out(32), complement2(31) => 
                           minus2A_out(31), complement2(30) => minus2A_out(30),
                           complement2(29) => minus2A_out(29), complement2(28) 
                           => minus2A_out(28), complement2(27) => 
                           minus2A_out(27), complement2(26) => minus2A_out(26),
                           complement2(25) => minus2A_out(25), complement2(24) 
                           => minus2A_out(24), complement2(23) => 
                           minus2A_out(23), complement2(22) => minus2A_out(22),
                           complement2(21) => minus2A_out(21), complement2(20) 
                           => minus2A_out(20), complement2(19) => 
                           minus2A_out(19), complement2(18) => minus2A_out(18),
                           complement2(17) => minus2A_out(17), complement2(16) 
                           => minus2A_out(16), complement2(15) => 
                           minus2A_out(15), complement2(14) => minus2A_out(14),
                           complement2(13) => minus2A_out(13), complement2(12) 
                           => minus2A_out(12), complement2(11) => 
                           minus2A_out(11), complement2(10) => minus2A_out(10),
                           complement2(9) => minus2A_out(9), complement2(8) => 
                           minus2A_out(8), complement2(7) => minus2A_out(7), 
                           complement2(6) => minus2A_out(6), complement2(5) => 
                           minus2A_out(5), complement2(4) => minus2A_out(4), 
                           complement2(3) => minus2A_out(3), complement2(2) => 
                           minus2A_out(2), complement2(1) => minus2A_out(1), 
                           complement2(0) => minus2A_out(0));
   complementer_2 : complementer_N64_9 port map( input(63) => 
                           plus4A_out_63_port, input(62) => plus4A_out_62_port,
                           input(61) => plus4A_out_61_port, input(60) => 
                           plus4A_out_60_port, input(59) => plus4A_out_59_port,
                           input(58) => plus4A_out_58_port, input(57) => 
                           plus4A_out_57_port, input(56) => plus4A_out_56_port,
                           input(55) => plus4A_out_55_port, input(54) => 
                           plus4A_out_54_port, input(53) => plus4A_out_53_port,
                           input(52) => plus4A_out_52_port, input(51) => 
                           plus4A_out_51_port, input(50) => plus4A_out_50_port,
                           input(49) => plus4A_out_49_port, input(48) => 
                           plus4A_out_48_port, input(47) => plus4A_out_47_port,
                           input(46) => plus4A_out_46_port, input(45) => 
                           plus4A_out_45_port, input(44) => plus4A_out_44_port,
                           input(43) => plus4A_out_43_port, input(42) => 
                           plus4A_out_42_port, input(41) => plus4A_out_41_port,
                           input(40) => plus4A_out_40_port, input(39) => 
                           plus4A_out_39_port, input(38) => plus4A_out_38_port,
                           input(37) => plus4A_out_37_port, input(36) => 
                           plus4A_out_36_port, input(35) => plus4A_out_35_port,
                           input(34) => plus4A_out_34_port, input(33) => 
                           plus4A_out_33_port, input(32) => plus4A_out_32_port,
                           input(31) => plus4A_out_31_port, input(30) => 
                           plus4A_out_30_port, input(29) => plus4A_out_29_port,
                           input(28) => plus4A_out_28_port, input(27) => 
                           plus4A_out_27_port, input(26) => plus4A_out_26_port,
                           input(25) => plus4A_out_25_port, input(24) => 
                           plus4A_out_24_port, input(23) => plus4A_out_23_port,
                           input(22) => plus4A_out_22_port, input(21) => 
                           plus4A_out_21_port, input(20) => plus4A_out_20_port,
                           input(19) => plus4A_out_19_port, input(18) => 
                           plus4A_out_18_port, input(17) => plus4A_out_17_port,
                           input(16) => plus4A_out_16_port, input(15) => 
                           plus4A_out_15_port, input(14) => plus4A_out_14_port,
                           input(13) => plus4A_out_13_port, input(12) => 
                           plus4A_out_12_port, input(11) => plus4A_out_11_port,
                           input(10) => plus4A_out_10_port, input(9) => 
                           plus4A_out_9_port, input(8) => plus4A_out_8_port, 
                           input(7) => plus4A_out_7_port, input(6) => 
                           plus4A_out_6_port, input(5) => plus4A_out_5_port, 
                           input(4) => plus4A_out_4_port, input(3) => 
                           plus4A_out_3_port, input(2) => plus4A_out_2_port, 
                           input(1) => plus4A_out_1_port, input(0) => 
                           plus4A_out_0_port, complement2(63) => 
                           minus4A_out(63), complement2(62) => minus4A_out(62),
                           complement2(61) => minus4A_out(61), complement2(60) 
                           => minus4A_out(60), complement2(59) => 
                           minus4A_out(59), complement2(58) => minus4A_out(58),
                           complement2(57) => minus4A_out(57), complement2(56) 
                           => minus4A_out(56), complement2(55) => 
                           minus4A_out(55), complement2(54) => minus4A_out(54),
                           complement2(53) => minus4A_out(53), complement2(52) 
                           => minus4A_out(52), complement2(51) => 
                           minus4A_out(51), complement2(50) => minus4A_out(50),
                           complement2(49) => minus4A_out(49), complement2(48) 
                           => minus4A_out(48), complement2(47) => 
                           minus4A_out(47), complement2(46) => minus4A_out(46),
                           complement2(45) => minus4A_out(45), complement2(44) 
                           => minus4A_out(44), complement2(43) => 
                           minus4A_out(43), complement2(42) => minus4A_out(42),
                           complement2(41) => minus4A_out(41), complement2(40) 
                           => minus4A_out(40), complement2(39) => 
                           minus4A_out(39), complement2(38) => minus4A_out(38),
                           complement2(37) => minus4A_out(37), complement2(36) 
                           => minus4A_out(36), complement2(35) => 
                           minus4A_out(35), complement2(34) => minus4A_out(34),
                           complement2(33) => minus4A_out(33), complement2(32) 
                           => minus4A_out(32), complement2(31) => 
                           minus4A_out(31), complement2(30) => minus4A_out(30),
                           complement2(29) => minus4A_out(29), complement2(28) 
                           => minus4A_out(28), complement2(27) => 
                           minus4A_out(27), complement2(26) => minus4A_out(26),
                           complement2(25) => minus4A_out(25), complement2(24) 
                           => minus4A_out(24), complement2(23) => 
                           minus4A_out(23), complement2(22) => minus4A_out(22),
                           complement2(21) => minus4A_out(21), complement2(20) 
                           => minus4A_out(20), complement2(19) => 
                           minus4A_out(19), complement2(18) => minus4A_out(18),
                           complement2(17) => minus4A_out(17), complement2(16) 
                           => minus4A_out(16), complement2(15) => 
                           minus4A_out(15), complement2(14) => minus4A_out(14),
                           complement2(13) => minus4A_out(13), complement2(12) 
                           => minus4A_out(12), complement2(11) => 
                           minus4A_out(11), complement2(10) => minus4A_out(10),
                           complement2(9) => minus4A_out(9), complement2(8) => 
                           minus4A_out(8), complement2(7) => minus4A_out(7), 
                           complement2(6) => minus4A_out(6), complement2(5) => 
                           minus4A_out(5), complement2(4) => minus4A_out(4), 
                           complement2(3) => minus4A_out(3), complement2(2) => 
                           minus4A_out(2), complement2(1) => minus4A_out(1), 
                           complement2(0) => minus4A_out(0));
   U3 : BUF_X1 port map( A => n32, Z => plus2A_out_57_port);
   U4 : BUF_X1 port map( A => n61, Z => plus2A_out_23_port);
   U5 : BUF_X1 port map( A => n59, Z => plus2A_out_25_port);
   U6 : BUF_X1 port map( A => n60, Z => plus2A_out_24_port);
   U7 : BUF_X1 port map( A => n58, Z => plus2A_out_26_port);
   U8 : BUF_X1 port map( A => n62, Z => plus2A_out_22_port);
   U9 : BUF_X1 port map( A => n49, Z => plus2A_out_35_port);
   U10 : BUF_X1 port map( A => n53, Z => plus2A_out_31_port);
   U11 : BUF_X1 port map( A => n57, Z => plus2A_out_27_port);
   U12 : BUF_X1 port map( A => n47, Z => plus2A_out_37_port);
   U13 : BUF_X1 port map( A => n51, Z => plus2A_out_33_port);
   U14 : BUF_X1 port map( A => n55, Z => plus2A_out_29_port);
   U15 : BUF_X1 port map( A => n48, Z => plus2A_out_36_port);
   U16 : BUF_X1 port map( A => n52, Z => plus2A_out_32_port);
   U17 : BUF_X1 port map( A => n56, Z => plus2A_out_28_port);
   U18 : BUF_X1 port map( A => n50, Z => plus2A_out_34_port);
   U19 : BUF_X1 port map( A => n54, Z => plus2A_out_30_port);
   U20 : BUF_X1 port map( A => n37, Z => plus2A_out_47_port);
   U21 : BUF_X1 port map( A => n41, Z => plus2A_out_43_port);
   U22 : BUF_X1 port map( A => n45, Z => plus2A_out_39_port);
   U23 : BUF_X1 port map( A => n39, Z => plus2A_out_45_port);
   U24 : BUF_X1 port map( A => n43, Z => plus2A_out_41_port);
   U25 : BUF_X1 port map( A => n36, Z => plus2A_out_48_port);
   U26 : BUF_X1 port map( A => n40, Z => plus2A_out_44_port);
   U27 : BUF_X1 port map( A => n44, Z => plus2A_out_40_port);
   U28 : BUF_X1 port map( A => n38, Z => plus2A_out_46_port);
   U29 : BUF_X1 port map( A => n42, Z => plus2A_out_42_port);
   U30 : BUF_X1 port map( A => n46, Z => plus2A_out_38_port);
   U31 : BUF_X1 port map( A => n33, Z => plus2A_out_51_port);
   U32 : BUF_X1 port map( A => n35, Z => plus2A_out_49_port);
   U33 : BUF_X1 port map( A => n34, Z => plus2A_out_50_port);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity ShiftnCompl_N64_6 is

   port( plusA : in std_logic_vector (63 downto 0);  plus2A_out, minus2A_out, 
         plus4A_out, minus4A_out : out std_logic_vector (63 downto 0));

end ShiftnCompl_N64_6;

architecture SYN_struct of ShiftnCompl_N64_6 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component complementer_N64_11
      port( input : in std_logic_vector (63 downto 0);  complement2 : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component complementer_N64_12
      port( input : in std_logic_vector (63 downto 0);  complement2 : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component shifter_N64_11
      port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component shifter_N64_12
      port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
            std_logic_vector (63 downto 0));
   end component;
   
   signal plus2A_out_63_port, plus2A_out_62_port, plus2A_out_61_port, 
      plus2A_out_60_port, plus2A_out_59_port, plus2A_out_58_port, n5, 
      plus2A_out_56_port, plus2A_out_55_port, plus2A_out_54_port, 
      plus2A_out_53_port, plus2A_out_52_port, plus2A_out_51_port, 
      plus2A_out_50_port, plus2A_out_49_port, plus2A_out_48_port, 
      plus2A_out_47_port, plus2A_out_46_port, plus2A_out_45_port, 
      plus2A_out_44_port, plus2A_out_43_port, plus2A_out_42_port, 
      plus2A_out_41_port, plus2A_out_40_port, plus2A_out_39_port, 
      plus2A_out_38_port, plus2A_out_37_port, plus2A_out_36_port, 
      plus2A_out_35_port, plus2A_out_34_port, plus2A_out_33_port, 
      plus2A_out_32_port, plus2A_out_31_port, plus2A_out_30_port, 
      plus2A_out_29_port, plus2A_out_28_port, plus2A_out_27_port, 
      plus2A_out_26_port, plus2A_out_25_port, plus2A_out_24_port, 
      plus2A_out_23_port, plus2A_out_22_port, plus2A_out_21_port, 
      plus2A_out_20_port, plus2A_out_19_port, plus2A_out_18_port, 
      plus2A_out_17_port, plus2A_out_16_port, plus2A_out_15_port, 
      plus2A_out_14_port, plus2A_out_13_port, plus2A_out_12_port, 
      plus2A_out_11_port, plus2A_out_10_port, plus2A_out_9_port, 
      plus2A_out_8_port, plus2A_out_7_port, plus2A_out_6_port, 
      plus2A_out_5_port, plus2A_out_4_port, plus2A_out_3_port, 
      plus2A_out_2_port, plus2A_out_1_port, plus2A_out_0_port, 
      plus4A_out_63_port, plus4A_out_62_port, plus4A_out_61_port, 
      plus4A_out_60_port, plus4A_out_59_port, plus4A_out_58_port, 
      plus4A_out_57_port, plus4A_out_56_port, plus4A_out_55_port, 
      plus4A_out_54_port, n6, n7, n8, plus4A_out_50_port, plus4A_out_49_port, 
      plus4A_out_48_port, plus4A_out_47_port, plus4A_out_46_port, 
      plus4A_out_45_port, plus4A_out_44_port, plus4A_out_43_port, 
      plus4A_out_42_port, plus4A_out_41_port, plus4A_out_40_port, 
      plus4A_out_39_port, plus4A_out_38_port, plus4A_out_37_port, 
      plus4A_out_36_port, plus4A_out_35_port, plus4A_out_34_port, 
      plus4A_out_33_port, plus4A_out_32_port, plus4A_out_31_port, 
      plus4A_out_30_port, plus4A_out_29_port, plus4A_out_28_port, 
      plus4A_out_27_port, plus4A_out_26_port, plus4A_out_25_port, 
      plus4A_out_24_port, plus4A_out_23_port, plus4A_out_22_port, 
      plus4A_out_21_port, plus4A_out_20_port, plus4A_out_19_port, 
      plus4A_out_18_port, plus4A_out_17_port, plus4A_out_16_port, 
      plus4A_out_15_port, plus4A_out_14_port, plus4A_out_13_port, 
      plus4A_out_12_port, plus4A_out_11_port, plus4A_out_10_port, 
      plus4A_out_9_port, plus4A_out_8_port, plus4A_out_7_port, 
      plus4A_out_6_port, plus4A_out_5_port, plus4A_out_4_port, 
      plus4A_out_3_port, plus4A_out_2_port, plus4A_out_1_port, 
      plus4A_out_0_port, plus4A_out_51_port, plus4A_out_52_port, 
      plus4A_out_53_port, plus2A_out_57_port, n_3154, n_3155 : std_logic;

begin
   plus2A_out <= ( plus2A_out_63_port, plus2A_out_62_port, plus2A_out_61_port, 
      plus2A_out_60_port, plus2A_out_59_port, plus2A_out_58_port, 
      plus2A_out_57_port, plus2A_out_56_port, plus2A_out_55_port, 
      plus2A_out_54_port, plus2A_out_53_port, plus2A_out_52_port, 
      plus2A_out_51_port, plus2A_out_50_port, plus2A_out_49_port, 
      plus2A_out_48_port, plus2A_out_47_port, plus2A_out_46_port, 
      plus2A_out_45_port, plus2A_out_44_port, plus2A_out_43_port, 
      plus2A_out_42_port, plus2A_out_41_port, plus2A_out_40_port, 
      plus2A_out_39_port, plus2A_out_38_port, plus2A_out_37_port, 
      plus2A_out_36_port, plus2A_out_35_port, plus2A_out_34_port, 
      plus2A_out_33_port, plus2A_out_32_port, plus2A_out_31_port, 
      plus2A_out_30_port, plus2A_out_29_port, plus2A_out_28_port, 
      plus2A_out_27_port, plus2A_out_26_port, plus2A_out_25_port, 
      plus2A_out_24_port, plus2A_out_23_port, plus2A_out_22_port, 
      plus2A_out_21_port, plus2A_out_20_port, plus2A_out_19_port, 
      plus2A_out_18_port, plus2A_out_17_port, plus2A_out_16_port, 
      plus2A_out_15_port, plus2A_out_14_port, plus2A_out_13_port, 
      plus2A_out_12_port, plus2A_out_11_port, plus2A_out_10_port, 
      plus2A_out_9_port, plus2A_out_8_port, plus2A_out_7_port, 
      plus2A_out_6_port, plus2A_out_5_port, plus2A_out_4_port, 
      plus2A_out_3_port, plus2A_out_2_port, plus2A_out_1_port, 
      plus2A_out_0_port );
   plus4A_out <= ( plus4A_out_63_port, plus4A_out_62_port, plus4A_out_61_port, 
      plus4A_out_60_port, plus4A_out_59_port, plus4A_out_58_port, 
      plus4A_out_57_port, plus4A_out_56_port, plus4A_out_55_port, 
      plus4A_out_54_port, plus4A_out_53_port, plus4A_out_52_port, 
      plus4A_out_51_port, plus4A_out_50_port, plus4A_out_49_port, 
      plus4A_out_48_port, plus4A_out_47_port, plus4A_out_46_port, 
      plus4A_out_45_port, plus4A_out_44_port, plus4A_out_43_port, 
      plus4A_out_42_port, plus4A_out_41_port, plus4A_out_40_port, 
      plus4A_out_39_port, plus4A_out_38_port, plus4A_out_37_port, 
      plus4A_out_36_port, plus4A_out_35_port, plus4A_out_34_port, 
      plus4A_out_33_port, plus4A_out_32_port, plus4A_out_31_port, 
      plus4A_out_30_port, plus4A_out_29_port, plus4A_out_28_port, 
      plus4A_out_27_port, plus4A_out_26_port, plus4A_out_25_port, 
      plus4A_out_24_port, plus4A_out_23_port, plus4A_out_22_port, 
      plus4A_out_21_port, plus4A_out_20_port, plus4A_out_19_port, 
      plus4A_out_18_port, plus4A_out_17_port, plus4A_out_16_port, 
      plus4A_out_15_port, plus4A_out_14_port, plus4A_out_13_port, 
      plus4A_out_12_port, plus4A_out_11_port, plus4A_out_10_port, 
      plus4A_out_9_port, plus4A_out_8_port, plus4A_out_7_port, 
      plus4A_out_6_port, plus4A_out_5_port, plus4A_out_4_port, 
      plus4A_out_3_port, plus4A_out_2_port, plus4A_out_1_port, 
      plus4A_out_0_port );
   
   plus2A_out_0_port <= '0';
   plus4A_out_0_port <= '0';
   shifter_1 : shifter_N64_12 port map( input(63) => plusA(63), input(62) => 
                           plusA(62), input(61) => plusA(61), input(60) => 
                           plusA(60), input(59) => plusA(59), input(58) => 
                           plusA(58), input(57) => plusA(57), input(56) => 
                           plusA(56), input(55) => plusA(55), input(54) => 
                           plusA(54), input(53) => plusA(53), input(52) => 
                           plusA(52), input(51) => plusA(51), input(50) => 
                           plusA(50), input(49) => plusA(49), input(48) => 
                           plusA(48), input(47) => plusA(47), input(46) => 
                           plusA(46), input(45) => plusA(45), input(44) => 
                           plusA(44), input(43) => plusA(43), input(42) => 
                           plusA(42), input(41) => plusA(41), input(40) => 
                           plusA(40), input(39) => plusA(39), input(38) => 
                           plusA(38), input(37) => plusA(37), input(36) => 
                           plusA(36), input(35) => plusA(35), input(34) => 
                           plusA(34), input(33) => plusA(33), input(32) => 
                           plusA(32), input(31) => plusA(31), input(30) => 
                           plusA(30), input(29) => plusA(29), input(28) => 
                           plusA(28), input(27) => plusA(27), input(26) => 
                           plusA(26), input(25) => plusA(25), input(24) => 
                           plusA(24), input(23) => plusA(23), input(22) => 
                           plusA(22), input(21) => plusA(21), input(20) => 
                           plusA(20), input(19) => plusA(19), input(18) => 
                           plusA(18), input(17) => plusA(17), input(16) => 
                           plusA(16), input(15) => plusA(15), input(14) => 
                           plusA(14), input(13) => plusA(13), input(12) => 
                           plusA(12), input(11) => plusA(11), input(10) => 
                           plusA(10), input(9) => plusA(9), input(8) => 
                           plusA(8), input(7) => plusA(7), input(6) => plusA(6)
                           , input(5) => plusA(5), input(4) => plusA(4), 
                           input(3) => plusA(3), input(2) => plusA(2), input(1)
                           => plusA(1), input(0) => plusA(0), 
                           shiftLeftOnePos(63) => plus2A_out_63_port, 
                           shiftLeftOnePos(62) => plus2A_out_62_port, 
                           shiftLeftOnePos(61) => plus2A_out_61_port, 
                           shiftLeftOnePos(60) => plus2A_out_60_port, 
                           shiftLeftOnePos(59) => plus2A_out_59_port, 
                           shiftLeftOnePos(58) => plus2A_out_58_port, 
                           shiftLeftOnePos(57) => n5, shiftLeftOnePos(56) => 
                           plus2A_out_56_port, shiftLeftOnePos(55) => 
                           plus2A_out_55_port, shiftLeftOnePos(54) => 
                           plus2A_out_54_port, shiftLeftOnePos(53) => 
                           plus2A_out_53_port, shiftLeftOnePos(52) => 
                           plus2A_out_52_port, shiftLeftOnePos(51) => 
                           plus2A_out_51_port, shiftLeftOnePos(50) => 
                           plus2A_out_50_port, shiftLeftOnePos(49) => 
                           plus2A_out_49_port, shiftLeftOnePos(48) => 
                           plus2A_out_48_port, shiftLeftOnePos(47) => 
                           plus2A_out_47_port, shiftLeftOnePos(46) => 
                           plus2A_out_46_port, shiftLeftOnePos(45) => 
                           plus2A_out_45_port, shiftLeftOnePos(44) => 
                           plus2A_out_44_port, shiftLeftOnePos(43) => 
                           plus2A_out_43_port, shiftLeftOnePos(42) => 
                           plus2A_out_42_port, shiftLeftOnePos(41) => 
                           plus2A_out_41_port, shiftLeftOnePos(40) => 
                           plus2A_out_40_port, shiftLeftOnePos(39) => 
                           plus2A_out_39_port, shiftLeftOnePos(38) => 
                           plus2A_out_38_port, shiftLeftOnePos(37) => 
                           plus2A_out_37_port, shiftLeftOnePos(36) => 
                           plus2A_out_36_port, shiftLeftOnePos(35) => 
                           plus2A_out_35_port, shiftLeftOnePos(34) => 
                           plus2A_out_34_port, shiftLeftOnePos(33) => 
                           plus2A_out_33_port, shiftLeftOnePos(32) => 
                           plus2A_out_32_port, shiftLeftOnePos(31) => 
                           plus2A_out_31_port, shiftLeftOnePos(30) => 
                           plus2A_out_30_port, shiftLeftOnePos(29) => 
                           plus2A_out_29_port, shiftLeftOnePos(28) => 
                           plus2A_out_28_port, shiftLeftOnePos(27) => 
                           plus2A_out_27_port, shiftLeftOnePos(26) => 
                           plus2A_out_26_port, shiftLeftOnePos(25) => 
                           plus2A_out_25_port, shiftLeftOnePos(24) => 
                           plus2A_out_24_port, shiftLeftOnePos(23) => 
                           plus2A_out_23_port, shiftLeftOnePos(22) => 
                           plus2A_out_22_port, shiftLeftOnePos(21) => 
                           plus2A_out_21_port, shiftLeftOnePos(20) => 
                           plus2A_out_20_port, shiftLeftOnePos(19) => 
                           plus2A_out_19_port, shiftLeftOnePos(18) => 
                           plus2A_out_18_port, shiftLeftOnePos(17) => 
                           plus2A_out_17_port, shiftLeftOnePos(16) => 
                           plus2A_out_16_port, shiftLeftOnePos(15) => 
                           plus2A_out_15_port, shiftLeftOnePos(14) => 
                           plus2A_out_14_port, shiftLeftOnePos(13) => 
                           plus2A_out_13_port, shiftLeftOnePos(12) => 
                           plus2A_out_12_port, shiftLeftOnePos(11) => 
                           plus2A_out_11_port, shiftLeftOnePos(10) => 
                           plus2A_out_10_port, shiftLeftOnePos(9) => 
                           plus2A_out_9_port, shiftLeftOnePos(8) => 
                           plus2A_out_8_port, shiftLeftOnePos(7) => 
                           plus2A_out_7_port, shiftLeftOnePos(6) => 
                           plus2A_out_6_port, shiftLeftOnePos(5) => 
                           plus2A_out_5_port, shiftLeftOnePos(4) => 
                           plus2A_out_4_port, shiftLeftOnePos(3) => 
                           plus2A_out_3_port, shiftLeftOnePos(2) => 
                           plus2A_out_2_port, shiftLeftOnePos(1) => 
                           plus2A_out_1_port, shiftLeftOnePos(0) => n_3154);
   shifter_2 : shifter_N64_11 port map( input(63) => plus2A_out_63_port, 
                           input(62) => plus2A_out_62_port, input(61) => 
                           plus2A_out_61_port, input(60) => plus2A_out_60_port,
                           input(59) => plus2A_out_59_port, input(58) => 
                           plus2A_out_58_port, input(57) => plus2A_out_57_port,
                           input(56) => plus2A_out_56_port, input(55) => 
                           plus2A_out_55_port, input(54) => plus2A_out_54_port,
                           input(53) => plus2A_out_53_port, input(52) => 
                           plus2A_out_52_port, input(51) => plus2A_out_51_port,
                           input(50) => plus2A_out_50_port, input(49) => 
                           plus2A_out_49_port, input(48) => plus2A_out_48_port,
                           input(47) => plus2A_out_47_port, input(46) => 
                           plus2A_out_46_port, input(45) => plus2A_out_45_port,
                           input(44) => plus2A_out_44_port, input(43) => 
                           plus2A_out_43_port, input(42) => plus2A_out_42_port,
                           input(41) => plus2A_out_41_port, input(40) => 
                           plus2A_out_40_port, input(39) => plus2A_out_39_port,
                           input(38) => plus2A_out_38_port, input(37) => 
                           plus2A_out_37_port, input(36) => plus2A_out_36_port,
                           input(35) => plus2A_out_35_port, input(34) => 
                           plus2A_out_34_port, input(33) => plus2A_out_33_port,
                           input(32) => plus2A_out_32_port, input(31) => 
                           plus2A_out_31_port, input(30) => plus2A_out_30_port,
                           input(29) => plus2A_out_29_port, input(28) => 
                           plus2A_out_28_port, input(27) => plus2A_out_27_port,
                           input(26) => plus2A_out_26_port, input(25) => 
                           plus2A_out_25_port, input(24) => plus2A_out_24_port,
                           input(23) => plus2A_out_23_port, input(22) => 
                           plus2A_out_22_port, input(21) => plus2A_out_21_port,
                           input(20) => plus2A_out_20_port, input(19) => 
                           plus2A_out_19_port, input(18) => plus2A_out_18_port,
                           input(17) => plus2A_out_17_port, input(16) => 
                           plus2A_out_16_port, input(15) => plus2A_out_15_port,
                           input(14) => plus2A_out_14_port, input(13) => 
                           plus2A_out_13_port, input(12) => plus2A_out_12_port,
                           input(11) => plus2A_out_11_port, input(10) => 
                           plus2A_out_10_port, input(9) => plus2A_out_9_port, 
                           input(8) => plus2A_out_8_port, input(7) => 
                           plus2A_out_7_port, input(6) => plus2A_out_6_port, 
                           input(5) => plus2A_out_5_port, input(4) => 
                           plus2A_out_4_port, input(3) => plus2A_out_3_port, 
                           input(2) => plus2A_out_2_port, input(1) => 
                           plus2A_out_1_port, input(0) => plus2A_out_0_port, 
                           shiftLeftOnePos(63) => plus4A_out_63_port, 
                           shiftLeftOnePos(62) => plus4A_out_62_port, 
                           shiftLeftOnePos(61) => plus4A_out_61_port, 
                           shiftLeftOnePos(60) => plus4A_out_60_port, 
                           shiftLeftOnePos(59) => plus4A_out_59_port, 
                           shiftLeftOnePos(58) => plus4A_out_58_port, 
                           shiftLeftOnePos(57) => plus4A_out_57_port, 
                           shiftLeftOnePos(56) => plus4A_out_56_port, 
                           shiftLeftOnePos(55) => plus4A_out_55_port, 
                           shiftLeftOnePos(54) => plus4A_out_54_port, 
                           shiftLeftOnePos(53) => n6, shiftLeftOnePos(52) => n7
                           , shiftLeftOnePos(51) => n8, shiftLeftOnePos(50) => 
                           plus4A_out_50_port, shiftLeftOnePos(49) => 
                           plus4A_out_49_port, shiftLeftOnePos(48) => 
                           plus4A_out_48_port, shiftLeftOnePos(47) => 
                           plus4A_out_47_port, shiftLeftOnePos(46) => 
                           plus4A_out_46_port, shiftLeftOnePos(45) => 
                           plus4A_out_45_port, shiftLeftOnePos(44) => 
                           plus4A_out_44_port, shiftLeftOnePos(43) => 
                           plus4A_out_43_port, shiftLeftOnePos(42) => 
                           plus4A_out_42_port, shiftLeftOnePos(41) => 
                           plus4A_out_41_port, shiftLeftOnePos(40) => 
                           plus4A_out_40_port, shiftLeftOnePos(39) => 
                           plus4A_out_39_port, shiftLeftOnePos(38) => 
                           plus4A_out_38_port, shiftLeftOnePos(37) => 
                           plus4A_out_37_port, shiftLeftOnePos(36) => 
                           plus4A_out_36_port, shiftLeftOnePos(35) => 
                           plus4A_out_35_port, shiftLeftOnePos(34) => 
                           plus4A_out_34_port, shiftLeftOnePos(33) => 
                           plus4A_out_33_port, shiftLeftOnePos(32) => 
                           plus4A_out_32_port, shiftLeftOnePos(31) => 
                           plus4A_out_31_port, shiftLeftOnePos(30) => 
                           plus4A_out_30_port, shiftLeftOnePos(29) => 
                           plus4A_out_29_port, shiftLeftOnePos(28) => 
                           plus4A_out_28_port, shiftLeftOnePos(27) => 
                           plus4A_out_27_port, shiftLeftOnePos(26) => 
                           plus4A_out_26_port, shiftLeftOnePos(25) => 
                           plus4A_out_25_port, shiftLeftOnePos(24) => 
                           plus4A_out_24_port, shiftLeftOnePos(23) => 
                           plus4A_out_23_port, shiftLeftOnePos(22) => 
                           plus4A_out_22_port, shiftLeftOnePos(21) => 
                           plus4A_out_21_port, shiftLeftOnePos(20) => 
                           plus4A_out_20_port, shiftLeftOnePos(19) => 
                           plus4A_out_19_port, shiftLeftOnePos(18) => 
                           plus4A_out_18_port, shiftLeftOnePos(17) => 
                           plus4A_out_17_port, shiftLeftOnePos(16) => 
                           plus4A_out_16_port, shiftLeftOnePos(15) => 
                           plus4A_out_15_port, shiftLeftOnePos(14) => 
                           plus4A_out_14_port, shiftLeftOnePos(13) => 
                           plus4A_out_13_port, shiftLeftOnePos(12) => 
                           plus4A_out_12_port, shiftLeftOnePos(11) => 
                           plus4A_out_11_port, shiftLeftOnePos(10) => 
                           plus4A_out_10_port, shiftLeftOnePos(9) => 
                           plus4A_out_9_port, shiftLeftOnePos(8) => 
                           plus4A_out_8_port, shiftLeftOnePos(7) => 
                           plus4A_out_7_port, shiftLeftOnePos(6) => 
                           plus4A_out_6_port, shiftLeftOnePos(5) => 
                           plus4A_out_5_port, shiftLeftOnePos(4) => 
                           plus4A_out_4_port, shiftLeftOnePos(3) => 
                           plus4A_out_3_port, shiftLeftOnePos(2) => 
                           plus4A_out_2_port, shiftLeftOnePos(1) => 
                           plus4A_out_1_port, shiftLeftOnePos(0) => n_3155);
   complementer_1 : complementer_N64_12 port map( input(63) => 
                           plus2A_out_63_port, input(62) => plus2A_out_62_port,
                           input(61) => plus2A_out_61_port, input(60) => 
                           plus2A_out_60_port, input(59) => plus2A_out_59_port,
                           input(58) => plus2A_out_58_port, input(57) => 
                           plus2A_out_57_port, input(56) => plus2A_out_56_port,
                           input(55) => plus2A_out_55_port, input(54) => 
                           plus2A_out_54_port, input(53) => plus2A_out_53_port,
                           input(52) => plus2A_out_52_port, input(51) => 
                           plus2A_out_51_port, input(50) => plus2A_out_50_port,
                           input(49) => plus2A_out_49_port, input(48) => 
                           plus2A_out_48_port, input(47) => plus2A_out_47_port,
                           input(46) => plus2A_out_46_port, input(45) => 
                           plus2A_out_45_port, input(44) => plus2A_out_44_port,
                           input(43) => plus2A_out_43_port, input(42) => 
                           plus2A_out_42_port, input(41) => plus2A_out_41_port,
                           input(40) => plus2A_out_40_port, input(39) => 
                           plus2A_out_39_port, input(38) => plus2A_out_38_port,
                           input(37) => plus2A_out_37_port, input(36) => 
                           plus2A_out_36_port, input(35) => plus2A_out_35_port,
                           input(34) => plus2A_out_34_port, input(33) => 
                           plus2A_out_33_port, input(32) => plus2A_out_32_port,
                           input(31) => plus2A_out_31_port, input(30) => 
                           plus2A_out_30_port, input(29) => plus2A_out_29_port,
                           input(28) => plus2A_out_28_port, input(27) => 
                           plus2A_out_27_port, input(26) => plus2A_out_26_port,
                           input(25) => plus2A_out_25_port, input(24) => 
                           plus2A_out_24_port, input(23) => plus2A_out_23_port,
                           input(22) => plus2A_out_22_port, input(21) => 
                           plus2A_out_21_port, input(20) => plus2A_out_20_port,
                           input(19) => plus2A_out_19_port, input(18) => 
                           plus2A_out_18_port, input(17) => plus2A_out_17_port,
                           input(16) => plus2A_out_16_port, input(15) => 
                           plus2A_out_15_port, input(14) => plus2A_out_14_port,
                           input(13) => plus2A_out_13_port, input(12) => 
                           plus2A_out_12_port, input(11) => plus2A_out_11_port,
                           input(10) => plus2A_out_10_port, input(9) => 
                           plus2A_out_9_port, input(8) => plus2A_out_8_port, 
                           input(7) => plus2A_out_7_port, input(6) => 
                           plus2A_out_6_port, input(5) => plus2A_out_5_port, 
                           input(4) => plus2A_out_4_port, input(3) => 
                           plus2A_out_3_port, input(2) => plus2A_out_2_port, 
                           input(1) => plus2A_out_1_port, input(0) => 
                           plus2A_out_0_port, complement2(63) => 
                           minus2A_out(63), complement2(62) => minus2A_out(62),
                           complement2(61) => minus2A_out(61), complement2(60) 
                           => minus2A_out(60), complement2(59) => 
                           minus2A_out(59), complement2(58) => minus2A_out(58),
                           complement2(57) => minus2A_out(57), complement2(56) 
                           => minus2A_out(56), complement2(55) => 
                           minus2A_out(55), complement2(54) => minus2A_out(54),
                           complement2(53) => minus2A_out(53), complement2(52) 
                           => minus2A_out(52), complement2(51) => 
                           minus2A_out(51), complement2(50) => minus2A_out(50),
                           complement2(49) => minus2A_out(49), complement2(48) 
                           => minus2A_out(48), complement2(47) => 
                           minus2A_out(47), complement2(46) => minus2A_out(46),
                           complement2(45) => minus2A_out(45), complement2(44) 
                           => minus2A_out(44), complement2(43) => 
                           minus2A_out(43), complement2(42) => minus2A_out(42),
                           complement2(41) => minus2A_out(41), complement2(40) 
                           => minus2A_out(40), complement2(39) => 
                           minus2A_out(39), complement2(38) => minus2A_out(38),
                           complement2(37) => minus2A_out(37), complement2(36) 
                           => minus2A_out(36), complement2(35) => 
                           minus2A_out(35), complement2(34) => minus2A_out(34),
                           complement2(33) => minus2A_out(33), complement2(32) 
                           => minus2A_out(32), complement2(31) => 
                           minus2A_out(31), complement2(30) => minus2A_out(30),
                           complement2(29) => minus2A_out(29), complement2(28) 
                           => minus2A_out(28), complement2(27) => 
                           minus2A_out(27), complement2(26) => minus2A_out(26),
                           complement2(25) => minus2A_out(25), complement2(24) 
                           => minus2A_out(24), complement2(23) => 
                           minus2A_out(23), complement2(22) => minus2A_out(22),
                           complement2(21) => minus2A_out(21), complement2(20) 
                           => minus2A_out(20), complement2(19) => 
                           minus2A_out(19), complement2(18) => minus2A_out(18),
                           complement2(17) => minus2A_out(17), complement2(16) 
                           => minus2A_out(16), complement2(15) => 
                           minus2A_out(15), complement2(14) => minus2A_out(14),
                           complement2(13) => minus2A_out(13), complement2(12) 
                           => minus2A_out(12), complement2(11) => 
                           minus2A_out(11), complement2(10) => minus2A_out(10),
                           complement2(9) => minus2A_out(9), complement2(8) => 
                           minus2A_out(8), complement2(7) => minus2A_out(7), 
                           complement2(6) => minus2A_out(6), complement2(5) => 
                           minus2A_out(5), complement2(4) => minus2A_out(4), 
                           complement2(3) => minus2A_out(3), complement2(2) => 
                           minus2A_out(2), complement2(1) => minus2A_out(1), 
                           complement2(0) => minus2A_out(0));
   complementer_2 : complementer_N64_11 port map( input(63) => 
                           plus4A_out_63_port, input(62) => plus4A_out_62_port,
                           input(61) => plus4A_out_61_port, input(60) => 
                           plus4A_out_60_port, input(59) => plus4A_out_59_port,
                           input(58) => plus4A_out_58_port, input(57) => 
                           plus4A_out_57_port, input(56) => plus4A_out_56_port,
                           input(55) => plus4A_out_55_port, input(54) => 
                           plus4A_out_54_port, input(53) => plus4A_out_53_port,
                           input(52) => plus4A_out_52_port, input(51) => 
                           plus4A_out_51_port, input(50) => plus4A_out_50_port,
                           input(49) => plus4A_out_49_port, input(48) => 
                           plus4A_out_48_port, input(47) => plus4A_out_47_port,
                           input(46) => plus4A_out_46_port, input(45) => 
                           plus4A_out_45_port, input(44) => plus4A_out_44_port,
                           input(43) => plus4A_out_43_port, input(42) => 
                           plus4A_out_42_port, input(41) => plus4A_out_41_port,
                           input(40) => plus4A_out_40_port, input(39) => 
                           plus4A_out_39_port, input(38) => plus4A_out_38_port,
                           input(37) => plus4A_out_37_port, input(36) => 
                           plus4A_out_36_port, input(35) => plus4A_out_35_port,
                           input(34) => plus4A_out_34_port, input(33) => 
                           plus4A_out_33_port, input(32) => plus4A_out_32_port,
                           input(31) => plus4A_out_31_port, input(30) => 
                           plus4A_out_30_port, input(29) => plus4A_out_29_port,
                           input(28) => plus4A_out_28_port, input(27) => 
                           plus4A_out_27_port, input(26) => plus4A_out_26_port,
                           input(25) => plus4A_out_25_port, input(24) => 
                           plus4A_out_24_port, input(23) => plus4A_out_23_port,
                           input(22) => plus4A_out_22_port, input(21) => 
                           plus4A_out_21_port, input(20) => plus4A_out_20_port,
                           input(19) => plus4A_out_19_port, input(18) => 
                           plus4A_out_18_port, input(17) => plus4A_out_17_port,
                           input(16) => plus4A_out_16_port, input(15) => 
                           plus4A_out_15_port, input(14) => plus4A_out_14_port,
                           input(13) => plus4A_out_13_port, input(12) => 
                           plus4A_out_12_port, input(11) => plus4A_out_11_port,
                           input(10) => plus4A_out_10_port, input(9) => 
                           plus4A_out_9_port, input(8) => plus4A_out_8_port, 
                           input(7) => plus4A_out_7_port, input(6) => 
                           plus4A_out_6_port, input(5) => plus4A_out_5_port, 
                           input(4) => plus4A_out_4_port, input(3) => 
                           plus4A_out_3_port, input(2) => plus4A_out_2_port, 
                           input(1) => plus4A_out_1_port, input(0) => 
                           plus4A_out_0_port, complement2(63) => 
                           minus4A_out(63), complement2(62) => minus4A_out(62),
                           complement2(61) => minus4A_out(61), complement2(60) 
                           => minus4A_out(60), complement2(59) => 
                           minus4A_out(59), complement2(58) => minus4A_out(58),
                           complement2(57) => minus4A_out(57), complement2(56) 
                           => minus4A_out(56), complement2(55) => 
                           minus4A_out(55), complement2(54) => minus4A_out(54),
                           complement2(53) => minus4A_out(53), complement2(52) 
                           => minus4A_out(52), complement2(51) => 
                           minus4A_out(51), complement2(50) => minus4A_out(50),
                           complement2(49) => minus4A_out(49), complement2(48) 
                           => minus4A_out(48), complement2(47) => 
                           minus4A_out(47), complement2(46) => minus4A_out(46),
                           complement2(45) => minus4A_out(45), complement2(44) 
                           => minus4A_out(44), complement2(43) => 
                           minus4A_out(43), complement2(42) => minus4A_out(42),
                           complement2(41) => minus4A_out(41), complement2(40) 
                           => minus4A_out(40), complement2(39) => 
                           minus4A_out(39), complement2(38) => minus4A_out(38),
                           complement2(37) => minus4A_out(37), complement2(36) 
                           => minus4A_out(36), complement2(35) => 
                           minus4A_out(35), complement2(34) => minus4A_out(34),
                           complement2(33) => minus4A_out(33), complement2(32) 
                           => minus4A_out(32), complement2(31) => 
                           minus4A_out(31), complement2(30) => minus4A_out(30),
                           complement2(29) => minus4A_out(29), complement2(28) 
                           => minus4A_out(28), complement2(27) => 
                           minus4A_out(27), complement2(26) => minus4A_out(26),
                           complement2(25) => minus4A_out(25), complement2(24) 
                           => minus4A_out(24), complement2(23) => 
                           minus4A_out(23), complement2(22) => minus4A_out(22),
                           complement2(21) => minus4A_out(21), complement2(20) 
                           => minus4A_out(20), complement2(19) => 
                           minus4A_out(19), complement2(18) => minus4A_out(18),
                           complement2(17) => minus4A_out(17), complement2(16) 
                           => minus4A_out(16), complement2(15) => 
                           minus4A_out(15), complement2(14) => minus4A_out(14),
                           complement2(13) => minus4A_out(13), complement2(12) 
                           => minus4A_out(12), complement2(11) => 
                           minus4A_out(11), complement2(10) => minus4A_out(10),
                           complement2(9) => minus4A_out(9), complement2(8) => 
                           minus4A_out(8), complement2(7) => minus4A_out(7), 
                           complement2(6) => minus4A_out(6), complement2(5) => 
                           minus4A_out(5), complement2(4) => minus4A_out(4), 
                           complement2(3) => minus4A_out(3), complement2(2) => 
                           minus4A_out(2), complement2(1) => minus4A_out(1), 
                           complement2(0) => minus4A_out(0));
   U3 : BUF_X1 port map( A => n5, Z => plus2A_out_57_port);
   U4 : BUF_X1 port map( A => n8, Z => plus4A_out_51_port);
   U5 : BUF_X1 port map( A => n7, Z => plus4A_out_52_port);
   U6 : BUF_X1 port map( A => n6, Z => plus4A_out_53_port);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity ShiftnCompl_N64_7 is

   port( plusA : in std_logic_vector (63 downto 0);  plus2A_out, minus2A_out, 
         plus4A_out, minus4A_out : out std_logic_vector (63 downto 0));

end ShiftnCompl_N64_7;

architecture SYN_struct of ShiftnCompl_N64_7 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component complementer_N64_13
      port( input : in std_logic_vector (63 downto 0);  complement2 : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component complementer_N64_14
      port( input : in std_logic_vector (63 downto 0);  complement2 : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component shifter_N64_13
      port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component shifter_N64_14
      port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
            std_logic_vector (63 downto 0));
   end component;
   
   signal plus2A_out_63_port, plus2A_out_62_port, plus2A_out_61_port, 
      plus2A_out_60_port, plus2A_out_59_port, plus2A_out_58_port, n4, 
      plus2A_out_56_port, plus2A_out_55_port, plus2A_out_54_port, 
      plus2A_out_53_port, plus2A_out_52_port, plus2A_out_51_port, 
      plus2A_out_50_port, plus2A_out_49_port, plus2A_out_48_port, 
      plus2A_out_47_port, plus2A_out_46_port, plus2A_out_45_port, 
      plus2A_out_44_port, plus2A_out_43_port, plus2A_out_42_port, 
      plus2A_out_41_port, plus2A_out_40_port, plus2A_out_39_port, 
      plus2A_out_38_port, plus2A_out_37_port, plus2A_out_36_port, 
      plus2A_out_35_port, plus2A_out_34_port, plus2A_out_33_port, 
      plus2A_out_32_port, plus2A_out_31_port, plus2A_out_30_port, 
      plus2A_out_29_port, plus2A_out_28_port, plus2A_out_27_port, 
      plus2A_out_26_port, plus2A_out_25_port, plus2A_out_24_port, 
      plus2A_out_23_port, plus2A_out_22_port, plus2A_out_21_port, 
      plus2A_out_20_port, plus2A_out_19_port, plus2A_out_18_port, 
      plus2A_out_17_port, plus2A_out_16_port, plus2A_out_15_port, 
      plus2A_out_14_port, plus2A_out_13_port, plus2A_out_12_port, 
      plus2A_out_11_port, plus2A_out_10_port, plus2A_out_9_port, 
      plus2A_out_8_port, plus2A_out_7_port, plus2A_out_6_port, 
      plus2A_out_5_port, plus2A_out_4_port, plus2A_out_3_port, 
      plus2A_out_2_port, plus2A_out_1_port, plus2A_out_0_port, 
      plus4A_out_63_port, plus4A_out_62_port, plus4A_out_61_port, 
      plus4A_out_60_port, plus4A_out_59_port, plus4A_out_58_port, 
      plus4A_out_57_port, plus4A_out_56_port, plus4A_out_55_port, 
      plus4A_out_54_port, n5, n6, plus4A_out_51_port, plus4A_out_50_port, 
      plus4A_out_49_port, plus4A_out_48_port, plus4A_out_47_port, 
      plus4A_out_46_port, plus4A_out_45_port, plus4A_out_44_port, 
      plus4A_out_43_port, plus4A_out_42_port, plus4A_out_41_port, 
      plus4A_out_40_port, plus4A_out_39_port, plus4A_out_38_port, 
      plus4A_out_37_port, plus4A_out_36_port, plus4A_out_35_port, 
      plus4A_out_34_port, plus4A_out_33_port, plus4A_out_32_port, 
      plus4A_out_31_port, plus4A_out_30_port, plus4A_out_29_port, 
      plus4A_out_28_port, plus4A_out_27_port, plus4A_out_26_port, 
      plus4A_out_25_port, plus4A_out_24_port, plus4A_out_23_port, 
      plus4A_out_22_port, plus4A_out_21_port, plus4A_out_20_port, 
      plus4A_out_19_port, plus4A_out_18_port, plus4A_out_17_port, 
      plus4A_out_16_port, plus4A_out_15_port, plus4A_out_14_port, 
      plus4A_out_13_port, plus4A_out_12_port, plus4A_out_11_port, 
      plus4A_out_10_port, plus4A_out_9_port, plus4A_out_8_port, 
      plus4A_out_7_port, plus4A_out_6_port, plus4A_out_5_port, 
      plus4A_out_4_port, plus4A_out_3_port, plus4A_out_2_port, 
      plus4A_out_1_port, plus4A_out_0_port, plus4A_out_52_port, 
      plus4A_out_53_port, plus2A_out_57_port, n_3156, n_3157 : std_logic;

begin
   plus2A_out <= ( plus2A_out_63_port, plus2A_out_62_port, plus2A_out_61_port, 
      plus2A_out_60_port, plus2A_out_59_port, plus2A_out_58_port, 
      plus2A_out_57_port, plus2A_out_56_port, plus2A_out_55_port, 
      plus2A_out_54_port, plus2A_out_53_port, plus2A_out_52_port, 
      plus2A_out_51_port, plus2A_out_50_port, plus2A_out_49_port, 
      plus2A_out_48_port, plus2A_out_47_port, plus2A_out_46_port, 
      plus2A_out_45_port, plus2A_out_44_port, plus2A_out_43_port, 
      plus2A_out_42_port, plus2A_out_41_port, plus2A_out_40_port, 
      plus2A_out_39_port, plus2A_out_38_port, plus2A_out_37_port, 
      plus2A_out_36_port, plus2A_out_35_port, plus2A_out_34_port, 
      plus2A_out_33_port, plus2A_out_32_port, plus2A_out_31_port, 
      plus2A_out_30_port, plus2A_out_29_port, plus2A_out_28_port, 
      plus2A_out_27_port, plus2A_out_26_port, plus2A_out_25_port, 
      plus2A_out_24_port, plus2A_out_23_port, plus2A_out_22_port, 
      plus2A_out_21_port, plus2A_out_20_port, plus2A_out_19_port, 
      plus2A_out_18_port, plus2A_out_17_port, plus2A_out_16_port, 
      plus2A_out_15_port, plus2A_out_14_port, plus2A_out_13_port, 
      plus2A_out_12_port, plus2A_out_11_port, plus2A_out_10_port, 
      plus2A_out_9_port, plus2A_out_8_port, plus2A_out_7_port, 
      plus2A_out_6_port, plus2A_out_5_port, plus2A_out_4_port, 
      plus2A_out_3_port, plus2A_out_2_port, plus2A_out_1_port, 
      plus2A_out_0_port );
   plus4A_out <= ( plus4A_out_63_port, plus4A_out_62_port, plus4A_out_61_port, 
      plus4A_out_60_port, plus4A_out_59_port, plus4A_out_58_port, 
      plus4A_out_57_port, plus4A_out_56_port, plus4A_out_55_port, 
      plus4A_out_54_port, plus4A_out_53_port, plus4A_out_52_port, 
      plus4A_out_51_port, plus4A_out_50_port, plus4A_out_49_port, 
      plus4A_out_48_port, plus4A_out_47_port, plus4A_out_46_port, 
      plus4A_out_45_port, plus4A_out_44_port, plus4A_out_43_port, 
      plus4A_out_42_port, plus4A_out_41_port, plus4A_out_40_port, 
      plus4A_out_39_port, plus4A_out_38_port, plus4A_out_37_port, 
      plus4A_out_36_port, plus4A_out_35_port, plus4A_out_34_port, 
      plus4A_out_33_port, plus4A_out_32_port, plus4A_out_31_port, 
      plus4A_out_30_port, plus4A_out_29_port, plus4A_out_28_port, 
      plus4A_out_27_port, plus4A_out_26_port, plus4A_out_25_port, 
      plus4A_out_24_port, plus4A_out_23_port, plus4A_out_22_port, 
      plus4A_out_21_port, plus4A_out_20_port, plus4A_out_19_port, 
      plus4A_out_18_port, plus4A_out_17_port, plus4A_out_16_port, 
      plus4A_out_15_port, plus4A_out_14_port, plus4A_out_13_port, 
      plus4A_out_12_port, plus4A_out_11_port, plus4A_out_10_port, 
      plus4A_out_9_port, plus4A_out_8_port, plus4A_out_7_port, 
      plus4A_out_6_port, plus4A_out_5_port, plus4A_out_4_port, 
      plus4A_out_3_port, plus4A_out_2_port, plus4A_out_1_port, 
      plus4A_out_0_port );
   
   plus2A_out_0_port <= '0';
   plus4A_out_0_port <= '0';
   shifter_1 : shifter_N64_14 port map( input(63) => plusA(63), input(62) => 
                           plusA(62), input(61) => plusA(61), input(60) => 
                           plusA(60), input(59) => plusA(59), input(58) => 
                           plusA(58), input(57) => plusA(57), input(56) => 
                           plusA(56), input(55) => plusA(55), input(54) => 
                           plusA(54), input(53) => plusA(53), input(52) => 
                           plusA(52), input(51) => plusA(51), input(50) => 
                           plusA(50), input(49) => plusA(49), input(48) => 
                           plusA(48), input(47) => plusA(47), input(46) => 
                           plusA(46), input(45) => plusA(45), input(44) => 
                           plusA(44), input(43) => plusA(43), input(42) => 
                           plusA(42), input(41) => plusA(41), input(40) => 
                           plusA(40), input(39) => plusA(39), input(38) => 
                           plusA(38), input(37) => plusA(37), input(36) => 
                           plusA(36), input(35) => plusA(35), input(34) => 
                           plusA(34), input(33) => plusA(33), input(32) => 
                           plusA(32), input(31) => plusA(31), input(30) => 
                           plusA(30), input(29) => plusA(29), input(28) => 
                           plusA(28), input(27) => plusA(27), input(26) => 
                           plusA(26), input(25) => plusA(25), input(24) => 
                           plusA(24), input(23) => plusA(23), input(22) => 
                           plusA(22), input(21) => plusA(21), input(20) => 
                           plusA(20), input(19) => plusA(19), input(18) => 
                           plusA(18), input(17) => plusA(17), input(16) => 
                           plusA(16), input(15) => plusA(15), input(14) => 
                           plusA(14), input(13) => plusA(13), input(12) => 
                           plusA(12), input(11) => plusA(11), input(10) => 
                           plusA(10), input(9) => plusA(9), input(8) => 
                           plusA(8), input(7) => plusA(7), input(6) => plusA(6)
                           , input(5) => plusA(5), input(4) => plusA(4), 
                           input(3) => plusA(3), input(2) => plusA(2), input(1)
                           => plusA(1), input(0) => plusA(0), 
                           shiftLeftOnePos(63) => plus2A_out_63_port, 
                           shiftLeftOnePos(62) => plus2A_out_62_port, 
                           shiftLeftOnePos(61) => plus2A_out_61_port, 
                           shiftLeftOnePos(60) => plus2A_out_60_port, 
                           shiftLeftOnePos(59) => plus2A_out_59_port, 
                           shiftLeftOnePos(58) => plus2A_out_58_port, 
                           shiftLeftOnePos(57) => n4, shiftLeftOnePos(56) => 
                           plus2A_out_56_port, shiftLeftOnePos(55) => 
                           plus2A_out_55_port, shiftLeftOnePos(54) => 
                           plus2A_out_54_port, shiftLeftOnePos(53) => 
                           plus2A_out_53_port, shiftLeftOnePos(52) => 
                           plus2A_out_52_port, shiftLeftOnePos(51) => 
                           plus2A_out_51_port, shiftLeftOnePos(50) => 
                           plus2A_out_50_port, shiftLeftOnePos(49) => 
                           plus2A_out_49_port, shiftLeftOnePos(48) => 
                           plus2A_out_48_port, shiftLeftOnePos(47) => 
                           plus2A_out_47_port, shiftLeftOnePos(46) => 
                           plus2A_out_46_port, shiftLeftOnePos(45) => 
                           plus2A_out_45_port, shiftLeftOnePos(44) => 
                           plus2A_out_44_port, shiftLeftOnePos(43) => 
                           plus2A_out_43_port, shiftLeftOnePos(42) => 
                           plus2A_out_42_port, shiftLeftOnePos(41) => 
                           plus2A_out_41_port, shiftLeftOnePos(40) => 
                           plus2A_out_40_port, shiftLeftOnePos(39) => 
                           plus2A_out_39_port, shiftLeftOnePos(38) => 
                           plus2A_out_38_port, shiftLeftOnePos(37) => 
                           plus2A_out_37_port, shiftLeftOnePos(36) => 
                           plus2A_out_36_port, shiftLeftOnePos(35) => 
                           plus2A_out_35_port, shiftLeftOnePos(34) => 
                           plus2A_out_34_port, shiftLeftOnePos(33) => 
                           plus2A_out_33_port, shiftLeftOnePos(32) => 
                           plus2A_out_32_port, shiftLeftOnePos(31) => 
                           plus2A_out_31_port, shiftLeftOnePos(30) => 
                           plus2A_out_30_port, shiftLeftOnePos(29) => 
                           plus2A_out_29_port, shiftLeftOnePos(28) => 
                           plus2A_out_28_port, shiftLeftOnePos(27) => 
                           plus2A_out_27_port, shiftLeftOnePos(26) => 
                           plus2A_out_26_port, shiftLeftOnePos(25) => 
                           plus2A_out_25_port, shiftLeftOnePos(24) => 
                           plus2A_out_24_port, shiftLeftOnePos(23) => 
                           plus2A_out_23_port, shiftLeftOnePos(22) => 
                           plus2A_out_22_port, shiftLeftOnePos(21) => 
                           plus2A_out_21_port, shiftLeftOnePos(20) => 
                           plus2A_out_20_port, shiftLeftOnePos(19) => 
                           plus2A_out_19_port, shiftLeftOnePos(18) => 
                           plus2A_out_18_port, shiftLeftOnePos(17) => 
                           plus2A_out_17_port, shiftLeftOnePos(16) => 
                           plus2A_out_16_port, shiftLeftOnePos(15) => 
                           plus2A_out_15_port, shiftLeftOnePos(14) => 
                           plus2A_out_14_port, shiftLeftOnePos(13) => 
                           plus2A_out_13_port, shiftLeftOnePos(12) => 
                           plus2A_out_12_port, shiftLeftOnePos(11) => 
                           plus2A_out_11_port, shiftLeftOnePos(10) => 
                           plus2A_out_10_port, shiftLeftOnePos(9) => 
                           plus2A_out_9_port, shiftLeftOnePos(8) => 
                           plus2A_out_8_port, shiftLeftOnePos(7) => 
                           plus2A_out_7_port, shiftLeftOnePos(6) => 
                           plus2A_out_6_port, shiftLeftOnePos(5) => 
                           plus2A_out_5_port, shiftLeftOnePos(4) => 
                           plus2A_out_4_port, shiftLeftOnePos(3) => 
                           plus2A_out_3_port, shiftLeftOnePos(2) => 
                           plus2A_out_2_port, shiftLeftOnePos(1) => 
                           plus2A_out_1_port, shiftLeftOnePos(0) => n_3156);
   shifter_2 : shifter_N64_13 port map( input(63) => plus2A_out_63_port, 
                           input(62) => plus2A_out_62_port, input(61) => 
                           plus2A_out_61_port, input(60) => plus2A_out_60_port,
                           input(59) => plus2A_out_59_port, input(58) => 
                           plus2A_out_58_port, input(57) => plus2A_out_57_port,
                           input(56) => plus2A_out_56_port, input(55) => 
                           plus2A_out_55_port, input(54) => plus2A_out_54_port,
                           input(53) => plus2A_out_53_port, input(52) => 
                           plus2A_out_52_port, input(51) => plus2A_out_51_port,
                           input(50) => plus2A_out_50_port, input(49) => 
                           plus2A_out_49_port, input(48) => plus2A_out_48_port,
                           input(47) => plus2A_out_47_port, input(46) => 
                           plus2A_out_46_port, input(45) => plus2A_out_45_port,
                           input(44) => plus2A_out_44_port, input(43) => 
                           plus2A_out_43_port, input(42) => plus2A_out_42_port,
                           input(41) => plus2A_out_41_port, input(40) => 
                           plus2A_out_40_port, input(39) => plus2A_out_39_port,
                           input(38) => plus2A_out_38_port, input(37) => 
                           plus2A_out_37_port, input(36) => plus2A_out_36_port,
                           input(35) => plus2A_out_35_port, input(34) => 
                           plus2A_out_34_port, input(33) => plus2A_out_33_port,
                           input(32) => plus2A_out_32_port, input(31) => 
                           plus2A_out_31_port, input(30) => plus2A_out_30_port,
                           input(29) => plus2A_out_29_port, input(28) => 
                           plus2A_out_28_port, input(27) => plus2A_out_27_port,
                           input(26) => plus2A_out_26_port, input(25) => 
                           plus2A_out_25_port, input(24) => plus2A_out_24_port,
                           input(23) => plus2A_out_23_port, input(22) => 
                           plus2A_out_22_port, input(21) => plus2A_out_21_port,
                           input(20) => plus2A_out_20_port, input(19) => 
                           plus2A_out_19_port, input(18) => plus2A_out_18_port,
                           input(17) => plus2A_out_17_port, input(16) => 
                           plus2A_out_16_port, input(15) => plus2A_out_15_port,
                           input(14) => plus2A_out_14_port, input(13) => 
                           plus2A_out_13_port, input(12) => plus2A_out_12_port,
                           input(11) => plus2A_out_11_port, input(10) => 
                           plus2A_out_10_port, input(9) => plus2A_out_9_port, 
                           input(8) => plus2A_out_8_port, input(7) => 
                           plus2A_out_7_port, input(6) => plus2A_out_6_port, 
                           input(5) => plus2A_out_5_port, input(4) => 
                           plus2A_out_4_port, input(3) => plus2A_out_3_port, 
                           input(2) => plus2A_out_2_port, input(1) => 
                           plus2A_out_1_port, input(0) => plus2A_out_0_port, 
                           shiftLeftOnePos(63) => plus4A_out_63_port, 
                           shiftLeftOnePos(62) => plus4A_out_62_port, 
                           shiftLeftOnePos(61) => plus4A_out_61_port, 
                           shiftLeftOnePos(60) => plus4A_out_60_port, 
                           shiftLeftOnePos(59) => plus4A_out_59_port, 
                           shiftLeftOnePos(58) => plus4A_out_58_port, 
                           shiftLeftOnePos(57) => plus4A_out_57_port, 
                           shiftLeftOnePos(56) => plus4A_out_56_port, 
                           shiftLeftOnePos(55) => plus4A_out_55_port, 
                           shiftLeftOnePos(54) => plus4A_out_54_port, 
                           shiftLeftOnePos(53) => n5, shiftLeftOnePos(52) => n6
                           , shiftLeftOnePos(51) => plus4A_out_51_port, 
                           shiftLeftOnePos(50) => plus4A_out_50_port, 
                           shiftLeftOnePos(49) => plus4A_out_49_port, 
                           shiftLeftOnePos(48) => plus4A_out_48_port, 
                           shiftLeftOnePos(47) => plus4A_out_47_port, 
                           shiftLeftOnePos(46) => plus4A_out_46_port, 
                           shiftLeftOnePos(45) => plus4A_out_45_port, 
                           shiftLeftOnePos(44) => plus4A_out_44_port, 
                           shiftLeftOnePos(43) => plus4A_out_43_port, 
                           shiftLeftOnePos(42) => plus4A_out_42_port, 
                           shiftLeftOnePos(41) => plus4A_out_41_port, 
                           shiftLeftOnePos(40) => plus4A_out_40_port, 
                           shiftLeftOnePos(39) => plus4A_out_39_port, 
                           shiftLeftOnePos(38) => plus4A_out_38_port, 
                           shiftLeftOnePos(37) => plus4A_out_37_port, 
                           shiftLeftOnePos(36) => plus4A_out_36_port, 
                           shiftLeftOnePos(35) => plus4A_out_35_port, 
                           shiftLeftOnePos(34) => plus4A_out_34_port, 
                           shiftLeftOnePos(33) => plus4A_out_33_port, 
                           shiftLeftOnePos(32) => plus4A_out_32_port, 
                           shiftLeftOnePos(31) => plus4A_out_31_port, 
                           shiftLeftOnePos(30) => plus4A_out_30_port, 
                           shiftLeftOnePos(29) => plus4A_out_29_port, 
                           shiftLeftOnePos(28) => plus4A_out_28_port, 
                           shiftLeftOnePos(27) => plus4A_out_27_port, 
                           shiftLeftOnePos(26) => plus4A_out_26_port, 
                           shiftLeftOnePos(25) => plus4A_out_25_port, 
                           shiftLeftOnePos(24) => plus4A_out_24_port, 
                           shiftLeftOnePos(23) => plus4A_out_23_port, 
                           shiftLeftOnePos(22) => plus4A_out_22_port, 
                           shiftLeftOnePos(21) => plus4A_out_21_port, 
                           shiftLeftOnePos(20) => plus4A_out_20_port, 
                           shiftLeftOnePos(19) => plus4A_out_19_port, 
                           shiftLeftOnePos(18) => plus4A_out_18_port, 
                           shiftLeftOnePos(17) => plus4A_out_17_port, 
                           shiftLeftOnePos(16) => plus4A_out_16_port, 
                           shiftLeftOnePos(15) => plus4A_out_15_port, 
                           shiftLeftOnePos(14) => plus4A_out_14_port, 
                           shiftLeftOnePos(13) => plus4A_out_13_port, 
                           shiftLeftOnePos(12) => plus4A_out_12_port, 
                           shiftLeftOnePos(11) => plus4A_out_11_port, 
                           shiftLeftOnePos(10) => plus4A_out_10_port, 
                           shiftLeftOnePos(9) => plus4A_out_9_port, 
                           shiftLeftOnePos(8) => plus4A_out_8_port, 
                           shiftLeftOnePos(7) => plus4A_out_7_port, 
                           shiftLeftOnePos(6) => plus4A_out_6_port, 
                           shiftLeftOnePos(5) => plus4A_out_5_port, 
                           shiftLeftOnePos(4) => plus4A_out_4_port, 
                           shiftLeftOnePos(3) => plus4A_out_3_port, 
                           shiftLeftOnePos(2) => plus4A_out_2_port, 
                           shiftLeftOnePos(1) => plus4A_out_1_port, 
                           shiftLeftOnePos(0) => n_3157);
   complementer_1 : complementer_N64_14 port map( input(63) => 
                           plus2A_out_63_port, input(62) => plus2A_out_62_port,
                           input(61) => plus2A_out_61_port, input(60) => 
                           plus2A_out_60_port, input(59) => plus2A_out_59_port,
                           input(58) => plus2A_out_58_port, input(57) => 
                           plus2A_out_57_port, input(56) => plus2A_out_56_port,
                           input(55) => plus2A_out_55_port, input(54) => 
                           plus2A_out_54_port, input(53) => plus2A_out_53_port,
                           input(52) => plus2A_out_52_port, input(51) => 
                           plus2A_out_51_port, input(50) => plus2A_out_50_port,
                           input(49) => plus2A_out_49_port, input(48) => 
                           plus2A_out_48_port, input(47) => plus2A_out_47_port,
                           input(46) => plus2A_out_46_port, input(45) => 
                           plus2A_out_45_port, input(44) => plus2A_out_44_port,
                           input(43) => plus2A_out_43_port, input(42) => 
                           plus2A_out_42_port, input(41) => plus2A_out_41_port,
                           input(40) => plus2A_out_40_port, input(39) => 
                           plus2A_out_39_port, input(38) => plus2A_out_38_port,
                           input(37) => plus2A_out_37_port, input(36) => 
                           plus2A_out_36_port, input(35) => plus2A_out_35_port,
                           input(34) => plus2A_out_34_port, input(33) => 
                           plus2A_out_33_port, input(32) => plus2A_out_32_port,
                           input(31) => plus2A_out_31_port, input(30) => 
                           plus2A_out_30_port, input(29) => plus2A_out_29_port,
                           input(28) => plus2A_out_28_port, input(27) => 
                           plus2A_out_27_port, input(26) => plus2A_out_26_port,
                           input(25) => plus2A_out_25_port, input(24) => 
                           plus2A_out_24_port, input(23) => plus2A_out_23_port,
                           input(22) => plus2A_out_22_port, input(21) => 
                           plus2A_out_21_port, input(20) => plus2A_out_20_port,
                           input(19) => plus2A_out_19_port, input(18) => 
                           plus2A_out_18_port, input(17) => plus2A_out_17_port,
                           input(16) => plus2A_out_16_port, input(15) => 
                           plus2A_out_15_port, input(14) => plus2A_out_14_port,
                           input(13) => plus2A_out_13_port, input(12) => 
                           plus2A_out_12_port, input(11) => plus2A_out_11_port,
                           input(10) => plus2A_out_10_port, input(9) => 
                           plus2A_out_9_port, input(8) => plus2A_out_8_port, 
                           input(7) => plus2A_out_7_port, input(6) => 
                           plus2A_out_6_port, input(5) => plus2A_out_5_port, 
                           input(4) => plus2A_out_4_port, input(3) => 
                           plus2A_out_3_port, input(2) => plus2A_out_2_port, 
                           input(1) => plus2A_out_1_port, input(0) => 
                           plus2A_out_0_port, complement2(63) => 
                           minus2A_out(63), complement2(62) => minus2A_out(62),
                           complement2(61) => minus2A_out(61), complement2(60) 
                           => minus2A_out(60), complement2(59) => 
                           minus2A_out(59), complement2(58) => minus2A_out(58),
                           complement2(57) => minus2A_out(57), complement2(56) 
                           => minus2A_out(56), complement2(55) => 
                           minus2A_out(55), complement2(54) => minus2A_out(54),
                           complement2(53) => minus2A_out(53), complement2(52) 
                           => minus2A_out(52), complement2(51) => 
                           minus2A_out(51), complement2(50) => minus2A_out(50),
                           complement2(49) => minus2A_out(49), complement2(48) 
                           => minus2A_out(48), complement2(47) => 
                           minus2A_out(47), complement2(46) => minus2A_out(46),
                           complement2(45) => minus2A_out(45), complement2(44) 
                           => minus2A_out(44), complement2(43) => 
                           minus2A_out(43), complement2(42) => minus2A_out(42),
                           complement2(41) => minus2A_out(41), complement2(40) 
                           => minus2A_out(40), complement2(39) => 
                           minus2A_out(39), complement2(38) => minus2A_out(38),
                           complement2(37) => minus2A_out(37), complement2(36) 
                           => minus2A_out(36), complement2(35) => 
                           minus2A_out(35), complement2(34) => minus2A_out(34),
                           complement2(33) => minus2A_out(33), complement2(32) 
                           => minus2A_out(32), complement2(31) => 
                           minus2A_out(31), complement2(30) => minus2A_out(30),
                           complement2(29) => minus2A_out(29), complement2(28) 
                           => minus2A_out(28), complement2(27) => 
                           minus2A_out(27), complement2(26) => minus2A_out(26),
                           complement2(25) => minus2A_out(25), complement2(24) 
                           => minus2A_out(24), complement2(23) => 
                           minus2A_out(23), complement2(22) => minus2A_out(22),
                           complement2(21) => minus2A_out(21), complement2(20) 
                           => minus2A_out(20), complement2(19) => 
                           minus2A_out(19), complement2(18) => minus2A_out(18),
                           complement2(17) => minus2A_out(17), complement2(16) 
                           => minus2A_out(16), complement2(15) => 
                           minus2A_out(15), complement2(14) => minus2A_out(14),
                           complement2(13) => minus2A_out(13), complement2(12) 
                           => minus2A_out(12), complement2(11) => 
                           minus2A_out(11), complement2(10) => minus2A_out(10),
                           complement2(9) => minus2A_out(9), complement2(8) => 
                           minus2A_out(8), complement2(7) => minus2A_out(7), 
                           complement2(6) => minus2A_out(6), complement2(5) => 
                           minus2A_out(5), complement2(4) => minus2A_out(4), 
                           complement2(3) => minus2A_out(3), complement2(2) => 
                           minus2A_out(2), complement2(1) => minus2A_out(1), 
                           complement2(0) => minus2A_out(0));
   complementer_2 : complementer_N64_13 port map( input(63) => 
                           plus4A_out_63_port, input(62) => plus4A_out_62_port,
                           input(61) => plus4A_out_61_port, input(60) => 
                           plus4A_out_60_port, input(59) => plus4A_out_59_port,
                           input(58) => plus4A_out_58_port, input(57) => 
                           plus4A_out_57_port, input(56) => plus4A_out_56_port,
                           input(55) => plus4A_out_55_port, input(54) => 
                           plus4A_out_54_port, input(53) => plus4A_out_53_port,
                           input(52) => plus4A_out_52_port, input(51) => 
                           plus4A_out_51_port, input(50) => plus4A_out_50_port,
                           input(49) => plus4A_out_49_port, input(48) => 
                           plus4A_out_48_port, input(47) => plus4A_out_47_port,
                           input(46) => plus4A_out_46_port, input(45) => 
                           plus4A_out_45_port, input(44) => plus4A_out_44_port,
                           input(43) => plus4A_out_43_port, input(42) => 
                           plus4A_out_42_port, input(41) => plus4A_out_41_port,
                           input(40) => plus4A_out_40_port, input(39) => 
                           plus4A_out_39_port, input(38) => plus4A_out_38_port,
                           input(37) => plus4A_out_37_port, input(36) => 
                           plus4A_out_36_port, input(35) => plus4A_out_35_port,
                           input(34) => plus4A_out_34_port, input(33) => 
                           plus4A_out_33_port, input(32) => plus4A_out_32_port,
                           input(31) => plus4A_out_31_port, input(30) => 
                           plus4A_out_30_port, input(29) => plus4A_out_29_port,
                           input(28) => plus4A_out_28_port, input(27) => 
                           plus4A_out_27_port, input(26) => plus4A_out_26_port,
                           input(25) => plus4A_out_25_port, input(24) => 
                           plus4A_out_24_port, input(23) => plus4A_out_23_port,
                           input(22) => plus4A_out_22_port, input(21) => 
                           plus4A_out_21_port, input(20) => plus4A_out_20_port,
                           input(19) => plus4A_out_19_port, input(18) => 
                           plus4A_out_18_port, input(17) => plus4A_out_17_port,
                           input(16) => plus4A_out_16_port, input(15) => 
                           plus4A_out_15_port, input(14) => plus4A_out_14_port,
                           input(13) => plus4A_out_13_port, input(12) => 
                           plus4A_out_12_port, input(11) => plus4A_out_11_port,
                           input(10) => plus4A_out_10_port, input(9) => 
                           plus4A_out_9_port, input(8) => plus4A_out_8_port, 
                           input(7) => plus4A_out_7_port, input(6) => 
                           plus4A_out_6_port, input(5) => plus4A_out_5_port, 
                           input(4) => plus4A_out_4_port, input(3) => 
                           plus4A_out_3_port, input(2) => plus4A_out_2_port, 
                           input(1) => plus4A_out_1_port, input(0) => 
                           plus4A_out_0_port, complement2(63) => 
                           minus4A_out(63), complement2(62) => minus4A_out(62),
                           complement2(61) => minus4A_out(61), complement2(60) 
                           => minus4A_out(60), complement2(59) => 
                           minus4A_out(59), complement2(58) => minus4A_out(58),
                           complement2(57) => minus4A_out(57), complement2(56) 
                           => minus4A_out(56), complement2(55) => 
                           minus4A_out(55), complement2(54) => minus4A_out(54),
                           complement2(53) => minus4A_out(53), complement2(52) 
                           => minus4A_out(52), complement2(51) => 
                           minus4A_out(51), complement2(50) => minus4A_out(50),
                           complement2(49) => minus4A_out(49), complement2(48) 
                           => minus4A_out(48), complement2(47) => 
                           minus4A_out(47), complement2(46) => minus4A_out(46),
                           complement2(45) => minus4A_out(45), complement2(44) 
                           => minus4A_out(44), complement2(43) => 
                           minus4A_out(43), complement2(42) => minus4A_out(42),
                           complement2(41) => minus4A_out(41), complement2(40) 
                           => minus4A_out(40), complement2(39) => 
                           minus4A_out(39), complement2(38) => minus4A_out(38),
                           complement2(37) => minus4A_out(37), complement2(36) 
                           => minus4A_out(36), complement2(35) => 
                           minus4A_out(35), complement2(34) => minus4A_out(34),
                           complement2(33) => minus4A_out(33), complement2(32) 
                           => minus4A_out(32), complement2(31) => 
                           minus4A_out(31), complement2(30) => minus4A_out(30),
                           complement2(29) => minus4A_out(29), complement2(28) 
                           => minus4A_out(28), complement2(27) => 
                           minus4A_out(27), complement2(26) => minus4A_out(26),
                           complement2(25) => minus4A_out(25), complement2(24) 
                           => minus4A_out(24), complement2(23) => 
                           minus4A_out(23), complement2(22) => minus4A_out(22),
                           complement2(21) => minus4A_out(21), complement2(20) 
                           => minus4A_out(20), complement2(19) => 
                           minus4A_out(19), complement2(18) => minus4A_out(18),
                           complement2(17) => minus4A_out(17), complement2(16) 
                           => minus4A_out(16), complement2(15) => 
                           minus4A_out(15), complement2(14) => minus4A_out(14),
                           complement2(13) => minus4A_out(13), complement2(12) 
                           => minus4A_out(12), complement2(11) => 
                           minus4A_out(11), complement2(10) => minus4A_out(10),
                           complement2(9) => minus4A_out(9), complement2(8) => 
                           minus4A_out(8), complement2(7) => minus4A_out(7), 
                           complement2(6) => minus4A_out(6), complement2(5) => 
                           minus4A_out(5), complement2(4) => minus4A_out(4), 
                           complement2(3) => minus4A_out(3), complement2(2) => 
                           minus4A_out(2), complement2(1) => minus4A_out(1), 
                           complement2(0) => minus4A_out(0));
   U3 : BUF_X1 port map( A => n4, Z => plus2A_out_57_port);
   U4 : BUF_X1 port map( A => n6, Z => plus4A_out_52_port);
   U5 : BUF_X1 port map( A => n5, Z => plus4A_out_53_port);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity ShiftnCompl_N64_8 is

   port( plusA : in std_logic_vector (63 downto 0);  plus2A_out, minus2A_out, 
         plus4A_out, minus4A_out : out std_logic_vector (63 downto 0));

end ShiftnCompl_N64_8;

architecture SYN_struct of ShiftnCompl_N64_8 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component complementer_N64_15
      port( input : in std_logic_vector (63 downto 0);  complement2 : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component complementer_N64_16
      port( input : in std_logic_vector (63 downto 0);  complement2 : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component shifter_N64_15
      port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component shifter_N64_16
      port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
            std_logic_vector (63 downto 0));
   end component;
   
   signal plus2A_out_63_port, plus2A_out_62_port, plus2A_out_61_port, 
      plus2A_out_60_port, plus2A_out_59_port, plus2A_out_58_port, n37, 
      plus2A_out_56_port, plus2A_out_55_port, plus2A_out_54_port, 
      plus2A_out_53_port, plus2A_out_52_port, plus2A_out_51_port, 
      plus2A_out_50_port, plus2A_out_49_port, n38, n39, n40, plus2A_out_45_port
      , plus2A_out_44_port, plus2A_out_43_port, plus2A_out_42_port, 
      plus2A_out_41_port, plus2A_out_40_port, plus2A_out_39_port, 
      plus2A_out_38_port, plus2A_out_37_port, plus2A_out_36_port, 
      plus2A_out_35_port, plus2A_out_34_port, plus2A_out_33_port, 
      plus2A_out_32_port, plus2A_out_31_port, plus2A_out_30_port, 
      plus2A_out_29_port, plus2A_out_28_port, plus2A_out_27_port, 
      plus2A_out_26_port, plus2A_out_25_port, plus2A_out_24_port, 
      plus2A_out_23_port, plus2A_out_22_port, plus2A_out_21_port, 
      plus2A_out_20_port, plus2A_out_19_port, plus2A_out_18_port, 
      plus2A_out_17_port, plus2A_out_16_port, plus2A_out_15_port, 
      plus2A_out_14_port, plus2A_out_13_port, plus2A_out_12_port, 
      plus2A_out_11_port, plus2A_out_10_port, plus2A_out_9_port, 
      plus2A_out_8_port, plus2A_out_7_port, plus2A_out_6_port, 
      plus2A_out_5_port, plus2A_out_4_port, plus2A_out_3_port, 
      plus2A_out_2_port, plus2A_out_1_port, plus2A_out_0_port, 
      plus4A_out_63_port, plus4A_out_62_port, plus4A_out_61_port, 
      plus4A_out_60_port, plus4A_out_59_port, plus4A_out_58_port, 
      plus4A_out_57_port, plus4A_out_56_port, plus4A_out_55_port, 
      plus4A_out_54_port, n41, n42, plus4A_out_51_port, plus4A_out_50_port, 
      plus4A_out_49_port, plus4A_out_48_port, plus4A_out_47_port, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, 
      plus4A_out_16_port, plus4A_out_15_port, plus4A_out_14_port, 
      plus4A_out_13_port, plus4A_out_12_port, plus4A_out_11_port, 
      plus4A_out_10_port, plus4A_out_9_port, plus4A_out_8_port, 
      plus4A_out_7_port, plus4A_out_6_port, plus4A_out_5_port, 
      plus4A_out_4_port, plus4A_out_3_port, plus4A_out_2_port, 
      plus4A_out_1_port, plus4A_out_0_port, plus4A_out_17_port, 
      plus4A_out_18_port, plus4A_out_19_port, plus4A_out_20_port, 
      plus4A_out_21_port, plus4A_out_22_port, plus4A_out_23_port, 
      plus4A_out_24_port, plus4A_out_25_port, plus4A_out_26_port, 
      plus4A_out_27_port, plus4A_out_28_port, plus4A_out_29_port, 
      plus4A_out_30_port, plus4A_out_31_port, plus4A_out_32_port, 
      plus4A_out_33_port, plus4A_out_34_port, plus4A_out_35_port, 
      plus4A_out_36_port, plus4A_out_37_port, plus4A_out_38_port, 
      plus4A_out_39_port, plus4A_out_40_port, plus4A_out_41_port, 
      plus4A_out_42_port, plus4A_out_43_port, plus4A_out_44_port, 
      plus4A_out_45_port, plus4A_out_46_port, plus2A_out_46_port, 
      plus2A_out_47_port, plus2A_out_48_port, plus4A_out_52_port, 
      plus4A_out_53_port, plus2A_out_57_port, n_3158, n_3159 : std_logic;

begin
   plus2A_out <= ( plus2A_out_63_port, plus2A_out_62_port, plus2A_out_61_port, 
      plus2A_out_60_port, plus2A_out_59_port, plus2A_out_58_port, 
      plus2A_out_57_port, plus2A_out_56_port, plus2A_out_55_port, 
      plus2A_out_54_port, plus2A_out_53_port, plus2A_out_52_port, 
      plus2A_out_51_port, plus2A_out_50_port, plus2A_out_49_port, 
      plus2A_out_48_port, plus2A_out_47_port, plus2A_out_46_port, 
      plus2A_out_45_port, plus2A_out_44_port, plus2A_out_43_port, 
      plus2A_out_42_port, plus2A_out_41_port, plus2A_out_40_port, 
      plus2A_out_39_port, plus2A_out_38_port, plus2A_out_37_port, 
      plus2A_out_36_port, plus2A_out_35_port, plus2A_out_34_port, 
      plus2A_out_33_port, plus2A_out_32_port, plus2A_out_31_port, 
      plus2A_out_30_port, plus2A_out_29_port, plus2A_out_28_port, 
      plus2A_out_27_port, plus2A_out_26_port, plus2A_out_25_port, 
      plus2A_out_24_port, plus2A_out_23_port, plus2A_out_22_port, 
      plus2A_out_21_port, plus2A_out_20_port, plus2A_out_19_port, 
      plus2A_out_18_port, plus2A_out_17_port, plus2A_out_16_port, 
      plus2A_out_15_port, plus2A_out_14_port, plus2A_out_13_port, 
      plus2A_out_12_port, plus2A_out_11_port, plus2A_out_10_port, 
      plus2A_out_9_port, plus2A_out_8_port, plus2A_out_7_port, 
      plus2A_out_6_port, plus2A_out_5_port, plus2A_out_4_port, 
      plus2A_out_3_port, plus2A_out_2_port, plus2A_out_1_port, 
      plus2A_out_0_port );
   plus4A_out <= ( plus4A_out_63_port, plus4A_out_62_port, plus4A_out_61_port, 
      plus4A_out_60_port, plus4A_out_59_port, plus4A_out_58_port, 
      plus4A_out_57_port, plus4A_out_56_port, plus4A_out_55_port, 
      plus4A_out_54_port, plus4A_out_53_port, plus4A_out_52_port, 
      plus4A_out_51_port, plus4A_out_50_port, plus4A_out_49_port, 
      plus4A_out_48_port, plus4A_out_47_port, plus4A_out_46_port, 
      plus4A_out_45_port, plus4A_out_44_port, plus4A_out_43_port, 
      plus4A_out_42_port, plus4A_out_41_port, plus4A_out_40_port, 
      plus4A_out_39_port, plus4A_out_38_port, plus4A_out_37_port, 
      plus4A_out_36_port, plus4A_out_35_port, plus4A_out_34_port, 
      plus4A_out_33_port, plus4A_out_32_port, plus4A_out_31_port, 
      plus4A_out_30_port, plus4A_out_29_port, plus4A_out_28_port, 
      plus4A_out_27_port, plus4A_out_26_port, plus4A_out_25_port, 
      plus4A_out_24_port, plus4A_out_23_port, plus4A_out_22_port, 
      plus4A_out_21_port, plus4A_out_20_port, plus4A_out_19_port, 
      plus4A_out_18_port, plus4A_out_17_port, plus4A_out_16_port, 
      plus4A_out_15_port, plus4A_out_14_port, plus4A_out_13_port, 
      plus4A_out_12_port, plus4A_out_11_port, plus4A_out_10_port, 
      plus4A_out_9_port, plus4A_out_8_port, plus4A_out_7_port, 
      plus4A_out_6_port, plus4A_out_5_port, plus4A_out_4_port, 
      plus4A_out_3_port, plus4A_out_2_port, plus4A_out_1_port, 
      plus4A_out_0_port );
   
   plus2A_out_0_port <= '0';
   plus4A_out_0_port <= '0';
   shifter_1 : shifter_N64_16 port map( input(63) => plusA(63), input(62) => 
                           plusA(62), input(61) => plusA(61), input(60) => 
                           plusA(60), input(59) => plusA(59), input(58) => 
                           plusA(58), input(57) => plusA(57), input(56) => 
                           plusA(56), input(55) => plusA(55), input(54) => 
                           plusA(54), input(53) => plusA(53), input(52) => 
                           plusA(52), input(51) => plusA(51), input(50) => 
                           plusA(50), input(49) => plusA(49), input(48) => 
                           plusA(48), input(47) => plusA(47), input(46) => 
                           plusA(46), input(45) => plusA(45), input(44) => 
                           plusA(44), input(43) => plusA(43), input(42) => 
                           plusA(42), input(41) => plusA(41), input(40) => 
                           plusA(40), input(39) => plusA(39), input(38) => 
                           plusA(38), input(37) => plusA(37), input(36) => 
                           plusA(36), input(35) => plusA(35), input(34) => 
                           plusA(34), input(33) => plusA(33), input(32) => 
                           plusA(32), input(31) => plusA(31), input(30) => 
                           plusA(30), input(29) => plusA(29), input(28) => 
                           plusA(28), input(27) => plusA(27), input(26) => 
                           plusA(26), input(25) => plusA(25), input(24) => 
                           plusA(24), input(23) => plusA(23), input(22) => 
                           plusA(22), input(21) => plusA(21), input(20) => 
                           plusA(20), input(19) => plusA(19), input(18) => 
                           plusA(18), input(17) => plusA(17), input(16) => 
                           plusA(16), input(15) => plusA(15), input(14) => 
                           plusA(14), input(13) => plusA(13), input(12) => 
                           plusA(12), input(11) => plusA(11), input(10) => 
                           plusA(10), input(9) => plusA(9), input(8) => 
                           plusA(8), input(7) => plusA(7), input(6) => plusA(6)
                           , input(5) => plusA(5), input(4) => plusA(4), 
                           input(3) => plusA(3), input(2) => plusA(2), input(1)
                           => plusA(1), input(0) => plusA(0), 
                           shiftLeftOnePos(63) => plus2A_out_63_port, 
                           shiftLeftOnePos(62) => plus2A_out_62_port, 
                           shiftLeftOnePos(61) => plus2A_out_61_port, 
                           shiftLeftOnePos(60) => plus2A_out_60_port, 
                           shiftLeftOnePos(59) => plus2A_out_59_port, 
                           shiftLeftOnePos(58) => plus2A_out_58_port, 
                           shiftLeftOnePos(57) => n37, shiftLeftOnePos(56) => 
                           plus2A_out_56_port, shiftLeftOnePos(55) => 
                           plus2A_out_55_port, shiftLeftOnePos(54) => 
                           plus2A_out_54_port, shiftLeftOnePos(53) => 
                           plus2A_out_53_port, shiftLeftOnePos(52) => 
                           plus2A_out_52_port, shiftLeftOnePos(51) => 
                           plus2A_out_51_port, shiftLeftOnePos(50) => 
                           plus2A_out_50_port, shiftLeftOnePos(49) => 
                           plus2A_out_49_port, shiftLeftOnePos(48) => n38, 
                           shiftLeftOnePos(47) => n39, shiftLeftOnePos(46) => 
                           n40, shiftLeftOnePos(45) => plus2A_out_45_port, 
                           shiftLeftOnePos(44) => plus2A_out_44_port, 
                           shiftLeftOnePos(43) => plus2A_out_43_port, 
                           shiftLeftOnePos(42) => plus2A_out_42_port, 
                           shiftLeftOnePos(41) => plus2A_out_41_port, 
                           shiftLeftOnePos(40) => plus2A_out_40_port, 
                           shiftLeftOnePos(39) => plus2A_out_39_port, 
                           shiftLeftOnePos(38) => plus2A_out_38_port, 
                           shiftLeftOnePos(37) => plus2A_out_37_port, 
                           shiftLeftOnePos(36) => plus2A_out_36_port, 
                           shiftLeftOnePos(35) => plus2A_out_35_port, 
                           shiftLeftOnePos(34) => plus2A_out_34_port, 
                           shiftLeftOnePos(33) => plus2A_out_33_port, 
                           shiftLeftOnePos(32) => plus2A_out_32_port, 
                           shiftLeftOnePos(31) => plus2A_out_31_port, 
                           shiftLeftOnePos(30) => plus2A_out_30_port, 
                           shiftLeftOnePos(29) => plus2A_out_29_port, 
                           shiftLeftOnePos(28) => plus2A_out_28_port, 
                           shiftLeftOnePos(27) => plus2A_out_27_port, 
                           shiftLeftOnePos(26) => plus2A_out_26_port, 
                           shiftLeftOnePos(25) => plus2A_out_25_port, 
                           shiftLeftOnePos(24) => plus2A_out_24_port, 
                           shiftLeftOnePos(23) => plus2A_out_23_port, 
                           shiftLeftOnePos(22) => plus2A_out_22_port, 
                           shiftLeftOnePos(21) => plus2A_out_21_port, 
                           shiftLeftOnePos(20) => plus2A_out_20_port, 
                           shiftLeftOnePos(19) => plus2A_out_19_port, 
                           shiftLeftOnePos(18) => plus2A_out_18_port, 
                           shiftLeftOnePos(17) => plus2A_out_17_port, 
                           shiftLeftOnePos(16) => plus2A_out_16_port, 
                           shiftLeftOnePos(15) => plus2A_out_15_port, 
                           shiftLeftOnePos(14) => plus2A_out_14_port, 
                           shiftLeftOnePos(13) => plus2A_out_13_port, 
                           shiftLeftOnePos(12) => plus2A_out_12_port, 
                           shiftLeftOnePos(11) => plus2A_out_11_port, 
                           shiftLeftOnePos(10) => plus2A_out_10_port, 
                           shiftLeftOnePos(9) => plus2A_out_9_port, 
                           shiftLeftOnePos(8) => plus2A_out_8_port, 
                           shiftLeftOnePos(7) => plus2A_out_7_port, 
                           shiftLeftOnePos(6) => plus2A_out_6_port, 
                           shiftLeftOnePos(5) => plus2A_out_5_port, 
                           shiftLeftOnePos(4) => plus2A_out_4_port, 
                           shiftLeftOnePos(3) => plus2A_out_3_port, 
                           shiftLeftOnePos(2) => plus2A_out_2_port, 
                           shiftLeftOnePos(1) => plus2A_out_1_port, 
                           shiftLeftOnePos(0) => n_3158);
   shifter_2 : shifter_N64_15 port map( input(63) => plus2A_out_63_port, 
                           input(62) => plus2A_out_62_port, input(61) => 
                           plus2A_out_61_port, input(60) => plus2A_out_60_port,
                           input(59) => plus2A_out_59_port, input(58) => 
                           plus2A_out_58_port, input(57) => plus2A_out_57_port,
                           input(56) => plus2A_out_56_port, input(55) => 
                           plus2A_out_55_port, input(54) => plus2A_out_54_port,
                           input(53) => plus2A_out_53_port, input(52) => 
                           plus2A_out_52_port, input(51) => plus2A_out_51_port,
                           input(50) => plus2A_out_50_port, input(49) => 
                           plus2A_out_49_port, input(48) => plus2A_out_48_port,
                           input(47) => plus2A_out_47_port, input(46) => 
                           plus2A_out_46_port, input(45) => plus2A_out_45_port,
                           input(44) => plus2A_out_44_port, input(43) => 
                           plus2A_out_43_port, input(42) => plus2A_out_42_port,
                           input(41) => plus2A_out_41_port, input(40) => 
                           plus2A_out_40_port, input(39) => plus2A_out_39_port,
                           input(38) => plus2A_out_38_port, input(37) => 
                           plus2A_out_37_port, input(36) => plus2A_out_36_port,
                           input(35) => plus2A_out_35_port, input(34) => 
                           plus2A_out_34_port, input(33) => plus2A_out_33_port,
                           input(32) => plus2A_out_32_port, input(31) => 
                           plus2A_out_31_port, input(30) => plus2A_out_30_port,
                           input(29) => plus2A_out_29_port, input(28) => 
                           plus2A_out_28_port, input(27) => plus2A_out_27_port,
                           input(26) => plus2A_out_26_port, input(25) => 
                           plus2A_out_25_port, input(24) => plus2A_out_24_port,
                           input(23) => plus2A_out_23_port, input(22) => 
                           plus2A_out_22_port, input(21) => plus2A_out_21_port,
                           input(20) => plus2A_out_20_port, input(19) => 
                           plus2A_out_19_port, input(18) => plus2A_out_18_port,
                           input(17) => plus2A_out_17_port, input(16) => 
                           plus2A_out_16_port, input(15) => plus2A_out_15_port,
                           input(14) => plus2A_out_14_port, input(13) => 
                           plus2A_out_13_port, input(12) => plus2A_out_12_port,
                           input(11) => plus2A_out_11_port, input(10) => 
                           plus2A_out_10_port, input(9) => plus2A_out_9_port, 
                           input(8) => plus2A_out_8_port, input(7) => 
                           plus2A_out_7_port, input(6) => plus2A_out_6_port, 
                           input(5) => plus2A_out_5_port, input(4) => 
                           plus2A_out_4_port, input(3) => plus2A_out_3_port, 
                           input(2) => plus2A_out_2_port, input(1) => 
                           plus2A_out_1_port, input(0) => plus2A_out_0_port, 
                           shiftLeftOnePos(63) => plus4A_out_63_port, 
                           shiftLeftOnePos(62) => plus4A_out_62_port, 
                           shiftLeftOnePos(61) => plus4A_out_61_port, 
                           shiftLeftOnePos(60) => plus4A_out_60_port, 
                           shiftLeftOnePos(59) => plus4A_out_59_port, 
                           shiftLeftOnePos(58) => plus4A_out_58_port, 
                           shiftLeftOnePos(57) => plus4A_out_57_port, 
                           shiftLeftOnePos(56) => plus4A_out_56_port, 
                           shiftLeftOnePos(55) => plus4A_out_55_port, 
                           shiftLeftOnePos(54) => plus4A_out_54_port, 
                           shiftLeftOnePos(53) => n41, shiftLeftOnePos(52) => 
                           n42, shiftLeftOnePos(51) => plus4A_out_51_port, 
                           shiftLeftOnePos(50) => plus4A_out_50_port, 
                           shiftLeftOnePos(49) => plus4A_out_49_port, 
                           shiftLeftOnePos(48) => plus4A_out_48_port, 
                           shiftLeftOnePos(47) => plus4A_out_47_port, 
                           shiftLeftOnePos(46) => n43, shiftLeftOnePos(45) => 
                           n44, shiftLeftOnePos(44) => n45, shiftLeftOnePos(43)
                           => n46, shiftLeftOnePos(42) => n47, 
                           shiftLeftOnePos(41) => n48, shiftLeftOnePos(40) => 
                           n49, shiftLeftOnePos(39) => n50, shiftLeftOnePos(38)
                           => n51, shiftLeftOnePos(37) => n52, 
                           shiftLeftOnePos(36) => n53, shiftLeftOnePos(35) => 
                           n54, shiftLeftOnePos(34) => n55, shiftLeftOnePos(33)
                           => n56, shiftLeftOnePos(32) => n57, 
                           shiftLeftOnePos(31) => n58, shiftLeftOnePos(30) => 
                           n59, shiftLeftOnePos(29) => n60, shiftLeftOnePos(28)
                           => n61, shiftLeftOnePos(27) => n62, 
                           shiftLeftOnePos(26) => n63, shiftLeftOnePos(25) => 
                           n64, shiftLeftOnePos(24) => n65, shiftLeftOnePos(23)
                           => n66, shiftLeftOnePos(22) => n67, 
                           shiftLeftOnePos(21) => n68, shiftLeftOnePos(20) => 
                           n69, shiftLeftOnePos(19) => n70, shiftLeftOnePos(18)
                           => n71, shiftLeftOnePos(17) => n72, 
                           shiftLeftOnePos(16) => plus4A_out_16_port, 
                           shiftLeftOnePos(15) => plus4A_out_15_port, 
                           shiftLeftOnePos(14) => plus4A_out_14_port, 
                           shiftLeftOnePos(13) => plus4A_out_13_port, 
                           shiftLeftOnePos(12) => plus4A_out_12_port, 
                           shiftLeftOnePos(11) => plus4A_out_11_port, 
                           shiftLeftOnePos(10) => plus4A_out_10_port, 
                           shiftLeftOnePos(9) => plus4A_out_9_port, 
                           shiftLeftOnePos(8) => plus4A_out_8_port, 
                           shiftLeftOnePos(7) => plus4A_out_7_port, 
                           shiftLeftOnePos(6) => plus4A_out_6_port, 
                           shiftLeftOnePos(5) => plus4A_out_5_port, 
                           shiftLeftOnePos(4) => plus4A_out_4_port, 
                           shiftLeftOnePos(3) => plus4A_out_3_port, 
                           shiftLeftOnePos(2) => plus4A_out_2_port, 
                           shiftLeftOnePos(1) => plus4A_out_1_port, 
                           shiftLeftOnePos(0) => n_3159);
   complementer_1 : complementer_N64_16 port map( input(63) => 
                           plus2A_out_63_port, input(62) => plus2A_out_62_port,
                           input(61) => plus2A_out_61_port, input(60) => 
                           plus2A_out_60_port, input(59) => plus2A_out_59_port,
                           input(58) => plus2A_out_58_port, input(57) => 
                           plus2A_out_57_port, input(56) => plus2A_out_56_port,
                           input(55) => plus2A_out_55_port, input(54) => 
                           plus2A_out_54_port, input(53) => plus2A_out_53_port,
                           input(52) => plus2A_out_52_port, input(51) => 
                           plus2A_out_51_port, input(50) => plus2A_out_50_port,
                           input(49) => plus2A_out_49_port, input(48) => 
                           plus2A_out_48_port, input(47) => plus2A_out_47_port,
                           input(46) => plus2A_out_46_port, input(45) => 
                           plus2A_out_45_port, input(44) => plus2A_out_44_port,
                           input(43) => plus2A_out_43_port, input(42) => 
                           plus2A_out_42_port, input(41) => plus2A_out_41_port,
                           input(40) => plus2A_out_40_port, input(39) => 
                           plus2A_out_39_port, input(38) => plus2A_out_38_port,
                           input(37) => plus2A_out_37_port, input(36) => 
                           plus2A_out_36_port, input(35) => plus2A_out_35_port,
                           input(34) => plus2A_out_34_port, input(33) => 
                           plus2A_out_33_port, input(32) => plus2A_out_32_port,
                           input(31) => plus2A_out_31_port, input(30) => 
                           plus2A_out_30_port, input(29) => plus2A_out_29_port,
                           input(28) => plus2A_out_28_port, input(27) => 
                           plus2A_out_27_port, input(26) => plus2A_out_26_port,
                           input(25) => plus2A_out_25_port, input(24) => 
                           plus2A_out_24_port, input(23) => plus2A_out_23_port,
                           input(22) => plus2A_out_22_port, input(21) => 
                           plus2A_out_21_port, input(20) => plus2A_out_20_port,
                           input(19) => plus2A_out_19_port, input(18) => 
                           plus2A_out_18_port, input(17) => plus2A_out_17_port,
                           input(16) => plus2A_out_16_port, input(15) => 
                           plus2A_out_15_port, input(14) => plus2A_out_14_port,
                           input(13) => plus2A_out_13_port, input(12) => 
                           plus2A_out_12_port, input(11) => plus2A_out_11_port,
                           input(10) => plus2A_out_10_port, input(9) => 
                           plus2A_out_9_port, input(8) => plus2A_out_8_port, 
                           input(7) => plus2A_out_7_port, input(6) => 
                           plus2A_out_6_port, input(5) => plus2A_out_5_port, 
                           input(4) => plus2A_out_4_port, input(3) => 
                           plus2A_out_3_port, input(2) => plus2A_out_2_port, 
                           input(1) => plus2A_out_1_port, input(0) => 
                           plus2A_out_0_port, complement2(63) => 
                           minus2A_out(63), complement2(62) => minus2A_out(62),
                           complement2(61) => minus2A_out(61), complement2(60) 
                           => minus2A_out(60), complement2(59) => 
                           minus2A_out(59), complement2(58) => minus2A_out(58),
                           complement2(57) => minus2A_out(57), complement2(56) 
                           => minus2A_out(56), complement2(55) => 
                           minus2A_out(55), complement2(54) => minus2A_out(54),
                           complement2(53) => minus2A_out(53), complement2(52) 
                           => minus2A_out(52), complement2(51) => 
                           minus2A_out(51), complement2(50) => minus2A_out(50),
                           complement2(49) => minus2A_out(49), complement2(48) 
                           => minus2A_out(48), complement2(47) => 
                           minus2A_out(47), complement2(46) => minus2A_out(46),
                           complement2(45) => minus2A_out(45), complement2(44) 
                           => minus2A_out(44), complement2(43) => 
                           minus2A_out(43), complement2(42) => minus2A_out(42),
                           complement2(41) => minus2A_out(41), complement2(40) 
                           => minus2A_out(40), complement2(39) => 
                           minus2A_out(39), complement2(38) => minus2A_out(38),
                           complement2(37) => minus2A_out(37), complement2(36) 
                           => minus2A_out(36), complement2(35) => 
                           minus2A_out(35), complement2(34) => minus2A_out(34),
                           complement2(33) => minus2A_out(33), complement2(32) 
                           => minus2A_out(32), complement2(31) => 
                           minus2A_out(31), complement2(30) => minus2A_out(30),
                           complement2(29) => minus2A_out(29), complement2(28) 
                           => minus2A_out(28), complement2(27) => 
                           minus2A_out(27), complement2(26) => minus2A_out(26),
                           complement2(25) => minus2A_out(25), complement2(24) 
                           => minus2A_out(24), complement2(23) => 
                           minus2A_out(23), complement2(22) => minus2A_out(22),
                           complement2(21) => minus2A_out(21), complement2(20) 
                           => minus2A_out(20), complement2(19) => 
                           minus2A_out(19), complement2(18) => minus2A_out(18),
                           complement2(17) => minus2A_out(17), complement2(16) 
                           => minus2A_out(16), complement2(15) => 
                           minus2A_out(15), complement2(14) => minus2A_out(14),
                           complement2(13) => minus2A_out(13), complement2(12) 
                           => minus2A_out(12), complement2(11) => 
                           minus2A_out(11), complement2(10) => minus2A_out(10),
                           complement2(9) => minus2A_out(9), complement2(8) => 
                           minus2A_out(8), complement2(7) => minus2A_out(7), 
                           complement2(6) => minus2A_out(6), complement2(5) => 
                           minus2A_out(5), complement2(4) => minus2A_out(4), 
                           complement2(3) => minus2A_out(3), complement2(2) => 
                           minus2A_out(2), complement2(1) => minus2A_out(1), 
                           complement2(0) => minus2A_out(0));
   complementer_2 : complementer_N64_15 port map( input(63) => 
                           plus4A_out_63_port, input(62) => plus4A_out_62_port,
                           input(61) => plus4A_out_61_port, input(60) => 
                           plus4A_out_60_port, input(59) => plus4A_out_59_port,
                           input(58) => plus4A_out_58_port, input(57) => 
                           plus4A_out_57_port, input(56) => plus4A_out_56_port,
                           input(55) => plus4A_out_55_port, input(54) => 
                           plus4A_out_54_port, input(53) => plus4A_out_53_port,
                           input(52) => plus4A_out_52_port, input(51) => 
                           plus4A_out_51_port, input(50) => plus4A_out_50_port,
                           input(49) => plus4A_out_49_port, input(48) => 
                           plus4A_out_48_port, input(47) => plus4A_out_47_port,
                           input(46) => plus4A_out_46_port, input(45) => 
                           plus4A_out_45_port, input(44) => plus4A_out_44_port,
                           input(43) => plus4A_out_43_port, input(42) => 
                           plus4A_out_42_port, input(41) => plus4A_out_41_port,
                           input(40) => plus4A_out_40_port, input(39) => 
                           plus4A_out_39_port, input(38) => plus4A_out_38_port,
                           input(37) => plus4A_out_37_port, input(36) => 
                           plus4A_out_36_port, input(35) => plus4A_out_35_port,
                           input(34) => plus4A_out_34_port, input(33) => 
                           plus4A_out_33_port, input(32) => plus4A_out_32_port,
                           input(31) => plus4A_out_31_port, input(30) => 
                           plus4A_out_30_port, input(29) => plus4A_out_29_port,
                           input(28) => plus4A_out_28_port, input(27) => 
                           plus4A_out_27_port, input(26) => plus4A_out_26_port,
                           input(25) => plus4A_out_25_port, input(24) => 
                           plus4A_out_24_port, input(23) => plus4A_out_23_port,
                           input(22) => plus4A_out_22_port, input(21) => 
                           plus4A_out_21_port, input(20) => plus4A_out_20_port,
                           input(19) => plus4A_out_19_port, input(18) => 
                           plus4A_out_18_port, input(17) => plus4A_out_17_port,
                           input(16) => plus4A_out_16_port, input(15) => 
                           plus4A_out_15_port, input(14) => plus4A_out_14_port,
                           input(13) => plus4A_out_13_port, input(12) => 
                           plus4A_out_12_port, input(11) => plus4A_out_11_port,
                           input(10) => plus4A_out_10_port, input(9) => 
                           plus4A_out_9_port, input(8) => plus4A_out_8_port, 
                           input(7) => plus4A_out_7_port, input(6) => 
                           plus4A_out_6_port, input(5) => plus4A_out_5_port, 
                           input(4) => plus4A_out_4_port, input(3) => 
                           plus4A_out_3_port, input(2) => plus4A_out_2_port, 
                           input(1) => plus4A_out_1_port, input(0) => 
                           plus4A_out_0_port, complement2(63) => 
                           minus4A_out(63), complement2(62) => minus4A_out(62),
                           complement2(61) => minus4A_out(61), complement2(60) 
                           => minus4A_out(60), complement2(59) => 
                           minus4A_out(59), complement2(58) => minus4A_out(58),
                           complement2(57) => minus4A_out(57), complement2(56) 
                           => minus4A_out(56), complement2(55) => 
                           minus4A_out(55), complement2(54) => minus4A_out(54),
                           complement2(53) => minus4A_out(53), complement2(52) 
                           => minus4A_out(52), complement2(51) => 
                           minus4A_out(51), complement2(50) => minus4A_out(50),
                           complement2(49) => minus4A_out(49), complement2(48) 
                           => minus4A_out(48), complement2(47) => 
                           minus4A_out(47), complement2(46) => minus4A_out(46),
                           complement2(45) => minus4A_out(45), complement2(44) 
                           => minus4A_out(44), complement2(43) => 
                           minus4A_out(43), complement2(42) => minus4A_out(42),
                           complement2(41) => minus4A_out(41), complement2(40) 
                           => minus4A_out(40), complement2(39) => 
                           minus4A_out(39), complement2(38) => minus4A_out(38),
                           complement2(37) => minus4A_out(37), complement2(36) 
                           => minus4A_out(36), complement2(35) => 
                           minus4A_out(35), complement2(34) => minus4A_out(34),
                           complement2(33) => minus4A_out(33), complement2(32) 
                           => minus4A_out(32), complement2(31) => 
                           minus4A_out(31), complement2(30) => minus4A_out(30),
                           complement2(29) => minus4A_out(29), complement2(28) 
                           => minus4A_out(28), complement2(27) => 
                           minus4A_out(27), complement2(26) => minus4A_out(26),
                           complement2(25) => minus4A_out(25), complement2(24) 
                           => minus4A_out(24), complement2(23) => 
                           minus4A_out(23), complement2(22) => minus4A_out(22),
                           complement2(21) => minus4A_out(21), complement2(20) 
                           => minus4A_out(20), complement2(19) => 
                           minus4A_out(19), complement2(18) => minus4A_out(18),
                           complement2(17) => minus4A_out(17), complement2(16) 
                           => minus4A_out(16), complement2(15) => 
                           minus4A_out(15), complement2(14) => minus4A_out(14),
                           complement2(13) => minus4A_out(13), complement2(12) 
                           => minus4A_out(12), complement2(11) => 
                           minus4A_out(11), complement2(10) => minus4A_out(10),
                           complement2(9) => minus4A_out(9), complement2(8) => 
                           minus4A_out(8), complement2(7) => minus4A_out(7), 
                           complement2(6) => minus4A_out(6), complement2(5) => 
                           minus4A_out(5), complement2(4) => minus4A_out(4), 
                           complement2(3) => minus4A_out(3), complement2(2) => 
                           minus4A_out(2), complement2(1) => minus4A_out(1), 
                           complement2(0) => minus4A_out(0));
   U3 : BUF_X1 port map( A => n50, Z => plus4A_out_39_port);
   U4 : BUF_X1 port map( A => n54, Z => plus4A_out_35_port);
   U5 : BUF_X1 port map( A => n58, Z => plus4A_out_31_port);
   U6 : BUF_X1 port map( A => n52, Z => plus4A_out_37_port);
   U7 : BUF_X1 port map( A => n56, Z => plus4A_out_33_port);
   U8 : BUF_X1 port map( A => n55, Z => plus4A_out_34_port);
   U9 : BUF_X1 port map( A => n57, Z => plus4A_out_32_port);
   U10 : BUF_X1 port map( A => n39, Z => plus2A_out_47_port);
   U11 : BUF_X1 port map( A => n46, Z => plus4A_out_43_port);
   U12 : BUF_X1 port map( A => n44, Z => plus4A_out_45_port);
   U13 : BUF_X1 port map( A => n48, Z => plus4A_out_41_port);
   U14 : BUF_X1 port map( A => n43, Z => plus4A_out_46_port);
   U15 : BUF_X1 port map( A => n47, Z => plus4A_out_42_port);
   U16 : BUF_X1 port map( A => n38, Z => plus2A_out_48_port);
   U17 : BUF_X1 port map( A => n45, Z => plus4A_out_44_port);
   U18 : BUF_X1 port map( A => n40, Z => plus2A_out_46_port);
   U19 : BUF_X1 port map( A => n37, Z => plus2A_out_57_port);
   U20 : BUF_X1 port map( A => n42, Z => plus4A_out_52_port);
   U21 : BUF_X1 port map( A => n41, Z => plus4A_out_53_port);
   U22 : BUF_X1 port map( A => n70, Z => plus4A_out_19_port);
   U23 : BUF_X1 port map( A => n72, Z => plus4A_out_17_port);
   U24 : BUF_X1 port map( A => n71, Z => plus4A_out_18_port);
   U25 : BUF_X1 port map( A => n62, Z => plus4A_out_27_port);
   U26 : BUF_X1 port map( A => n66, Z => plus4A_out_23_port);
   U27 : BUF_X1 port map( A => n60, Z => plus4A_out_29_port);
   U28 : BUF_X1 port map( A => n64, Z => plus4A_out_25_port);
   U29 : BUF_X1 port map( A => n68, Z => plus4A_out_21_port);
   U30 : BUF_X1 port map( A => n61, Z => plus4A_out_28_port);
   U31 : BUF_X1 port map( A => n65, Z => plus4A_out_24_port);
   U32 : BUF_X1 port map( A => n69, Z => plus4A_out_20_port);
   U33 : BUF_X1 port map( A => n59, Z => plus4A_out_30_port);
   U34 : BUF_X1 port map( A => n63, Z => plus4A_out_26_port);
   U35 : BUF_X1 port map( A => n67, Z => plus4A_out_22_port);
   U36 : BUF_X1 port map( A => n49, Z => plus4A_out_40_port);
   U37 : BUF_X1 port map( A => n53, Z => plus4A_out_36_port);
   U38 : BUF_X1 port map( A => n51, Z => plus4A_out_38_port);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity ShiftnCompl_N64_9 is

   port( plusA : in std_logic_vector (63 downto 0);  plus2A_out, minus2A_out, 
         plus4A_out, minus4A_out : out std_logic_vector (63 downto 0));

end ShiftnCompl_N64_9;

architecture SYN_struct of ShiftnCompl_N64_9 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component complementer_N64_17
      port( input : in std_logic_vector (63 downto 0);  complement2 : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component complementer_N64_18
      port( input : in std_logic_vector (63 downto 0);  complement2 : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component shifter_N64_17
      port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component shifter_N64_18
      port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
            std_logic_vector (63 downto 0));
   end component;
   
   signal plus2A_out_63_port, plus2A_out_62_port, plus2A_out_61_port, 
      plus2A_out_60_port, plus2A_out_59_port, plus2A_out_58_port, n6, 
      plus2A_out_56_port, plus2A_out_55_port, plus2A_out_54_port, 
      plus2A_out_53_port, plus2A_out_52_port, plus2A_out_51_port, 
      plus2A_out_50_port, plus2A_out_49_port, n7, n8, plus2A_out_46_port, 
      plus2A_out_45_port, plus2A_out_44_port, plus2A_out_43_port, 
      plus2A_out_42_port, plus2A_out_41_port, plus2A_out_40_port, 
      plus2A_out_39_port, plus2A_out_38_port, plus2A_out_37_port, 
      plus2A_out_36_port, plus2A_out_35_port, plus2A_out_34_port, 
      plus2A_out_33_port, plus2A_out_32_port, plus2A_out_31_port, 
      plus2A_out_30_port, plus2A_out_29_port, plus2A_out_28_port, 
      plus2A_out_27_port, plus2A_out_26_port, plus2A_out_25_port, 
      plus2A_out_24_port, plus2A_out_23_port, plus2A_out_22_port, 
      plus2A_out_21_port, plus2A_out_20_port, plus2A_out_19_port, 
      plus2A_out_18_port, plus2A_out_17_port, plus2A_out_16_port, 
      plus2A_out_15_port, plus2A_out_14_port, plus2A_out_13_port, 
      plus2A_out_12_port, plus2A_out_11_port, plus2A_out_10_port, 
      plus2A_out_9_port, plus2A_out_8_port, plus2A_out_7_port, 
      plus2A_out_6_port, plus2A_out_5_port, plus2A_out_4_port, 
      plus2A_out_3_port, plus2A_out_2_port, plus2A_out_1_port, 
      plus2A_out_0_port, plus4A_out_63_port, plus4A_out_62_port, 
      plus4A_out_61_port, plus4A_out_60_port, plus4A_out_59_port, 
      plus4A_out_58_port, plus4A_out_57_port, plus4A_out_56_port, 
      plus4A_out_55_port, plus4A_out_54_port, n9, n10, plus4A_out_51_port, 
      plus4A_out_50_port, plus4A_out_49_port, plus4A_out_48_port, 
      plus4A_out_47_port, plus4A_out_46_port, plus4A_out_45_port, 
      plus4A_out_44_port, plus4A_out_43_port, plus4A_out_42_port, 
      plus4A_out_41_port, plus4A_out_40_port, plus4A_out_39_port, 
      plus4A_out_38_port, plus4A_out_37_port, plus4A_out_36_port, 
      plus4A_out_35_port, plus4A_out_34_port, plus4A_out_33_port, 
      plus4A_out_32_port, plus4A_out_31_port, plus4A_out_30_port, 
      plus4A_out_29_port, plus4A_out_28_port, plus4A_out_27_port, 
      plus4A_out_26_port, plus4A_out_25_port, plus4A_out_24_port, 
      plus4A_out_23_port, plus4A_out_22_port, plus4A_out_21_port, 
      plus4A_out_20_port, plus4A_out_19_port, plus4A_out_18_port, 
      plus4A_out_17_port, plus4A_out_16_port, plus4A_out_15_port, 
      plus4A_out_14_port, plus4A_out_13_port, plus4A_out_12_port, 
      plus4A_out_11_port, plus4A_out_10_port, plus4A_out_9_port, 
      plus4A_out_8_port, plus4A_out_7_port, plus4A_out_6_port, 
      plus4A_out_5_port, plus4A_out_4_port, plus4A_out_3_port, 
      plus4A_out_2_port, plus4A_out_1_port, plus4A_out_0_port, 
      plus2A_out_47_port, plus2A_out_48_port, plus4A_out_52_port, 
      plus4A_out_53_port, plus2A_out_57_port, n_3160, n_3161 : std_logic;

begin
   plus2A_out <= ( plus2A_out_63_port, plus2A_out_62_port, plus2A_out_61_port, 
      plus2A_out_60_port, plus2A_out_59_port, plus2A_out_58_port, 
      plus2A_out_57_port, plus2A_out_56_port, plus2A_out_55_port, 
      plus2A_out_54_port, plus2A_out_53_port, plus2A_out_52_port, 
      plus2A_out_51_port, plus2A_out_50_port, plus2A_out_49_port, 
      plus2A_out_48_port, plus2A_out_47_port, plus2A_out_46_port, 
      plus2A_out_45_port, plus2A_out_44_port, plus2A_out_43_port, 
      plus2A_out_42_port, plus2A_out_41_port, plus2A_out_40_port, 
      plus2A_out_39_port, plus2A_out_38_port, plus2A_out_37_port, 
      plus2A_out_36_port, plus2A_out_35_port, plus2A_out_34_port, 
      plus2A_out_33_port, plus2A_out_32_port, plus2A_out_31_port, 
      plus2A_out_30_port, plus2A_out_29_port, plus2A_out_28_port, 
      plus2A_out_27_port, plus2A_out_26_port, plus2A_out_25_port, 
      plus2A_out_24_port, plus2A_out_23_port, plus2A_out_22_port, 
      plus2A_out_21_port, plus2A_out_20_port, plus2A_out_19_port, 
      plus2A_out_18_port, plus2A_out_17_port, plus2A_out_16_port, 
      plus2A_out_15_port, plus2A_out_14_port, plus2A_out_13_port, 
      plus2A_out_12_port, plus2A_out_11_port, plus2A_out_10_port, 
      plus2A_out_9_port, plus2A_out_8_port, plus2A_out_7_port, 
      plus2A_out_6_port, plus2A_out_5_port, plus2A_out_4_port, 
      plus2A_out_3_port, plus2A_out_2_port, plus2A_out_1_port, 
      plus2A_out_0_port );
   plus4A_out <= ( plus4A_out_63_port, plus4A_out_62_port, plus4A_out_61_port, 
      plus4A_out_60_port, plus4A_out_59_port, plus4A_out_58_port, 
      plus4A_out_57_port, plus4A_out_56_port, plus4A_out_55_port, 
      plus4A_out_54_port, plus4A_out_53_port, plus4A_out_52_port, 
      plus4A_out_51_port, plus4A_out_50_port, plus4A_out_49_port, 
      plus4A_out_48_port, plus4A_out_47_port, plus4A_out_46_port, 
      plus4A_out_45_port, plus4A_out_44_port, plus4A_out_43_port, 
      plus4A_out_42_port, plus4A_out_41_port, plus4A_out_40_port, 
      plus4A_out_39_port, plus4A_out_38_port, plus4A_out_37_port, 
      plus4A_out_36_port, plus4A_out_35_port, plus4A_out_34_port, 
      plus4A_out_33_port, plus4A_out_32_port, plus4A_out_31_port, 
      plus4A_out_30_port, plus4A_out_29_port, plus4A_out_28_port, 
      plus4A_out_27_port, plus4A_out_26_port, plus4A_out_25_port, 
      plus4A_out_24_port, plus4A_out_23_port, plus4A_out_22_port, 
      plus4A_out_21_port, plus4A_out_20_port, plus4A_out_19_port, 
      plus4A_out_18_port, plus4A_out_17_port, plus4A_out_16_port, 
      plus4A_out_15_port, plus4A_out_14_port, plus4A_out_13_port, 
      plus4A_out_12_port, plus4A_out_11_port, plus4A_out_10_port, 
      plus4A_out_9_port, plus4A_out_8_port, plus4A_out_7_port, 
      plus4A_out_6_port, plus4A_out_5_port, plus4A_out_4_port, 
      plus4A_out_3_port, plus4A_out_2_port, plus4A_out_1_port, 
      plus4A_out_0_port );
   
   plus2A_out_0_port <= '0';
   plus4A_out_0_port <= '0';
   shifter_1 : shifter_N64_18 port map( input(63) => plusA(63), input(62) => 
                           plusA(62), input(61) => plusA(61), input(60) => 
                           plusA(60), input(59) => plusA(59), input(58) => 
                           plusA(58), input(57) => plusA(57), input(56) => 
                           plusA(56), input(55) => plusA(55), input(54) => 
                           plusA(54), input(53) => plusA(53), input(52) => 
                           plusA(52), input(51) => plusA(51), input(50) => 
                           plusA(50), input(49) => plusA(49), input(48) => 
                           plusA(48), input(47) => plusA(47), input(46) => 
                           plusA(46), input(45) => plusA(45), input(44) => 
                           plusA(44), input(43) => plusA(43), input(42) => 
                           plusA(42), input(41) => plusA(41), input(40) => 
                           plusA(40), input(39) => plusA(39), input(38) => 
                           plusA(38), input(37) => plusA(37), input(36) => 
                           plusA(36), input(35) => plusA(35), input(34) => 
                           plusA(34), input(33) => plusA(33), input(32) => 
                           plusA(32), input(31) => plusA(31), input(30) => 
                           plusA(30), input(29) => plusA(29), input(28) => 
                           plusA(28), input(27) => plusA(27), input(26) => 
                           plusA(26), input(25) => plusA(25), input(24) => 
                           plusA(24), input(23) => plusA(23), input(22) => 
                           plusA(22), input(21) => plusA(21), input(20) => 
                           plusA(20), input(19) => plusA(19), input(18) => 
                           plusA(18), input(17) => plusA(17), input(16) => 
                           plusA(16), input(15) => plusA(15), input(14) => 
                           plusA(14), input(13) => plusA(13), input(12) => 
                           plusA(12), input(11) => plusA(11), input(10) => 
                           plusA(10), input(9) => plusA(9), input(8) => 
                           plusA(8), input(7) => plusA(7), input(6) => plusA(6)
                           , input(5) => plusA(5), input(4) => plusA(4), 
                           input(3) => plusA(3), input(2) => plusA(2), input(1)
                           => plusA(1), input(0) => plusA(0), 
                           shiftLeftOnePos(63) => plus2A_out_63_port, 
                           shiftLeftOnePos(62) => plus2A_out_62_port, 
                           shiftLeftOnePos(61) => plus2A_out_61_port, 
                           shiftLeftOnePos(60) => plus2A_out_60_port, 
                           shiftLeftOnePos(59) => plus2A_out_59_port, 
                           shiftLeftOnePos(58) => plus2A_out_58_port, 
                           shiftLeftOnePos(57) => n6, shiftLeftOnePos(56) => 
                           plus2A_out_56_port, shiftLeftOnePos(55) => 
                           plus2A_out_55_port, shiftLeftOnePos(54) => 
                           plus2A_out_54_port, shiftLeftOnePos(53) => 
                           plus2A_out_53_port, shiftLeftOnePos(52) => 
                           plus2A_out_52_port, shiftLeftOnePos(51) => 
                           plus2A_out_51_port, shiftLeftOnePos(50) => 
                           plus2A_out_50_port, shiftLeftOnePos(49) => 
                           plus2A_out_49_port, shiftLeftOnePos(48) => n7, 
                           shiftLeftOnePos(47) => n8, shiftLeftOnePos(46) => 
                           plus2A_out_46_port, shiftLeftOnePos(45) => 
                           plus2A_out_45_port, shiftLeftOnePos(44) => 
                           plus2A_out_44_port, shiftLeftOnePos(43) => 
                           plus2A_out_43_port, shiftLeftOnePos(42) => 
                           plus2A_out_42_port, shiftLeftOnePos(41) => 
                           plus2A_out_41_port, shiftLeftOnePos(40) => 
                           plus2A_out_40_port, shiftLeftOnePos(39) => 
                           plus2A_out_39_port, shiftLeftOnePos(38) => 
                           plus2A_out_38_port, shiftLeftOnePos(37) => 
                           plus2A_out_37_port, shiftLeftOnePos(36) => 
                           plus2A_out_36_port, shiftLeftOnePos(35) => 
                           plus2A_out_35_port, shiftLeftOnePos(34) => 
                           plus2A_out_34_port, shiftLeftOnePos(33) => 
                           plus2A_out_33_port, shiftLeftOnePos(32) => 
                           plus2A_out_32_port, shiftLeftOnePos(31) => 
                           plus2A_out_31_port, shiftLeftOnePos(30) => 
                           plus2A_out_30_port, shiftLeftOnePos(29) => 
                           plus2A_out_29_port, shiftLeftOnePos(28) => 
                           plus2A_out_28_port, shiftLeftOnePos(27) => 
                           plus2A_out_27_port, shiftLeftOnePos(26) => 
                           plus2A_out_26_port, shiftLeftOnePos(25) => 
                           plus2A_out_25_port, shiftLeftOnePos(24) => 
                           plus2A_out_24_port, shiftLeftOnePos(23) => 
                           plus2A_out_23_port, shiftLeftOnePos(22) => 
                           plus2A_out_22_port, shiftLeftOnePos(21) => 
                           plus2A_out_21_port, shiftLeftOnePos(20) => 
                           plus2A_out_20_port, shiftLeftOnePos(19) => 
                           plus2A_out_19_port, shiftLeftOnePos(18) => 
                           plus2A_out_18_port, shiftLeftOnePos(17) => 
                           plus2A_out_17_port, shiftLeftOnePos(16) => 
                           plus2A_out_16_port, shiftLeftOnePos(15) => 
                           plus2A_out_15_port, shiftLeftOnePos(14) => 
                           plus2A_out_14_port, shiftLeftOnePos(13) => 
                           plus2A_out_13_port, shiftLeftOnePos(12) => 
                           plus2A_out_12_port, shiftLeftOnePos(11) => 
                           plus2A_out_11_port, shiftLeftOnePos(10) => 
                           plus2A_out_10_port, shiftLeftOnePos(9) => 
                           plus2A_out_9_port, shiftLeftOnePos(8) => 
                           plus2A_out_8_port, shiftLeftOnePos(7) => 
                           plus2A_out_7_port, shiftLeftOnePos(6) => 
                           plus2A_out_6_port, shiftLeftOnePos(5) => 
                           plus2A_out_5_port, shiftLeftOnePos(4) => 
                           plus2A_out_4_port, shiftLeftOnePos(3) => 
                           plus2A_out_3_port, shiftLeftOnePos(2) => 
                           plus2A_out_2_port, shiftLeftOnePos(1) => 
                           plus2A_out_1_port, shiftLeftOnePos(0) => n_3160);
   shifter_2 : shifter_N64_17 port map( input(63) => plus2A_out_63_port, 
                           input(62) => plus2A_out_62_port, input(61) => 
                           plus2A_out_61_port, input(60) => plus2A_out_60_port,
                           input(59) => plus2A_out_59_port, input(58) => 
                           plus2A_out_58_port, input(57) => plus2A_out_57_port,
                           input(56) => plus2A_out_56_port, input(55) => 
                           plus2A_out_55_port, input(54) => plus2A_out_54_port,
                           input(53) => plus2A_out_53_port, input(52) => 
                           plus2A_out_52_port, input(51) => plus2A_out_51_port,
                           input(50) => plus2A_out_50_port, input(49) => 
                           plus2A_out_49_port, input(48) => plus2A_out_48_port,
                           input(47) => plus2A_out_47_port, input(46) => 
                           plus2A_out_46_port, input(45) => plus2A_out_45_port,
                           input(44) => plus2A_out_44_port, input(43) => 
                           plus2A_out_43_port, input(42) => plus2A_out_42_port,
                           input(41) => plus2A_out_41_port, input(40) => 
                           plus2A_out_40_port, input(39) => plus2A_out_39_port,
                           input(38) => plus2A_out_38_port, input(37) => 
                           plus2A_out_37_port, input(36) => plus2A_out_36_port,
                           input(35) => plus2A_out_35_port, input(34) => 
                           plus2A_out_34_port, input(33) => plus2A_out_33_port,
                           input(32) => plus2A_out_32_port, input(31) => 
                           plus2A_out_31_port, input(30) => plus2A_out_30_port,
                           input(29) => plus2A_out_29_port, input(28) => 
                           plus2A_out_28_port, input(27) => plus2A_out_27_port,
                           input(26) => plus2A_out_26_port, input(25) => 
                           plus2A_out_25_port, input(24) => plus2A_out_24_port,
                           input(23) => plus2A_out_23_port, input(22) => 
                           plus2A_out_22_port, input(21) => plus2A_out_21_port,
                           input(20) => plus2A_out_20_port, input(19) => 
                           plus2A_out_19_port, input(18) => plus2A_out_18_port,
                           input(17) => plus2A_out_17_port, input(16) => 
                           plus2A_out_16_port, input(15) => plus2A_out_15_port,
                           input(14) => plus2A_out_14_port, input(13) => 
                           plus2A_out_13_port, input(12) => plus2A_out_12_port,
                           input(11) => plus2A_out_11_port, input(10) => 
                           plus2A_out_10_port, input(9) => plus2A_out_9_port, 
                           input(8) => plus2A_out_8_port, input(7) => 
                           plus2A_out_7_port, input(6) => plus2A_out_6_port, 
                           input(5) => plus2A_out_5_port, input(4) => 
                           plus2A_out_4_port, input(3) => plus2A_out_3_port, 
                           input(2) => plus2A_out_2_port, input(1) => 
                           plus2A_out_1_port, input(0) => plus2A_out_0_port, 
                           shiftLeftOnePos(63) => plus4A_out_63_port, 
                           shiftLeftOnePos(62) => plus4A_out_62_port, 
                           shiftLeftOnePos(61) => plus4A_out_61_port, 
                           shiftLeftOnePos(60) => plus4A_out_60_port, 
                           shiftLeftOnePos(59) => plus4A_out_59_port, 
                           shiftLeftOnePos(58) => plus4A_out_58_port, 
                           shiftLeftOnePos(57) => plus4A_out_57_port, 
                           shiftLeftOnePos(56) => plus4A_out_56_port, 
                           shiftLeftOnePos(55) => plus4A_out_55_port, 
                           shiftLeftOnePos(54) => plus4A_out_54_port, 
                           shiftLeftOnePos(53) => n9, shiftLeftOnePos(52) => 
                           n10, shiftLeftOnePos(51) => plus4A_out_51_port, 
                           shiftLeftOnePos(50) => plus4A_out_50_port, 
                           shiftLeftOnePos(49) => plus4A_out_49_port, 
                           shiftLeftOnePos(48) => plus4A_out_48_port, 
                           shiftLeftOnePos(47) => plus4A_out_47_port, 
                           shiftLeftOnePos(46) => plus4A_out_46_port, 
                           shiftLeftOnePos(45) => plus4A_out_45_port, 
                           shiftLeftOnePos(44) => plus4A_out_44_port, 
                           shiftLeftOnePos(43) => plus4A_out_43_port, 
                           shiftLeftOnePos(42) => plus4A_out_42_port, 
                           shiftLeftOnePos(41) => plus4A_out_41_port, 
                           shiftLeftOnePos(40) => plus4A_out_40_port, 
                           shiftLeftOnePos(39) => plus4A_out_39_port, 
                           shiftLeftOnePos(38) => plus4A_out_38_port, 
                           shiftLeftOnePos(37) => plus4A_out_37_port, 
                           shiftLeftOnePos(36) => plus4A_out_36_port, 
                           shiftLeftOnePos(35) => plus4A_out_35_port, 
                           shiftLeftOnePos(34) => plus4A_out_34_port, 
                           shiftLeftOnePos(33) => plus4A_out_33_port, 
                           shiftLeftOnePos(32) => plus4A_out_32_port, 
                           shiftLeftOnePos(31) => plus4A_out_31_port, 
                           shiftLeftOnePos(30) => plus4A_out_30_port, 
                           shiftLeftOnePos(29) => plus4A_out_29_port, 
                           shiftLeftOnePos(28) => plus4A_out_28_port, 
                           shiftLeftOnePos(27) => plus4A_out_27_port, 
                           shiftLeftOnePos(26) => plus4A_out_26_port, 
                           shiftLeftOnePos(25) => plus4A_out_25_port, 
                           shiftLeftOnePos(24) => plus4A_out_24_port, 
                           shiftLeftOnePos(23) => plus4A_out_23_port, 
                           shiftLeftOnePos(22) => plus4A_out_22_port, 
                           shiftLeftOnePos(21) => plus4A_out_21_port, 
                           shiftLeftOnePos(20) => plus4A_out_20_port, 
                           shiftLeftOnePos(19) => plus4A_out_19_port, 
                           shiftLeftOnePos(18) => plus4A_out_18_port, 
                           shiftLeftOnePos(17) => plus4A_out_17_port, 
                           shiftLeftOnePos(16) => plus4A_out_16_port, 
                           shiftLeftOnePos(15) => plus4A_out_15_port, 
                           shiftLeftOnePos(14) => plus4A_out_14_port, 
                           shiftLeftOnePos(13) => plus4A_out_13_port, 
                           shiftLeftOnePos(12) => plus4A_out_12_port, 
                           shiftLeftOnePos(11) => plus4A_out_11_port, 
                           shiftLeftOnePos(10) => plus4A_out_10_port, 
                           shiftLeftOnePos(9) => plus4A_out_9_port, 
                           shiftLeftOnePos(8) => plus4A_out_8_port, 
                           shiftLeftOnePos(7) => plus4A_out_7_port, 
                           shiftLeftOnePos(6) => plus4A_out_6_port, 
                           shiftLeftOnePos(5) => plus4A_out_5_port, 
                           shiftLeftOnePos(4) => plus4A_out_4_port, 
                           shiftLeftOnePos(3) => plus4A_out_3_port, 
                           shiftLeftOnePos(2) => plus4A_out_2_port, 
                           shiftLeftOnePos(1) => plus4A_out_1_port, 
                           shiftLeftOnePos(0) => n_3161);
   complementer_1 : complementer_N64_18 port map( input(63) => 
                           plus2A_out_63_port, input(62) => plus2A_out_62_port,
                           input(61) => plus2A_out_61_port, input(60) => 
                           plus2A_out_60_port, input(59) => plus2A_out_59_port,
                           input(58) => plus2A_out_58_port, input(57) => 
                           plus2A_out_57_port, input(56) => plus2A_out_56_port,
                           input(55) => plus2A_out_55_port, input(54) => 
                           plus2A_out_54_port, input(53) => plus2A_out_53_port,
                           input(52) => plus2A_out_52_port, input(51) => 
                           plus2A_out_51_port, input(50) => plus2A_out_50_port,
                           input(49) => plus2A_out_49_port, input(48) => 
                           plus2A_out_48_port, input(47) => plus2A_out_47_port,
                           input(46) => plus2A_out_46_port, input(45) => 
                           plus2A_out_45_port, input(44) => plus2A_out_44_port,
                           input(43) => plus2A_out_43_port, input(42) => 
                           plus2A_out_42_port, input(41) => plus2A_out_41_port,
                           input(40) => plus2A_out_40_port, input(39) => 
                           plus2A_out_39_port, input(38) => plus2A_out_38_port,
                           input(37) => plus2A_out_37_port, input(36) => 
                           plus2A_out_36_port, input(35) => plus2A_out_35_port,
                           input(34) => plus2A_out_34_port, input(33) => 
                           plus2A_out_33_port, input(32) => plus2A_out_32_port,
                           input(31) => plus2A_out_31_port, input(30) => 
                           plus2A_out_30_port, input(29) => plus2A_out_29_port,
                           input(28) => plus2A_out_28_port, input(27) => 
                           plus2A_out_27_port, input(26) => plus2A_out_26_port,
                           input(25) => plus2A_out_25_port, input(24) => 
                           plus2A_out_24_port, input(23) => plus2A_out_23_port,
                           input(22) => plus2A_out_22_port, input(21) => 
                           plus2A_out_21_port, input(20) => plus2A_out_20_port,
                           input(19) => plus2A_out_19_port, input(18) => 
                           plus2A_out_18_port, input(17) => plus2A_out_17_port,
                           input(16) => plus2A_out_16_port, input(15) => 
                           plus2A_out_15_port, input(14) => plus2A_out_14_port,
                           input(13) => plus2A_out_13_port, input(12) => 
                           plus2A_out_12_port, input(11) => plus2A_out_11_port,
                           input(10) => plus2A_out_10_port, input(9) => 
                           plus2A_out_9_port, input(8) => plus2A_out_8_port, 
                           input(7) => plus2A_out_7_port, input(6) => 
                           plus2A_out_6_port, input(5) => plus2A_out_5_port, 
                           input(4) => plus2A_out_4_port, input(3) => 
                           plus2A_out_3_port, input(2) => plus2A_out_2_port, 
                           input(1) => plus2A_out_1_port, input(0) => 
                           plus2A_out_0_port, complement2(63) => 
                           minus2A_out(63), complement2(62) => minus2A_out(62),
                           complement2(61) => minus2A_out(61), complement2(60) 
                           => minus2A_out(60), complement2(59) => 
                           minus2A_out(59), complement2(58) => minus2A_out(58),
                           complement2(57) => minus2A_out(57), complement2(56) 
                           => minus2A_out(56), complement2(55) => 
                           minus2A_out(55), complement2(54) => minus2A_out(54),
                           complement2(53) => minus2A_out(53), complement2(52) 
                           => minus2A_out(52), complement2(51) => 
                           minus2A_out(51), complement2(50) => minus2A_out(50),
                           complement2(49) => minus2A_out(49), complement2(48) 
                           => minus2A_out(48), complement2(47) => 
                           minus2A_out(47), complement2(46) => minus2A_out(46),
                           complement2(45) => minus2A_out(45), complement2(44) 
                           => minus2A_out(44), complement2(43) => 
                           minus2A_out(43), complement2(42) => minus2A_out(42),
                           complement2(41) => minus2A_out(41), complement2(40) 
                           => minus2A_out(40), complement2(39) => 
                           minus2A_out(39), complement2(38) => minus2A_out(38),
                           complement2(37) => minus2A_out(37), complement2(36) 
                           => minus2A_out(36), complement2(35) => 
                           minus2A_out(35), complement2(34) => minus2A_out(34),
                           complement2(33) => minus2A_out(33), complement2(32) 
                           => minus2A_out(32), complement2(31) => 
                           minus2A_out(31), complement2(30) => minus2A_out(30),
                           complement2(29) => minus2A_out(29), complement2(28) 
                           => minus2A_out(28), complement2(27) => 
                           minus2A_out(27), complement2(26) => minus2A_out(26),
                           complement2(25) => minus2A_out(25), complement2(24) 
                           => minus2A_out(24), complement2(23) => 
                           minus2A_out(23), complement2(22) => minus2A_out(22),
                           complement2(21) => minus2A_out(21), complement2(20) 
                           => minus2A_out(20), complement2(19) => 
                           minus2A_out(19), complement2(18) => minus2A_out(18),
                           complement2(17) => minus2A_out(17), complement2(16) 
                           => minus2A_out(16), complement2(15) => 
                           minus2A_out(15), complement2(14) => minus2A_out(14),
                           complement2(13) => minus2A_out(13), complement2(12) 
                           => minus2A_out(12), complement2(11) => 
                           minus2A_out(11), complement2(10) => minus2A_out(10),
                           complement2(9) => minus2A_out(9), complement2(8) => 
                           minus2A_out(8), complement2(7) => minus2A_out(7), 
                           complement2(6) => minus2A_out(6), complement2(5) => 
                           minus2A_out(5), complement2(4) => minus2A_out(4), 
                           complement2(3) => minus2A_out(3), complement2(2) => 
                           minus2A_out(2), complement2(1) => minus2A_out(1), 
                           complement2(0) => minus2A_out(0));
   complementer_2 : complementer_N64_17 port map( input(63) => 
                           plus4A_out_63_port, input(62) => plus4A_out_62_port,
                           input(61) => plus4A_out_61_port, input(60) => 
                           plus4A_out_60_port, input(59) => plus4A_out_59_port,
                           input(58) => plus4A_out_58_port, input(57) => 
                           plus4A_out_57_port, input(56) => plus4A_out_56_port,
                           input(55) => plus4A_out_55_port, input(54) => 
                           plus4A_out_54_port, input(53) => plus4A_out_53_port,
                           input(52) => plus4A_out_52_port, input(51) => 
                           plus4A_out_51_port, input(50) => plus4A_out_50_port,
                           input(49) => plus4A_out_49_port, input(48) => 
                           plus4A_out_48_port, input(47) => plus4A_out_47_port,
                           input(46) => plus4A_out_46_port, input(45) => 
                           plus4A_out_45_port, input(44) => plus4A_out_44_port,
                           input(43) => plus4A_out_43_port, input(42) => 
                           plus4A_out_42_port, input(41) => plus4A_out_41_port,
                           input(40) => plus4A_out_40_port, input(39) => 
                           plus4A_out_39_port, input(38) => plus4A_out_38_port,
                           input(37) => plus4A_out_37_port, input(36) => 
                           plus4A_out_36_port, input(35) => plus4A_out_35_port,
                           input(34) => plus4A_out_34_port, input(33) => 
                           plus4A_out_33_port, input(32) => plus4A_out_32_port,
                           input(31) => plus4A_out_31_port, input(30) => 
                           plus4A_out_30_port, input(29) => plus4A_out_29_port,
                           input(28) => plus4A_out_28_port, input(27) => 
                           plus4A_out_27_port, input(26) => plus4A_out_26_port,
                           input(25) => plus4A_out_25_port, input(24) => 
                           plus4A_out_24_port, input(23) => plus4A_out_23_port,
                           input(22) => plus4A_out_22_port, input(21) => 
                           plus4A_out_21_port, input(20) => plus4A_out_20_port,
                           input(19) => plus4A_out_19_port, input(18) => 
                           plus4A_out_18_port, input(17) => plus4A_out_17_port,
                           input(16) => plus4A_out_16_port, input(15) => 
                           plus4A_out_15_port, input(14) => plus4A_out_14_port,
                           input(13) => plus4A_out_13_port, input(12) => 
                           plus4A_out_12_port, input(11) => plus4A_out_11_port,
                           input(10) => plus4A_out_10_port, input(9) => 
                           plus4A_out_9_port, input(8) => plus4A_out_8_port, 
                           input(7) => plus4A_out_7_port, input(6) => 
                           plus4A_out_6_port, input(5) => plus4A_out_5_port, 
                           input(4) => plus4A_out_4_port, input(3) => 
                           plus4A_out_3_port, input(2) => plus4A_out_2_port, 
                           input(1) => plus4A_out_1_port, input(0) => 
                           plus4A_out_0_port, complement2(63) => 
                           minus4A_out(63), complement2(62) => minus4A_out(62),
                           complement2(61) => minus4A_out(61), complement2(60) 
                           => minus4A_out(60), complement2(59) => 
                           minus4A_out(59), complement2(58) => minus4A_out(58),
                           complement2(57) => minus4A_out(57), complement2(56) 
                           => minus4A_out(56), complement2(55) => 
                           minus4A_out(55), complement2(54) => minus4A_out(54),
                           complement2(53) => minus4A_out(53), complement2(52) 
                           => minus4A_out(52), complement2(51) => 
                           minus4A_out(51), complement2(50) => minus4A_out(50),
                           complement2(49) => minus4A_out(49), complement2(48) 
                           => minus4A_out(48), complement2(47) => 
                           minus4A_out(47), complement2(46) => minus4A_out(46),
                           complement2(45) => minus4A_out(45), complement2(44) 
                           => minus4A_out(44), complement2(43) => 
                           minus4A_out(43), complement2(42) => minus4A_out(42),
                           complement2(41) => minus4A_out(41), complement2(40) 
                           => minus4A_out(40), complement2(39) => 
                           minus4A_out(39), complement2(38) => minus4A_out(38),
                           complement2(37) => minus4A_out(37), complement2(36) 
                           => minus4A_out(36), complement2(35) => 
                           minus4A_out(35), complement2(34) => minus4A_out(34),
                           complement2(33) => minus4A_out(33), complement2(32) 
                           => minus4A_out(32), complement2(31) => 
                           minus4A_out(31), complement2(30) => minus4A_out(30),
                           complement2(29) => minus4A_out(29), complement2(28) 
                           => minus4A_out(28), complement2(27) => 
                           minus4A_out(27), complement2(26) => minus4A_out(26),
                           complement2(25) => minus4A_out(25), complement2(24) 
                           => minus4A_out(24), complement2(23) => 
                           minus4A_out(23), complement2(22) => minus4A_out(22),
                           complement2(21) => minus4A_out(21), complement2(20) 
                           => minus4A_out(20), complement2(19) => 
                           minus4A_out(19), complement2(18) => minus4A_out(18),
                           complement2(17) => minus4A_out(17), complement2(16) 
                           => minus4A_out(16), complement2(15) => 
                           minus4A_out(15), complement2(14) => minus4A_out(14),
                           complement2(13) => minus4A_out(13), complement2(12) 
                           => minus4A_out(12), complement2(11) => 
                           minus4A_out(11), complement2(10) => minus4A_out(10),
                           complement2(9) => minus4A_out(9), complement2(8) => 
                           minus4A_out(8), complement2(7) => minus4A_out(7), 
                           complement2(6) => minus4A_out(6), complement2(5) => 
                           minus4A_out(5), complement2(4) => minus4A_out(4), 
                           complement2(3) => minus4A_out(3), complement2(2) => 
                           minus4A_out(2), complement2(1) => minus4A_out(1), 
                           complement2(0) => minus4A_out(0));
   U3 : BUF_X1 port map( A => n10, Z => plus4A_out_52_port);
   U4 : BUF_X1 port map( A => n9, Z => plus4A_out_53_port);
   U5 : BUF_X1 port map( A => n8, Z => plus2A_out_47_port);
   U6 : BUF_X1 port map( A => n7, Z => plus2A_out_48_port);
   U7 : BUF_X1 port map( A => n6, Z => plus2A_out_57_port);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity ShiftnCompl_N64_10 is

   port( plusA : in std_logic_vector (63 downto 0);  plus2A_out, minus2A_out, 
         plus4A_out, minus4A_out : out std_logic_vector (63 downto 0));

end ShiftnCompl_N64_10;

architecture SYN_struct of ShiftnCompl_N64_10 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component complementer_N64_19
      port( input : in std_logic_vector (63 downto 0);  complement2 : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component complementer_N64_20
      port( input : in std_logic_vector (63 downto 0);  complement2 : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component shifter_N64_19
      port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component shifter_N64_20
      port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
            std_logic_vector (63 downto 0));
   end component;
   
   signal plus2A_out_63_port, plus2A_out_62_port, plus2A_out_61_port, 
      plus2A_out_60_port, plus2A_out_59_port, plus2A_out_58_port, n36, 
      plus2A_out_56_port, plus2A_out_55_port, plus2A_out_54_port, 
      plus2A_out_53_port, plus2A_out_52_port, plus2A_out_51_port, 
      plus2A_out_50_port, plus2A_out_49_port, n37, n38, plus2A_out_46_port, 
      plus2A_out_45_port, plus2A_out_44_port, plus2A_out_43_port, 
      plus2A_out_42_port, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49
      , n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, 
      n64, n65, n66, n67, n68, plus2A_out_11_port, plus2A_out_10_port, 
      plus2A_out_9_port, plus2A_out_8_port, plus2A_out_7_port, 
      plus2A_out_6_port, plus2A_out_5_port, plus2A_out_4_port, 
      plus2A_out_3_port, plus2A_out_2_port, plus2A_out_1_port, 
      plus2A_out_0_port, plus4A_out_63_port, plus4A_out_62_port, 
      plus4A_out_61_port, plus4A_out_60_port, plus4A_out_59_port, 
      plus4A_out_58_port, plus4A_out_57_port, plus4A_out_56_port, 
      plus4A_out_55_port, plus4A_out_54_port, n69, n70, plus4A_out_51_port, 
      plus4A_out_50_port, plus4A_out_49_port, plus4A_out_48_port, 
      plus4A_out_47_port, plus4A_out_46_port, plus4A_out_45_port, 
      plus4A_out_44_port, plus4A_out_43_port, plus4A_out_42_port, 
      plus4A_out_41_port, plus4A_out_40_port, plus4A_out_39_port, 
      plus4A_out_38_port, plus4A_out_37_port, plus4A_out_36_port, 
      plus4A_out_35_port, plus4A_out_34_port, plus4A_out_33_port, 
      plus4A_out_32_port, plus4A_out_31_port, plus4A_out_30_port, 
      plus4A_out_29_port, plus4A_out_28_port, plus4A_out_27_port, 
      plus4A_out_26_port, plus4A_out_25_port, plus4A_out_24_port, 
      plus4A_out_23_port, plus4A_out_22_port, plus4A_out_21_port, 
      plus4A_out_20_port, plus4A_out_19_port, plus4A_out_18_port, 
      plus4A_out_17_port, plus4A_out_16_port, plus4A_out_15_port, 
      plus4A_out_14_port, plus4A_out_13_port, plus4A_out_12_port, 
      plus4A_out_11_port, plus4A_out_10_port, plus4A_out_9_port, 
      plus4A_out_8_port, plus4A_out_7_port, plus4A_out_6_port, 
      plus4A_out_5_port, plus4A_out_4_port, plus4A_out_3_port, 
      plus4A_out_2_port, plus4A_out_1_port, plus4A_out_0_port, 
      plus2A_out_12_port, plus2A_out_13_port, plus2A_out_14_port, 
      plus2A_out_15_port, plus2A_out_16_port, plus2A_out_17_port, 
      plus2A_out_18_port, plus2A_out_19_port, plus2A_out_20_port, 
      plus2A_out_21_port, plus2A_out_22_port, plus2A_out_23_port, 
      plus2A_out_24_port, plus2A_out_25_port, plus2A_out_26_port, 
      plus2A_out_27_port, plus2A_out_28_port, plus2A_out_29_port, 
      plus2A_out_30_port, plus2A_out_31_port, plus2A_out_32_port, 
      plus2A_out_33_port, plus2A_out_34_port, plus2A_out_35_port, 
      plus2A_out_36_port, plus2A_out_37_port, plus2A_out_38_port, 
      plus2A_out_39_port, plus2A_out_40_port, plus2A_out_41_port, 
      plus2A_out_47_port, plus2A_out_48_port, plus4A_out_52_port, 
      plus4A_out_53_port, plus2A_out_57_port, n_3162, n_3163 : std_logic;

begin
   plus2A_out <= ( plus2A_out_63_port, plus2A_out_62_port, plus2A_out_61_port, 
      plus2A_out_60_port, plus2A_out_59_port, plus2A_out_58_port, 
      plus2A_out_57_port, plus2A_out_56_port, plus2A_out_55_port, 
      plus2A_out_54_port, plus2A_out_53_port, plus2A_out_52_port, 
      plus2A_out_51_port, plus2A_out_50_port, plus2A_out_49_port, 
      plus2A_out_48_port, plus2A_out_47_port, plus2A_out_46_port, 
      plus2A_out_45_port, plus2A_out_44_port, plus2A_out_43_port, 
      plus2A_out_42_port, plus2A_out_41_port, plus2A_out_40_port, 
      plus2A_out_39_port, plus2A_out_38_port, plus2A_out_37_port, 
      plus2A_out_36_port, plus2A_out_35_port, plus2A_out_34_port, 
      plus2A_out_33_port, plus2A_out_32_port, plus2A_out_31_port, 
      plus2A_out_30_port, plus2A_out_29_port, plus2A_out_28_port, 
      plus2A_out_27_port, plus2A_out_26_port, plus2A_out_25_port, 
      plus2A_out_24_port, plus2A_out_23_port, plus2A_out_22_port, 
      plus2A_out_21_port, plus2A_out_20_port, plus2A_out_19_port, 
      plus2A_out_18_port, plus2A_out_17_port, plus2A_out_16_port, 
      plus2A_out_15_port, plus2A_out_14_port, plus2A_out_13_port, 
      plus2A_out_12_port, plus2A_out_11_port, plus2A_out_10_port, 
      plus2A_out_9_port, plus2A_out_8_port, plus2A_out_7_port, 
      plus2A_out_6_port, plus2A_out_5_port, plus2A_out_4_port, 
      plus2A_out_3_port, plus2A_out_2_port, plus2A_out_1_port, 
      plus2A_out_0_port );
   plus4A_out <= ( plus4A_out_63_port, plus4A_out_62_port, plus4A_out_61_port, 
      plus4A_out_60_port, plus4A_out_59_port, plus4A_out_58_port, 
      plus4A_out_57_port, plus4A_out_56_port, plus4A_out_55_port, 
      plus4A_out_54_port, plus4A_out_53_port, plus4A_out_52_port, 
      plus4A_out_51_port, plus4A_out_50_port, plus4A_out_49_port, 
      plus4A_out_48_port, plus4A_out_47_port, plus4A_out_46_port, 
      plus4A_out_45_port, plus4A_out_44_port, plus4A_out_43_port, 
      plus4A_out_42_port, plus4A_out_41_port, plus4A_out_40_port, 
      plus4A_out_39_port, plus4A_out_38_port, plus4A_out_37_port, 
      plus4A_out_36_port, plus4A_out_35_port, plus4A_out_34_port, 
      plus4A_out_33_port, plus4A_out_32_port, plus4A_out_31_port, 
      plus4A_out_30_port, plus4A_out_29_port, plus4A_out_28_port, 
      plus4A_out_27_port, plus4A_out_26_port, plus4A_out_25_port, 
      plus4A_out_24_port, plus4A_out_23_port, plus4A_out_22_port, 
      plus4A_out_21_port, plus4A_out_20_port, plus4A_out_19_port, 
      plus4A_out_18_port, plus4A_out_17_port, plus4A_out_16_port, 
      plus4A_out_15_port, plus4A_out_14_port, plus4A_out_13_port, 
      plus4A_out_12_port, plus4A_out_11_port, plus4A_out_10_port, 
      plus4A_out_9_port, plus4A_out_8_port, plus4A_out_7_port, 
      plus4A_out_6_port, plus4A_out_5_port, plus4A_out_4_port, 
      plus4A_out_3_port, plus4A_out_2_port, plus4A_out_1_port, 
      plus4A_out_0_port );
   
   plus2A_out_0_port <= '0';
   plus4A_out_0_port <= '0';
   shifter_1 : shifter_N64_20 port map( input(63) => plusA(63), input(62) => 
                           plusA(62), input(61) => plusA(61), input(60) => 
                           plusA(60), input(59) => plusA(59), input(58) => 
                           plusA(58), input(57) => plusA(57), input(56) => 
                           plusA(56), input(55) => plusA(55), input(54) => 
                           plusA(54), input(53) => plusA(53), input(52) => 
                           plusA(52), input(51) => plusA(51), input(50) => 
                           plusA(50), input(49) => plusA(49), input(48) => 
                           plusA(48), input(47) => plusA(47), input(46) => 
                           plusA(46), input(45) => plusA(45), input(44) => 
                           plusA(44), input(43) => plusA(43), input(42) => 
                           plusA(42), input(41) => plusA(41), input(40) => 
                           plusA(40), input(39) => plusA(39), input(38) => 
                           plusA(38), input(37) => plusA(37), input(36) => 
                           plusA(36), input(35) => plusA(35), input(34) => 
                           plusA(34), input(33) => plusA(33), input(32) => 
                           plusA(32), input(31) => plusA(31), input(30) => 
                           plusA(30), input(29) => plusA(29), input(28) => 
                           plusA(28), input(27) => plusA(27), input(26) => 
                           plusA(26), input(25) => plusA(25), input(24) => 
                           plusA(24), input(23) => plusA(23), input(22) => 
                           plusA(22), input(21) => plusA(21), input(20) => 
                           plusA(20), input(19) => plusA(19), input(18) => 
                           plusA(18), input(17) => plusA(17), input(16) => 
                           plusA(16), input(15) => plusA(15), input(14) => 
                           plusA(14), input(13) => plusA(13), input(12) => 
                           plusA(12), input(11) => plusA(11), input(10) => 
                           plusA(10), input(9) => plusA(9), input(8) => 
                           plusA(8), input(7) => plusA(7), input(6) => plusA(6)
                           , input(5) => plusA(5), input(4) => plusA(4), 
                           input(3) => plusA(3), input(2) => plusA(2), input(1)
                           => plusA(1), input(0) => plusA(0), 
                           shiftLeftOnePos(63) => plus2A_out_63_port, 
                           shiftLeftOnePos(62) => plus2A_out_62_port, 
                           shiftLeftOnePos(61) => plus2A_out_61_port, 
                           shiftLeftOnePos(60) => plus2A_out_60_port, 
                           shiftLeftOnePos(59) => plus2A_out_59_port, 
                           shiftLeftOnePos(58) => plus2A_out_58_port, 
                           shiftLeftOnePos(57) => n36, shiftLeftOnePos(56) => 
                           plus2A_out_56_port, shiftLeftOnePos(55) => 
                           plus2A_out_55_port, shiftLeftOnePos(54) => 
                           plus2A_out_54_port, shiftLeftOnePos(53) => 
                           plus2A_out_53_port, shiftLeftOnePos(52) => 
                           plus2A_out_52_port, shiftLeftOnePos(51) => 
                           plus2A_out_51_port, shiftLeftOnePos(50) => 
                           plus2A_out_50_port, shiftLeftOnePos(49) => 
                           plus2A_out_49_port, shiftLeftOnePos(48) => n37, 
                           shiftLeftOnePos(47) => n38, shiftLeftOnePos(46) => 
                           plus2A_out_46_port, shiftLeftOnePos(45) => 
                           plus2A_out_45_port, shiftLeftOnePos(44) => 
                           plus2A_out_44_port, shiftLeftOnePos(43) => 
                           plus2A_out_43_port, shiftLeftOnePos(42) => 
                           plus2A_out_42_port, shiftLeftOnePos(41) => n39, 
                           shiftLeftOnePos(40) => n40, shiftLeftOnePos(39) => 
                           n41, shiftLeftOnePos(38) => n42, shiftLeftOnePos(37)
                           => n43, shiftLeftOnePos(36) => n44, 
                           shiftLeftOnePos(35) => n45, shiftLeftOnePos(34) => 
                           n46, shiftLeftOnePos(33) => n47, shiftLeftOnePos(32)
                           => n48, shiftLeftOnePos(31) => n49, 
                           shiftLeftOnePos(30) => n50, shiftLeftOnePos(29) => 
                           n51, shiftLeftOnePos(28) => n52, shiftLeftOnePos(27)
                           => n53, shiftLeftOnePos(26) => n54, 
                           shiftLeftOnePos(25) => n55, shiftLeftOnePos(24) => 
                           n56, shiftLeftOnePos(23) => n57, shiftLeftOnePos(22)
                           => n58, shiftLeftOnePos(21) => n59, 
                           shiftLeftOnePos(20) => n60, shiftLeftOnePos(19) => 
                           n61, shiftLeftOnePos(18) => n62, shiftLeftOnePos(17)
                           => n63, shiftLeftOnePos(16) => n64, 
                           shiftLeftOnePos(15) => n65, shiftLeftOnePos(14) => 
                           n66, shiftLeftOnePos(13) => n67, shiftLeftOnePos(12)
                           => n68, shiftLeftOnePos(11) => plus2A_out_11_port, 
                           shiftLeftOnePos(10) => plus2A_out_10_port, 
                           shiftLeftOnePos(9) => plus2A_out_9_port, 
                           shiftLeftOnePos(8) => plus2A_out_8_port, 
                           shiftLeftOnePos(7) => plus2A_out_7_port, 
                           shiftLeftOnePos(6) => plus2A_out_6_port, 
                           shiftLeftOnePos(5) => plus2A_out_5_port, 
                           shiftLeftOnePos(4) => plus2A_out_4_port, 
                           shiftLeftOnePos(3) => plus2A_out_3_port, 
                           shiftLeftOnePos(2) => plus2A_out_2_port, 
                           shiftLeftOnePos(1) => plus2A_out_1_port, 
                           shiftLeftOnePos(0) => n_3162);
   shifter_2 : shifter_N64_19 port map( input(63) => plus2A_out_63_port, 
                           input(62) => plus2A_out_62_port, input(61) => 
                           plus2A_out_61_port, input(60) => plus2A_out_60_port,
                           input(59) => plus2A_out_59_port, input(58) => 
                           plus2A_out_58_port, input(57) => plus2A_out_57_port,
                           input(56) => plus2A_out_56_port, input(55) => 
                           plus2A_out_55_port, input(54) => plus2A_out_54_port,
                           input(53) => plus2A_out_53_port, input(52) => 
                           plus2A_out_52_port, input(51) => plus2A_out_51_port,
                           input(50) => plus2A_out_50_port, input(49) => 
                           plus2A_out_49_port, input(48) => plus2A_out_48_port,
                           input(47) => plus2A_out_47_port, input(46) => 
                           plus2A_out_46_port, input(45) => plus2A_out_45_port,
                           input(44) => plus2A_out_44_port, input(43) => 
                           plus2A_out_43_port, input(42) => plus2A_out_42_port,
                           input(41) => plus2A_out_41_port, input(40) => 
                           plus2A_out_40_port, input(39) => plus2A_out_39_port,
                           input(38) => plus2A_out_38_port, input(37) => 
                           plus2A_out_37_port, input(36) => plus2A_out_36_port,
                           input(35) => plus2A_out_35_port, input(34) => 
                           plus2A_out_34_port, input(33) => plus2A_out_33_port,
                           input(32) => plus2A_out_32_port, input(31) => 
                           plus2A_out_31_port, input(30) => plus2A_out_30_port,
                           input(29) => plus2A_out_29_port, input(28) => 
                           plus2A_out_28_port, input(27) => plus2A_out_27_port,
                           input(26) => plus2A_out_26_port, input(25) => 
                           plus2A_out_25_port, input(24) => plus2A_out_24_port,
                           input(23) => plus2A_out_23_port, input(22) => 
                           plus2A_out_22_port, input(21) => plus2A_out_21_port,
                           input(20) => plus2A_out_20_port, input(19) => 
                           plus2A_out_19_port, input(18) => plus2A_out_18_port,
                           input(17) => plus2A_out_17_port, input(16) => 
                           plus2A_out_16_port, input(15) => plus2A_out_15_port,
                           input(14) => plus2A_out_14_port, input(13) => 
                           plus2A_out_13_port, input(12) => plus2A_out_12_port,
                           input(11) => plus2A_out_11_port, input(10) => 
                           plus2A_out_10_port, input(9) => plus2A_out_9_port, 
                           input(8) => plus2A_out_8_port, input(7) => 
                           plus2A_out_7_port, input(6) => plus2A_out_6_port, 
                           input(5) => plus2A_out_5_port, input(4) => 
                           plus2A_out_4_port, input(3) => plus2A_out_3_port, 
                           input(2) => plus2A_out_2_port, input(1) => 
                           plus2A_out_1_port, input(0) => plus2A_out_0_port, 
                           shiftLeftOnePos(63) => plus4A_out_63_port, 
                           shiftLeftOnePos(62) => plus4A_out_62_port, 
                           shiftLeftOnePos(61) => plus4A_out_61_port, 
                           shiftLeftOnePos(60) => plus4A_out_60_port, 
                           shiftLeftOnePos(59) => plus4A_out_59_port, 
                           shiftLeftOnePos(58) => plus4A_out_58_port, 
                           shiftLeftOnePos(57) => plus4A_out_57_port, 
                           shiftLeftOnePos(56) => plus4A_out_56_port, 
                           shiftLeftOnePos(55) => plus4A_out_55_port, 
                           shiftLeftOnePos(54) => plus4A_out_54_port, 
                           shiftLeftOnePos(53) => n69, shiftLeftOnePos(52) => 
                           n70, shiftLeftOnePos(51) => plus4A_out_51_port, 
                           shiftLeftOnePos(50) => plus4A_out_50_port, 
                           shiftLeftOnePos(49) => plus4A_out_49_port, 
                           shiftLeftOnePos(48) => plus4A_out_48_port, 
                           shiftLeftOnePos(47) => plus4A_out_47_port, 
                           shiftLeftOnePos(46) => plus4A_out_46_port, 
                           shiftLeftOnePos(45) => plus4A_out_45_port, 
                           shiftLeftOnePos(44) => plus4A_out_44_port, 
                           shiftLeftOnePos(43) => plus4A_out_43_port, 
                           shiftLeftOnePos(42) => plus4A_out_42_port, 
                           shiftLeftOnePos(41) => plus4A_out_41_port, 
                           shiftLeftOnePos(40) => plus4A_out_40_port, 
                           shiftLeftOnePos(39) => plus4A_out_39_port, 
                           shiftLeftOnePos(38) => plus4A_out_38_port, 
                           shiftLeftOnePos(37) => plus4A_out_37_port, 
                           shiftLeftOnePos(36) => plus4A_out_36_port, 
                           shiftLeftOnePos(35) => plus4A_out_35_port, 
                           shiftLeftOnePos(34) => plus4A_out_34_port, 
                           shiftLeftOnePos(33) => plus4A_out_33_port, 
                           shiftLeftOnePos(32) => plus4A_out_32_port, 
                           shiftLeftOnePos(31) => plus4A_out_31_port, 
                           shiftLeftOnePos(30) => plus4A_out_30_port, 
                           shiftLeftOnePos(29) => plus4A_out_29_port, 
                           shiftLeftOnePos(28) => plus4A_out_28_port, 
                           shiftLeftOnePos(27) => plus4A_out_27_port, 
                           shiftLeftOnePos(26) => plus4A_out_26_port, 
                           shiftLeftOnePos(25) => plus4A_out_25_port, 
                           shiftLeftOnePos(24) => plus4A_out_24_port, 
                           shiftLeftOnePos(23) => plus4A_out_23_port, 
                           shiftLeftOnePos(22) => plus4A_out_22_port, 
                           shiftLeftOnePos(21) => plus4A_out_21_port, 
                           shiftLeftOnePos(20) => plus4A_out_20_port, 
                           shiftLeftOnePos(19) => plus4A_out_19_port, 
                           shiftLeftOnePos(18) => plus4A_out_18_port, 
                           shiftLeftOnePos(17) => plus4A_out_17_port, 
                           shiftLeftOnePos(16) => plus4A_out_16_port, 
                           shiftLeftOnePos(15) => plus4A_out_15_port, 
                           shiftLeftOnePos(14) => plus4A_out_14_port, 
                           shiftLeftOnePos(13) => plus4A_out_13_port, 
                           shiftLeftOnePos(12) => plus4A_out_12_port, 
                           shiftLeftOnePos(11) => plus4A_out_11_port, 
                           shiftLeftOnePos(10) => plus4A_out_10_port, 
                           shiftLeftOnePos(9) => plus4A_out_9_port, 
                           shiftLeftOnePos(8) => plus4A_out_8_port, 
                           shiftLeftOnePos(7) => plus4A_out_7_port, 
                           shiftLeftOnePos(6) => plus4A_out_6_port, 
                           shiftLeftOnePos(5) => plus4A_out_5_port, 
                           shiftLeftOnePos(4) => plus4A_out_4_port, 
                           shiftLeftOnePos(3) => plus4A_out_3_port, 
                           shiftLeftOnePos(2) => plus4A_out_2_port, 
                           shiftLeftOnePos(1) => plus4A_out_1_port, 
                           shiftLeftOnePos(0) => n_3163);
   complementer_1 : complementer_N64_20 port map( input(63) => 
                           plus2A_out_63_port, input(62) => plus2A_out_62_port,
                           input(61) => plus2A_out_61_port, input(60) => 
                           plus2A_out_60_port, input(59) => plus2A_out_59_port,
                           input(58) => plus2A_out_58_port, input(57) => 
                           plus2A_out_57_port, input(56) => plus2A_out_56_port,
                           input(55) => plus2A_out_55_port, input(54) => 
                           plus2A_out_54_port, input(53) => plus2A_out_53_port,
                           input(52) => plus2A_out_52_port, input(51) => 
                           plus2A_out_51_port, input(50) => plus2A_out_50_port,
                           input(49) => plus2A_out_49_port, input(48) => 
                           plus2A_out_48_port, input(47) => plus2A_out_47_port,
                           input(46) => plus2A_out_46_port, input(45) => 
                           plus2A_out_45_port, input(44) => plus2A_out_44_port,
                           input(43) => plus2A_out_43_port, input(42) => 
                           plus2A_out_42_port, input(41) => plus2A_out_41_port,
                           input(40) => plus2A_out_40_port, input(39) => 
                           plus2A_out_39_port, input(38) => plus2A_out_38_port,
                           input(37) => plus2A_out_37_port, input(36) => 
                           plus2A_out_36_port, input(35) => plus2A_out_35_port,
                           input(34) => plus2A_out_34_port, input(33) => 
                           plus2A_out_33_port, input(32) => plus2A_out_32_port,
                           input(31) => plus2A_out_31_port, input(30) => 
                           plus2A_out_30_port, input(29) => plus2A_out_29_port,
                           input(28) => plus2A_out_28_port, input(27) => 
                           plus2A_out_27_port, input(26) => plus2A_out_26_port,
                           input(25) => plus2A_out_25_port, input(24) => 
                           plus2A_out_24_port, input(23) => plus2A_out_23_port,
                           input(22) => plus2A_out_22_port, input(21) => 
                           plus2A_out_21_port, input(20) => plus2A_out_20_port,
                           input(19) => plus2A_out_19_port, input(18) => 
                           plus2A_out_18_port, input(17) => plus2A_out_17_port,
                           input(16) => plus2A_out_16_port, input(15) => 
                           plus2A_out_15_port, input(14) => plus2A_out_14_port,
                           input(13) => plus2A_out_13_port, input(12) => 
                           plus2A_out_12_port, input(11) => plus2A_out_11_port,
                           input(10) => plus2A_out_10_port, input(9) => 
                           plus2A_out_9_port, input(8) => plus2A_out_8_port, 
                           input(7) => plus2A_out_7_port, input(6) => 
                           plus2A_out_6_port, input(5) => plus2A_out_5_port, 
                           input(4) => plus2A_out_4_port, input(3) => 
                           plus2A_out_3_port, input(2) => plus2A_out_2_port, 
                           input(1) => plus2A_out_1_port, input(0) => 
                           plus2A_out_0_port, complement2(63) => 
                           minus2A_out(63), complement2(62) => minus2A_out(62),
                           complement2(61) => minus2A_out(61), complement2(60) 
                           => minus2A_out(60), complement2(59) => 
                           minus2A_out(59), complement2(58) => minus2A_out(58),
                           complement2(57) => minus2A_out(57), complement2(56) 
                           => minus2A_out(56), complement2(55) => 
                           minus2A_out(55), complement2(54) => minus2A_out(54),
                           complement2(53) => minus2A_out(53), complement2(52) 
                           => minus2A_out(52), complement2(51) => 
                           minus2A_out(51), complement2(50) => minus2A_out(50),
                           complement2(49) => minus2A_out(49), complement2(48) 
                           => minus2A_out(48), complement2(47) => 
                           minus2A_out(47), complement2(46) => minus2A_out(46),
                           complement2(45) => minus2A_out(45), complement2(44) 
                           => minus2A_out(44), complement2(43) => 
                           minus2A_out(43), complement2(42) => minus2A_out(42),
                           complement2(41) => minus2A_out(41), complement2(40) 
                           => minus2A_out(40), complement2(39) => 
                           minus2A_out(39), complement2(38) => minus2A_out(38),
                           complement2(37) => minus2A_out(37), complement2(36) 
                           => minus2A_out(36), complement2(35) => 
                           minus2A_out(35), complement2(34) => minus2A_out(34),
                           complement2(33) => minus2A_out(33), complement2(32) 
                           => minus2A_out(32), complement2(31) => 
                           minus2A_out(31), complement2(30) => minus2A_out(30),
                           complement2(29) => minus2A_out(29), complement2(28) 
                           => minus2A_out(28), complement2(27) => 
                           minus2A_out(27), complement2(26) => minus2A_out(26),
                           complement2(25) => minus2A_out(25), complement2(24) 
                           => minus2A_out(24), complement2(23) => 
                           minus2A_out(23), complement2(22) => minus2A_out(22),
                           complement2(21) => minus2A_out(21), complement2(20) 
                           => minus2A_out(20), complement2(19) => 
                           minus2A_out(19), complement2(18) => minus2A_out(18),
                           complement2(17) => minus2A_out(17), complement2(16) 
                           => minus2A_out(16), complement2(15) => 
                           minus2A_out(15), complement2(14) => minus2A_out(14),
                           complement2(13) => minus2A_out(13), complement2(12) 
                           => minus2A_out(12), complement2(11) => 
                           minus2A_out(11), complement2(10) => minus2A_out(10),
                           complement2(9) => minus2A_out(9), complement2(8) => 
                           minus2A_out(8), complement2(7) => minus2A_out(7), 
                           complement2(6) => minus2A_out(6), complement2(5) => 
                           minus2A_out(5), complement2(4) => minus2A_out(4), 
                           complement2(3) => minus2A_out(3), complement2(2) => 
                           minus2A_out(2), complement2(1) => minus2A_out(1), 
                           complement2(0) => minus2A_out(0));
   complementer_2 : complementer_N64_19 port map( input(63) => 
                           plus4A_out_63_port, input(62) => plus4A_out_62_port,
                           input(61) => plus4A_out_61_port, input(60) => 
                           plus4A_out_60_port, input(59) => plus4A_out_59_port,
                           input(58) => plus4A_out_58_port, input(57) => 
                           plus4A_out_57_port, input(56) => plus4A_out_56_port,
                           input(55) => plus4A_out_55_port, input(54) => 
                           plus4A_out_54_port, input(53) => plus4A_out_53_port,
                           input(52) => plus4A_out_52_port, input(51) => 
                           plus4A_out_51_port, input(50) => plus4A_out_50_port,
                           input(49) => plus4A_out_49_port, input(48) => 
                           plus4A_out_48_port, input(47) => plus4A_out_47_port,
                           input(46) => plus4A_out_46_port, input(45) => 
                           plus4A_out_45_port, input(44) => plus4A_out_44_port,
                           input(43) => plus4A_out_43_port, input(42) => 
                           plus4A_out_42_port, input(41) => plus4A_out_41_port,
                           input(40) => plus4A_out_40_port, input(39) => 
                           plus4A_out_39_port, input(38) => plus4A_out_38_port,
                           input(37) => plus4A_out_37_port, input(36) => 
                           plus4A_out_36_port, input(35) => plus4A_out_35_port,
                           input(34) => plus4A_out_34_port, input(33) => 
                           plus4A_out_33_port, input(32) => plus4A_out_32_port,
                           input(31) => plus4A_out_31_port, input(30) => 
                           plus4A_out_30_port, input(29) => plus4A_out_29_port,
                           input(28) => plus4A_out_28_port, input(27) => 
                           plus4A_out_27_port, input(26) => plus4A_out_26_port,
                           input(25) => plus4A_out_25_port, input(24) => 
                           plus4A_out_24_port, input(23) => plus4A_out_23_port,
                           input(22) => plus4A_out_22_port, input(21) => 
                           plus4A_out_21_port, input(20) => plus4A_out_20_port,
                           input(19) => plus4A_out_19_port, input(18) => 
                           plus4A_out_18_port, input(17) => plus4A_out_17_port,
                           input(16) => plus4A_out_16_port, input(15) => 
                           plus4A_out_15_port, input(14) => plus4A_out_14_port,
                           input(13) => plus4A_out_13_port, input(12) => 
                           plus4A_out_12_port, input(11) => plus4A_out_11_port,
                           input(10) => plus4A_out_10_port, input(9) => 
                           plus4A_out_9_port, input(8) => plus4A_out_8_port, 
                           input(7) => plus4A_out_7_port, input(6) => 
                           plus4A_out_6_port, input(5) => plus4A_out_5_port, 
                           input(4) => plus4A_out_4_port, input(3) => 
                           plus4A_out_3_port, input(2) => plus4A_out_2_port, 
                           input(1) => plus4A_out_1_port, input(0) => 
                           plus4A_out_0_port, complement2(63) => 
                           minus4A_out(63), complement2(62) => minus4A_out(62),
                           complement2(61) => minus4A_out(61), complement2(60) 
                           => minus4A_out(60), complement2(59) => 
                           minus4A_out(59), complement2(58) => minus4A_out(58),
                           complement2(57) => minus4A_out(57), complement2(56) 
                           => minus4A_out(56), complement2(55) => 
                           minus4A_out(55), complement2(54) => minus4A_out(54),
                           complement2(53) => minus4A_out(53), complement2(52) 
                           => minus4A_out(52), complement2(51) => 
                           minus4A_out(51), complement2(50) => minus4A_out(50),
                           complement2(49) => minus4A_out(49), complement2(48) 
                           => minus4A_out(48), complement2(47) => 
                           minus4A_out(47), complement2(46) => minus4A_out(46),
                           complement2(45) => minus4A_out(45), complement2(44) 
                           => minus4A_out(44), complement2(43) => 
                           minus4A_out(43), complement2(42) => minus4A_out(42),
                           complement2(41) => minus4A_out(41), complement2(40) 
                           => minus4A_out(40), complement2(39) => 
                           minus4A_out(39), complement2(38) => minus4A_out(38),
                           complement2(37) => minus4A_out(37), complement2(36) 
                           => minus4A_out(36), complement2(35) => 
                           minus4A_out(35), complement2(34) => minus4A_out(34),
                           complement2(33) => minus4A_out(33), complement2(32) 
                           => minus4A_out(32), complement2(31) => 
                           minus4A_out(31), complement2(30) => minus4A_out(30),
                           complement2(29) => minus4A_out(29), complement2(28) 
                           => minus4A_out(28), complement2(27) => 
                           minus4A_out(27), complement2(26) => minus4A_out(26),
                           complement2(25) => minus4A_out(25), complement2(24) 
                           => minus4A_out(24), complement2(23) => 
                           minus4A_out(23), complement2(22) => minus4A_out(22),
                           complement2(21) => minus4A_out(21), complement2(20) 
                           => minus4A_out(20), complement2(19) => 
                           minus4A_out(19), complement2(18) => minus4A_out(18),
                           complement2(17) => minus4A_out(17), complement2(16) 
                           => minus4A_out(16), complement2(15) => 
                           minus4A_out(15), complement2(14) => minus4A_out(14),
                           complement2(13) => minus4A_out(13), complement2(12) 
                           => minus4A_out(12), complement2(11) => 
                           minus4A_out(11), complement2(10) => minus4A_out(10),
                           complement2(9) => minus4A_out(9), complement2(8) => 
                           minus4A_out(8), complement2(7) => minus4A_out(7), 
                           complement2(6) => minus4A_out(6), complement2(5) => 
                           minus4A_out(5), complement2(4) => minus4A_out(4), 
                           complement2(3) => minus4A_out(3), complement2(2) => 
                           minus4A_out(2), complement2(1) => minus4A_out(1), 
                           complement2(0) => minus4A_out(0));
   U3 : CLKBUF_X1 port map( A => n65, Z => plus2A_out_15_port);
   U4 : CLKBUF_X1 port map( A => n63, Z => plus2A_out_17_port);
   U5 : CLKBUF_X1 port map( A => n67, Z => plus2A_out_13_port);
   U6 : CLKBUF_X1 port map( A => n66, Z => plus2A_out_14_port);
   U7 : BUF_X1 port map( A => n61, Z => plus2A_out_19_port);
   U8 : BUF_X1 port map( A => n62, Z => plus2A_out_18_port);
   U9 : BUF_X1 port map( A => n53, Z => plus2A_out_27_port);
   U10 : BUF_X1 port map( A => n51, Z => plus2A_out_29_port);
   U11 : BUF_X1 port map( A => n49, Z => plus2A_out_31_port);
   U12 : BUF_X1 port map( A => n57, Z => plus2A_out_23_port);
   U13 : BUF_X1 port map( A => n55, Z => plus2A_out_25_port);
   U14 : BUF_X1 port map( A => n59, Z => plus2A_out_21_port);
   U15 : BUF_X1 port map( A => n50, Z => plus2A_out_30_port);
   U16 : BUF_X1 port map( A => n54, Z => plus2A_out_26_port);
   U17 : BUF_X1 port map( A => n52, Z => plus2A_out_28_port);
   U18 : BUF_X1 port map( A => n58, Z => plus2A_out_22_port);
   U19 : BUF_X1 port map( A => n56, Z => plus2A_out_24_port);
   U20 : BUF_X1 port map( A => n60, Z => plus2A_out_20_port);
   U21 : BUF_X1 port map( A => n41, Z => plus2A_out_39_port);
   U22 : BUF_X1 port map( A => n39, Z => plus2A_out_41_port);
   U23 : BUF_X1 port map( A => n43, Z => plus2A_out_37_port);
   U24 : BUF_X1 port map( A => n45, Z => plus2A_out_35_port);
   U25 : BUF_X1 port map( A => n47, Z => plus2A_out_33_port);
   U26 : BUF_X1 port map( A => n42, Z => plus2A_out_38_port);
   U27 : BUF_X1 port map( A => n46, Z => plus2A_out_34_port);
   U28 : BUF_X1 port map( A => n40, Z => plus2A_out_40_port);
   U29 : BUF_X1 port map( A => n44, Z => plus2A_out_36_port);
   U30 : BUF_X1 port map( A => n48, Z => plus2A_out_32_port);
   U31 : BUF_X1 port map( A => n38, Z => plus2A_out_47_port);
   U32 : BUF_X1 port map( A => n70, Z => plus4A_out_52_port);
   U33 : BUF_X1 port map( A => n69, Z => plus4A_out_53_port);
   U34 : BUF_X1 port map( A => n37, Z => plus2A_out_48_port);
   U35 : BUF_X1 port map( A => n36, Z => plus2A_out_57_port);
   U36 : BUF_X1 port map( A => n68, Z => plus2A_out_12_port);
   U37 : BUF_X1 port map( A => n64, Z => plus2A_out_16_port);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity ShiftnCompl_N64_11 is

   port( plusA : in std_logic_vector (63 downto 0);  plus2A_out, minus2A_out, 
         plus4A_out, minus4A_out : out std_logic_vector (63 downto 0));

end ShiftnCompl_N64_11;

architecture SYN_struct of ShiftnCompl_N64_11 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component complementer_N64_21
      port( input : in std_logic_vector (63 downto 0);  complement2 : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component complementer_N64_22
      port( input : in std_logic_vector (63 downto 0);  complement2 : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component shifter_N64_21
      port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component shifter_N64_22
      port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
            std_logic_vector (63 downto 0));
   end component;
   
   signal plus2A_out_63_port, plus2A_out_62_port, plus2A_out_61_port, 
      plus2A_out_60_port, plus2A_out_59_port, plus2A_out_58_port, n9, 
      plus2A_out_56_port, plus2A_out_55_port, plus2A_out_54_port, 
      plus2A_out_53_port, plus2A_out_52_port, plus2A_out_51_port, 
      plus2A_out_50_port, plus2A_out_49_port, n10, n11, plus2A_out_46_port, 
      plus2A_out_45_port, plus2A_out_44_port, plus2A_out_43_port, 
      plus2A_out_42_port, plus2A_out_41_port, plus2A_out_40_port, 
      plus2A_out_39_port, plus2A_out_38_port, plus2A_out_37_port, 
      plus2A_out_36_port, plus2A_out_35_port, plus2A_out_34_port, 
      plus2A_out_33_port, plus2A_out_32_port, plus2A_out_31_port, 
      plus2A_out_30_port, plus2A_out_29_port, plus2A_out_28_port, 
      plus2A_out_27_port, plus2A_out_26_port, plus2A_out_25_port, 
      plus2A_out_24_port, plus2A_out_23_port, plus2A_out_22_port, 
      plus2A_out_21_port, plus2A_out_20_port, plus2A_out_19_port, 
      plus2A_out_18_port, plus2A_out_17_port, plus2A_out_16_port, 
      plus2A_out_15_port, plus2A_out_14_port, plus2A_out_13_port, 
      plus2A_out_12_port, plus2A_out_11_port, plus2A_out_10_port, 
      plus2A_out_9_port, plus2A_out_8_port, plus2A_out_7_port, 
      plus2A_out_6_port, plus2A_out_5_port, plus2A_out_4_port, 
      plus2A_out_3_port, plus2A_out_2_port, plus2A_out_1_port, 
      plus2A_out_0_port, plus4A_out_63_port, plus4A_out_62_port, 
      plus4A_out_61_port, plus4A_out_60_port, plus4A_out_59_port, 
      plus4A_out_58_port, plus4A_out_57_port, plus4A_out_56_port, 
      plus4A_out_55_port, plus4A_out_54_port, n12, n13, plus4A_out_51_port, 
      plus4A_out_50_port, plus4A_out_49_port, plus4A_out_48_port, 
      plus4A_out_47_port, plus4A_out_46_port, plus4A_out_45_port, 
      plus4A_out_44_port, n14, n15, n16, plus4A_out_40_port, plus4A_out_39_port
      , plus4A_out_38_port, plus4A_out_37_port, plus4A_out_36_port, 
      plus4A_out_35_port, plus4A_out_34_port, plus4A_out_33_port, 
      plus4A_out_32_port, plus4A_out_31_port, plus4A_out_30_port, 
      plus4A_out_29_port, plus4A_out_28_port, plus4A_out_27_port, 
      plus4A_out_26_port, plus4A_out_25_port, plus4A_out_24_port, 
      plus4A_out_23_port, plus4A_out_22_port, plus4A_out_21_port, 
      plus4A_out_20_port, plus4A_out_19_port, plus4A_out_18_port, 
      plus4A_out_17_port, plus4A_out_16_port, plus4A_out_15_port, 
      plus4A_out_14_port, plus4A_out_13_port, plus4A_out_12_port, 
      plus4A_out_11_port, plus4A_out_10_port, plus4A_out_9_port, 
      plus4A_out_8_port, plus4A_out_7_port, plus4A_out_6_port, 
      plus4A_out_5_port, plus4A_out_4_port, plus4A_out_3_port, 
      plus4A_out_2_port, plus4A_out_1_port, plus4A_out_0_port, 
      plus4A_out_41_port, plus4A_out_42_port, plus4A_out_43_port, 
      plus2A_out_47_port, plus2A_out_48_port, plus4A_out_52_port, 
      plus4A_out_53_port, plus2A_out_57_port, n_3164, n_3165 : std_logic;

begin
   plus2A_out <= ( plus2A_out_63_port, plus2A_out_62_port, plus2A_out_61_port, 
      plus2A_out_60_port, plus2A_out_59_port, plus2A_out_58_port, 
      plus2A_out_57_port, plus2A_out_56_port, plus2A_out_55_port, 
      plus2A_out_54_port, plus2A_out_53_port, plus2A_out_52_port, 
      plus2A_out_51_port, plus2A_out_50_port, plus2A_out_49_port, 
      plus2A_out_48_port, plus2A_out_47_port, plus2A_out_46_port, 
      plus2A_out_45_port, plus2A_out_44_port, plus2A_out_43_port, 
      plus2A_out_42_port, plus2A_out_41_port, plus2A_out_40_port, 
      plus2A_out_39_port, plus2A_out_38_port, plus2A_out_37_port, 
      plus2A_out_36_port, plus2A_out_35_port, plus2A_out_34_port, 
      plus2A_out_33_port, plus2A_out_32_port, plus2A_out_31_port, 
      plus2A_out_30_port, plus2A_out_29_port, plus2A_out_28_port, 
      plus2A_out_27_port, plus2A_out_26_port, plus2A_out_25_port, 
      plus2A_out_24_port, plus2A_out_23_port, plus2A_out_22_port, 
      plus2A_out_21_port, plus2A_out_20_port, plus2A_out_19_port, 
      plus2A_out_18_port, plus2A_out_17_port, plus2A_out_16_port, 
      plus2A_out_15_port, plus2A_out_14_port, plus2A_out_13_port, 
      plus2A_out_12_port, plus2A_out_11_port, plus2A_out_10_port, 
      plus2A_out_9_port, plus2A_out_8_port, plus2A_out_7_port, 
      plus2A_out_6_port, plus2A_out_5_port, plus2A_out_4_port, 
      plus2A_out_3_port, plus2A_out_2_port, plus2A_out_1_port, 
      plus2A_out_0_port );
   plus4A_out <= ( plus4A_out_63_port, plus4A_out_62_port, plus4A_out_61_port, 
      plus4A_out_60_port, plus4A_out_59_port, plus4A_out_58_port, 
      plus4A_out_57_port, plus4A_out_56_port, plus4A_out_55_port, 
      plus4A_out_54_port, plus4A_out_53_port, plus4A_out_52_port, 
      plus4A_out_51_port, plus4A_out_50_port, plus4A_out_49_port, 
      plus4A_out_48_port, plus4A_out_47_port, plus4A_out_46_port, 
      plus4A_out_45_port, plus4A_out_44_port, plus4A_out_43_port, 
      plus4A_out_42_port, plus4A_out_41_port, plus4A_out_40_port, 
      plus4A_out_39_port, plus4A_out_38_port, plus4A_out_37_port, 
      plus4A_out_36_port, plus4A_out_35_port, plus4A_out_34_port, 
      plus4A_out_33_port, plus4A_out_32_port, plus4A_out_31_port, 
      plus4A_out_30_port, plus4A_out_29_port, plus4A_out_28_port, 
      plus4A_out_27_port, plus4A_out_26_port, plus4A_out_25_port, 
      plus4A_out_24_port, plus4A_out_23_port, plus4A_out_22_port, 
      plus4A_out_21_port, plus4A_out_20_port, plus4A_out_19_port, 
      plus4A_out_18_port, plus4A_out_17_port, plus4A_out_16_port, 
      plus4A_out_15_port, plus4A_out_14_port, plus4A_out_13_port, 
      plus4A_out_12_port, plus4A_out_11_port, plus4A_out_10_port, 
      plus4A_out_9_port, plus4A_out_8_port, plus4A_out_7_port, 
      plus4A_out_6_port, plus4A_out_5_port, plus4A_out_4_port, 
      plus4A_out_3_port, plus4A_out_2_port, plus4A_out_1_port, 
      plus4A_out_0_port );
   
   plus2A_out_0_port <= '0';
   plus4A_out_0_port <= '0';
   shifter_1 : shifter_N64_22 port map( input(63) => plusA(63), input(62) => 
                           plusA(62), input(61) => plusA(61), input(60) => 
                           plusA(60), input(59) => plusA(59), input(58) => 
                           plusA(58), input(57) => plusA(57), input(56) => 
                           plusA(56), input(55) => plusA(55), input(54) => 
                           plusA(54), input(53) => plusA(53), input(52) => 
                           plusA(52), input(51) => plusA(51), input(50) => 
                           plusA(50), input(49) => plusA(49), input(48) => 
                           plusA(48), input(47) => plusA(47), input(46) => 
                           plusA(46), input(45) => plusA(45), input(44) => 
                           plusA(44), input(43) => plusA(43), input(42) => 
                           plusA(42), input(41) => plusA(41), input(40) => 
                           plusA(40), input(39) => plusA(39), input(38) => 
                           plusA(38), input(37) => plusA(37), input(36) => 
                           plusA(36), input(35) => plusA(35), input(34) => 
                           plusA(34), input(33) => plusA(33), input(32) => 
                           plusA(32), input(31) => plusA(31), input(30) => 
                           plusA(30), input(29) => plusA(29), input(28) => 
                           plusA(28), input(27) => plusA(27), input(26) => 
                           plusA(26), input(25) => plusA(25), input(24) => 
                           plusA(24), input(23) => plusA(23), input(22) => 
                           plusA(22), input(21) => plusA(21), input(20) => 
                           plusA(20), input(19) => plusA(19), input(18) => 
                           plusA(18), input(17) => plusA(17), input(16) => 
                           plusA(16), input(15) => plusA(15), input(14) => 
                           plusA(14), input(13) => plusA(13), input(12) => 
                           plusA(12), input(11) => plusA(11), input(10) => 
                           plusA(10), input(9) => plusA(9), input(8) => 
                           plusA(8), input(7) => plusA(7), input(6) => plusA(6)
                           , input(5) => plusA(5), input(4) => plusA(4), 
                           input(3) => plusA(3), input(2) => plusA(2), input(1)
                           => plusA(1), input(0) => plusA(0), 
                           shiftLeftOnePos(63) => plus2A_out_63_port, 
                           shiftLeftOnePos(62) => plus2A_out_62_port, 
                           shiftLeftOnePos(61) => plus2A_out_61_port, 
                           shiftLeftOnePos(60) => plus2A_out_60_port, 
                           shiftLeftOnePos(59) => plus2A_out_59_port, 
                           shiftLeftOnePos(58) => plus2A_out_58_port, 
                           shiftLeftOnePos(57) => n9, shiftLeftOnePos(56) => 
                           plus2A_out_56_port, shiftLeftOnePos(55) => 
                           plus2A_out_55_port, shiftLeftOnePos(54) => 
                           plus2A_out_54_port, shiftLeftOnePos(53) => 
                           plus2A_out_53_port, shiftLeftOnePos(52) => 
                           plus2A_out_52_port, shiftLeftOnePos(51) => 
                           plus2A_out_51_port, shiftLeftOnePos(50) => 
                           plus2A_out_50_port, shiftLeftOnePos(49) => 
                           plus2A_out_49_port, shiftLeftOnePos(48) => n10, 
                           shiftLeftOnePos(47) => n11, shiftLeftOnePos(46) => 
                           plus2A_out_46_port, shiftLeftOnePos(45) => 
                           plus2A_out_45_port, shiftLeftOnePos(44) => 
                           plus2A_out_44_port, shiftLeftOnePos(43) => 
                           plus2A_out_43_port, shiftLeftOnePos(42) => 
                           plus2A_out_42_port, shiftLeftOnePos(41) => 
                           plus2A_out_41_port, shiftLeftOnePos(40) => 
                           plus2A_out_40_port, shiftLeftOnePos(39) => 
                           plus2A_out_39_port, shiftLeftOnePos(38) => 
                           plus2A_out_38_port, shiftLeftOnePos(37) => 
                           plus2A_out_37_port, shiftLeftOnePos(36) => 
                           plus2A_out_36_port, shiftLeftOnePos(35) => 
                           plus2A_out_35_port, shiftLeftOnePos(34) => 
                           plus2A_out_34_port, shiftLeftOnePos(33) => 
                           plus2A_out_33_port, shiftLeftOnePos(32) => 
                           plus2A_out_32_port, shiftLeftOnePos(31) => 
                           plus2A_out_31_port, shiftLeftOnePos(30) => 
                           plus2A_out_30_port, shiftLeftOnePos(29) => 
                           plus2A_out_29_port, shiftLeftOnePos(28) => 
                           plus2A_out_28_port, shiftLeftOnePos(27) => 
                           plus2A_out_27_port, shiftLeftOnePos(26) => 
                           plus2A_out_26_port, shiftLeftOnePos(25) => 
                           plus2A_out_25_port, shiftLeftOnePos(24) => 
                           plus2A_out_24_port, shiftLeftOnePos(23) => 
                           plus2A_out_23_port, shiftLeftOnePos(22) => 
                           plus2A_out_22_port, shiftLeftOnePos(21) => 
                           plus2A_out_21_port, shiftLeftOnePos(20) => 
                           plus2A_out_20_port, shiftLeftOnePos(19) => 
                           plus2A_out_19_port, shiftLeftOnePos(18) => 
                           plus2A_out_18_port, shiftLeftOnePos(17) => 
                           plus2A_out_17_port, shiftLeftOnePos(16) => 
                           plus2A_out_16_port, shiftLeftOnePos(15) => 
                           plus2A_out_15_port, shiftLeftOnePos(14) => 
                           plus2A_out_14_port, shiftLeftOnePos(13) => 
                           plus2A_out_13_port, shiftLeftOnePos(12) => 
                           plus2A_out_12_port, shiftLeftOnePos(11) => 
                           plus2A_out_11_port, shiftLeftOnePos(10) => 
                           plus2A_out_10_port, shiftLeftOnePos(9) => 
                           plus2A_out_9_port, shiftLeftOnePos(8) => 
                           plus2A_out_8_port, shiftLeftOnePos(7) => 
                           plus2A_out_7_port, shiftLeftOnePos(6) => 
                           plus2A_out_6_port, shiftLeftOnePos(5) => 
                           plus2A_out_5_port, shiftLeftOnePos(4) => 
                           plus2A_out_4_port, shiftLeftOnePos(3) => 
                           plus2A_out_3_port, shiftLeftOnePos(2) => 
                           plus2A_out_2_port, shiftLeftOnePos(1) => 
                           plus2A_out_1_port, shiftLeftOnePos(0) => n_3164);
   shifter_2 : shifter_N64_21 port map( input(63) => plus2A_out_63_port, 
                           input(62) => plus2A_out_62_port, input(61) => 
                           plus2A_out_61_port, input(60) => plus2A_out_60_port,
                           input(59) => plus2A_out_59_port, input(58) => 
                           plus2A_out_58_port, input(57) => plus2A_out_57_port,
                           input(56) => plus2A_out_56_port, input(55) => 
                           plus2A_out_55_port, input(54) => plus2A_out_54_port,
                           input(53) => plus2A_out_53_port, input(52) => 
                           plus2A_out_52_port, input(51) => plus2A_out_51_port,
                           input(50) => plus2A_out_50_port, input(49) => 
                           plus2A_out_49_port, input(48) => plus2A_out_48_port,
                           input(47) => plus2A_out_47_port, input(46) => 
                           plus2A_out_46_port, input(45) => plus2A_out_45_port,
                           input(44) => plus2A_out_44_port, input(43) => 
                           plus2A_out_43_port, input(42) => plus2A_out_42_port,
                           input(41) => plus2A_out_41_port, input(40) => 
                           plus2A_out_40_port, input(39) => plus2A_out_39_port,
                           input(38) => plus2A_out_38_port, input(37) => 
                           plus2A_out_37_port, input(36) => plus2A_out_36_port,
                           input(35) => plus2A_out_35_port, input(34) => 
                           plus2A_out_34_port, input(33) => plus2A_out_33_port,
                           input(32) => plus2A_out_32_port, input(31) => 
                           plus2A_out_31_port, input(30) => plus2A_out_30_port,
                           input(29) => plus2A_out_29_port, input(28) => 
                           plus2A_out_28_port, input(27) => plus2A_out_27_port,
                           input(26) => plus2A_out_26_port, input(25) => 
                           plus2A_out_25_port, input(24) => plus2A_out_24_port,
                           input(23) => plus2A_out_23_port, input(22) => 
                           plus2A_out_22_port, input(21) => plus2A_out_21_port,
                           input(20) => plus2A_out_20_port, input(19) => 
                           plus2A_out_19_port, input(18) => plus2A_out_18_port,
                           input(17) => plus2A_out_17_port, input(16) => 
                           plus2A_out_16_port, input(15) => plus2A_out_15_port,
                           input(14) => plus2A_out_14_port, input(13) => 
                           plus2A_out_13_port, input(12) => plus2A_out_12_port,
                           input(11) => plus2A_out_11_port, input(10) => 
                           plus2A_out_10_port, input(9) => plus2A_out_9_port, 
                           input(8) => plus2A_out_8_port, input(7) => 
                           plus2A_out_7_port, input(6) => plus2A_out_6_port, 
                           input(5) => plus2A_out_5_port, input(4) => 
                           plus2A_out_4_port, input(3) => plus2A_out_3_port, 
                           input(2) => plus2A_out_2_port, input(1) => 
                           plus2A_out_1_port, input(0) => plus2A_out_0_port, 
                           shiftLeftOnePos(63) => plus4A_out_63_port, 
                           shiftLeftOnePos(62) => plus4A_out_62_port, 
                           shiftLeftOnePos(61) => plus4A_out_61_port, 
                           shiftLeftOnePos(60) => plus4A_out_60_port, 
                           shiftLeftOnePos(59) => plus4A_out_59_port, 
                           shiftLeftOnePos(58) => plus4A_out_58_port, 
                           shiftLeftOnePos(57) => plus4A_out_57_port, 
                           shiftLeftOnePos(56) => plus4A_out_56_port, 
                           shiftLeftOnePos(55) => plus4A_out_55_port, 
                           shiftLeftOnePos(54) => plus4A_out_54_port, 
                           shiftLeftOnePos(53) => n12, shiftLeftOnePos(52) => 
                           n13, shiftLeftOnePos(51) => plus4A_out_51_port, 
                           shiftLeftOnePos(50) => plus4A_out_50_port, 
                           shiftLeftOnePos(49) => plus4A_out_49_port, 
                           shiftLeftOnePos(48) => plus4A_out_48_port, 
                           shiftLeftOnePos(47) => plus4A_out_47_port, 
                           shiftLeftOnePos(46) => plus4A_out_46_port, 
                           shiftLeftOnePos(45) => plus4A_out_45_port, 
                           shiftLeftOnePos(44) => plus4A_out_44_port, 
                           shiftLeftOnePos(43) => n14, shiftLeftOnePos(42) => 
                           n15, shiftLeftOnePos(41) => n16, shiftLeftOnePos(40)
                           => plus4A_out_40_port, shiftLeftOnePos(39) => 
                           plus4A_out_39_port, shiftLeftOnePos(38) => 
                           plus4A_out_38_port, shiftLeftOnePos(37) => 
                           plus4A_out_37_port, shiftLeftOnePos(36) => 
                           plus4A_out_36_port, shiftLeftOnePos(35) => 
                           plus4A_out_35_port, shiftLeftOnePos(34) => 
                           plus4A_out_34_port, shiftLeftOnePos(33) => 
                           plus4A_out_33_port, shiftLeftOnePos(32) => 
                           plus4A_out_32_port, shiftLeftOnePos(31) => 
                           plus4A_out_31_port, shiftLeftOnePos(30) => 
                           plus4A_out_30_port, shiftLeftOnePos(29) => 
                           plus4A_out_29_port, shiftLeftOnePos(28) => 
                           plus4A_out_28_port, shiftLeftOnePos(27) => 
                           plus4A_out_27_port, shiftLeftOnePos(26) => 
                           plus4A_out_26_port, shiftLeftOnePos(25) => 
                           plus4A_out_25_port, shiftLeftOnePos(24) => 
                           plus4A_out_24_port, shiftLeftOnePos(23) => 
                           plus4A_out_23_port, shiftLeftOnePos(22) => 
                           plus4A_out_22_port, shiftLeftOnePos(21) => 
                           plus4A_out_21_port, shiftLeftOnePos(20) => 
                           plus4A_out_20_port, shiftLeftOnePos(19) => 
                           plus4A_out_19_port, shiftLeftOnePos(18) => 
                           plus4A_out_18_port, shiftLeftOnePos(17) => 
                           plus4A_out_17_port, shiftLeftOnePos(16) => 
                           plus4A_out_16_port, shiftLeftOnePos(15) => 
                           plus4A_out_15_port, shiftLeftOnePos(14) => 
                           plus4A_out_14_port, shiftLeftOnePos(13) => 
                           plus4A_out_13_port, shiftLeftOnePos(12) => 
                           plus4A_out_12_port, shiftLeftOnePos(11) => 
                           plus4A_out_11_port, shiftLeftOnePos(10) => 
                           plus4A_out_10_port, shiftLeftOnePos(9) => 
                           plus4A_out_9_port, shiftLeftOnePos(8) => 
                           plus4A_out_8_port, shiftLeftOnePos(7) => 
                           plus4A_out_7_port, shiftLeftOnePos(6) => 
                           plus4A_out_6_port, shiftLeftOnePos(5) => 
                           plus4A_out_5_port, shiftLeftOnePos(4) => 
                           plus4A_out_4_port, shiftLeftOnePos(3) => 
                           plus4A_out_3_port, shiftLeftOnePos(2) => 
                           plus4A_out_2_port, shiftLeftOnePos(1) => 
                           plus4A_out_1_port, shiftLeftOnePos(0) => n_3165);
   complementer_1 : complementer_N64_22 port map( input(63) => 
                           plus2A_out_63_port, input(62) => plus2A_out_62_port,
                           input(61) => plus2A_out_61_port, input(60) => 
                           plus2A_out_60_port, input(59) => plus2A_out_59_port,
                           input(58) => plus2A_out_58_port, input(57) => 
                           plus2A_out_57_port, input(56) => plus2A_out_56_port,
                           input(55) => plus2A_out_55_port, input(54) => 
                           plus2A_out_54_port, input(53) => plus2A_out_53_port,
                           input(52) => plus2A_out_52_port, input(51) => 
                           plus2A_out_51_port, input(50) => plus2A_out_50_port,
                           input(49) => plus2A_out_49_port, input(48) => 
                           plus2A_out_48_port, input(47) => plus2A_out_47_port,
                           input(46) => plus2A_out_46_port, input(45) => 
                           plus2A_out_45_port, input(44) => plus2A_out_44_port,
                           input(43) => plus2A_out_43_port, input(42) => 
                           plus2A_out_42_port, input(41) => plus2A_out_41_port,
                           input(40) => plus2A_out_40_port, input(39) => 
                           plus2A_out_39_port, input(38) => plus2A_out_38_port,
                           input(37) => plus2A_out_37_port, input(36) => 
                           plus2A_out_36_port, input(35) => plus2A_out_35_port,
                           input(34) => plus2A_out_34_port, input(33) => 
                           plus2A_out_33_port, input(32) => plus2A_out_32_port,
                           input(31) => plus2A_out_31_port, input(30) => 
                           plus2A_out_30_port, input(29) => plus2A_out_29_port,
                           input(28) => plus2A_out_28_port, input(27) => 
                           plus2A_out_27_port, input(26) => plus2A_out_26_port,
                           input(25) => plus2A_out_25_port, input(24) => 
                           plus2A_out_24_port, input(23) => plus2A_out_23_port,
                           input(22) => plus2A_out_22_port, input(21) => 
                           plus2A_out_21_port, input(20) => plus2A_out_20_port,
                           input(19) => plus2A_out_19_port, input(18) => 
                           plus2A_out_18_port, input(17) => plus2A_out_17_port,
                           input(16) => plus2A_out_16_port, input(15) => 
                           plus2A_out_15_port, input(14) => plus2A_out_14_port,
                           input(13) => plus2A_out_13_port, input(12) => 
                           plus2A_out_12_port, input(11) => plus2A_out_11_port,
                           input(10) => plus2A_out_10_port, input(9) => 
                           plus2A_out_9_port, input(8) => plus2A_out_8_port, 
                           input(7) => plus2A_out_7_port, input(6) => 
                           plus2A_out_6_port, input(5) => plus2A_out_5_port, 
                           input(4) => plus2A_out_4_port, input(3) => 
                           plus2A_out_3_port, input(2) => plus2A_out_2_port, 
                           input(1) => plus2A_out_1_port, input(0) => 
                           plus2A_out_0_port, complement2(63) => 
                           minus2A_out(63), complement2(62) => minus2A_out(62),
                           complement2(61) => minus2A_out(61), complement2(60) 
                           => minus2A_out(60), complement2(59) => 
                           minus2A_out(59), complement2(58) => minus2A_out(58),
                           complement2(57) => minus2A_out(57), complement2(56) 
                           => minus2A_out(56), complement2(55) => 
                           minus2A_out(55), complement2(54) => minus2A_out(54),
                           complement2(53) => minus2A_out(53), complement2(52) 
                           => minus2A_out(52), complement2(51) => 
                           minus2A_out(51), complement2(50) => minus2A_out(50),
                           complement2(49) => minus2A_out(49), complement2(48) 
                           => minus2A_out(48), complement2(47) => 
                           minus2A_out(47), complement2(46) => minus2A_out(46),
                           complement2(45) => minus2A_out(45), complement2(44) 
                           => minus2A_out(44), complement2(43) => 
                           minus2A_out(43), complement2(42) => minus2A_out(42),
                           complement2(41) => minus2A_out(41), complement2(40) 
                           => minus2A_out(40), complement2(39) => 
                           minus2A_out(39), complement2(38) => minus2A_out(38),
                           complement2(37) => minus2A_out(37), complement2(36) 
                           => minus2A_out(36), complement2(35) => 
                           minus2A_out(35), complement2(34) => minus2A_out(34),
                           complement2(33) => minus2A_out(33), complement2(32) 
                           => minus2A_out(32), complement2(31) => 
                           minus2A_out(31), complement2(30) => minus2A_out(30),
                           complement2(29) => minus2A_out(29), complement2(28) 
                           => minus2A_out(28), complement2(27) => 
                           minus2A_out(27), complement2(26) => minus2A_out(26),
                           complement2(25) => minus2A_out(25), complement2(24) 
                           => minus2A_out(24), complement2(23) => 
                           minus2A_out(23), complement2(22) => minus2A_out(22),
                           complement2(21) => minus2A_out(21), complement2(20) 
                           => minus2A_out(20), complement2(19) => 
                           minus2A_out(19), complement2(18) => minus2A_out(18),
                           complement2(17) => minus2A_out(17), complement2(16) 
                           => minus2A_out(16), complement2(15) => 
                           minus2A_out(15), complement2(14) => minus2A_out(14),
                           complement2(13) => minus2A_out(13), complement2(12) 
                           => minus2A_out(12), complement2(11) => 
                           minus2A_out(11), complement2(10) => minus2A_out(10),
                           complement2(9) => minus2A_out(9), complement2(8) => 
                           minus2A_out(8), complement2(7) => minus2A_out(7), 
                           complement2(6) => minus2A_out(6), complement2(5) => 
                           minus2A_out(5), complement2(4) => minus2A_out(4), 
                           complement2(3) => minus2A_out(3), complement2(2) => 
                           minus2A_out(2), complement2(1) => minus2A_out(1), 
                           complement2(0) => minus2A_out(0));
   complementer_2 : complementer_N64_21 port map( input(63) => 
                           plus4A_out_63_port, input(62) => plus4A_out_62_port,
                           input(61) => plus4A_out_61_port, input(60) => 
                           plus4A_out_60_port, input(59) => plus4A_out_59_port,
                           input(58) => plus4A_out_58_port, input(57) => 
                           plus4A_out_57_port, input(56) => plus4A_out_56_port,
                           input(55) => plus4A_out_55_port, input(54) => 
                           plus4A_out_54_port, input(53) => plus4A_out_53_port,
                           input(52) => plus4A_out_52_port, input(51) => 
                           plus4A_out_51_port, input(50) => plus4A_out_50_port,
                           input(49) => plus4A_out_49_port, input(48) => 
                           plus4A_out_48_port, input(47) => plus4A_out_47_port,
                           input(46) => plus4A_out_46_port, input(45) => 
                           plus4A_out_45_port, input(44) => plus4A_out_44_port,
                           input(43) => plus4A_out_43_port, input(42) => 
                           plus4A_out_42_port, input(41) => plus4A_out_41_port,
                           input(40) => plus4A_out_40_port, input(39) => 
                           plus4A_out_39_port, input(38) => plus4A_out_38_port,
                           input(37) => plus4A_out_37_port, input(36) => 
                           plus4A_out_36_port, input(35) => plus4A_out_35_port,
                           input(34) => plus4A_out_34_port, input(33) => 
                           plus4A_out_33_port, input(32) => plus4A_out_32_port,
                           input(31) => plus4A_out_31_port, input(30) => 
                           plus4A_out_30_port, input(29) => plus4A_out_29_port,
                           input(28) => plus4A_out_28_port, input(27) => 
                           plus4A_out_27_port, input(26) => plus4A_out_26_port,
                           input(25) => plus4A_out_25_port, input(24) => 
                           plus4A_out_24_port, input(23) => plus4A_out_23_port,
                           input(22) => plus4A_out_22_port, input(21) => 
                           plus4A_out_21_port, input(20) => plus4A_out_20_port,
                           input(19) => plus4A_out_19_port, input(18) => 
                           plus4A_out_18_port, input(17) => plus4A_out_17_port,
                           input(16) => plus4A_out_16_port, input(15) => 
                           plus4A_out_15_port, input(14) => plus4A_out_14_port,
                           input(13) => plus4A_out_13_port, input(12) => 
                           plus4A_out_12_port, input(11) => plus4A_out_11_port,
                           input(10) => plus4A_out_10_port, input(9) => 
                           plus4A_out_9_port, input(8) => plus4A_out_8_port, 
                           input(7) => plus4A_out_7_port, input(6) => 
                           plus4A_out_6_port, input(5) => plus4A_out_5_port, 
                           input(4) => plus4A_out_4_port, input(3) => 
                           plus4A_out_3_port, input(2) => plus4A_out_2_port, 
                           input(1) => plus4A_out_1_port, input(0) => 
                           plus4A_out_0_port, complement2(63) => 
                           minus4A_out(63), complement2(62) => minus4A_out(62),
                           complement2(61) => minus4A_out(61), complement2(60) 
                           => minus4A_out(60), complement2(59) => 
                           minus4A_out(59), complement2(58) => minus4A_out(58),
                           complement2(57) => minus4A_out(57), complement2(56) 
                           => minus4A_out(56), complement2(55) => 
                           minus4A_out(55), complement2(54) => minus4A_out(54),
                           complement2(53) => minus4A_out(53), complement2(52) 
                           => minus4A_out(52), complement2(51) => 
                           minus4A_out(51), complement2(50) => minus4A_out(50),
                           complement2(49) => minus4A_out(49), complement2(48) 
                           => minus4A_out(48), complement2(47) => 
                           minus4A_out(47), complement2(46) => minus4A_out(46),
                           complement2(45) => minus4A_out(45), complement2(44) 
                           => minus4A_out(44), complement2(43) => 
                           minus4A_out(43), complement2(42) => minus4A_out(42),
                           complement2(41) => minus4A_out(41), complement2(40) 
                           => minus4A_out(40), complement2(39) => 
                           minus4A_out(39), complement2(38) => minus4A_out(38),
                           complement2(37) => minus4A_out(37), complement2(36) 
                           => minus4A_out(36), complement2(35) => 
                           minus4A_out(35), complement2(34) => minus4A_out(34),
                           complement2(33) => minus4A_out(33), complement2(32) 
                           => minus4A_out(32), complement2(31) => 
                           minus4A_out(31), complement2(30) => minus4A_out(30),
                           complement2(29) => minus4A_out(29), complement2(28) 
                           => minus4A_out(28), complement2(27) => 
                           minus4A_out(27), complement2(26) => minus4A_out(26),
                           complement2(25) => minus4A_out(25), complement2(24) 
                           => minus4A_out(24), complement2(23) => 
                           minus4A_out(23), complement2(22) => minus4A_out(22),
                           complement2(21) => minus4A_out(21), complement2(20) 
                           => minus4A_out(20), complement2(19) => 
                           minus4A_out(19), complement2(18) => minus4A_out(18),
                           complement2(17) => minus4A_out(17), complement2(16) 
                           => minus4A_out(16), complement2(15) => 
                           minus4A_out(15), complement2(14) => minus4A_out(14),
                           complement2(13) => minus4A_out(13), complement2(12) 
                           => minus4A_out(12), complement2(11) => 
                           minus4A_out(11), complement2(10) => minus4A_out(10),
                           complement2(9) => minus4A_out(9), complement2(8) => 
                           minus4A_out(8), complement2(7) => minus4A_out(7), 
                           complement2(6) => minus4A_out(6), complement2(5) => 
                           minus4A_out(5), complement2(4) => minus4A_out(4), 
                           complement2(3) => minus4A_out(3), complement2(2) => 
                           minus4A_out(2), complement2(1) => minus4A_out(1), 
                           complement2(0) => minus4A_out(0));
   U3 : BUF_X1 port map( A => n14, Z => plus4A_out_43_port);
   U4 : BUF_X1 port map( A => n16, Z => plus4A_out_41_port);
   U5 : BUF_X1 port map( A => n15, Z => plus4A_out_42_port);
   U6 : BUF_X1 port map( A => n11, Z => plus2A_out_47_port);
   U7 : BUF_X1 port map( A => n13, Z => plus4A_out_52_port);
   U8 : BUF_X1 port map( A => n10, Z => plus2A_out_48_port);
   U9 : BUF_X1 port map( A => n12, Z => plus4A_out_53_port);
   U10 : BUF_X1 port map( A => n9, Z => plus2A_out_57_port);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity MUX_GENERIC_N64_RADIX3_12 is

   port( plusA, minusA, plus2A, minus2A : in std_logic_vector (63 downto 0);  
         SEL : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (63 
         downto 0));

end MUX_GENERIC_N64_RADIX3_12;

architecture SYN_beh of MUX_GENERIC_N64_RADIX3_12 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component TBUF_X1
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   signal n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, 
      n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, 
      n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, 
      n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, 
      n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, 
      n266, n267, n268, n269, n270, n271, n4, n5, n6, n7, n8, n9, n10, n11, n12
      , n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, 
      n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41
      , n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, 
      n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70
      , n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, 
      n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99
      , n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
      n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, 
      n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, 
      n136, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, 
      n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, 
      n295, n296, n297, n298, n299, n300, n301, n302, n303, n304 : std_logic;

begin
   
   Y_tri_60_inst : TBUF_X1 port map( A => n268, EN => n301, Z => Y(60));
   Y_tri_61_inst : TBUF_X1 port map( A => n269, EN => n301, Z => Y(61));
   Y_tri_62_inst : TBUF_X1 port map( A => n270, EN => n301, Z => Y(62));
   Y_tri_63_inst : TBUF_X1 port map( A => n271, EN => n301, Z => Y(63));
   Y_tri_48_inst : TBUF_X1 port map( A => n256, EN => n300, Z => Y(48));
   Y_tri_49_inst : TBUF_X1 port map( A => n257, EN => n300, Z => Y(49));
   Y_tri_50_inst : TBUF_X1 port map( A => n258, EN => n300, Z => Y(50));
   Y_tri_51_inst : TBUF_X1 port map( A => n259, EN => n300, Z => Y(51));
   Y_tri_52_inst : TBUF_X1 port map( A => n260, EN => n300, Z => Y(52));
   Y_tri_53_inst : TBUF_X1 port map( A => n261, EN => n300, Z => Y(53));
   Y_tri_54_inst : TBUF_X1 port map( A => n262, EN => n300, Z => Y(54));
   Y_tri_55_inst : TBUF_X1 port map( A => n263, EN => n300, Z => Y(55));
   Y_tri_56_inst : TBUF_X1 port map( A => n264, EN => n300, Z => Y(56));
   Y_tri_57_inst : TBUF_X1 port map( A => n265, EN => n300, Z => Y(57));
   Y_tri_58_inst : TBUF_X1 port map( A => n266, EN => n300, Z => Y(58));
   Y_tri_59_inst : TBUF_X1 port map( A => n267, EN => n300, Z => Y(59));
   Y_tri_27_inst : TBUF_X1 port map( A => n235, EN => n298, Z => Y(27));
   Y_tri_28_inst : TBUF_X1 port map( A => n236, EN => n298, Z => Y(28));
   Y_tri_29_inst : TBUF_X1 port map( A => n237, EN => n298, Z => Y(29));
   Y_tri_30_inst : TBUF_X1 port map( A => n238, EN => n298, Z => Y(30));
   Y_tri_31_inst : TBUF_X1 port map( A => n239, EN => n298, Z => Y(31));
   Y_tri_32_inst : TBUF_X1 port map( A => n240, EN => n298, Z => Y(32));
   Y_tri_33_inst : TBUF_X1 port map( A => n241, EN => n298, Z => Y(33));
   Y_tri_34_inst : TBUF_X1 port map( A => n242, EN => n298, Z => Y(34));
   Y_tri_35_inst : TBUF_X1 port map( A => n243, EN => n298, Z => Y(35));
   Y_tri_36_inst : TBUF_X1 port map( A => n244, EN => n299, Z => Y(36));
   Y_tri_37_inst : TBUF_X1 port map( A => n245, EN => n299, Z => Y(37));
   Y_tri_38_inst : TBUF_X1 port map( A => n246, EN => n299, Z => Y(38));
   Y_tri_39_inst : TBUF_X1 port map( A => n247, EN => n299, Z => Y(39));
   Y_tri_40_inst : TBUF_X1 port map( A => n248, EN => n299, Z => Y(40));
   Y_tri_41_inst : TBUF_X1 port map( A => n249, EN => n299, Z => Y(41));
   Y_tri_42_inst : TBUF_X1 port map( A => n250, EN => n299, Z => Y(42));
   Y_tri_43_inst : TBUF_X1 port map( A => n251, EN => n299, Z => Y(43));
   Y_tri_44_inst : TBUF_X1 port map( A => n252, EN => n299, Z => Y(44));
   Y_tri_45_inst : TBUF_X1 port map( A => n253, EN => n299, Z => Y(45));
   Y_tri_46_inst : TBUF_X1 port map( A => n254, EN => n299, Z => Y(46));
   Y_tri_47_inst : TBUF_X1 port map( A => n255, EN => n299, Z => Y(47));
   Y_tri_20_inst : TBUF_X1 port map( A => n228, EN => n297, Z => Y(20));
   Y_tri_18_inst : TBUF_X1 port map( A => n226, EN => n297, Z => Y(18));
   Y_tri_17_inst : TBUF_X1 port map( A => n225, EN => n297, Z => Y(17));
   Y_tri_16_inst : TBUF_X1 port map( A => n224, EN => n297, Z => Y(16));
   Y_tri_11_inst : TBUF_X1 port map( A => n219, EN => n296, Z => Y(11));
   Y_tri_15_inst : TBUF_X1 port map( A => n223, EN => n297, Z => Y(15));
   Y_tri_14_inst : TBUF_X1 port map( A => n222, EN => n297, Z => Y(14));
   Y_tri_13_inst : TBUF_X1 port map( A => n221, EN => n297, Z => Y(13));
   Y_tri_25_inst : TBUF_X1 port map( A => n233, EN => n298, Z => Y(25));
   Y_tri_26_inst : TBUF_X1 port map( A => n234, EN => n298, Z => Y(26));
   Y_tri_24_inst : TBUF_X1 port map( A => n232, EN => n298, Z => Y(24));
   Y_tri_21_inst : TBUF_X1 port map( A => n229, EN => n297, Z => Y(21));
   Y_tri_23_inst : TBUF_X1 port map( A => n231, EN => n297, Z => Y(23));
   Y_tri_22_inst : TBUF_X1 port map( A => n230, EN => n297, Z => Y(22));
   Y_tri_12_inst : TBUF_X1 port map( A => n220, EN => n297, Z => Y(12));
   Y_tri_10_inst : TBUF_X1 port map( A => n218, EN => n296, Z => Y(10));
   Y_tri_9_inst : TBUF_X1 port map( A => n217, EN => n296, Z => Y(9));
   Y_tri_8_inst : TBUF_X1 port map( A => n215, EN => n296, Z => Y(8));
   Y_tri_7_inst : TBUF_X1 port map( A => n214, EN => n296, Z => Y(7));
   Y_tri_6_inst : TBUF_X1 port map( A => n213, EN => n296, Z => Y(6));
   Y_tri_5_inst : TBUF_X1 port map( A => n212, EN => n296, Z => Y(5));
   Y_tri_4_inst : TBUF_X1 port map( A => n211, EN => n296, Z => Y(4));
   Y_tri_3_inst : TBUF_X1 port map( A => n210, EN => n296, Z => Y(3));
   Y_tri_19_inst : TBUF_X1 port map( A => n227, EN => n297, Z => Y(19));
   Y_tri_2_inst : TBUF_X1 port map( A => n209, EN => n296, Z => Y(2));
   Y_tri_1_inst : TBUF_X1 port map( A => n208, EN => n296, Z => Y(1));
   Y_tri_0_inst : TBUF_X1 port map( A => n207, EN => n296, Z => Y(0));
   U2 : NOR3_X1 port map( A1 => SEL(0), A2 => SEL(2), A3 => n302, ZN => n7);
   U3 : NOR3_X1 port map( A1 => n302, A2 => SEL(2), A3 => n303, ZN => n9);
   U4 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => n303, ZN => n8);
   U5 : BUF_X2 port map( A => n216, Z => n296);
   U6 : CLKBUF_X1 port map( A => n6, Z => n292);
   U7 : CLKBUF_X1 port map( A => n6, Z => n293);
   U8 : CLKBUF_X1 port map( A => n6, Z => n294);
   U9 : CLKBUF_X1 port map( A => n216, Z => n297);
   U10 : CLKBUF_X1 port map( A => n216, Z => n298);
   U11 : CLKBUF_X1 port map( A => n6, Z => n291);
   U12 : CLKBUF_X1 port map( A => n216, Z => n299);
   U13 : CLKBUF_X1 port map( A => n216, Z => n300);
   U14 : BUF_X1 port map( A => n8, Z => n278);
   U15 : CLKBUF_X1 port map( A => n8, Z => n279);
   U16 : CLKBUF_X1 port map( A => n8, Z => n280);
   U17 : BUF_X1 port map( A => n7, Z => n284);
   U18 : BUF_X1 port map( A => n9, Z => n272);
   U19 : CLKBUF_X1 port map( A => n7, Z => n285);
   U20 : CLKBUF_X1 port map( A => n9, Z => n273);
   U21 : CLKBUF_X1 port map( A => n7, Z => n286);
   U22 : CLKBUF_X1 port map( A => n9, Z => n274);
   U23 : BUF_X1 port map( A => n6, Z => n290);
   U24 : NAND2_X1 port map( A1 => n62, A2 => n63, ZN => n244);
   U25 : AOI22_X1 port map( A1 => plusA(36), A2 => n281, B1 => plus2A(36), B2 
                           => n275, ZN => n62);
   U26 : AOI22_X1 port map( A1 => minus2A(36), A2 => n293, B1 => minusA(36), B2
                           => n287, ZN => n63);
   U27 : NAND2_X1 port map( A1 => n70, A2 => n71, ZN => n240);
   U28 : AOI22_X1 port map( A1 => plusA(32), A2 => n280, B1 => plus2A(32), B2 
                           => n274, ZN => n70);
   U29 : AOI22_X1 port map( A1 => minus2A(32), A2 => n292, B1 => minusA(32), B2
                           => n286, ZN => n71);
   U30 : NAND2_X1 port map( A1 => n84, A2 => n85, ZN => n233);
   U31 : AOI22_X1 port map( A1 => plusA(25), A2 => n280, B1 => plus2A(25), B2 
                           => n274, ZN => n84);
   U32 : AOI22_X1 port map( A1 => minus2A(25), A2 => n292, B1 => minusA(25), B2
                           => n286, ZN => n85);
   U33 : NAND2_X1 port map( A1 => n92, A2 => n93, ZN => n229);
   U34 : AOI22_X1 port map( A1 => plusA(21), A2 => n279, B1 => plus2A(21), B2 
                           => n273, ZN => n92);
   U35 : AOI22_X1 port map( A1 => minus2A(21), A2 => n291, B1 => minusA(21), B2
                           => n285, ZN => n93);
   U36 : NAND2_X1 port map( A1 => n108, A2 => n109, ZN => n221);
   U37 : AOI22_X1 port map( A1 => plusA(13), A2 => n279, B1 => plus2A(13), B2 
                           => n273, ZN => n108);
   U38 : AOI22_X1 port map( A1 => minus2A(13), A2 => n291, B1 => minusA(13), B2
                           => n285, ZN => n109);
   U39 : NAND2_X1 port map( A1 => n100, A2 => n101, ZN => n225);
   U40 : AOI22_X1 port map( A1 => plusA(17), A2 => n279, B1 => plus2A(17), B2 
                           => n273, ZN => n100);
   U41 : AOI22_X1 port map( A1 => minus2A(17), A2 => n291, B1 => minusA(17), B2
                           => n285, ZN => n101);
   U42 : NAND2_X1 port map( A1 => n40, A2 => n41, ZN => n255);
   U43 : AOI22_X1 port map( A1 => plusA(47), A2 => n281, B1 => plus2A(47), B2 
                           => n275, ZN => n40);
   U44 : AOI22_X1 port map( A1 => minus2A(47), A2 => n293, B1 => minusA(47), B2
                           => n287, ZN => n41);
   U45 : NAND2_X1 port map( A1 => n44, A2 => n45, ZN => n253);
   U46 : AOI22_X1 port map( A1 => plusA(45), A2 => n281, B1 => plus2A(45), B2 
                           => n275, ZN => n44);
   U47 : AOI22_X1 port map( A1 => minus2A(45), A2 => n293, B1 => minusA(45), B2
                           => n287, ZN => n45);
   U48 : NAND2_X1 port map( A1 => n48, A2 => n49, ZN => n251);
   U49 : AOI22_X1 port map( A1 => plusA(43), A2 => n281, B1 => plus2A(43), B2 
                           => n275, ZN => n48);
   U50 : AOI22_X1 port map( A1 => minus2A(43), A2 => n293, B1 => minusA(43), B2
                           => n287, ZN => n49);
   U51 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => n245);
   U52 : AOI22_X1 port map( A1 => plusA(37), A2 => n281, B1 => plus2A(37), B2 
                           => n275, ZN => n60);
   U53 : AOI22_X1 port map( A1 => minus2A(37), A2 => n293, B1 => minusA(37), B2
                           => n287, ZN => n61);
   U54 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => n241);
   U55 : AOI22_X1 port map( A1 => plusA(33), A2 => n280, B1 => plus2A(33), B2 
                           => n274, ZN => n68);
   U56 : AOI22_X1 port map( A1 => minus2A(33), A2 => n292, B1 => minusA(33), B2
                           => n286, ZN => n69);
   U57 : NAND2_X1 port map( A1 => n76, A2 => n77, ZN => n237);
   U58 : AOI22_X1 port map( A1 => plusA(29), A2 => n280, B1 => plus2A(29), B2 
                           => n274, ZN => n76);
   U59 : AOI22_X1 port map( A1 => minus2A(29), A2 => n292, B1 => minusA(29), B2
                           => n286, ZN => n77);
   U60 : NAND2_X1 port map( A1 => n54, A2 => n55, ZN => n248);
   U61 : AOI22_X1 port map( A1 => plusA(40), A2 => n281, B1 => plus2A(40), B2 
                           => n275, ZN => n54);
   U62 : AOI22_X1 port map( A1 => minus2A(40), A2 => n293, B1 => minusA(40), B2
                           => n287, ZN => n55);
   U63 : NAND2_X1 port map( A1 => n112, A2 => n113, ZN => n219);
   U64 : AOI22_X1 port map( A1 => plusA(11), A2 => n278, B1 => plus2A(11), B2 
                           => n272, ZN => n112);
   U65 : AOI22_X1 port map( A1 => minus2A(11), A2 => n290, B1 => minusA(11), B2
                           => n284, ZN => n113);
   U66 : NAND2_X1 port map( A1 => n88, A2 => n89, ZN => n231);
   U67 : AOI22_X1 port map( A1 => plusA(23), A2 => n279, B1 => plus2A(23), B2 
                           => n273, ZN => n88);
   U68 : AOI22_X1 port map( A1 => minus2A(23), A2 => n291, B1 => minusA(23), B2
                           => n285, ZN => n89);
   U69 : NAND2_X1 port map( A1 => n104, A2 => n105, ZN => n223);
   U70 : AOI22_X1 port map( A1 => plusA(15), A2 => n279, B1 => plus2A(15), B2 
                           => n273, ZN => n104);
   U71 : AOI22_X1 port map( A1 => minus2A(15), A2 => n291, B1 => minusA(15), B2
                           => n285, ZN => n105);
   U72 : NAND2_X1 port map( A1 => n96, A2 => n97, ZN => n227);
   U73 : AOI22_X1 port map( A1 => plusA(19), A2 => n279, B1 => plus2A(19), B2 
                           => n273, ZN => n96);
   U74 : AOI22_X1 port map( A1 => minus2A(19), A2 => n291, B1 => minusA(19), B2
                           => n285, ZN => n97);
   U75 : NAND2_X1 port map( A1 => n64, A2 => n65, ZN => n243);
   U76 : AOI22_X1 port map( A1 => plusA(35), A2 => n280, B1 => plus2A(35), B2 
                           => n274, ZN => n64);
   U77 : AOI22_X1 port map( A1 => minus2A(35), A2 => n292, B1 => minusA(35), B2
                           => n286, ZN => n65);
   U78 : NAND2_X1 port map( A1 => n72, A2 => n73, ZN => n239);
   U79 : AOI22_X1 port map( A1 => plusA(31), A2 => n280, B1 => plus2A(31), B2 
                           => n274, ZN => n72);
   U80 : AOI22_X1 port map( A1 => minus2A(31), A2 => n292, B1 => minusA(31), B2
                           => n286, ZN => n73);
   U81 : NAND2_X1 port map( A1 => n80, A2 => n81, ZN => n235);
   U82 : AOI22_X1 port map( A1 => plusA(27), A2 => n280, B1 => plus2A(27), B2 
                           => n274, ZN => n80);
   U83 : AOI22_X1 port map( A1 => minus2A(27), A2 => n292, B1 => minusA(27), B2
                           => n286, ZN => n81);
   U84 : NAND2_X1 port map( A1 => n56, A2 => n57, ZN => n247);
   U85 : AOI22_X1 port map( A1 => plusA(39), A2 => n281, B1 => plus2A(39), B2 
                           => n275, ZN => n56);
   U86 : AOI22_X1 port map( A1 => minus2A(39), A2 => n293, B1 => minusA(39), B2
                           => n287, ZN => n57);
   U87 : NAND2_X1 port map( A1 => n114, A2 => n115, ZN => n218);
   U88 : AOI22_X1 port map( A1 => plusA(10), A2 => n278, B1 => plus2A(10), B2 
                           => n272, ZN => n114);
   U89 : AOI22_X1 port map( A1 => minus2A(10), A2 => n290, B1 => minusA(10), B2
                           => n284, ZN => n115);
   U90 : NAND2_X1 port map( A1 => n82, A2 => n83, ZN => n234);
   U91 : AOI22_X1 port map( A1 => plusA(26), A2 => n280, B1 => plus2A(26), B2 
                           => n274, ZN => n82);
   U92 : AOI22_X1 port map( A1 => minus2A(26), A2 => n292, B1 => minusA(26), B2
                           => n286, ZN => n83);
   U93 : NAND2_X1 port map( A1 => n90, A2 => n91, ZN => n230);
   U94 : AOI22_X1 port map( A1 => plusA(22), A2 => n279, B1 => plus2A(22), B2 
                           => n273, ZN => n90);
   U95 : AOI22_X1 port map( A1 => minus2A(22), A2 => n291, B1 => minusA(22), B2
                           => n285, ZN => n91);
   U96 : NAND2_X1 port map( A1 => n106, A2 => n107, ZN => n222);
   U97 : AOI22_X1 port map( A1 => plusA(14), A2 => n279, B1 => plus2A(14), B2 
                           => n273, ZN => n106);
   U98 : AOI22_X1 port map( A1 => minus2A(14), A2 => n291, B1 => minusA(14), B2
                           => n285, ZN => n107);
   U99 : NAND2_X1 port map( A1 => n98, A2 => n99, ZN => n226);
   U100 : AOI22_X1 port map( A1 => plusA(18), A2 => n279, B1 => plus2A(18), B2 
                           => n273, ZN => n98);
   U101 : AOI22_X1 port map( A1 => minus2A(18), A2 => n291, B1 => minusA(18), 
                           B2 => n285, ZN => n99);
   U102 : NAND2_X1 port map( A1 => n58, A2 => n59, ZN => n246);
   U103 : AOI22_X1 port map( A1 => plusA(38), A2 => n281, B1 => plus2A(38), B2 
                           => n275, ZN => n58);
   U104 : AOI22_X1 port map( A1 => minus2A(38), A2 => n293, B1 => minusA(38), 
                           B2 => n287, ZN => n59);
   U105 : NAND2_X1 port map( A1 => n66, A2 => n67, ZN => n242);
   U106 : AOI22_X1 port map( A1 => plusA(34), A2 => n280, B1 => plus2A(34), B2 
                           => n274, ZN => n66);
   U107 : AOI22_X1 port map( A1 => minus2A(34), A2 => n292, B1 => minusA(34), 
                           B2 => n286, ZN => n67);
   U108 : NAND2_X1 port map( A1 => n74, A2 => n75, ZN => n238);
   U109 : AOI22_X1 port map( A1 => plusA(30), A2 => n280, B1 => plus2A(30), B2 
                           => n274, ZN => n74);
   U110 : AOI22_X1 port map( A1 => minus2A(30), A2 => n292, B1 => minusA(30), 
                           B2 => n286, ZN => n75);
   U111 : NAND2_X1 port map( A1 => n110, A2 => n111, ZN => n220);
   U112 : AOI22_X1 port map( A1 => plusA(12), A2 => n279, B1 => plus2A(12), B2 
                           => n273, ZN => n110);
   U113 : AOI22_X1 port map( A1 => minus2A(12), A2 => n291, B1 => minusA(12), 
                           B2 => n285, ZN => n111);
   U114 : NAND2_X1 port map( A1 => n86, A2 => n87, ZN => n232);
   U115 : AOI22_X1 port map( A1 => plusA(24), A2 => n280, B1 => plus2A(24), B2 
                           => n274, ZN => n86);
   U116 : AOI22_X1 port map( A1 => minus2A(24), A2 => n292, B1 => minusA(24), 
                           B2 => n286, ZN => n87);
   U117 : NAND2_X1 port map( A1 => n102, A2 => n103, ZN => n224);
   U118 : AOI22_X1 port map( A1 => plusA(16), A2 => n279, B1 => plus2A(16), B2 
                           => n273, ZN => n102);
   U119 : AOI22_X1 port map( A1 => minus2A(16), A2 => n291, B1 => minusA(16), 
                           B2 => n285, ZN => n103);
   U120 : NAND2_X1 port map( A1 => n94, A2 => n95, ZN => n228);
   U121 : AOI22_X1 port map( A1 => plusA(20), A2 => n279, B1 => plus2A(20), B2 
                           => n273, ZN => n94);
   U122 : AOI22_X1 port map( A1 => minus2A(20), A2 => n291, B1 => minusA(20), 
                           B2 => n285, ZN => n95);
   U123 : NAND2_X1 port map( A1 => n42, A2 => n43, ZN => n254);
   U124 : AOI22_X1 port map( A1 => plusA(46), A2 => n281, B1 => plus2A(46), B2 
                           => n275, ZN => n42);
   U125 : AOI22_X1 port map( A1 => minus2A(46), A2 => n293, B1 => minusA(46), 
                           B2 => n287, ZN => n43);
   U126 : NAND2_X1 port map( A1 => n46, A2 => n47, ZN => n252);
   U127 : AOI22_X1 port map( A1 => plusA(44), A2 => n281, B1 => plus2A(44), B2 
                           => n275, ZN => n46);
   U128 : AOI22_X1 port map( A1 => minus2A(44), A2 => n293, B1 => minusA(44), 
                           B2 => n287, ZN => n47);
   U129 : NAND2_X1 port map( A1 => n78, A2 => n79, ZN => n236);
   U130 : AOI22_X1 port map( A1 => plusA(28), A2 => n280, B1 => plus2A(28), B2 
                           => n274, ZN => n78);
   U131 : AOI22_X1 port map( A1 => minus2A(28), A2 => n292, B1 => minusA(28), 
                           B2 => n286, ZN => n79);
   U132 : CLKBUF_X1 port map( A => n8, Z => n281);
   U133 : CLKBUF_X1 port map( A => n7, Z => n287);
   U134 : CLKBUF_X1 port map( A => n9, Z => n275);
   U135 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => n268);
   U136 : AOI22_X1 port map( A1 => plusA(60), A2 => n283, B1 => plus2A(60), B2 
                           => n277, ZN => n14);
   U137 : AOI22_X1 port map( A1 => minus2A(60), A2 => n295, B1 => minusA(60), 
                           B2 => n289, ZN => n15);
   U138 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => n267);
   U139 : AOI22_X1 port map( A1 => plusA(59), A2 => n282, B1 => plus2A(59), B2 
                           => n276, ZN => n16);
   U140 : AOI22_X1 port map( A1 => minus2A(59), A2 => n294, B1 => minusA(59), 
                           B2 => n288, ZN => n17);
   U141 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => n266);
   U142 : AOI22_X1 port map( A1 => plusA(58), A2 => n282, B1 => plus2A(58), B2 
                           => n276, ZN => n18);
   U143 : AOI22_X1 port map( A1 => minus2A(58), A2 => n294, B1 => minusA(58), 
                           B2 => n288, ZN => n19);
   U144 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => n265);
   U145 : AOI22_X1 port map( A1 => plusA(57), A2 => n282, B1 => plus2A(57), B2 
                           => n276, ZN => n20);
   U146 : AOI22_X1 port map( A1 => minus2A(57), A2 => n294, B1 => minusA(57), 
                           B2 => n288, ZN => n21);
   U147 : NAND2_X1 port map( A1 => n24, A2 => n25, ZN => n263);
   U148 : AOI22_X1 port map( A1 => plusA(55), A2 => n282, B1 => plus2A(55), B2 
                           => n276, ZN => n24);
   U149 : AOI22_X1 port map( A1 => minus2A(55), A2 => n294, B1 => minusA(55), 
                           B2 => n288, ZN => n25);
   U150 : NAND2_X1 port map( A1 => n26, A2 => n27, ZN => n262);
   U151 : AOI22_X1 port map( A1 => plusA(54), A2 => n282, B1 => plus2A(54), B2 
                           => n276, ZN => n26);
   U152 : AOI22_X1 port map( A1 => minus2A(54), A2 => n294, B1 => minusA(54), 
                           B2 => n288, ZN => n27);
   U153 : NAND2_X1 port map( A1 => n28, A2 => n29, ZN => n261);
   U154 : AOI22_X1 port map( A1 => plusA(53), A2 => n282, B1 => plus2A(53), B2 
                           => n276, ZN => n28);
   U155 : AOI22_X1 port map( A1 => minus2A(53), A2 => n294, B1 => minusA(53), 
                           B2 => n288, ZN => n29);
   U156 : NAND2_X1 port map( A1 => n34, A2 => n35, ZN => n258);
   U157 : AOI22_X1 port map( A1 => plusA(50), A2 => n282, B1 => plus2A(50), B2 
                           => n276, ZN => n34);
   U158 : AOI22_X1 port map( A1 => minus2A(50), A2 => n294, B1 => minusA(50), 
                           B2 => n288, ZN => n35);
   U159 : NAND2_X1 port map( A1 => n38, A2 => n39, ZN => n256);
   U160 : AOI22_X1 port map( A1 => plusA(48), A2 => n282, B1 => plus2A(48), B2 
                           => n276, ZN => n38);
   U161 : AOI22_X1 port map( A1 => minus2A(48), A2 => n294, B1 => minusA(48), 
                           B2 => n288, ZN => n39);
   U162 : NAND2_X1 port map( A1 => n36, A2 => n37, ZN => n257);
   U163 : AOI22_X1 port map( A1 => plusA(49), A2 => n282, B1 => plus2A(49), B2 
                           => n276, ZN => n36);
   U164 : AOI22_X1 port map( A1 => minus2A(49), A2 => n294, B1 => minusA(49), 
                           B2 => n288, ZN => n37);
   U165 : NAND2_X1 port map( A1 => n22, A2 => n23, ZN => n264);
   U166 : AOI22_X1 port map( A1 => plusA(56), A2 => n282, B1 => plus2A(56), B2 
                           => n276, ZN => n22);
   U167 : AOI22_X1 port map( A1 => minus2A(56), A2 => n294, B1 => minusA(56), 
                           B2 => n288, ZN => n23);
   U168 : CLKBUF_X1 port map( A => n8, Z => n282);
   U169 : CLKBUF_X1 port map( A => n7, Z => n288);
   U170 : CLKBUF_X1 port map( A => n9, Z => n276);
   U171 : NOR2_X1 port map( A1 => n118, A2 => n304, ZN => n216);
   U172 : INV_X1 port map( A => SEL(2), ZN => n304);
   U173 : NOR2_X1 port map( A1 => SEL(1), A2 => SEL(0), ZN => n118);
   U174 : AND2_X1 port map( A1 => SEL(2), A2 => n118, ZN => n6);
   U175 : NAND2_X1 port map( A1 => n116, A2 => n117, ZN => n217);
   U176 : AOI22_X1 port map( A1 => plusA(9), A2 => n278, B1 => plus2A(9), B2 =>
                           n272, ZN => n116);
   U177 : AOI22_X1 port map( A1 => minus2A(9), A2 => n290, B1 => minusA(9), B2 
                           => n284, ZN => n117);
   U178 : INV_X1 port map( A => SEL(1), ZN => n302);
   U179 : INV_X1 port map( A => SEL(0), ZN => n303);
   U180 : NAND2_X1 port map( A1 => n52, A2 => n53, ZN => n249);
   U181 : AOI22_X1 port map( A1 => plusA(41), A2 => n281, B1 => plus2A(41), B2 
                           => n275, ZN => n52);
   U182 : AOI22_X1 port map( A1 => minus2A(41), A2 => n293, B1 => minusA(41), 
                           B2 => n287, ZN => n53);
   U183 : NAND2_X1 port map( A1 => n50, A2 => n51, ZN => n250);
   U184 : AOI22_X1 port map( A1 => plusA(42), A2 => n281, B1 => plus2A(42), B2 
                           => n275, ZN => n50);
   U185 : AOI22_X1 port map( A1 => minus2A(42), A2 => n293, B1 => minusA(42), 
                           B2 => n287, ZN => n51);
   U186 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => n271);
   U187 : AOI22_X1 port map( A1 => plusA(63), A2 => n283, B1 => plus2A(63), B2 
                           => n277, ZN => n4);
   U188 : AOI22_X1 port map( A1 => minus2A(63), A2 => n295, B1 => minusA(63), 
                           B2 => n289, ZN => n5);
   U189 : NAND2_X1 port map( A1 => n10, A2 => n11, ZN => n270);
   U190 : AOI22_X1 port map( A1 => plusA(62), A2 => n283, B1 => plus2A(62), B2 
                           => n277, ZN => n10);
   U191 : AOI22_X1 port map( A1 => minus2A(62), A2 => n295, B1 => minusA(62), 
                           B2 => n289, ZN => n11);
   U192 : NAND2_X1 port map( A1 => n12, A2 => n13, ZN => n269);
   U193 : AOI22_X1 port map( A1 => plusA(61), A2 => n283, B1 => plus2A(61), B2 
                           => n277, ZN => n12);
   U194 : AOI22_X1 port map( A1 => minus2A(61), A2 => n295, B1 => minusA(61), 
                           B2 => n289, ZN => n13);
   U195 : NAND2_X1 port map( A1 => n32, A2 => n33, ZN => n259);
   U196 : AOI22_X1 port map( A1 => plusA(51), A2 => n282, B1 => plus2A(51), B2 
                           => n276, ZN => n32);
   U197 : AOI22_X1 port map( A1 => minus2A(51), A2 => n294, B1 => minusA(51), 
                           B2 => n288, ZN => n33);
   U198 : NAND2_X1 port map( A1 => n30, A2 => n31, ZN => n260);
   U199 : AOI22_X1 port map( A1 => plusA(52), A2 => n282, B1 => plus2A(52), B2 
                           => n276, ZN => n30);
   U200 : AOI22_X1 port map( A1 => minus2A(52), A2 => n294, B1 => minusA(52), 
                           B2 => n288, ZN => n31);
   U201 : NAND2_X1 port map( A1 => n119, A2 => n120, ZN => n215);
   U202 : AOI22_X1 port map( A1 => plusA(8), A2 => n278, B1 => plus2A(8), B2 =>
                           n272, ZN => n119);
   U203 : AOI22_X1 port map( A1 => minus2A(8), A2 => n290, B1 => minusA(8), B2 
                           => n284, ZN => n120);
   U204 : NAND2_X1 port map( A1 => n121, A2 => n122, ZN => n214);
   U205 : AOI22_X1 port map( A1 => plusA(7), A2 => n278, B1 => plus2A(7), B2 =>
                           n272, ZN => n121);
   U206 : AOI22_X1 port map( A1 => minus2A(7), A2 => n290, B1 => minusA(7), B2 
                           => n284, ZN => n122);
   U207 : NAND2_X1 port map( A1 => n123, A2 => n124, ZN => n213);
   U208 : AOI22_X1 port map( A1 => plusA(6), A2 => n278, B1 => plus2A(6), B2 =>
                           n272, ZN => n123);
   U209 : AOI22_X1 port map( A1 => minus2A(6), A2 => n290, B1 => minusA(6), B2 
                           => n284, ZN => n124);
   U210 : NAND2_X1 port map( A1 => n125, A2 => n126, ZN => n212);
   U211 : AOI22_X1 port map( A1 => plusA(5), A2 => n278, B1 => plus2A(5), B2 =>
                           n272, ZN => n125);
   U212 : AOI22_X1 port map( A1 => minus2A(5), A2 => n290, B1 => minusA(5), B2 
                           => n284, ZN => n126);
   U213 : NAND2_X1 port map( A1 => n129, A2 => n130, ZN => n210);
   U214 : AOI22_X1 port map( A1 => plusA(3), A2 => n278, B1 => plus2A(3), B2 =>
                           n272, ZN => n129);
   U215 : AOI22_X1 port map( A1 => minus2A(3), A2 => n290, B1 => minusA(3), B2 
                           => n284, ZN => n130);
   U216 : NAND2_X1 port map( A1 => n127, A2 => n128, ZN => n211);
   U217 : AOI22_X1 port map( A1 => plusA(4), A2 => n278, B1 => plus2A(4), B2 =>
                           n272, ZN => n127);
   U218 : AOI22_X1 port map( A1 => minus2A(4), A2 => n290, B1 => minusA(4), B2 
                           => n284, ZN => n128);
   U219 : NAND2_X1 port map( A1 => n131, A2 => n132, ZN => n209);
   U220 : AOI22_X1 port map( A1 => plusA(2), A2 => n278, B1 => plus2A(2), B2 =>
                           n272, ZN => n131);
   U221 : AOI22_X1 port map( A1 => minus2A(2), A2 => n290, B1 => minusA(2), B2 
                           => n284, ZN => n132);
   U222 : NAND2_X1 port map( A1 => n133, A2 => n134, ZN => n208);
   U223 : AOI22_X1 port map( A1 => plusA(1), A2 => n278, B1 => plus2A(1), B2 =>
                           n272, ZN => n133);
   U224 : AOI22_X1 port map( A1 => minus2A(1), A2 => n290, B1 => minusA(1), B2 
                           => n284, ZN => n134);
   U225 : NAND2_X1 port map( A1 => n135, A2 => n136, ZN => n207);
   U226 : AOI22_X1 port map( A1 => plusA(0), A2 => n278, B1 => plus2A(0), B2 =>
                           n272, ZN => n135);
   U227 : AOI22_X1 port map( A1 => minus2A(0), A2 => n290, B1 => minusA(0), B2 
                           => n284, ZN => n136);
   U228 : CLKBUF_X1 port map( A => n9, Z => n277);
   U229 : CLKBUF_X1 port map( A => n8, Z => n283);
   U230 : CLKBUF_X1 port map( A => n7, Z => n289);
   U231 : CLKBUF_X1 port map( A => n6, Z => n295);
   U232 : CLKBUF_X1 port map( A => n216, Z => n301);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity ShiftnCompl_N64_12 is

   port( plusA : in std_logic_vector (63 downto 0);  plus2A_out, minus2A_out, 
         plus4A_out, minus4A_out : out std_logic_vector (63 downto 0));

end ShiftnCompl_N64_12;

architecture SYN_struct of ShiftnCompl_N64_12 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component complementer_N64_23
      port( input : in std_logic_vector (63 downto 0);  complement2 : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component complementer_N64_24
      port( input : in std_logic_vector (63 downto 0);  complement2 : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component shifter_N64_23
      port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component shifter_N64_24
      port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
            std_logic_vector (63 downto 0));
   end component;
   
   signal plus2A_out_63_port, plus2A_out_62_port, plus2A_out_61_port, 
      plus2A_out_60_port, plus2A_out_59_port, plus2A_out_58_port, n8, 
      plus2A_out_56_port, plus2A_out_55_port, plus2A_out_54_port, 
      plus2A_out_53_port, plus2A_out_52_port, plus2A_out_51_port, 
      plus2A_out_50_port, plus2A_out_49_port, n9, n10, plus2A_out_46_port, 
      plus2A_out_45_port, plus2A_out_44_port, plus2A_out_43_port, 
      plus2A_out_42_port, plus2A_out_41_port, plus2A_out_40_port, 
      plus2A_out_39_port, plus2A_out_38_port, plus2A_out_37_port, 
      plus2A_out_36_port, plus2A_out_35_port, plus2A_out_34_port, 
      plus2A_out_33_port, plus2A_out_32_port, plus2A_out_31_port, 
      plus2A_out_30_port, plus2A_out_29_port, plus2A_out_28_port, 
      plus2A_out_27_port, plus2A_out_26_port, plus2A_out_25_port, 
      plus2A_out_24_port, plus2A_out_23_port, plus2A_out_22_port, 
      plus2A_out_21_port, plus2A_out_20_port, plus2A_out_19_port, 
      plus2A_out_18_port, plus2A_out_17_port, plus2A_out_16_port, 
      plus2A_out_15_port, plus2A_out_14_port, plus2A_out_13_port, 
      plus2A_out_12_port, plus2A_out_11_port, plus2A_out_10_port, 
      plus2A_out_9_port, plus2A_out_8_port, plus2A_out_7_port, 
      plus2A_out_6_port, plus2A_out_5_port, plus2A_out_4_port, 
      plus2A_out_3_port, plus2A_out_2_port, plus2A_out_1_port, 
      plus2A_out_0_port, plus4A_out_63_port, plus4A_out_62_port, 
      plus4A_out_61_port, plus4A_out_60_port, plus4A_out_59_port, 
      plus4A_out_58_port, plus4A_out_57_port, plus4A_out_56_port, 
      plus4A_out_55_port, plus4A_out_54_port, n11, n12, plus4A_out_51_port, 
      plus4A_out_50_port, plus4A_out_49_port, plus4A_out_48_port, 
      plus4A_out_47_port, plus4A_out_46_port, plus4A_out_45_port, 
      plus4A_out_44_port, n13, n14, plus4A_out_41_port, plus4A_out_40_port, 
      plus4A_out_39_port, plus4A_out_38_port, plus4A_out_37_port, 
      plus4A_out_36_port, plus4A_out_35_port, plus4A_out_34_port, 
      plus4A_out_33_port, plus4A_out_32_port, plus4A_out_31_port, 
      plus4A_out_30_port, plus4A_out_29_port, plus4A_out_28_port, 
      plus4A_out_27_port, plus4A_out_26_port, plus4A_out_25_port, 
      plus4A_out_24_port, plus4A_out_23_port, plus4A_out_22_port, 
      plus4A_out_21_port, plus4A_out_20_port, plus4A_out_19_port, 
      plus4A_out_18_port, plus4A_out_17_port, plus4A_out_16_port, 
      plus4A_out_15_port, plus4A_out_14_port, plus4A_out_13_port, 
      plus4A_out_12_port, plus4A_out_11_port, plus4A_out_10_port, 
      plus4A_out_9_port, plus4A_out_8_port, plus4A_out_7_port, 
      plus4A_out_6_port, plus4A_out_5_port, plus4A_out_4_port, 
      plus4A_out_3_port, plus4A_out_2_port, plus4A_out_1_port, 
      plus4A_out_0_port, plus4A_out_42_port, plus4A_out_43_port, 
      plus2A_out_47_port, plus2A_out_48_port, plus4A_out_52_port, 
      plus4A_out_53_port, plus2A_out_57_port, n_3166, n_3167 : std_logic;

begin
   plus2A_out <= ( plus2A_out_63_port, plus2A_out_62_port, plus2A_out_61_port, 
      plus2A_out_60_port, plus2A_out_59_port, plus2A_out_58_port, 
      plus2A_out_57_port, plus2A_out_56_port, plus2A_out_55_port, 
      plus2A_out_54_port, plus2A_out_53_port, plus2A_out_52_port, 
      plus2A_out_51_port, plus2A_out_50_port, plus2A_out_49_port, 
      plus2A_out_48_port, plus2A_out_47_port, plus2A_out_46_port, 
      plus2A_out_45_port, plus2A_out_44_port, plus2A_out_43_port, 
      plus2A_out_42_port, plus2A_out_41_port, plus2A_out_40_port, 
      plus2A_out_39_port, plus2A_out_38_port, plus2A_out_37_port, 
      plus2A_out_36_port, plus2A_out_35_port, plus2A_out_34_port, 
      plus2A_out_33_port, plus2A_out_32_port, plus2A_out_31_port, 
      plus2A_out_30_port, plus2A_out_29_port, plus2A_out_28_port, 
      plus2A_out_27_port, plus2A_out_26_port, plus2A_out_25_port, 
      plus2A_out_24_port, plus2A_out_23_port, plus2A_out_22_port, 
      plus2A_out_21_port, plus2A_out_20_port, plus2A_out_19_port, 
      plus2A_out_18_port, plus2A_out_17_port, plus2A_out_16_port, 
      plus2A_out_15_port, plus2A_out_14_port, plus2A_out_13_port, 
      plus2A_out_12_port, plus2A_out_11_port, plus2A_out_10_port, 
      plus2A_out_9_port, plus2A_out_8_port, plus2A_out_7_port, 
      plus2A_out_6_port, plus2A_out_5_port, plus2A_out_4_port, 
      plus2A_out_3_port, plus2A_out_2_port, plus2A_out_1_port, 
      plus2A_out_0_port );
   plus4A_out <= ( plus4A_out_63_port, plus4A_out_62_port, plus4A_out_61_port, 
      plus4A_out_60_port, plus4A_out_59_port, plus4A_out_58_port, 
      plus4A_out_57_port, plus4A_out_56_port, plus4A_out_55_port, 
      plus4A_out_54_port, plus4A_out_53_port, plus4A_out_52_port, 
      plus4A_out_51_port, plus4A_out_50_port, plus4A_out_49_port, 
      plus4A_out_48_port, plus4A_out_47_port, plus4A_out_46_port, 
      plus4A_out_45_port, plus4A_out_44_port, plus4A_out_43_port, 
      plus4A_out_42_port, plus4A_out_41_port, plus4A_out_40_port, 
      plus4A_out_39_port, plus4A_out_38_port, plus4A_out_37_port, 
      plus4A_out_36_port, plus4A_out_35_port, plus4A_out_34_port, 
      plus4A_out_33_port, plus4A_out_32_port, plus4A_out_31_port, 
      plus4A_out_30_port, plus4A_out_29_port, plus4A_out_28_port, 
      plus4A_out_27_port, plus4A_out_26_port, plus4A_out_25_port, 
      plus4A_out_24_port, plus4A_out_23_port, plus4A_out_22_port, 
      plus4A_out_21_port, plus4A_out_20_port, plus4A_out_19_port, 
      plus4A_out_18_port, plus4A_out_17_port, plus4A_out_16_port, 
      plus4A_out_15_port, plus4A_out_14_port, plus4A_out_13_port, 
      plus4A_out_12_port, plus4A_out_11_port, plus4A_out_10_port, 
      plus4A_out_9_port, plus4A_out_8_port, plus4A_out_7_port, 
      plus4A_out_6_port, plus4A_out_5_port, plus4A_out_4_port, 
      plus4A_out_3_port, plus4A_out_2_port, plus4A_out_1_port, 
      plus4A_out_0_port );
   
   plus2A_out_0_port <= '0';
   plus4A_out_0_port <= '0';
   shifter_1 : shifter_N64_24 port map( input(63) => plusA(63), input(62) => 
                           plusA(62), input(61) => plusA(61), input(60) => 
                           plusA(60), input(59) => plusA(59), input(58) => 
                           plusA(58), input(57) => plusA(57), input(56) => 
                           plusA(56), input(55) => plusA(55), input(54) => 
                           plusA(54), input(53) => plusA(53), input(52) => 
                           plusA(52), input(51) => plusA(51), input(50) => 
                           plusA(50), input(49) => plusA(49), input(48) => 
                           plusA(48), input(47) => plusA(47), input(46) => 
                           plusA(46), input(45) => plusA(45), input(44) => 
                           plusA(44), input(43) => plusA(43), input(42) => 
                           plusA(42), input(41) => plusA(41), input(40) => 
                           plusA(40), input(39) => plusA(39), input(38) => 
                           plusA(38), input(37) => plusA(37), input(36) => 
                           plusA(36), input(35) => plusA(35), input(34) => 
                           plusA(34), input(33) => plusA(33), input(32) => 
                           plusA(32), input(31) => plusA(31), input(30) => 
                           plusA(30), input(29) => plusA(29), input(28) => 
                           plusA(28), input(27) => plusA(27), input(26) => 
                           plusA(26), input(25) => plusA(25), input(24) => 
                           plusA(24), input(23) => plusA(23), input(22) => 
                           plusA(22), input(21) => plusA(21), input(20) => 
                           plusA(20), input(19) => plusA(19), input(18) => 
                           plusA(18), input(17) => plusA(17), input(16) => 
                           plusA(16), input(15) => plusA(15), input(14) => 
                           plusA(14), input(13) => plusA(13), input(12) => 
                           plusA(12), input(11) => plusA(11), input(10) => 
                           plusA(10), input(9) => plusA(9), input(8) => 
                           plusA(8), input(7) => plusA(7), input(6) => plusA(6)
                           , input(5) => plusA(5), input(4) => plusA(4), 
                           input(3) => plusA(3), input(2) => plusA(2), input(1)
                           => plusA(1), input(0) => plusA(0), 
                           shiftLeftOnePos(63) => plus2A_out_63_port, 
                           shiftLeftOnePos(62) => plus2A_out_62_port, 
                           shiftLeftOnePos(61) => plus2A_out_61_port, 
                           shiftLeftOnePos(60) => plus2A_out_60_port, 
                           shiftLeftOnePos(59) => plus2A_out_59_port, 
                           shiftLeftOnePos(58) => plus2A_out_58_port, 
                           shiftLeftOnePos(57) => n8, shiftLeftOnePos(56) => 
                           plus2A_out_56_port, shiftLeftOnePos(55) => 
                           plus2A_out_55_port, shiftLeftOnePos(54) => 
                           plus2A_out_54_port, shiftLeftOnePos(53) => 
                           plus2A_out_53_port, shiftLeftOnePos(52) => 
                           plus2A_out_52_port, shiftLeftOnePos(51) => 
                           plus2A_out_51_port, shiftLeftOnePos(50) => 
                           plus2A_out_50_port, shiftLeftOnePos(49) => 
                           plus2A_out_49_port, shiftLeftOnePos(48) => n9, 
                           shiftLeftOnePos(47) => n10, shiftLeftOnePos(46) => 
                           plus2A_out_46_port, shiftLeftOnePos(45) => 
                           plus2A_out_45_port, shiftLeftOnePos(44) => 
                           plus2A_out_44_port, shiftLeftOnePos(43) => 
                           plus2A_out_43_port, shiftLeftOnePos(42) => 
                           plus2A_out_42_port, shiftLeftOnePos(41) => 
                           plus2A_out_41_port, shiftLeftOnePos(40) => 
                           plus2A_out_40_port, shiftLeftOnePos(39) => 
                           plus2A_out_39_port, shiftLeftOnePos(38) => 
                           plus2A_out_38_port, shiftLeftOnePos(37) => 
                           plus2A_out_37_port, shiftLeftOnePos(36) => 
                           plus2A_out_36_port, shiftLeftOnePos(35) => 
                           plus2A_out_35_port, shiftLeftOnePos(34) => 
                           plus2A_out_34_port, shiftLeftOnePos(33) => 
                           plus2A_out_33_port, shiftLeftOnePos(32) => 
                           plus2A_out_32_port, shiftLeftOnePos(31) => 
                           plus2A_out_31_port, shiftLeftOnePos(30) => 
                           plus2A_out_30_port, shiftLeftOnePos(29) => 
                           plus2A_out_29_port, shiftLeftOnePos(28) => 
                           plus2A_out_28_port, shiftLeftOnePos(27) => 
                           plus2A_out_27_port, shiftLeftOnePos(26) => 
                           plus2A_out_26_port, shiftLeftOnePos(25) => 
                           plus2A_out_25_port, shiftLeftOnePos(24) => 
                           plus2A_out_24_port, shiftLeftOnePos(23) => 
                           plus2A_out_23_port, shiftLeftOnePos(22) => 
                           plus2A_out_22_port, shiftLeftOnePos(21) => 
                           plus2A_out_21_port, shiftLeftOnePos(20) => 
                           plus2A_out_20_port, shiftLeftOnePos(19) => 
                           plus2A_out_19_port, shiftLeftOnePos(18) => 
                           plus2A_out_18_port, shiftLeftOnePos(17) => 
                           plus2A_out_17_port, shiftLeftOnePos(16) => 
                           plus2A_out_16_port, shiftLeftOnePos(15) => 
                           plus2A_out_15_port, shiftLeftOnePos(14) => 
                           plus2A_out_14_port, shiftLeftOnePos(13) => 
                           plus2A_out_13_port, shiftLeftOnePos(12) => 
                           plus2A_out_12_port, shiftLeftOnePos(11) => 
                           plus2A_out_11_port, shiftLeftOnePos(10) => 
                           plus2A_out_10_port, shiftLeftOnePos(9) => 
                           plus2A_out_9_port, shiftLeftOnePos(8) => 
                           plus2A_out_8_port, shiftLeftOnePos(7) => 
                           plus2A_out_7_port, shiftLeftOnePos(6) => 
                           plus2A_out_6_port, shiftLeftOnePos(5) => 
                           plus2A_out_5_port, shiftLeftOnePos(4) => 
                           plus2A_out_4_port, shiftLeftOnePos(3) => 
                           plus2A_out_3_port, shiftLeftOnePos(2) => 
                           plus2A_out_2_port, shiftLeftOnePos(1) => 
                           plus2A_out_1_port, shiftLeftOnePos(0) => n_3166);
   shifter_2 : shifter_N64_23 port map( input(63) => plus2A_out_63_port, 
                           input(62) => plus2A_out_62_port, input(61) => 
                           plus2A_out_61_port, input(60) => plus2A_out_60_port,
                           input(59) => plus2A_out_59_port, input(58) => 
                           plus2A_out_58_port, input(57) => plus2A_out_57_port,
                           input(56) => plus2A_out_56_port, input(55) => 
                           plus2A_out_55_port, input(54) => plus2A_out_54_port,
                           input(53) => plus2A_out_53_port, input(52) => 
                           plus2A_out_52_port, input(51) => plus2A_out_51_port,
                           input(50) => plus2A_out_50_port, input(49) => 
                           plus2A_out_49_port, input(48) => plus2A_out_48_port,
                           input(47) => plus2A_out_47_port, input(46) => 
                           plus2A_out_46_port, input(45) => plus2A_out_45_port,
                           input(44) => plus2A_out_44_port, input(43) => 
                           plus2A_out_43_port, input(42) => plus2A_out_42_port,
                           input(41) => plus2A_out_41_port, input(40) => 
                           plus2A_out_40_port, input(39) => plus2A_out_39_port,
                           input(38) => plus2A_out_38_port, input(37) => 
                           plus2A_out_37_port, input(36) => plus2A_out_36_port,
                           input(35) => plus2A_out_35_port, input(34) => 
                           plus2A_out_34_port, input(33) => plus2A_out_33_port,
                           input(32) => plus2A_out_32_port, input(31) => 
                           plus2A_out_31_port, input(30) => plus2A_out_30_port,
                           input(29) => plus2A_out_29_port, input(28) => 
                           plus2A_out_28_port, input(27) => plus2A_out_27_port,
                           input(26) => plus2A_out_26_port, input(25) => 
                           plus2A_out_25_port, input(24) => plus2A_out_24_port,
                           input(23) => plus2A_out_23_port, input(22) => 
                           plus2A_out_22_port, input(21) => plus2A_out_21_port,
                           input(20) => plus2A_out_20_port, input(19) => 
                           plus2A_out_19_port, input(18) => plus2A_out_18_port,
                           input(17) => plus2A_out_17_port, input(16) => 
                           plus2A_out_16_port, input(15) => plus2A_out_15_port,
                           input(14) => plus2A_out_14_port, input(13) => 
                           plus2A_out_13_port, input(12) => plus2A_out_12_port,
                           input(11) => plus2A_out_11_port, input(10) => 
                           plus2A_out_10_port, input(9) => plus2A_out_9_port, 
                           input(8) => plus2A_out_8_port, input(7) => 
                           plus2A_out_7_port, input(6) => plus2A_out_6_port, 
                           input(5) => plus2A_out_5_port, input(4) => 
                           plus2A_out_4_port, input(3) => plus2A_out_3_port, 
                           input(2) => plus2A_out_2_port, input(1) => 
                           plus2A_out_1_port, input(0) => plus2A_out_0_port, 
                           shiftLeftOnePos(63) => plus4A_out_63_port, 
                           shiftLeftOnePos(62) => plus4A_out_62_port, 
                           shiftLeftOnePos(61) => plus4A_out_61_port, 
                           shiftLeftOnePos(60) => plus4A_out_60_port, 
                           shiftLeftOnePos(59) => plus4A_out_59_port, 
                           shiftLeftOnePos(58) => plus4A_out_58_port, 
                           shiftLeftOnePos(57) => plus4A_out_57_port, 
                           shiftLeftOnePos(56) => plus4A_out_56_port, 
                           shiftLeftOnePos(55) => plus4A_out_55_port, 
                           shiftLeftOnePos(54) => plus4A_out_54_port, 
                           shiftLeftOnePos(53) => n11, shiftLeftOnePos(52) => 
                           n12, shiftLeftOnePos(51) => plus4A_out_51_port, 
                           shiftLeftOnePos(50) => plus4A_out_50_port, 
                           shiftLeftOnePos(49) => plus4A_out_49_port, 
                           shiftLeftOnePos(48) => plus4A_out_48_port, 
                           shiftLeftOnePos(47) => plus4A_out_47_port, 
                           shiftLeftOnePos(46) => plus4A_out_46_port, 
                           shiftLeftOnePos(45) => plus4A_out_45_port, 
                           shiftLeftOnePos(44) => plus4A_out_44_port, 
                           shiftLeftOnePos(43) => n13, shiftLeftOnePos(42) => 
                           n14, shiftLeftOnePos(41) => plus4A_out_41_port, 
                           shiftLeftOnePos(40) => plus4A_out_40_port, 
                           shiftLeftOnePos(39) => plus4A_out_39_port, 
                           shiftLeftOnePos(38) => plus4A_out_38_port, 
                           shiftLeftOnePos(37) => plus4A_out_37_port, 
                           shiftLeftOnePos(36) => plus4A_out_36_port, 
                           shiftLeftOnePos(35) => plus4A_out_35_port, 
                           shiftLeftOnePos(34) => plus4A_out_34_port, 
                           shiftLeftOnePos(33) => plus4A_out_33_port, 
                           shiftLeftOnePos(32) => plus4A_out_32_port, 
                           shiftLeftOnePos(31) => plus4A_out_31_port, 
                           shiftLeftOnePos(30) => plus4A_out_30_port, 
                           shiftLeftOnePos(29) => plus4A_out_29_port, 
                           shiftLeftOnePos(28) => plus4A_out_28_port, 
                           shiftLeftOnePos(27) => plus4A_out_27_port, 
                           shiftLeftOnePos(26) => plus4A_out_26_port, 
                           shiftLeftOnePos(25) => plus4A_out_25_port, 
                           shiftLeftOnePos(24) => plus4A_out_24_port, 
                           shiftLeftOnePos(23) => plus4A_out_23_port, 
                           shiftLeftOnePos(22) => plus4A_out_22_port, 
                           shiftLeftOnePos(21) => plus4A_out_21_port, 
                           shiftLeftOnePos(20) => plus4A_out_20_port, 
                           shiftLeftOnePos(19) => plus4A_out_19_port, 
                           shiftLeftOnePos(18) => plus4A_out_18_port, 
                           shiftLeftOnePos(17) => plus4A_out_17_port, 
                           shiftLeftOnePos(16) => plus4A_out_16_port, 
                           shiftLeftOnePos(15) => plus4A_out_15_port, 
                           shiftLeftOnePos(14) => plus4A_out_14_port, 
                           shiftLeftOnePos(13) => plus4A_out_13_port, 
                           shiftLeftOnePos(12) => plus4A_out_12_port, 
                           shiftLeftOnePos(11) => plus4A_out_11_port, 
                           shiftLeftOnePos(10) => plus4A_out_10_port, 
                           shiftLeftOnePos(9) => plus4A_out_9_port, 
                           shiftLeftOnePos(8) => plus4A_out_8_port, 
                           shiftLeftOnePos(7) => plus4A_out_7_port, 
                           shiftLeftOnePos(6) => plus4A_out_6_port, 
                           shiftLeftOnePos(5) => plus4A_out_5_port, 
                           shiftLeftOnePos(4) => plus4A_out_4_port, 
                           shiftLeftOnePos(3) => plus4A_out_3_port, 
                           shiftLeftOnePos(2) => plus4A_out_2_port, 
                           shiftLeftOnePos(1) => plus4A_out_1_port, 
                           shiftLeftOnePos(0) => n_3167);
   complementer_1 : complementer_N64_24 port map( input(63) => 
                           plus2A_out_63_port, input(62) => plus2A_out_62_port,
                           input(61) => plus2A_out_61_port, input(60) => 
                           plus2A_out_60_port, input(59) => plus2A_out_59_port,
                           input(58) => plus2A_out_58_port, input(57) => 
                           plus2A_out_57_port, input(56) => plus2A_out_56_port,
                           input(55) => plus2A_out_55_port, input(54) => 
                           plus2A_out_54_port, input(53) => plus2A_out_53_port,
                           input(52) => plus2A_out_52_port, input(51) => 
                           plus2A_out_51_port, input(50) => plus2A_out_50_port,
                           input(49) => plus2A_out_49_port, input(48) => 
                           plus2A_out_48_port, input(47) => plus2A_out_47_port,
                           input(46) => plus2A_out_46_port, input(45) => 
                           plus2A_out_45_port, input(44) => plus2A_out_44_port,
                           input(43) => plus2A_out_43_port, input(42) => 
                           plus2A_out_42_port, input(41) => plus2A_out_41_port,
                           input(40) => plus2A_out_40_port, input(39) => 
                           plus2A_out_39_port, input(38) => plus2A_out_38_port,
                           input(37) => plus2A_out_37_port, input(36) => 
                           plus2A_out_36_port, input(35) => plus2A_out_35_port,
                           input(34) => plus2A_out_34_port, input(33) => 
                           plus2A_out_33_port, input(32) => plus2A_out_32_port,
                           input(31) => plus2A_out_31_port, input(30) => 
                           plus2A_out_30_port, input(29) => plus2A_out_29_port,
                           input(28) => plus2A_out_28_port, input(27) => 
                           plus2A_out_27_port, input(26) => plus2A_out_26_port,
                           input(25) => plus2A_out_25_port, input(24) => 
                           plus2A_out_24_port, input(23) => plus2A_out_23_port,
                           input(22) => plus2A_out_22_port, input(21) => 
                           plus2A_out_21_port, input(20) => plus2A_out_20_port,
                           input(19) => plus2A_out_19_port, input(18) => 
                           plus2A_out_18_port, input(17) => plus2A_out_17_port,
                           input(16) => plus2A_out_16_port, input(15) => 
                           plus2A_out_15_port, input(14) => plus2A_out_14_port,
                           input(13) => plus2A_out_13_port, input(12) => 
                           plus2A_out_12_port, input(11) => plus2A_out_11_port,
                           input(10) => plus2A_out_10_port, input(9) => 
                           plus2A_out_9_port, input(8) => plus2A_out_8_port, 
                           input(7) => plus2A_out_7_port, input(6) => 
                           plus2A_out_6_port, input(5) => plus2A_out_5_port, 
                           input(4) => plus2A_out_4_port, input(3) => 
                           plus2A_out_3_port, input(2) => plus2A_out_2_port, 
                           input(1) => plus2A_out_1_port, input(0) => 
                           plus2A_out_0_port, complement2(63) => 
                           minus2A_out(63), complement2(62) => minus2A_out(62),
                           complement2(61) => minus2A_out(61), complement2(60) 
                           => minus2A_out(60), complement2(59) => 
                           minus2A_out(59), complement2(58) => minus2A_out(58),
                           complement2(57) => minus2A_out(57), complement2(56) 
                           => minus2A_out(56), complement2(55) => 
                           minus2A_out(55), complement2(54) => minus2A_out(54),
                           complement2(53) => minus2A_out(53), complement2(52) 
                           => minus2A_out(52), complement2(51) => 
                           minus2A_out(51), complement2(50) => minus2A_out(50),
                           complement2(49) => minus2A_out(49), complement2(48) 
                           => minus2A_out(48), complement2(47) => 
                           minus2A_out(47), complement2(46) => minus2A_out(46),
                           complement2(45) => minus2A_out(45), complement2(44) 
                           => minus2A_out(44), complement2(43) => 
                           minus2A_out(43), complement2(42) => minus2A_out(42),
                           complement2(41) => minus2A_out(41), complement2(40) 
                           => minus2A_out(40), complement2(39) => 
                           minus2A_out(39), complement2(38) => minus2A_out(38),
                           complement2(37) => minus2A_out(37), complement2(36) 
                           => minus2A_out(36), complement2(35) => 
                           minus2A_out(35), complement2(34) => minus2A_out(34),
                           complement2(33) => minus2A_out(33), complement2(32) 
                           => minus2A_out(32), complement2(31) => 
                           minus2A_out(31), complement2(30) => minus2A_out(30),
                           complement2(29) => minus2A_out(29), complement2(28) 
                           => minus2A_out(28), complement2(27) => 
                           minus2A_out(27), complement2(26) => minus2A_out(26),
                           complement2(25) => minus2A_out(25), complement2(24) 
                           => minus2A_out(24), complement2(23) => 
                           minus2A_out(23), complement2(22) => minus2A_out(22),
                           complement2(21) => minus2A_out(21), complement2(20) 
                           => minus2A_out(20), complement2(19) => 
                           minus2A_out(19), complement2(18) => minus2A_out(18),
                           complement2(17) => minus2A_out(17), complement2(16) 
                           => minus2A_out(16), complement2(15) => 
                           minus2A_out(15), complement2(14) => minus2A_out(14),
                           complement2(13) => minus2A_out(13), complement2(12) 
                           => minus2A_out(12), complement2(11) => 
                           minus2A_out(11), complement2(10) => minus2A_out(10),
                           complement2(9) => minus2A_out(9), complement2(8) => 
                           minus2A_out(8), complement2(7) => minus2A_out(7), 
                           complement2(6) => minus2A_out(6), complement2(5) => 
                           minus2A_out(5), complement2(4) => minus2A_out(4), 
                           complement2(3) => minus2A_out(3), complement2(2) => 
                           minus2A_out(2), complement2(1) => minus2A_out(1), 
                           complement2(0) => minus2A_out(0));
   complementer_2 : complementer_N64_23 port map( input(63) => 
                           plus4A_out_63_port, input(62) => plus4A_out_62_port,
                           input(61) => plus4A_out_61_port, input(60) => 
                           plus4A_out_60_port, input(59) => plus4A_out_59_port,
                           input(58) => plus4A_out_58_port, input(57) => 
                           plus4A_out_57_port, input(56) => plus4A_out_56_port,
                           input(55) => plus4A_out_55_port, input(54) => 
                           plus4A_out_54_port, input(53) => plus4A_out_53_port,
                           input(52) => plus4A_out_52_port, input(51) => 
                           plus4A_out_51_port, input(50) => plus4A_out_50_port,
                           input(49) => plus4A_out_49_port, input(48) => 
                           plus4A_out_48_port, input(47) => plus4A_out_47_port,
                           input(46) => plus4A_out_46_port, input(45) => 
                           plus4A_out_45_port, input(44) => plus4A_out_44_port,
                           input(43) => plus4A_out_43_port, input(42) => 
                           plus4A_out_42_port, input(41) => plus4A_out_41_port,
                           input(40) => plus4A_out_40_port, input(39) => 
                           plus4A_out_39_port, input(38) => plus4A_out_38_port,
                           input(37) => plus4A_out_37_port, input(36) => 
                           plus4A_out_36_port, input(35) => plus4A_out_35_port,
                           input(34) => plus4A_out_34_port, input(33) => 
                           plus4A_out_33_port, input(32) => plus4A_out_32_port,
                           input(31) => plus4A_out_31_port, input(30) => 
                           plus4A_out_30_port, input(29) => plus4A_out_29_port,
                           input(28) => plus4A_out_28_port, input(27) => 
                           plus4A_out_27_port, input(26) => plus4A_out_26_port,
                           input(25) => plus4A_out_25_port, input(24) => 
                           plus4A_out_24_port, input(23) => plus4A_out_23_port,
                           input(22) => plus4A_out_22_port, input(21) => 
                           plus4A_out_21_port, input(20) => plus4A_out_20_port,
                           input(19) => plus4A_out_19_port, input(18) => 
                           plus4A_out_18_port, input(17) => plus4A_out_17_port,
                           input(16) => plus4A_out_16_port, input(15) => 
                           plus4A_out_15_port, input(14) => plus4A_out_14_port,
                           input(13) => plus4A_out_13_port, input(12) => 
                           plus4A_out_12_port, input(11) => plus4A_out_11_port,
                           input(10) => plus4A_out_10_port, input(9) => 
                           plus4A_out_9_port, input(8) => plus4A_out_8_port, 
                           input(7) => plus4A_out_7_port, input(6) => 
                           plus4A_out_6_port, input(5) => plus4A_out_5_port, 
                           input(4) => plus4A_out_4_port, input(3) => 
                           plus4A_out_3_port, input(2) => plus4A_out_2_port, 
                           input(1) => plus4A_out_1_port, input(0) => 
                           plus4A_out_0_port, complement2(63) => 
                           minus4A_out(63), complement2(62) => minus4A_out(62),
                           complement2(61) => minus4A_out(61), complement2(60) 
                           => minus4A_out(60), complement2(59) => 
                           minus4A_out(59), complement2(58) => minus4A_out(58),
                           complement2(57) => minus4A_out(57), complement2(56) 
                           => minus4A_out(56), complement2(55) => 
                           minus4A_out(55), complement2(54) => minus4A_out(54),
                           complement2(53) => minus4A_out(53), complement2(52) 
                           => minus4A_out(52), complement2(51) => 
                           minus4A_out(51), complement2(50) => minus4A_out(50),
                           complement2(49) => minus4A_out(49), complement2(48) 
                           => minus4A_out(48), complement2(47) => 
                           minus4A_out(47), complement2(46) => minus4A_out(46),
                           complement2(45) => minus4A_out(45), complement2(44) 
                           => minus4A_out(44), complement2(43) => 
                           minus4A_out(43), complement2(42) => minus4A_out(42),
                           complement2(41) => minus4A_out(41), complement2(40) 
                           => minus4A_out(40), complement2(39) => 
                           minus4A_out(39), complement2(38) => minus4A_out(38),
                           complement2(37) => minus4A_out(37), complement2(36) 
                           => minus4A_out(36), complement2(35) => 
                           minus4A_out(35), complement2(34) => minus4A_out(34),
                           complement2(33) => minus4A_out(33), complement2(32) 
                           => minus4A_out(32), complement2(31) => 
                           minus4A_out(31), complement2(30) => minus4A_out(30),
                           complement2(29) => minus4A_out(29), complement2(28) 
                           => minus4A_out(28), complement2(27) => 
                           minus4A_out(27), complement2(26) => minus4A_out(26),
                           complement2(25) => minus4A_out(25), complement2(24) 
                           => minus4A_out(24), complement2(23) => 
                           minus4A_out(23), complement2(22) => minus4A_out(22),
                           complement2(21) => minus4A_out(21), complement2(20) 
                           => minus4A_out(20), complement2(19) => 
                           minus4A_out(19), complement2(18) => minus4A_out(18),
                           complement2(17) => minus4A_out(17), complement2(16) 
                           => minus4A_out(16), complement2(15) => 
                           minus4A_out(15), complement2(14) => minus4A_out(14),
                           complement2(13) => minus4A_out(13), complement2(12) 
                           => minus4A_out(12), complement2(11) => 
                           minus4A_out(11), complement2(10) => minus4A_out(10),
                           complement2(9) => minus4A_out(9), complement2(8) => 
                           minus4A_out(8), complement2(7) => minus4A_out(7), 
                           complement2(6) => minus4A_out(6), complement2(5) => 
                           minus4A_out(5), complement2(4) => minus4A_out(4), 
                           complement2(3) => minus4A_out(3), complement2(2) => 
                           minus4A_out(2), complement2(1) => minus4A_out(1), 
                           complement2(0) => minus4A_out(0));
   U3 : BUF_X1 port map( A => n13, Z => plus4A_out_43_port);
   U4 : BUF_X1 port map( A => n14, Z => plus4A_out_42_port);
   U5 : BUF_X1 port map( A => n10, Z => plus2A_out_47_port);
   U6 : BUF_X1 port map( A => n12, Z => plus4A_out_52_port);
   U7 : BUF_X1 port map( A => n9, Z => plus2A_out_48_port);
   U8 : BUF_X1 port map( A => n11, Z => plus4A_out_53_port);
   U9 : BUF_X1 port map( A => n8, Z => plus2A_out_57_port);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity ShiftnCompl_N64_13 is

   port( plusA : in std_logic_vector (63 downto 0);  plus2A_out, minus2A_out, 
         plus4A_out, minus4A_out : out std_logic_vector (63 downto 0));

end ShiftnCompl_N64_13;

architecture SYN_struct of ShiftnCompl_N64_13 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component complementer_N64_25
      port( input : in std_logic_vector (63 downto 0);  complement2 : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component complementer_N64_26
      port( input : in std_logic_vector (63 downto 0);  complement2 : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component shifter_N64_25
      port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component shifter_N64_26
      port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
            std_logic_vector (63 downto 0));
   end component;
   
   signal plus2A_out_63_port, plus2A_out_62_port, plus2A_out_61_port, 
      plus2A_out_60_port, plus2A_out_59_port, plus2A_out_58_port, n41, 
      plus2A_out_56_port, plus2A_out_55_port, plus2A_out_54_port, 
      plus2A_out_53_port, plus2A_out_52_port, plus2A_out_51_port, 
      plus2A_out_50_port, plus2A_out_49_port, n42, n43, plus2A_out_46_port, 
      plus2A_out_45_port, plus2A_out_44_port, plus2A_out_43_port, 
      plus2A_out_42_port, plus2A_out_41_port, plus2A_out_40_port, 
      plus2A_out_39_port, n44, n45, n46, plus2A_out_35_port, plus2A_out_34_port
      , plus2A_out_33_port, plus2A_out_32_port, plus2A_out_31_port, 
      plus2A_out_30_port, plus2A_out_29_port, plus2A_out_28_port, 
      plus2A_out_27_port, plus2A_out_26_port, plus2A_out_25_port, 
      plus2A_out_24_port, plus2A_out_23_port, plus2A_out_22_port, 
      plus2A_out_21_port, plus2A_out_20_port, plus2A_out_19_port, 
      plus2A_out_18_port, plus2A_out_17_port, plus2A_out_16_port, 
      plus2A_out_15_port, plus2A_out_14_port, plus2A_out_13_port, 
      plus2A_out_12_port, plus2A_out_11_port, plus2A_out_10_port, 
      plus2A_out_9_port, plus2A_out_8_port, plus2A_out_7_port, 
      plus2A_out_6_port, plus2A_out_5_port, plus2A_out_4_port, 
      plus2A_out_3_port, plus2A_out_2_port, plus2A_out_1_port, 
      plus2A_out_0_port, plus4A_out_63_port, plus4A_out_62_port, 
      plus4A_out_61_port, plus4A_out_60_port, plus4A_out_59_port, 
      plus4A_out_58_port, plus4A_out_57_port, plus4A_out_56_port, 
      plus4A_out_55_port, plus4A_out_54_port, n47, n48, plus4A_out_51_port, 
      plus4A_out_50_port, plus4A_out_49_port, plus4A_out_48_port, 
      plus4A_out_47_port, plus4A_out_46_port, plus4A_out_45_port, 
      plus4A_out_44_port, n49, n50, plus4A_out_41_port, plus4A_out_40_port, 
      plus4A_out_39_port, plus4A_out_38_port, plus4A_out_37_port, n51, n52, n53
      , n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, 
      n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, 
      plus4A_out_6_port, plus4A_out_5_port, plus4A_out_4_port, 
      plus4A_out_3_port, plus4A_out_2_port, plus4A_out_1_port, 
      plus4A_out_0_port, plus4A_out_7_port, plus4A_out_8_port, 
      plus4A_out_9_port, plus4A_out_10_port, plus4A_out_11_port, 
      plus4A_out_12_port, plus4A_out_13_port, plus4A_out_14_port, 
      plus4A_out_15_port, plus4A_out_16_port, plus4A_out_17_port, 
      plus4A_out_18_port, plus4A_out_19_port, plus4A_out_20_port, 
      plus4A_out_21_port, plus4A_out_22_port, plus4A_out_23_port, 
      plus4A_out_24_port, plus4A_out_25_port, plus4A_out_26_port, 
      plus4A_out_27_port, plus4A_out_28_port, plus4A_out_29_port, 
      plus4A_out_30_port, plus4A_out_31_port, plus4A_out_32_port, 
      plus4A_out_33_port, plus4A_out_34_port, plus4A_out_35_port, 
      plus4A_out_36_port, plus2A_out_36_port, plus2A_out_37_port, 
      plus2A_out_38_port, plus4A_out_42_port, plus4A_out_43_port, 
      plus2A_out_47_port, plus2A_out_48_port, plus4A_out_52_port, 
      plus4A_out_53_port, plus2A_out_57_port, n_3168, n_3169 : std_logic;

begin
   plus2A_out <= ( plus2A_out_63_port, plus2A_out_62_port, plus2A_out_61_port, 
      plus2A_out_60_port, plus2A_out_59_port, plus2A_out_58_port, 
      plus2A_out_57_port, plus2A_out_56_port, plus2A_out_55_port, 
      plus2A_out_54_port, plus2A_out_53_port, plus2A_out_52_port, 
      plus2A_out_51_port, plus2A_out_50_port, plus2A_out_49_port, 
      plus2A_out_48_port, plus2A_out_47_port, plus2A_out_46_port, 
      plus2A_out_45_port, plus2A_out_44_port, plus2A_out_43_port, 
      plus2A_out_42_port, plus2A_out_41_port, plus2A_out_40_port, 
      plus2A_out_39_port, plus2A_out_38_port, plus2A_out_37_port, 
      plus2A_out_36_port, plus2A_out_35_port, plus2A_out_34_port, 
      plus2A_out_33_port, plus2A_out_32_port, plus2A_out_31_port, 
      plus2A_out_30_port, plus2A_out_29_port, plus2A_out_28_port, 
      plus2A_out_27_port, plus2A_out_26_port, plus2A_out_25_port, 
      plus2A_out_24_port, plus2A_out_23_port, plus2A_out_22_port, 
      plus2A_out_21_port, plus2A_out_20_port, plus2A_out_19_port, 
      plus2A_out_18_port, plus2A_out_17_port, plus2A_out_16_port, 
      plus2A_out_15_port, plus2A_out_14_port, plus2A_out_13_port, 
      plus2A_out_12_port, plus2A_out_11_port, plus2A_out_10_port, 
      plus2A_out_9_port, plus2A_out_8_port, plus2A_out_7_port, 
      plus2A_out_6_port, plus2A_out_5_port, plus2A_out_4_port, 
      plus2A_out_3_port, plus2A_out_2_port, plus2A_out_1_port, 
      plus2A_out_0_port );
   plus4A_out <= ( plus4A_out_63_port, plus4A_out_62_port, plus4A_out_61_port, 
      plus4A_out_60_port, plus4A_out_59_port, plus4A_out_58_port, 
      plus4A_out_57_port, plus4A_out_56_port, plus4A_out_55_port, 
      plus4A_out_54_port, plus4A_out_53_port, plus4A_out_52_port, 
      plus4A_out_51_port, plus4A_out_50_port, plus4A_out_49_port, 
      plus4A_out_48_port, plus4A_out_47_port, plus4A_out_46_port, 
      plus4A_out_45_port, plus4A_out_44_port, plus4A_out_43_port, 
      plus4A_out_42_port, plus4A_out_41_port, plus4A_out_40_port, 
      plus4A_out_39_port, plus4A_out_38_port, plus4A_out_37_port, 
      plus4A_out_36_port, plus4A_out_35_port, plus4A_out_34_port, 
      plus4A_out_33_port, plus4A_out_32_port, plus4A_out_31_port, 
      plus4A_out_30_port, plus4A_out_29_port, plus4A_out_28_port, 
      plus4A_out_27_port, plus4A_out_26_port, plus4A_out_25_port, 
      plus4A_out_24_port, plus4A_out_23_port, plus4A_out_22_port, 
      plus4A_out_21_port, plus4A_out_20_port, plus4A_out_19_port, 
      plus4A_out_18_port, plus4A_out_17_port, plus4A_out_16_port, 
      plus4A_out_15_port, plus4A_out_14_port, plus4A_out_13_port, 
      plus4A_out_12_port, plus4A_out_11_port, plus4A_out_10_port, 
      plus4A_out_9_port, plus4A_out_8_port, plus4A_out_7_port, 
      plus4A_out_6_port, plus4A_out_5_port, plus4A_out_4_port, 
      plus4A_out_3_port, plus4A_out_2_port, plus4A_out_1_port, 
      plus4A_out_0_port );
   
   plus2A_out_0_port <= '0';
   plus4A_out_0_port <= '0';
   shifter_1 : shifter_N64_26 port map( input(63) => plusA(63), input(62) => 
                           plusA(62), input(61) => plusA(61), input(60) => 
                           plusA(60), input(59) => plusA(59), input(58) => 
                           plusA(58), input(57) => plusA(57), input(56) => 
                           plusA(56), input(55) => plusA(55), input(54) => 
                           plusA(54), input(53) => plusA(53), input(52) => 
                           plusA(52), input(51) => plusA(51), input(50) => 
                           plusA(50), input(49) => plusA(49), input(48) => 
                           plusA(48), input(47) => plusA(47), input(46) => 
                           plusA(46), input(45) => plusA(45), input(44) => 
                           plusA(44), input(43) => plusA(43), input(42) => 
                           plusA(42), input(41) => plusA(41), input(40) => 
                           plusA(40), input(39) => plusA(39), input(38) => 
                           plusA(38), input(37) => plusA(37), input(36) => 
                           plusA(36), input(35) => plusA(35), input(34) => 
                           plusA(34), input(33) => plusA(33), input(32) => 
                           plusA(32), input(31) => plusA(31), input(30) => 
                           plusA(30), input(29) => plusA(29), input(28) => 
                           plusA(28), input(27) => plusA(27), input(26) => 
                           plusA(26), input(25) => plusA(25), input(24) => 
                           plusA(24), input(23) => plusA(23), input(22) => 
                           plusA(22), input(21) => plusA(21), input(20) => 
                           plusA(20), input(19) => plusA(19), input(18) => 
                           plusA(18), input(17) => plusA(17), input(16) => 
                           plusA(16), input(15) => plusA(15), input(14) => 
                           plusA(14), input(13) => plusA(13), input(12) => 
                           plusA(12), input(11) => plusA(11), input(10) => 
                           plusA(10), input(9) => plusA(9), input(8) => 
                           plusA(8), input(7) => plusA(7), input(6) => plusA(6)
                           , input(5) => plusA(5), input(4) => plusA(4), 
                           input(3) => plusA(3), input(2) => plusA(2), input(1)
                           => plusA(1), input(0) => plusA(0), 
                           shiftLeftOnePos(63) => plus2A_out_63_port, 
                           shiftLeftOnePos(62) => plus2A_out_62_port, 
                           shiftLeftOnePos(61) => plus2A_out_61_port, 
                           shiftLeftOnePos(60) => plus2A_out_60_port, 
                           shiftLeftOnePos(59) => plus2A_out_59_port, 
                           shiftLeftOnePos(58) => plus2A_out_58_port, 
                           shiftLeftOnePos(57) => n41, shiftLeftOnePos(56) => 
                           plus2A_out_56_port, shiftLeftOnePos(55) => 
                           plus2A_out_55_port, shiftLeftOnePos(54) => 
                           plus2A_out_54_port, shiftLeftOnePos(53) => 
                           plus2A_out_53_port, shiftLeftOnePos(52) => 
                           plus2A_out_52_port, shiftLeftOnePos(51) => 
                           plus2A_out_51_port, shiftLeftOnePos(50) => 
                           plus2A_out_50_port, shiftLeftOnePos(49) => 
                           plus2A_out_49_port, shiftLeftOnePos(48) => n42, 
                           shiftLeftOnePos(47) => n43, shiftLeftOnePos(46) => 
                           plus2A_out_46_port, shiftLeftOnePos(45) => 
                           plus2A_out_45_port, shiftLeftOnePos(44) => 
                           plus2A_out_44_port, shiftLeftOnePos(43) => 
                           plus2A_out_43_port, shiftLeftOnePos(42) => 
                           plus2A_out_42_port, shiftLeftOnePos(41) => 
                           plus2A_out_41_port, shiftLeftOnePos(40) => 
                           plus2A_out_40_port, shiftLeftOnePos(39) => 
                           plus2A_out_39_port, shiftLeftOnePos(38) => n44, 
                           shiftLeftOnePos(37) => n45, shiftLeftOnePos(36) => 
                           n46, shiftLeftOnePos(35) => plus2A_out_35_port, 
                           shiftLeftOnePos(34) => plus2A_out_34_port, 
                           shiftLeftOnePos(33) => plus2A_out_33_port, 
                           shiftLeftOnePos(32) => plus2A_out_32_port, 
                           shiftLeftOnePos(31) => plus2A_out_31_port, 
                           shiftLeftOnePos(30) => plus2A_out_30_port, 
                           shiftLeftOnePos(29) => plus2A_out_29_port, 
                           shiftLeftOnePos(28) => plus2A_out_28_port, 
                           shiftLeftOnePos(27) => plus2A_out_27_port, 
                           shiftLeftOnePos(26) => plus2A_out_26_port, 
                           shiftLeftOnePos(25) => plus2A_out_25_port, 
                           shiftLeftOnePos(24) => plus2A_out_24_port, 
                           shiftLeftOnePos(23) => plus2A_out_23_port, 
                           shiftLeftOnePos(22) => plus2A_out_22_port, 
                           shiftLeftOnePos(21) => plus2A_out_21_port, 
                           shiftLeftOnePos(20) => plus2A_out_20_port, 
                           shiftLeftOnePos(19) => plus2A_out_19_port, 
                           shiftLeftOnePos(18) => plus2A_out_18_port, 
                           shiftLeftOnePos(17) => plus2A_out_17_port, 
                           shiftLeftOnePos(16) => plus2A_out_16_port, 
                           shiftLeftOnePos(15) => plus2A_out_15_port, 
                           shiftLeftOnePos(14) => plus2A_out_14_port, 
                           shiftLeftOnePos(13) => plus2A_out_13_port, 
                           shiftLeftOnePos(12) => plus2A_out_12_port, 
                           shiftLeftOnePos(11) => plus2A_out_11_port, 
                           shiftLeftOnePos(10) => plus2A_out_10_port, 
                           shiftLeftOnePos(9) => plus2A_out_9_port, 
                           shiftLeftOnePos(8) => plus2A_out_8_port, 
                           shiftLeftOnePos(7) => plus2A_out_7_port, 
                           shiftLeftOnePos(6) => plus2A_out_6_port, 
                           shiftLeftOnePos(5) => plus2A_out_5_port, 
                           shiftLeftOnePos(4) => plus2A_out_4_port, 
                           shiftLeftOnePos(3) => plus2A_out_3_port, 
                           shiftLeftOnePos(2) => plus2A_out_2_port, 
                           shiftLeftOnePos(1) => plus2A_out_1_port, 
                           shiftLeftOnePos(0) => n_3168);
   shifter_2 : shifter_N64_25 port map( input(63) => plus2A_out_63_port, 
                           input(62) => plus2A_out_62_port, input(61) => 
                           plus2A_out_61_port, input(60) => plus2A_out_60_port,
                           input(59) => plus2A_out_59_port, input(58) => 
                           plus2A_out_58_port, input(57) => plus2A_out_57_port,
                           input(56) => plus2A_out_56_port, input(55) => 
                           plus2A_out_55_port, input(54) => plus2A_out_54_port,
                           input(53) => plus2A_out_53_port, input(52) => 
                           plus2A_out_52_port, input(51) => plus2A_out_51_port,
                           input(50) => plus2A_out_50_port, input(49) => 
                           plus2A_out_49_port, input(48) => plus2A_out_48_port,
                           input(47) => plus2A_out_47_port, input(46) => 
                           plus2A_out_46_port, input(45) => plus2A_out_45_port,
                           input(44) => plus2A_out_44_port, input(43) => 
                           plus2A_out_43_port, input(42) => plus2A_out_42_port,
                           input(41) => plus2A_out_41_port, input(40) => 
                           plus2A_out_40_port, input(39) => plus2A_out_39_port,
                           input(38) => plus2A_out_38_port, input(37) => 
                           plus2A_out_37_port, input(36) => plus2A_out_36_port,
                           input(35) => plus2A_out_35_port, input(34) => 
                           plus2A_out_34_port, input(33) => plus2A_out_33_port,
                           input(32) => plus2A_out_32_port, input(31) => 
                           plus2A_out_31_port, input(30) => plus2A_out_30_port,
                           input(29) => plus2A_out_29_port, input(28) => 
                           plus2A_out_28_port, input(27) => plus2A_out_27_port,
                           input(26) => plus2A_out_26_port, input(25) => 
                           plus2A_out_25_port, input(24) => plus2A_out_24_port,
                           input(23) => plus2A_out_23_port, input(22) => 
                           plus2A_out_22_port, input(21) => plus2A_out_21_port,
                           input(20) => plus2A_out_20_port, input(19) => 
                           plus2A_out_19_port, input(18) => plus2A_out_18_port,
                           input(17) => plus2A_out_17_port, input(16) => 
                           plus2A_out_16_port, input(15) => plus2A_out_15_port,
                           input(14) => plus2A_out_14_port, input(13) => 
                           plus2A_out_13_port, input(12) => plus2A_out_12_port,
                           input(11) => plus2A_out_11_port, input(10) => 
                           plus2A_out_10_port, input(9) => plus2A_out_9_port, 
                           input(8) => plus2A_out_8_port, input(7) => 
                           plus2A_out_7_port, input(6) => plus2A_out_6_port, 
                           input(5) => plus2A_out_5_port, input(4) => 
                           plus2A_out_4_port, input(3) => plus2A_out_3_port, 
                           input(2) => plus2A_out_2_port, input(1) => 
                           plus2A_out_1_port, input(0) => plus2A_out_0_port, 
                           shiftLeftOnePos(63) => plus4A_out_63_port, 
                           shiftLeftOnePos(62) => plus4A_out_62_port, 
                           shiftLeftOnePos(61) => plus4A_out_61_port, 
                           shiftLeftOnePos(60) => plus4A_out_60_port, 
                           shiftLeftOnePos(59) => plus4A_out_59_port, 
                           shiftLeftOnePos(58) => plus4A_out_58_port, 
                           shiftLeftOnePos(57) => plus4A_out_57_port, 
                           shiftLeftOnePos(56) => plus4A_out_56_port, 
                           shiftLeftOnePos(55) => plus4A_out_55_port, 
                           shiftLeftOnePos(54) => plus4A_out_54_port, 
                           shiftLeftOnePos(53) => n47, shiftLeftOnePos(52) => 
                           n48, shiftLeftOnePos(51) => plus4A_out_51_port, 
                           shiftLeftOnePos(50) => plus4A_out_50_port, 
                           shiftLeftOnePos(49) => plus4A_out_49_port, 
                           shiftLeftOnePos(48) => plus4A_out_48_port, 
                           shiftLeftOnePos(47) => plus4A_out_47_port, 
                           shiftLeftOnePos(46) => plus4A_out_46_port, 
                           shiftLeftOnePos(45) => plus4A_out_45_port, 
                           shiftLeftOnePos(44) => plus4A_out_44_port, 
                           shiftLeftOnePos(43) => n49, shiftLeftOnePos(42) => 
                           n50, shiftLeftOnePos(41) => plus4A_out_41_port, 
                           shiftLeftOnePos(40) => plus4A_out_40_port, 
                           shiftLeftOnePos(39) => plus4A_out_39_port, 
                           shiftLeftOnePos(38) => plus4A_out_38_port, 
                           shiftLeftOnePos(37) => plus4A_out_37_port, 
                           shiftLeftOnePos(36) => n51, shiftLeftOnePos(35) => 
                           n52, shiftLeftOnePos(34) => n53, shiftLeftOnePos(33)
                           => n54, shiftLeftOnePos(32) => n55, 
                           shiftLeftOnePos(31) => n56, shiftLeftOnePos(30) => 
                           n57, shiftLeftOnePos(29) => n58, shiftLeftOnePos(28)
                           => n59, shiftLeftOnePos(27) => n60, 
                           shiftLeftOnePos(26) => n61, shiftLeftOnePos(25) => 
                           n62, shiftLeftOnePos(24) => n63, shiftLeftOnePos(23)
                           => n64, shiftLeftOnePos(22) => n65, 
                           shiftLeftOnePos(21) => n66, shiftLeftOnePos(20) => 
                           n67, shiftLeftOnePos(19) => n68, shiftLeftOnePos(18)
                           => n69, shiftLeftOnePos(17) => n70, 
                           shiftLeftOnePos(16) => n71, shiftLeftOnePos(15) => 
                           n72, shiftLeftOnePos(14) => n73, shiftLeftOnePos(13)
                           => n74, shiftLeftOnePos(12) => n75, 
                           shiftLeftOnePos(11) => n76, shiftLeftOnePos(10) => 
                           n77, shiftLeftOnePos(9) => n78, shiftLeftOnePos(8) 
                           => n79, shiftLeftOnePos(7) => n80, 
                           shiftLeftOnePos(6) => plus4A_out_6_port, 
                           shiftLeftOnePos(5) => plus4A_out_5_port, 
                           shiftLeftOnePos(4) => plus4A_out_4_port, 
                           shiftLeftOnePos(3) => plus4A_out_3_port, 
                           shiftLeftOnePos(2) => plus4A_out_2_port, 
                           shiftLeftOnePos(1) => plus4A_out_1_port, 
                           shiftLeftOnePos(0) => n_3169);
   complementer_1 : complementer_N64_26 port map( input(63) => 
                           plus2A_out_63_port, input(62) => plus2A_out_62_port,
                           input(61) => plus2A_out_61_port, input(60) => 
                           plus2A_out_60_port, input(59) => plus2A_out_59_port,
                           input(58) => plus2A_out_58_port, input(57) => 
                           plus2A_out_57_port, input(56) => plus2A_out_56_port,
                           input(55) => plus2A_out_55_port, input(54) => 
                           plus2A_out_54_port, input(53) => plus2A_out_53_port,
                           input(52) => plus2A_out_52_port, input(51) => 
                           plus2A_out_51_port, input(50) => plus2A_out_50_port,
                           input(49) => plus2A_out_49_port, input(48) => 
                           plus2A_out_48_port, input(47) => plus2A_out_47_port,
                           input(46) => plus2A_out_46_port, input(45) => 
                           plus2A_out_45_port, input(44) => plus2A_out_44_port,
                           input(43) => plus2A_out_43_port, input(42) => 
                           plus2A_out_42_port, input(41) => plus2A_out_41_port,
                           input(40) => plus2A_out_40_port, input(39) => 
                           plus2A_out_39_port, input(38) => plus2A_out_38_port,
                           input(37) => plus2A_out_37_port, input(36) => 
                           plus2A_out_36_port, input(35) => plus2A_out_35_port,
                           input(34) => plus2A_out_34_port, input(33) => 
                           plus2A_out_33_port, input(32) => plus2A_out_32_port,
                           input(31) => plus2A_out_31_port, input(30) => 
                           plus2A_out_30_port, input(29) => plus2A_out_29_port,
                           input(28) => plus2A_out_28_port, input(27) => 
                           plus2A_out_27_port, input(26) => plus2A_out_26_port,
                           input(25) => plus2A_out_25_port, input(24) => 
                           plus2A_out_24_port, input(23) => plus2A_out_23_port,
                           input(22) => plus2A_out_22_port, input(21) => 
                           plus2A_out_21_port, input(20) => plus2A_out_20_port,
                           input(19) => plus2A_out_19_port, input(18) => 
                           plus2A_out_18_port, input(17) => plus2A_out_17_port,
                           input(16) => plus2A_out_16_port, input(15) => 
                           plus2A_out_15_port, input(14) => plus2A_out_14_port,
                           input(13) => plus2A_out_13_port, input(12) => 
                           plus2A_out_12_port, input(11) => plus2A_out_11_port,
                           input(10) => plus2A_out_10_port, input(9) => 
                           plus2A_out_9_port, input(8) => plus2A_out_8_port, 
                           input(7) => plus2A_out_7_port, input(6) => 
                           plus2A_out_6_port, input(5) => plus2A_out_5_port, 
                           input(4) => plus2A_out_4_port, input(3) => 
                           plus2A_out_3_port, input(2) => plus2A_out_2_port, 
                           input(1) => plus2A_out_1_port, input(0) => 
                           plus2A_out_0_port, complement2(63) => 
                           minus2A_out(63), complement2(62) => minus2A_out(62),
                           complement2(61) => minus2A_out(61), complement2(60) 
                           => minus2A_out(60), complement2(59) => 
                           minus2A_out(59), complement2(58) => minus2A_out(58),
                           complement2(57) => minus2A_out(57), complement2(56) 
                           => minus2A_out(56), complement2(55) => 
                           minus2A_out(55), complement2(54) => minus2A_out(54),
                           complement2(53) => minus2A_out(53), complement2(52) 
                           => minus2A_out(52), complement2(51) => 
                           minus2A_out(51), complement2(50) => minus2A_out(50),
                           complement2(49) => minus2A_out(49), complement2(48) 
                           => minus2A_out(48), complement2(47) => 
                           minus2A_out(47), complement2(46) => minus2A_out(46),
                           complement2(45) => minus2A_out(45), complement2(44) 
                           => minus2A_out(44), complement2(43) => 
                           minus2A_out(43), complement2(42) => minus2A_out(42),
                           complement2(41) => minus2A_out(41), complement2(40) 
                           => minus2A_out(40), complement2(39) => 
                           minus2A_out(39), complement2(38) => minus2A_out(38),
                           complement2(37) => minus2A_out(37), complement2(36) 
                           => minus2A_out(36), complement2(35) => 
                           minus2A_out(35), complement2(34) => minus2A_out(34),
                           complement2(33) => minus2A_out(33), complement2(32) 
                           => minus2A_out(32), complement2(31) => 
                           minus2A_out(31), complement2(30) => minus2A_out(30),
                           complement2(29) => minus2A_out(29), complement2(28) 
                           => minus2A_out(28), complement2(27) => 
                           minus2A_out(27), complement2(26) => minus2A_out(26),
                           complement2(25) => minus2A_out(25), complement2(24) 
                           => minus2A_out(24), complement2(23) => 
                           minus2A_out(23), complement2(22) => minus2A_out(22),
                           complement2(21) => minus2A_out(21), complement2(20) 
                           => minus2A_out(20), complement2(19) => 
                           minus2A_out(19), complement2(18) => minus2A_out(18),
                           complement2(17) => minus2A_out(17), complement2(16) 
                           => minus2A_out(16), complement2(15) => 
                           minus2A_out(15), complement2(14) => minus2A_out(14),
                           complement2(13) => minus2A_out(13), complement2(12) 
                           => minus2A_out(12), complement2(11) => 
                           minus2A_out(11), complement2(10) => minus2A_out(10),
                           complement2(9) => minus2A_out(9), complement2(8) => 
                           minus2A_out(8), complement2(7) => minus2A_out(7), 
                           complement2(6) => minus2A_out(6), complement2(5) => 
                           minus2A_out(5), complement2(4) => minus2A_out(4), 
                           complement2(3) => minus2A_out(3), complement2(2) => 
                           minus2A_out(2), complement2(1) => minus2A_out(1), 
                           complement2(0) => minus2A_out(0));
   complementer_2 : complementer_N64_25 port map( input(63) => 
                           plus4A_out_63_port, input(62) => plus4A_out_62_port,
                           input(61) => plus4A_out_61_port, input(60) => 
                           plus4A_out_60_port, input(59) => plus4A_out_59_port,
                           input(58) => plus4A_out_58_port, input(57) => 
                           plus4A_out_57_port, input(56) => plus4A_out_56_port,
                           input(55) => plus4A_out_55_port, input(54) => 
                           plus4A_out_54_port, input(53) => plus4A_out_53_port,
                           input(52) => plus4A_out_52_port, input(51) => 
                           plus4A_out_51_port, input(50) => plus4A_out_50_port,
                           input(49) => plus4A_out_49_port, input(48) => 
                           plus4A_out_48_port, input(47) => plus4A_out_47_port,
                           input(46) => plus4A_out_46_port, input(45) => 
                           plus4A_out_45_port, input(44) => plus4A_out_44_port,
                           input(43) => plus4A_out_43_port, input(42) => 
                           plus4A_out_42_port, input(41) => plus4A_out_41_port,
                           input(40) => plus4A_out_40_port, input(39) => 
                           plus4A_out_39_port, input(38) => plus4A_out_38_port,
                           input(37) => plus4A_out_37_port, input(36) => 
                           plus4A_out_36_port, input(35) => plus4A_out_35_port,
                           input(34) => plus4A_out_34_port, input(33) => 
                           plus4A_out_33_port, input(32) => plus4A_out_32_port,
                           input(31) => plus4A_out_31_port, input(30) => 
                           plus4A_out_30_port, input(29) => plus4A_out_29_port,
                           input(28) => plus4A_out_28_port, input(27) => 
                           plus4A_out_27_port, input(26) => plus4A_out_26_port,
                           input(25) => plus4A_out_25_port, input(24) => 
                           plus4A_out_24_port, input(23) => plus4A_out_23_port,
                           input(22) => plus4A_out_22_port, input(21) => 
                           plus4A_out_21_port, input(20) => plus4A_out_20_port,
                           input(19) => plus4A_out_19_port, input(18) => 
                           plus4A_out_18_port, input(17) => plus4A_out_17_port,
                           input(16) => plus4A_out_16_port, input(15) => 
                           plus4A_out_15_port, input(14) => plus4A_out_14_port,
                           input(13) => plus4A_out_13_port, input(12) => 
                           plus4A_out_12_port, input(11) => plus4A_out_11_port,
                           input(10) => plus4A_out_10_port, input(9) => 
                           plus4A_out_9_port, input(8) => plus4A_out_8_port, 
                           input(7) => plus4A_out_7_port, input(6) => 
                           plus4A_out_6_port, input(5) => plus4A_out_5_port, 
                           input(4) => plus4A_out_4_port, input(3) => 
                           plus4A_out_3_port, input(2) => plus4A_out_2_port, 
                           input(1) => plus4A_out_1_port, input(0) => 
                           plus4A_out_0_port, complement2(63) => 
                           minus4A_out(63), complement2(62) => minus4A_out(62),
                           complement2(61) => minus4A_out(61), complement2(60) 
                           => minus4A_out(60), complement2(59) => 
                           minus4A_out(59), complement2(58) => minus4A_out(58),
                           complement2(57) => minus4A_out(57), complement2(56) 
                           => minus4A_out(56), complement2(55) => 
                           minus4A_out(55), complement2(54) => minus4A_out(54),
                           complement2(53) => minus4A_out(53), complement2(52) 
                           => minus4A_out(52), complement2(51) => 
                           minus4A_out(51), complement2(50) => minus4A_out(50),
                           complement2(49) => minus4A_out(49), complement2(48) 
                           => minus4A_out(48), complement2(47) => 
                           minus4A_out(47), complement2(46) => minus4A_out(46),
                           complement2(45) => minus4A_out(45), complement2(44) 
                           => minus4A_out(44), complement2(43) => 
                           minus4A_out(43), complement2(42) => minus4A_out(42),
                           complement2(41) => minus4A_out(41), complement2(40) 
                           => minus4A_out(40), complement2(39) => 
                           minus4A_out(39), complement2(38) => minus4A_out(38),
                           complement2(37) => minus4A_out(37), complement2(36) 
                           => minus4A_out(36), complement2(35) => 
                           minus4A_out(35), complement2(34) => minus4A_out(34),
                           complement2(33) => minus4A_out(33), complement2(32) 
                           => minus4A_out(32), complement2(31) => 
                           minus4A_out(31), complement2(30) => minus4A_out(30),
                           complement2(29) => minus4A_out(29), complement2(28) 
                           => minus4A_out(28), complement2(27) => 
                           minus4A_out(27), complement2(26) => minus4A_out(26),
                           complement2(25) => minus4A_out(25), complement2(24) 
                           => minus4A_out(24), complement2(23) => 
                           minus4A_out(23), complement2(22) => minus4A_out(22),
                           complement2(21) => minus4A_out(21), complement2(20) 
                           => minus4A_out(20), complement2(19) => 
                           minus4A_out(19), complement2(18) => minus4A_out(18),
                           complement2(17) => minus4A_out(17), complement2(16) 
                           => minus4A_out(16), complement2(15) => 
                           minus4A_out(15), complement2(14) => minus4A_out(14),
                           complement2(13) => minus4A_out(13), complement2(12) 
                           => minus4A_out(12), complement2(11) => 
                           minus4A_out(11), complement2(10) => minus4A_out(10),
                           complement2(9) => minus4A_out(9), complement2(8) => 
                           minus4A_out(8), complement2(7) => minus4A_out(7), 
                           complement2(6) => minus4A_out(6), complement2(5) => 
                           minus4A_out(5), complement2(4) => minus4A_out(4), 
                           complement2(3) => minus4A_out(3), complement2(2) => 
                           minus4A_out(2), complement2(1) => minus4A_out(1), 
                           complement2(0) => minus4A_out(0));
   U3 : CLKBUF_X1 port map( A => n68, Z => plus4A_out_19_port);
   U4 : CLKBUF_X1 port map( A => n76, Z => plus4A_out_11_port);
   U5 : CLKBUF_X1 port map( A => n66, Z => plus4A_out_21_port);
   U6 : CLKBUF_X1 port map( A => n70, Z => plus4A_out_17_port);
   U7 : CLKBUF_X1 port map( A => n74, Z => plus4A_out_13_port);
   U8 : CLKBUF_X1 port map( A => n69, Z => plus4A_out_18_port);
   U9 : CLKBUF_X1 port map( A => n73, Z => plus4A_out_14_port);
   U10 : CLKBUF_X1 port map( A => n67, Z => plus4A_out_20_port);
   U11 : CLKBUF_X1 port map( A => n80, Z => plus4A_out_7_port);
   U12 : CLKBUF_X1 port map( A => n79, Z => plus4A_out_8_port);
   U13 : CLKBUF_X1 port map( A => n72, Z => plus4A_out_15_port);
   U14 : BUF_X1 port map( A => n64, Z => plus4A_out_23_port);
   U15 : BUF_X1 port map( A => n65, Z => plus4A_out_22_port);
   U16 : CLKBUF_X1 port map( A => n71, Z => plus4A_out_16_port);
   U17 : CLKBUF_X1 port map( A => n75, Z => plus4A_out_12_port);
   U18 : BUF_X1 port map( A => n63, Z => plus4A_out_24_port);
   U19 : CLKBUF_X1 port map( A => n77, Z => plus4A_out_10_port);
   U20 : BUF_X1 port map( A => n52, Z => plus4A_out_35_port);
   U21 : BUF_X1 port map( A => n56, Z => plus4A_out_31_port);
   U22 : BUF_X1 port map( A => n60, Z => plus4A_out_27_port);
   U23 : BUF_X1 port map( A => n54, Z => plus4A_out_33_port);
   U24 : BUF_X1 port map( A => n58, Z => plus4A_out_29_port);
   U25 : BUF_X1 port map( A => n62, Z => plus4A_out_25_port);
   U26 : BUF_X1 port map( A => n53, Z => plus4A_out_34_port);
   U27 : BUF_X1 port map( A => n57, Z => plus4A_out_30_port);
   U28 : BUF_X1 port map( A => n61, Z => plus4A_out_26_port);
   U29 : BUF_X1 port map( A => n55, Z => plus4A_out_32_port);
   U30 : BUF_X1 port map( A => n59, Z => plus4A_out_28_port);
   U31 : BUF_X1 port map( A => n43, Z => plus2A_out_47_port);
   U32 : BUF_X1 port map( A => n45, Z => plus2A_out_37_port);
   U33 : BUF_X1 port map( A => n49, Z => plus4A_out_43_port);
   U34 : BUF_X1 port map( A => n50, Z => plus4A_out_42_port);
   U35 : BUF_X1 port map( A => n46, Z => plus2A_out_36_port);
   U36 : BUF_X1 port map( A => n51, Z => plus4A_out_36_port);
   U37 : BUF_X1 port map( A => n44, Z => plus2A_out_38_port);
   U38 : BUF_X1 port map( A => n41, Z => plus2A_out_57_port);
   U39 : BUF_X1 port map( A => n42, Z => plus2A_out_48_port);
   U40 : BUF_X1 port map( A => n48, Z => plus4A_out_52_port);
   U41 : BUF_X1 port map( A => n47, Z => plus4A_out_53_port);
   U42 : BUF_X1 port map( A => n78, Z => plus4A_out_9_port);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity ShiftnCompl_N64_14 is

   port( plusA : in std_logic_vector (63 downto 0);  plus2A_out, minus2A_out, 
         plus4A_out, minus4A_out : out std_logic_vector (63 downto 0));

end ShiftnCompl_N64_14;

architecture SYN_struct of ShiftnCompl_N64_14 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component complementer_N64_27
      port( input : in std_logic_vector (63 downto 0);  complement2 : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component complementer_N64_28
      port( input : in std_logic_vector (63 downto 0);  complement2 : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component shifter_N64_27
      port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component shifter_N64_28
      port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
            std_logic_vector (63 downto 0));
   end component;
   
   signal plus2A_out_63_port, plus2A_out_62_port, plus2A_out_61_port, 
      plus2A_out_60_port, plus2A_out_59_port, plus2A_out_58_port, n10, 
      plus2A_out_56_port, plus2A_out_55_port, plus2A_out_54_port, 
      plus2A_out_53_port, plus2A_out_52_port, plus2A_out_51_port, 
      plus2A_out_50_port, plus2A_out_49_port, n11, n12, plus2A_out_46_port, 
      plus2A_out_45_port, plus2A_out_44_port, plus2A_out_43_port, 
      plus2A_out_42_port, plus2A_out_41_port, plus2A_out_40_port, 
      plus2A_out_39_port, n13, n14, plus2A_out_36_port, plus2A_out_35_port, 
      plus2A_out_34_port, plus2A_out_33_port, plus2A_out_32_port, 
      plus2A_out_31_port, plus2A_out_30_port, plus2A_out_29_port, 
      plus2A_out_28_port, plus2A_out_27_port, plus2A_out_26_port, 
      plus2A_out_25_port, plus2A_out_24_port, plus2A_out_23_port, 
      plus2A_out_22_port, plus2A_out_21_port, plus2A_out_20_port, 
      plus2A_out_19_port, plus2A_out_18_port, plus2A_out_17_port, 
      plus2A_out_16_port, plus2A_out_15_port, plus2A_out_14_port, 
      plus2A_out_13_port, plus2A_out_12_port, plus2A_out_11_port, 
      plus2A_out_10_port, plus2A_out_9_port, plus2A_out_8_port, 
      plus2A_out_7_port, plus2A_out_6_port, plus2A_out_5_port, 
      plus2A_out_4_port, plus2A_out_3_port, plus2A_out_2_port, 
      plus2A_out_1_port, plus2A_out_0_port, plus4A_out_63_port, 
      plus4A_out_62_port, plus4A_out_61_port, plus4A_out_60_port, 
      plus4A_out_59_port, plus4A_out_58_port, plus4A_out_57_port, 
      plus4A_out_56_port, plus4A_out_55_port, plus4A_out_54_port, n15, n16, 
      plus4A_out_51_port, plus4A_out_50_port, plus4A_out_49_port, 
      plus4A_out_48_port, plus4A_out_47_port, plus4A_out_46_port, 
      plus4A_out_45_port, plus4A_out_44_port, n17, n18, plus4A_out_41_port, 
      plus4A_out_40_port, plus4A_out_39_port, plus4A_out_38_port, 
      plus4A_out_37_port, plus4A_out_36_port, plus4A_out_35_port, 
      plus4A_out_34_port, plus4A_out_33_port, plus4A_out_32_port, 
      plus4A_out_31_port, plus4A_out_30_port, plus4A_out_29_port, 
      plus4A_out_28_port, plus4A_out_27_port, plus4A_out_26_port, 
      plus4A_out_25_port, plus4A_out_24_port, plus4A_out_23_port, 
      plus4A_out_22_port, plus4A_out_21_port, plus4A_out_20_port, 
      plus4A_out_19_port, plus4A_out_18_port, plus4A_out_17_port, 
      plus4A_out_16_port, plus4A_out_15_port, plus4A_out_14_port, 
      plus4A_out_13_port, plus4A_out_12_port, plus4A_out_11_port, 
      plus4A_out_10_port, plus4A_out_9_port, plus4A_out_8_port, 
      plus4A_out_7_port, plus4A_out_6_port, plus4A_out_5_port, 
      plus4A_out_4_port, plus4A_out_3_port, plus4A_out_2_port, 
      plus4A_out_1_port, plus4A_out_0_port, plus2A_out_37_port, 
      plus2A_out_38_port, plus4A_out_42_port, plus4A_out_43_port, 
      plus2A_out_47_port, plus2A_out_48_port, plus4A_out_52_port, 
      plus4A_out_53_port, plus2A_out_57_port, n_3170, n_3171 : std_logic;

begin
   plus2A_out <= ( plus2A_out_63_port, plus2A_out_62_port, plus2A_out_61_port, 
      plus2A_out_60_port, plus2A_out_59_port, plus2A_out_58_port, 
      plus2A_out_57_port, plus2A_out_56_port, plus2A_out_55_port, 
      plus2A_out_54_port, plus2A_out_53_port, plus2A_out_52_port, 
      plus2A_out_51_port, plus2A_out_50_port, plus2A_out_49_port, 
      plus2A_out_48_port, plus2A_out_47_port, plus2A_out_46_port, 
      plus2A_out_45_port, plus2A_out_44_port, plus2A_out_43_port, 
      plus2A_out_42_port, plus2A_out_41_port, plus2A_out_40_port, 
      plus2A_out_39_port, plus2A_out_38_port, plus2A_out_37_port, 
      plus2A_out_36_port, plus2A_out_35_port, plus2A_out_34_port, 
      plus2A_out_33_port, plus2A_out_32_port, plus2A_out_31_port, 
      plus2A_out_30_port, plus2A_out_29_port, plus2A_out_28_port, 
      plus2A_out_27_port, plus2A_out_26_port, plus2A_out_25_port, 
      plus2A_out_24_port, plus2A_out_23_port, plus2A_out_22_port, 
      plus2A_out_21_port, plus2A_out_20_port, plus2A_out_19_port, 
      plus2A_out_18_port, plus2A_out_17_port, plus2A_out_16_port, 
      plus2A_out_15_port, plus2A_out_14_port, plus2A_out_13_port, 
      plus2A_out_12_port, plus2A_out_11_port, plus2A_out_10_port, 
      plus2A_out_9_port, plus2A_out_8_port, plus2A_out_7_port, 
      plus2A_out_6_port, plus2A_out_5_port, plus2A_out_4_port, 
      plus2A_out_3_port, plus2A_out_2_port, plus2A_out_1_port, 
      plus2A_out_0_port );
   plus4A_out <= ( plus4A_out_63_port, plus4A_out_62_port, plus4A_out_61_port, 
      plus4A_out_60_port, plus4A_out_59_port, plus4A_out_58_port, 
      plus4A_out_57_port, plus4A_out_56_port, plus4A_out_55_port, 
      plus4A_out_54_port, plus4A_out_53_port, plus4A_out_52_port, 
      plus4A_out_51_port, plus4A_out_50_port, plus4A_out_49_port, 
      plus4A_out_48_port, plus4A_out_47_port, plus4A_out_46_port, 
      plus4A_out_45_port, plus4A_out_44_port, plus4A_out_43_port, 
      plus4A_out_42_port, plus4A_out_41_port, plus4A_out_40_port, 
      plus4A_out_39_port, plus4A_out_38_port, plus4A_out_37_port, 
      plus4A_out_36_port, plus4A_out_35_port, plus4A_out_34_port, 
      plus4A_out_33_port, plus4A_out_32_port, plus4A_out_31_port, 
      plus4A_out_30_port, plus4A_out_29_port, plus4A_out_28_port, 
      plus4A_out_27_port, plus4A_out_26_port, plus4A_out_25_port, 
      plus4A_out_24_port, plus4A_out_23_port, plus4A_out_22_port, 
      plus4A_out_21_port, plus4A_out_20_port, plus4A_out_19_port, 
      plus4A_out_18_port, plus4A_out_17_port, plus4A_out_16_port, 
      plus4A_out_15_port, plus4A_out_14_port, plus4A_out_13_port, 
      plus4A_out_12_port, plus4A_out_11_port, plus4A_out_10_port, 
      plus4A_out_9_port, plus4A_out_8_port, plus4A_out_7_port, 
      plus4A_out_6_port, plus4A_out_5_port, plus4A_out_4_port, 
      plus4A_out_3_port, plus4A_out_2_port, plus4A_out_1_port, 
      plus4A_out_0_port );
   
   plus2A_out_0_port <= '0';
   plus4A_out_0_port <= '0';
   shifter_1 : shifter_N64_28 port map( input(63) => plusA(63), input(62) => 
                           plusA(62), input(61) => plusA(61), input(60) => 
                           plusA(60), input(59) => plusA(59), input(58) => 
                           plusA(58), input(57) => plusA(57), input(56) => 
                           plusA(56), input(55) => plusA(55), input(54) => 
                           plusA(54), input(53) => plusA(53), input(52) => 
                           plusA(52), input(51) => plusA(51), input(50) => 
                           plusA(50), input(49) => plusA(49), input(48) => 
                           plusA(48), input(47) => plusA(47), input(46) => 
                           plusA(46), input(45) => plusA(45), input(44) => 
                           plusA(44), input(43) => plusA(43), input(42) => 
                           plusA(42), input(41) => plusA(41), input(40) => 
                           plusA(40), input(39) => plusA(39), input(38) => 
                           plusA(38), input(37) => plusA(37), input(36) => 
                           plusA(36), input(35) => plusA(35), input(34) => 
                           plusA(34), input(33) => plusA(33), input(32) => 
                           plusA(32), input(31) => plusA(31), input(30) => 
                           plusA(30), input(29) => plusA(29), input(28) => 
                           plusA(28), input(27) => plusA(27), input(26) => 
                           plusA(26), input(25) => plusA(25), input(24) => 
                           plusA(24), input(23) => plusA(23), input(22) => 
                           plusA(22), input(21) => plusA(21), input(20) => 
                           plusA(20), input(19) => plusA(19), input(18) => 
                           plusA(18), input(17) => plusA(17), input(16) => 
                           plusA(16), input(15) => plusA(15), input(14) => 
                           plusA(14), input(13) => plusA(13), input(12) => 
                           plusA(12), input(11) => plusA(11), input(10) => 
                           plusA(10), input(9) => plusA(9), input(8) => 
                           plusA(8), input(7) => plusA(7), input(6) => plusA(6)
                           , input(5) => plusA(5), input(4) => plusA(4), 
                           input(3) => plusA(3), input(2) => plusA(2), input(1)
                           => plusA(1), input(0) => plusA(0), 
                           shiftLeftOnePos(63) => plus2A_out_63_port, 
                           shiftLeftOnePos(62) => plus2A_out_62_port, 
                           shiftLeftOnePos(61) => plus2A_out_61_port, 
                           shiftLeftOnePos(60) => plus2A_out_60_port, 
                           shiftLeftOnePos(59) => plus2A_out_59_port, 
                           shiftLeftOnePos(58) => plus2A_out_58_port, 
                           shiftLeftOnePos(57) => n10, shiftLeftOnePos(56) => 
                           plus2A_out_56_port, shiftLeftOnePos(55) => 
                           plus2A_out_55_port, shiftLeftOnePos(54) => 
                           plus2A_out_54_port, shiftLeftOnePos(53) => 
                           plus2A_out_53_port, shiftLeftOnePos(52) => 
                           plus2A_out_52_port, shiftLeftOnePos(51) => 
                           plus2A_out_51_port, shiftLeftOnePos(50) => 
                           plus2A_out_50_port, shiftLeftOnePos(49) => 
                           plus2A_out_49_port, shiftLeftOnePos(48) => n11, 
                           shiftLeftOnePos(47) => n12, shiftLeftOnePos(46) => 
                           plus2A_out_46_port, shiftLeftOnePos(45) => 
                           plus2A_out_45_port, shiftLeftOnePos(44) => 
                           plus2A_out_44_port, shiftLeftOnePos(43) => 
                           plus2A_out_43_port, shiftLeftOnePos(42) => 
                           plus2A_out_42_port, shiftLeftOnePos(41) => 
                           plus2A_out_41_port, shiftLeftOnePos(40) => 
                           plus2A_out_40_port, shiftLeftOnePos(39) => 
                           plus2A_out_39_port, shiftLeftOnePos(38) => n13, 
                           shiftLeftOnePos(37) => n14, shiftLeftOnePos(36) => 
                           plus2A_out_36_port, shiftLeftOnePos(35) => 
                           plus2A_out_35_port, shiftLeftOnePos(34) => 
                           plus2A_out_34_port, shiftLeftOnePos(33) => 
                           plus2A_out_33_port, shiftLeftOnePos(32) => 
                           plus2A_out_32_port, shiftLeftOnePos(31) => 
                           plus2A_out_31_port, shiftLeftOnePos(30) => 
                           plus2A_out_30_port, shiftLeftOnePos(29) => 
                           plus2A_out_29_port, shiftLeftOnePos(28) => 
                           plus2A_out_28_port, shiftLeftOnePos(27) => 
                           plus2A_out_27_port, shiftLeftOnePos(26) => 
                           plus2A_out_26_port, shiftLeftOnePos(25) => 
                           plus2A_out_25_port, shiftLeftOnePos(24) => 
                           plus2A_out_24_port, shiftLeftOnePos(23) => 
                           plus2A_out_23_port, shiftLeftOnePos(22) => 
                           plus2A_out_22_port, shiftLeftOnePos(21) => 
                           plus2A_out_21_port, shiftLeftOnePos(20) => 
                           plus2A_out_20_port, shiftLeftOnePos(19) => 
                           plus2A_out_19_port, shiftLeftOnePos(18) => 
                           plus2A_out_18_port, shiftLeftOnePos(17) => 
                           plus2A_out_17_port, shiftLeftOnePos(16) => 
                           plus2A_out_16_port, shiftLeftOnePos(15) => 
                           plus2A_out_15_port, shiftLeftOnePos(14) => 
                           plus2A_out_14_port, shiftLeftOnePos(13) => 
                           plus2A_out_13_port, shiftLeftOnePos(12) => 
                           plus2A_out_12_port, shiftLeftOnePos(11) => 
                           plus2A_out_11_port, shiftLeftOnePos(10) => 
                           plus2A_out_10_port, shiftLeftOnePos(9) => 
                           plus2A_out_9_port, shiftLeftOnePos(8) => 
                           plus2A_out_8_port, shiftLeftOnePos(7) => 
                           plus2A_out_7_port, shiftLeftOnePos(6) => 
                           plus2A_out_6_port, shiftLeftOnePos(5) => 
                           plus2A_out_5_port, shiftLeftOnePos(4) => 
                           plus2A_out_4_port, shiftLeftOnePos(3) => 
                           plus2A_out_3_port, shiftLeftOnePos(2) => 
                           plus2A_out_2_port, shiftLeftOnePos(1) => 
                           plus2A_out_1_port, shiftLeftOnePos(0) => n_3170);
   shifter_2 : shifter_N64_27 port map( input(63) => plus2A_out_63_port, 
                           input(62) => plus2A_out_62_port, input(61) => 
                           plus2A_out_61_port, input(60) => plus2A_out_60_port,
                           input(59) => plus2A_out_59_port, input(58) => 
                           plus2A_out_58_port, input(57) => plus2A_out_57_port,
                           input(56) => plus2A_out_56_port, input(55) => 
                           plus2A_out_55_port, input(54) => plus2A_out_54_port,
                           input(53) => plus2A_out_53_port, input(52) => 
                           plus2A_out_52_port, input(51) => plus2A_out_51_port,
                           input(50) => plus2A_out_50_port, input(49) => 
                           plus2A_out_49_port, input(48) => plus2A_out_48_port,
                           input(47) => plus2A_out_47_port, input(46) => 
                           plus2A_out_46_port, input(45) => plus2A_out_45_port,
                           input(44) => plus2A_out_44_port, input(43) => 
                           plus2A_out_43_port, input(42) => plus2A_out_42_port,
                           input(41) => plus2A_out_41_port, input(40) => 
                           plus2A_out_40_port, input(39) => plus2A_out_39_port,
                           input(38) => plus2A_out_38_port, input(37) => 
                           plus2A_out_37_port, input(36) => plus2A_out_36_port,
                           input(35) => plus2A_out_35_port, input(34) => 
                           plus2A_out_34_port, input(33) => plus2A_out_33_port,
                           input(32) => plus2A_out_32_port, input(31) => 
                           plus2A_out_31_port, input(30) => plus2A_out_30_port,
                           input(29) => plus2A_out_29_port, input(28) => 
                           plus2A_out_28_port, input(27) => plus2A_out_27_port,
                           input(26) => plus2A_out_26_port, input(25) => 
                           plus2A_out_25_port, input(24) => plus2A_out_24_port,
                           input(23) => plus2A_out_23_port, input(22) => 
                           plus2A_out_22_port, input(21) => plus2A_out_21_port,
                           input(20) => plus2A_out_20_port, input(19) => 
                           plus2A_out_19_port, input(18) => plus2A_out_18_port,
                           input(17) => plus2A_out_17_port, input(16) => 
                           plus2A_out_16_port, input(15) => plus2A_out_15_port,
                           input(14) => plus2A_out_14_port, input(13) => 
                           plus2A_out_13_port, input(12) => plus2A_out_12_port,
                           input(11) => plus2A_out_11_port, input(10) => 
                           plus2A_out_10_port, input(9) => plus2A_out_9_port, 
                           input(8) => plus2A_out_8_port, input(7) => 
                           plus2A_out_7_port, input(6) => plus2A_out_6_port, 
                           input(5) => plus2A_out_5_port, input(4) => 
                           plus2A_out_4_port, input(3) => plus2A_out_3_port, 
                           input(2) => plus2A_out_2_port, input(1) => 
                           plus2A_out_1_port, input(0) => plus2A_out_0_port, 
                           shiftLeftOnePos(63) => plus4A_out_63_port, 
                           shiftLeftOnePos(62) => plus4A_out_62_port, 
                           shiftLeftOnePos(61) => plus4A_out_61_port, 
                           shiftLeftOnePos(60) => plus4A_out_60_port, 
                           shiftLeftOnePos(59) => plus4A_out_59_port, 
                           shiftLeftOnePos(58) => plus4A_out_58_port, 
                           shiftLeftOnePos(57) => plus4A_out_57_port, 
                           shiftLeftOnePos(56) => plus4A_out_56_port, 
                           shiftLeftOnePos(55) => plus4A_out_55_port, 
                           shiftLeftOnePos(54) => plus4A_out_54_port, 
                           shiftLeftOnePos(53) => n15, shiftLeftOnePos(52) => 
                           n16, shiftLeftOnePos(51) => plus4A_out_51_port, 
                           shiftLeftOnePos(50) => plus4A_out_50_port, 
                           shiftLeftOnePos(49) => plus4A_out_49_port, 
                           shiftLeftOnePos(48) => plus4A_out_48_port, 
                           shiftLeftOnePos(47) => plus4A_out_47_port, 
                           shiftLeftOnePos(46) => plus4A_out_46_port, 
                           shiftLeftOnePos(45) => plus4A_out_45_port, 
                           shiftLeftOnePos(44) => plus4A_out_44_port, 
                           shiftLeftOnePos(43) => n17, shiftLeftOnePos(42) => 
                           n18, shiftLeftOnePos(41) => plus4A_out_41_port, 
                           shiftLeftOnePos(40) => plus4A_out_40_port, 
                           shiftLeftOnePos(39) => plus4A_out_39_port, 
                           shiftLeftOnePos(38) => plus4A_out_38_port, 
                           shiftLeftOnePos(37) => plus4A_out_37_port, 
                           shiftLeftOnePos(36) => plus4A_out_36_port, 
                           shiftLeftOnePos(35) => plus4A_out_35_port, 
                           shiftLeftOnePos(34) => plus4A_out_34_port, 
                           shiftLeftOnePos(33) => plus4A_out_33_port, 
                           shiftLeftOnePos(32) => plus4A_out_32_port, 
                           shiftLeftOnePos(31) => plus4A_out_31_port, 
                           shiftLeftOnePos(30) => plus4A_out_30_port, 
                           shiftLeftOnePos(29) => plus4A_out_29_port, 
                           shiftLeftOnePos(28) => plus4A_out_28_port, 
                           shiftLeftOnePos(27) => plus4A_out_27_port, 
                           shiftLeftOnePos(26) => plus4A_out_26_port, 
                           shiftLeftOnePos(25) => plus4A_out_25_port, 
                           shiftLeftOnePos(24) => plus4A_out_24_port, 
                           shiftLeftOnePos(23) => plus4A_out_23_port, 
                           shiftLeftOnePos(22) => plus4A_out_22_port, 
                           shiftLeftOnePos(21) => plus4A_out_21_port, 
                           shiftLeftOnePos(20) => plus4A_out_20_port, 
                           shiftLeftOnePos(19) => plus4A_out_19_port, 
                           shiftLeftOnePos(18) => plus4A_out_18_port, 
                           shiftLeftOnePos(17) => plus4A_out_17_port, 
                           shiftLeftOnePos(16) => plus4A_out_16_port, 
                           shiftLeftOnePos(15) => plus4A_out_15_port, 
                           shiftLeftOnePos(14) => plus4A_out_14_port, 
                           shiftLeftOnePos(13) => plus4A_out_13_port, 
                           shiftLeftOnePos(12) => plus4A_out_12_port, 
                           shiftLeftOnePos(11) => plus4A_out_11_port, 
                           shiftLeftOnePos(10) => plus4A_out_10_port, 
                           shiftLeftOnePos(9) => plus4A_out_9_port, 
                           shiftLeftOnePos(8) => plus4A_out_8_port, 
                           shiftLeftOnePos(7) => plus4A_out_7_port, 
                           shiftLeftOnePos(6) => plus4A_out_6_port, 
                           shiftLeftOnePos(5) => plus4A_out_5_port, 
                           shiftLeftOnePos(4) => plus4A_out_4_port, 
                           shiftLeftOnePos(3) => plus4A_out_3_port, 
                           shiftLeftOnePos(2) => plus4A_out_2_port, 
                           shiftLeftOnePos(1) => plus4A_out_1_port, 
                           shiftLeftOnePos(0) => n_3171);
   complementer_1 : complementer_N64_28 port map( input(63) => 
                           plus2A_out_63_port, input(62) => plus2A_out_62_port,
                           input(61) => plus2A_out_61_port, input(60) => 
                           plus2A_out_60_port, input(59) => plus2A_out_59_port,
                           input(58) => plus2A_out_58_port, input(57) => 
                           plus2A_out_57_port, input(56) => plus2A_out_56_port,
                           input(55) => plus2A_out_55_port, input(54) => 
                           plus2A_out_54_port, input(53) => plus2A_out_53_port,
                           input(52) => plus2A_out_52_port, input(51) => 
                           plus2A_out_51_port, input(50) => plus2A_out_50_port,
                           input(49) => plus2A_out_49_port, input(48) => 
                           plus2A_out_48_port, input(47) => plus2A_out_47_port,
                           input(46) => plus2A_out_46_port, input(45) => 
                           plus2A_out_45_port, input(44) => plus2A_out_44_port,
                           input(43) => plus2A_out_43_port, input(42) => 
                           plus2A_out_42_port, input(41) => plus2A_out_41_port,
                           input(40) => plus2A_out_40_port, input(39) => 
                           plus2A_out_39_port, input(38) => plus2A_out_38_port,
                           input(37) => plus2A_out_37_port, input(36) => 
                           plus2A_out_36_port, input(35) => plus2A_out_35_port,
                           input(34) => plus2A_out_34_port, input(33) => 
                           plus2A_out_33_port, input(32) => plus2A_out_32_port,
                           input(31) => plus2A_out_31_port, input(30) => 
                           plus2A_out_30_port, input(29) => plus2A_out_29_port,
                           input(28) => plus2A_out_28_port, input(27) => 
                           plus2A_out_27_port, input(26) => plus2A_out_26_port,
                           input(25) => plus2A_out_25_port, input(24) => 
                           plus2A_out_24_port, input(23) => plus2A_out_23_port,
                           input(22) => plus2A_out_22_port, input(21) => 
                           plus2A_out_21_port, input(20) => plus2A_out_20_port,
                           input(19) => plus2A_out_19_port, input(18) => 
                           plus2A_out_18_port, input(17) => plus2A_out_17_port,
                           input(16) => plus2A_out_16_port, input(15) => 
                           plus2A_out_15_port, input(14) => plus2A_out_14_port,
                           input(13) => plus2A_out_13_port, input(12) => 
                           plus2A_out_12_port, input(11) => plus2A_out_11_port,
                           input(10) => plus2A_out_10_port, input(9) => 
                           plus2A_out_9_port, input(8) => plus2A_out_8_port, 
                           input(7) => plus2A_out_7_port, input(6) => 
                           plus2A_out_6_port, input(5) => plus2A_out_5_port, 
                           input(4) => plus2A_out_4_port, input(3) => 
                           plus2A_out_3_port, input(2) => plus2A_out_2_port, 
                           input(1) => plus2A_out_1_port, input(0) => 
                           plus2A_out_0_port, complement2(63) => 
                           minus2A_out(63), complement2(62) => minus2A_out(62),
                           complement2(61) => minus2A_out(61), complement2(60) 
                           => minus2A_out(60), complement2(59) => 
                           minus2A_out(59), complement2(58) => minus2A_out(58),
                           complement2(57) => minus2A_out(57), complement2(56) 
                           => minus2A_out(56), complement2(55) => 
                           minus2A_out(55), complement2(54) => minus2A_out(54),
                           complement2(53) => minus2A_out(53), complement2(52) 
                           => minus2A_out(52), complement2(51) => 
                           minus2A_out(51), complement2(50) => minus2A_out(50),
                           complement2(49) => minus2A_out(49), complement2(48) 
                           => minus2A_out(48), complement2(47) => 
                           minus2A_out(47), complement2(46) => minus2A_out(46),
                           complement2(45) => minus2A_out(45), complement2(44) 
                           => minus2A_out(44), complement2(43) => 
                           minus2A_out(43), complement2(42) => minus2A_out(42),
                           complement2(41) => minus2A_out(41), complement2(40) 
                           => minus2A_out(40), complement2(39) => 
                           minus2A_out(39), complement2(38) => minus2A_out(38),
                           complement2(37) => minus2A_out(37), complement2(36) 
                           => minus2A_out(36), complement2(35) => 
                           minus2A_out(35), complement2(34) => minus2A_out(34),
                           complement2(33) => minus2A_out(33), complement2(32) 
                           => minus2A_out(32), complement2(31) => 
                           minus2A_out(31), complement2(30) => minus2A_out(30),
                           complement2(29) => minus2A_out(29), complement2(28) 
                           => minus2A_out(28), complement2(27) => 
                           minus2A_out(27), complement2(26) => minus2A_out(26),
                           complement2(25) => minus2A_out(25), complement2(24) 
                           => minus2A_out(24), complement2(23) => 
                           minus2A_out(23), complement2(22) => minus2A_out(22),
                           complement2(21) => minus2A_out(21), complement2(20) 
                           => minus2A_out(20), complement2(19) => 
                           minus2A_out(19), complement2(18) => minus2A_out(18),
                           complement2(17) => minus2A_out(17), complement2(16) 
                           => minus2A_out(16), complement2(15) => 
                           minus2A_out(15), complement2(14) => minus2A_out(14),
                           complement2(13) => minus2A_out(13), complement2(12) 
                           => minus2A_out(12), complement2(11) => 
                           minus2A_out(11), complement2(10) => minus2A_out(10),
                           complement2(9) => minus2A_out(9), complement2(8) => 
                           minus2A_out(8), complement2(7) => minus2A_out(7), 
                           complement2(6) => minus2A_out(6), complement2(5) => 
                           minus2A_out(5), complement2(4) => minus2A_out(4), 
                           complement2(3) => minus2A_out(3), complement2(2) => 
                           minus2A_out(2), complement2(1) => minus2A_out(1), 
                           complement2(0) => minus2A_out(0));
   complementer_2 : complementer_N64_27 port map( input(63) => 
                           plus4A_out_63_port, input(62) => plus4A_out_62_port,
                           input(61) => plus4A_out_61_port, input(60) => 
                           plus4A_out_60_port, input(59) => plus4A_out_59_port,
                           input(58) => plus4A_out_58_port, input(57) => 
                           plus4A_out_57_port, input(56) => plus4A_out_56_port,
                           input(55) => plus4A_out_55_port, input(54) => 
                           plus4A_out_54_port, input(53) => plus4A_out_53_port,
                           input(52) => plus4A_out_52_port, input(51) => 
                           plus4A_out_51_port, input(50) => plus4A_out_50_port,
                           input(49) => plus4A_out_49_port, input(48) => 
                           plus4A_out_48_port, input(47) => plus4A_out_47_port,
                           input(46) => plus4A_out_46_port, input(45) => 
                           plus4A_out_45_port, input(44) => plus4A_out_44_port,
                           input(43) => plus4A_out_43_port, input(42) => 
                           plus4A_out_42_port, input(41) => plus4A_out_41_port,
                           input(40) => plus4A_out_40_port, input(39) => 
                           plus4A_out_39_port, input(38) => plus4A_out_38_port,
                           input(37) => plus4A_out_37_port, input(36) => 
                           plus4A_out_36_port, input(35) => plus4A_out_35_port,
                           input(34) => plus4A_out_34_port, input(33) => 
                           plus4A_out_33_port, input(32) => plus4A_out_32_port,
                           input(31) => plus4A_out_31_port, input(30) => 
                           plus4A_out_30_port, input(29) => plus4A_out_29_port,
                           input(28) => plus4A_out_28_port, input(27) => 
                           plus4A_out_27_port, input(26) => plus4A_out_26_port,
                           input(25) => plus4A_out_25_port, input(24) => 
                           plus4A_out_24_port, input(23) => plus4A_out_23_port,
                           input(22) => plus4A_out_22_port, input(21) => 
                           plus4A_out_21_port, input(20) => plus4A_out_20_port,
                           input(19) => plus4A_out_19_port, input(18) => 
                           plus4A_out_18_port, input(17) => plus4A_out_17_port,
                           input(16) => plus4A_out_16_port, input(15) => 
                           plus4A_out_15_port, input(14) => plus4A_out_14_port,
                           input(13) => plus4A_out_13_port, input(12) => 
                           plus4A_out_12_port, input(11) => plus4A_out_11_port,
                           input(10) => plus4A_out_10_port, input(9) => 
                           plus4A_out_9_port, input(8) => plus4A_out_8_port, 
                           input(7) => plus4A_out_7_port, input(6) => 
                           plus4A_out_6_port, input(5) => plus4A_out_5_port, 
                           input(4) => plus4A_out_4_port, input(3) => 
                           plus4A_out_3_port, input(2) => plus4A_out_2_port, 
                           input(1) => plus4A_out_1_port, input(0) => 
                           plus4A_out_0_port, complement2(63) => 
                           minus4A_out(63), complement2(62) => minus4A_out(62),
                           complement2(61) => minus4A_out(61), complement2(60) 
                           => minus4A_out(60), complement2(59) => 
                           minus4A_out(59), complement2(58) => minus4A_out(58),
                           complement2(57) => minus4A_out(57), complement2(56) 
                           => minus4A_out(56), complement2(55) => 
                           minus4A_out(55), complement2(54) => minus4A_out(54),
                           complement2(53) => minus4A_out(53), complement2(52) 
                           => minus4A_out(52), complement2(51) => 
                           minus4A_out(51), complement2(50) => minus4A_out(50),
                           complement2(49) => minus4A_out(49), complement2(48) 
                           => minus4A_out(48), complement2(47) => 
                           minus4A_out(47), complement2(46) => minus4A_out(46),
                           complement2(45) => minus4A_out(45), complement2(44) 
                           => minus4A_out(44), complement2(43) => 
                           minus4A_out(43), complement2(42) => minus4A_out(42),
                           complement2(41) => minus4A_out(41), complement2(40) 
                           => minus4A_out(40), complement2(39) => 
                           minus4A_out(39), complement2(38) => minus4A_out(38),
                           complement2(37) => minus4A_out(37), complement2(36) 
                           => minus4A_out(36), complement2(35) => 
                           minus4A_out(35), complement2(34) => minus4A_out(34),
                           complement2(33) => minus4A_out(33), complement2(32) 
                           => minus4A_out(32), complement2(31) => 
                           minus4A_out(31), complement2(30) => minus4A_out(30),
                           complement2(29) => minus4A_out(29), complement2(28) 
                           => minus4A_out(28), complement2(27) => 
                           minus4A_out(27), complement2(26) => minus4A_out(26),
                           complement2(25) => minus4A_out(25), complement2(24) 
                           => minus4A_out(24), complement2(23) => 
                           minus4A_out(23), complement2(22) => minus4A_out(22),
                           complement2(21) => minus4A_out(21), complement2(20) 
                           => minus4A_out(20), complement2(19) => 
                           minus4A_out(19), complement2(18) => minus4A_out(18),
                           complement2(17) => minus4A_out(17), complement2(16) 
                           => minus4A_out(16), complement2(15) => 
                           minus4A_out(15), complement2(14) => minus4A_out(14),
                           complement2(13) => minus4A_out(13), complement2(12) 
                           => minus4A_out(12), complement2(11) => 
                           minus4A_out(11), complement2(10) => minus4A_out(10),
                           complement2(9) => minus4A_out(9), complement2(8) => 
                           minus4A_out(8), complement2(7) => minus4A_out(7), 
                           complement2(6) => minus4A_out(6), complement2(5) => 
                           minus4A_out(5), complement2(4) => minus4A_out(4), 
                           complement2(3) => minus4A_out(3), complement2(2) => 
                           minus4A_out(2), complement2(1) => minus4A_out(1), 
                           complement2(0) => minus4A_out(0));
   U3 : BUF_X1 port map( A => n17, Z => plus4A_out_43_port);
   U4 : BUF_X1 port map( A => n18, Z => plus4A_out_42_port);
   U5 : BUF_X1 port map( A => n16, Z => plus4A_out_52_port);
   U6 : BUF_X1 port map( A => n15, Z => plus4A_out_53_port);
   U7 : BUF_X1 port map( A => n14, Z => plus2A_out_37_port);
   U8 : BUF_X1 port map( A => n12, Z => plus2A_out_47_port);
   U9 : BUF_X1 port map( A => n13, Z => plus2A_out_38_port);
   U10 : BUF_X1 port map( A => n10, Z => plus2A_out_57_port);
   U11 : BUF_X1 port map( A => n11, Z => plus2A_out_48_port);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity RCA_N64_0 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_N64_0;

architecture SYN_STRUCTURAL of RCA_N64_0 is

   component FA_897
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_898
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_899
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_900
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_901
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_902
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_903
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_904
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_905
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_906
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_907
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_908
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_909
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_910
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_911
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_912
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_913
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_914
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_915
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_916
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_917
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_918
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_919
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_920
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_921
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_922
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_923
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_924
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_925
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_926
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_927
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_928
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_929
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_930
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_931
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_932
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_933
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_934
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_935
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_936
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_937
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_938
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_939
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_940
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_941
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_942
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_943
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_944
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_945
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_946
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_947
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_948
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_949
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_950
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_951
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_952
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_953
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_954
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_955
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_956
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_957
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_958
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_959
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_0
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_0 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_959 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_958 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_957 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_956 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_955 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_954 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_953 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_952 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_951 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_950 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_949 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_948 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_947 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_946 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_945 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_944 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_943 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_942 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_941 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_940 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_939 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_938 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_937 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_936 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_935 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_934 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_933 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_932 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_931 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_930 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_929 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_928 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_927 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_926 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_925 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_924 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_923 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_922 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_921 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_920 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_919 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_918 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_917 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_916 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_915 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_914 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_913 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_912 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_911 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_910 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_909 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_908 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_907 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_906 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_905 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_904 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_903 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_902 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_901 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_900 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_899 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_898 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_897 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity ShiftnCompl_N64_0 is

   port( plusA : in std_logic_vector (63 downto 0);  plus2A_out, minus2A_out, 
         plus4A_out, minus4A_out : out std_logic_vector (63 downto 0));

end ShiftnCompl_N64_0;

architecture SYN_struct of ShiftnCompl_N64_0 is

   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component complementer_N64_29
      port( input : in std_logic_vector (63 downto 0);  complement2 : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component complementer_N64_30
      port( input : in std_logic_vector (63 downto 0);  complement2 : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component shifter_N64_29
      port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component shifter_N64_30
      port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
            std_logic_vector (63 downto 0));
   end component;
   
   signal plus2A_out_63_port, plus2A_out_62_port, plus2A_out_61_port, 
      plus2A_out_60_port, plus2A_out_59_port, plus2A_out_58_port, n40, 
      plus2A_out_56_port, plus2A_out_55_port, plus2A_out_54_port, 
      plus2A_out_53_port, plus2A_out_52_port, plus2A_out_51_port, 
      plus2A_out_50_port, plus2A_out_49_port, n41, n42, plus2A_out_46_port, 
      plus2A_out_45_port, plus2A_out_44_port, plus2A_out_43_port, 
      plus2A_out_42_port, plus2A_out_41_port, plus2A_out_40_port, 
      plus2A_out_39_port, n43, n44, plus2A_out_36_port, plus2A_out_35_port, 
      plus2A_out_34_port, plus2A_out_33_port, plus2A_out_32_port, n45, n46, n47
      , n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, 
      n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, 
      plus2A_out_1_port, plus2A_out_0_port, plus4A_out_63_port, 
      plus4A_out_62_port, plus4A_out_61_port, plus4A_out_60_port, 
      plus4A_out_59_port, plus4A_out_58_port, plus4A_out_57_port, 
      plus4A_out_56_port, plus4A_out_55_port, plus4A_out_54_port, n75, n76, 
      plus4A_out_51_port, plus4A_out_50_port, plus4A_out_49_port, 
      plus4A_out_48_port, plus4A_out_47_port, plus4A_out_46_port, 
      plus4A_out_45_port, plus4A_out_44_port, n77, n78, plus4A_out_41_port, 
      plus4A_out_40_port, plus4A_out_39_port, plus4A_out_38_port, 
      plus4A_out_37_port, plus4A_out_36_port, plus4A_out_35_port, 
      plus4A_out_34_port, plus4A_out_33_port, plus4A_out_32_port, 
      plus4A_out_31_port, plus4A_out_30_port, plus4A_out_29_port, 
      plus4A_out_28_port, plus4A_out_27_port, plus4A_out_26_port, 
      plus4A_out_25_port, plus4A_out_24_port, plus4A_out_23_port, 
      plus4A_out_22_port, plus4A_out_21_port, plus4A_out_20_port, 
      plus4A_out_19_port, plus4A_out_18_port, plus4A_out_17_port, 
      plus4A_out_16_port, plus4A_out_15_port, plus4A_out_14_port, 
      plus4A_out_13_port, plus4A_out_12_port, plus4A_out_11_port, 
      plus4A_out_10_port, plus4A_out_9_port, plus4A_out_8_port, 
      plus4A_out_7_port, plus4A_out_6_port, plus4A_out_5_port, 
      plus4A_out_4_port, plus4A_out_3_port, plus4A_out_2_port, 
      plus4A_out_1_port, plus4A_out_0_port, plus2A_out_2_port, 
      plus2A_out_3_port, plus2A_out_4_port, plus2A_out_5_port, 
      plus2A_out_6_port, plus2A_out_7_port, plus2A_out_8_port, 
      plus2A_out_9_port, plus2A_out_10_port, plus2A_out_11_port, 
      plus2A_out_12_port, plus2A_out_13_port, plus2A_out_14_port, 
      plus2A_out_15_port, plus2A_out_16_port, plus2A_out_17_port, 
      plus2A_out_18_port, plus2A_out_19_port, plus2A_out_20_port, 
      plus2A_out_21_port, plus2A_out_22_port, plus2A_out_23_port, 
      plus2A_out_24_port, plus2A_out_25_port, plus2A_out_26_port, 
      plus2A_out_27_port, plus2A_out_28_port, plus2A_out_29_port, 
      plus2A_out_30_port, plus2A_out_31_port, plus2A_out_37_port, 
      plus2A_out_38_port, plus4A_out_42_port, plus4A_out_43_port, 
      plus2A_out_47_port, plus2A_out_48_port, plus4A_out_52_port, 
      plus4A_out_53_port, plus2A_out_57_port, n_3172, n_3173 : std_logic;

begin
   plus2A_out <= ( plus2A_out_63_port, plus2A_out_62_port, plus2A_out_61_port, 
      plus2A_out_60_port, plus2A_out_59_port, plus2A_out_58_port, 
      plus2A_out_57_port, plus2A_out_56_port, plus2A_out_55_port, 
      plus2A_out_54_port, plus2A_out_53_port, plus2A_out_52_port, 
      plus2A_out_51_port, plus2A_out_50_port, plus2A_out_49_port, 
      plus2A_out_48_port, plus2A_out_47_port, plus2A_out_46_port, 
      plus2A_out_45_port, plus2A_out_44_port, plus2A_out_43_port, 
      plus2A_out_42_port, plus2A_out_41_port, plus2A_out_40_port, 
      plus2A_out_39_port, plus2A_out_38_port, plus2A_out_37_port, 
      plus2A_out_36_port, plus2A_out_35_port, plus2A_out_34_port, 
      plus2A_out_33_port, plus2A_out_32_port, plus2A_out_31_port, 
      plus2A_out_30_port, plus2A_out_29_port, plus2A_out_28_port, 
      plus2A_out_27_port, plus2A_out_26_port, plus2A_out_25_port, 
      plus2A_out_24_port, plus2A_out_23_port, plus2A_out_22_port, 
      plus2A_out_21_port, plus2A_out_20_port, plus2A_out_19_port, 
      plus2A_out_18_port, plus2A_out_17_port, plus2A_out_16_port, 
      plus2A_out_15_port, plus2A_out_14_port, plus2A_out_13_port, 
      plus2A_out_12_port, plus2A_out_11_port, plus2A_out_10_port, 
      plus2A_out_9_port, plus2A_out_8_port, plus2A_out_7_port, 
      plus2A_out_6_port, plus2A_out_5_port, plus2A_out_4_port, 
      plus2A_out_3_port, plus2A_out_2_port, plus2A_out_1_port, 
      plus2A_out_0_port );
   plus4A_out <= ( plus4A_out_63_port, plus4A_out_62_port, plus4A_out_61_port, 
      plus4A_out_60_port, plus4A_out_59_port, plus4A_out_58_port, 
      plus4A_out_57_port, plus4A_out_56_port, plus4A_out_55_port, 
      plus4A_out_54_port, plus4A_out_53_port, plus4A_out_52_port, 
      plus4A_out_51_port, plus4A_out_50_port, plus4A_out_49_port, 
      plus4A_out_48_port, plus4A_out_47_port, plus4A_out_46_port, 
      plus4A_out_45_port, plus4A_out_44_port, plus4A_out_43_port, 
      plus4A_out_42_port, plus4A_out_41_port, plus4A_out_40_port, 
      plus4A_out_39_port, plus4A_out_38_port, plus4A_out_37_port, 
      plus4A_out_36_port, plus4A_out_35_port, plus4A_out_34_port, 
      plus4A_out_33_port, plus4A_out_32_port, plus4A_out_31_port, 
      plus4A_out_30_port, plus4A_out_29_port, plus4A_out_28_port, 
      plus4A_out_27_port, plus4A_out_26_port, plus4A_out_25_port, 
      plus4A_out_24_port, plus4A_out_23_port, plus4A_out_22_port, 
      plus4A_out_21_port, plus4A_out_20_port, plus4A_out_19_port, 
      plus4A_out_18_port, plus4A_out_17_port, plus4A_out_16_port, 
      plus4A_out_15_port, plus4A_out_14_port, plus4A_out_13_port, 
      plus4A_out_12_port, plus4A_out_11_port, plus4A_out_10_port, 
      plus4A_out_9_port, plus4A_out_8_port, plus4A_out_7_port, 
      plus4A_out_6_port, plus4A_out_5_port, plus4A_out_4_port, 
      plus4A_out_3_port, plus4A_out_2_port, plus4A_out_1_port, 
      plus4A_out_0_port );
   
   plus2A_out_0_port <= '0';
   plus4A_out_0_port <= '0';
   shifter_1 : shifter_N64_30 port map( input(63) => plusA(63), input(62) => 
                           plusA(62), input(61) => plusA(61), input(60) => 
                           plusA(60), input(59) => plusA(59), input(58) => 
                           plusA(58), input(57) => plusA(57), input(56) => 
                           plusA(56), input(55) => plusA(55), input(54) => 
                           plusA(54), input(53) => plusA(53), input(52) => 
                           plusA(52), input(51) => plusA(51), input(50) => 
                           plusA(50), input(49) => plusA(49), input(48) => 
                           plusA(48), input(47) => plusA(47), input(46) => 
                           plusA(46), input(45) => plusA(45), input(44) => 
                           plusA(44), input(43) => plusA(43), input(42) => 
                           plusA(42), input(41) => plusA(41), input(40) => 
                           plusA(40), input(39) => plusA(39), input(38) => 
                           plusA(38), input(37) => plusA(37), input(36) => 
                           plusA(36), input(35) => plusA(35), input(34) => 
                           plusA(34), input(33) => plusA(33), input(32) => 
                           plusA(32), input(31) => plusA(31), input(30) => 
                           plusA(30), input(29) => plusA(29), input(28) => 
                           plusA(28), input(27) => plusA(27), input(26) => 
                           plusA(26), input(25) => plusA(25), input(24) => 
                           plusA(24), input(23) => plusA(23), input(22) => 
                           plusA(22), input(21) => plusA(21), input(20) => 
                           plusA(20), input(19) => plusA(19), input(18) => 
                           plusA(18), input(17) => plusA(17), input(16) => 
                           plusA(16), input(15) => plusA(15), input(14) => 
                           plusA(14), input(13) => plusA(13), input(12) => 
                           plusA(12), input(11) => plusA(11), input(10) => 
                           plusA(10), input(9) => plusA(9), input(8) => 
                           plusA(8), input(7) => plusA(7), input(6) => plusA(6)
                           , input(5) => plusA(5), input(4) => plusA(4), 
                           input(3) => plusA(3), input(2) => plusA(2), input(1)
                           => plusA(1), input(0) => plusA(0), 
                           shiftLeftOnePos(63) => plus2A_out_63_port, 
                           shiftLeftOnePos(62) => plus2A_out_62_port, 
                           shiftLeftOnePos(61) => plus2A_out_61_port, 
                           shiftLeftOnePos(60) => plus2A_out_60_port, 
                           shiftLeftOnePos(59) => plus2A_out_59_port, 
                           shiftLeftOnePos(58) => plus2A_out_58_port, 
                           shiftLeftOnePos(57) => n40, shiftLeftOnePos(56) => 
                           plus2A_out_56_port, shiftLeftOnePos(55) => 
                           plus2A_out_55_port, shiftLeftOnePos(54) => 
                           plus2A_out_54_port, shiftLeftOnePos(53) => 
                           plus2A_out_53_port, shiftLeftOnePos(52) => 
                           plus2A_out_52_port, shiftLeftOnePos(51) => 
                           plus2A_out_51_port, shiftLeftOnePos(50) => 
                           plus2A_out_50_port, shiftLeftOnePos(49) => 
                           plus2A_out_49_port, shiftLeftOnePos(48) => n41, 
                           shiftLeftOnePos(47) => n42, shiftLeftOnePos(46) => 
                           plus2A_out_46_port, shiftLeftOnePos(45) => 
                           plus2A_out_45_port, shiftLeftOnePos(44) => 
                           plus2A_out_44_port, shiftLeftOnePos(43) => 
                           plus2A_out_43_port, shiftLeftOnePos(42) => 
                           plus2A_out_42_port, shiftLeftOnePos(41) => 
                           plus2A_out_41_port, shiftLeftOnePos(40) => 
                           plus2A_out_40_port, shiftLeftOnePos(39) => 
                           plus2A_out_39_port, shiftLeftOnePos(38) => n43, 
                           shiftLeftOnePos(37) => n44, shiftLeftOnePos(36) => 
                           plus2A_out_36_port, shiftLeftOnePos(35) => 
                           plus2A_out_35_port, shiftLeftOnePos(34) => 
                           plus2A_out_34_port, shiftLeftOnePos(33) => 
                           plus2A_out_33_port, shiftLeftOnePos(32) => 
                           plus2A_out_32_port, shiftLeftOnePos(31) => n45, 
                           shiftLeftOnePos(30) => n46, shiftLeftOnePos(29) => 
                           n47, shiftLeftOnePos(28) => n48, shiftLeftOnePos(27)
                           => n49, shiftLeftOnePos(26) => n50, 
                           shiftLeftOnePos(25) => n51, shiftLeftOnePos(24) => 
                           n52, shiftLeftOnePos(23) => n53, shiftLeftOnePos(22)
                           => n54, shiftLeftOnePos(21) => n55, 
                           shiftLeftOnePos(20) => n56, shiftLeftOnePos(19) => 
                           n57, shiftLeftOnePos(18) => n58, shiftLeftOnePos(17)
                           => n59, shiftLeftOnePos(16) => n60, 
                           shiftLeftOnePos(15) => n61, shiftLeftOnePos(14) => 
                           n62, shiftLeftOnePos(13) => n63, shiftLeftOnePos(12)
                           => n64, shiftLeftOnePos(11) => n65, 
                           shiftLeftOnePos(10) => n66, shiftLeftOnePos(9) => 
                           n67, shiftLeftOnePos(8) => n68, shiftLeftOnePos(7) 
                           => n69, shiftLeftOnePos(6) => n70, 
                           shiftLeftOnePos(5) => n71, shiftLeftOnePos(4) => n72
                           , shiftLeftOnePos(3) => n73, shiftLeftOnePos(2) => 
                           n74, shiftLeftOnePos(1) => plus2A_out_1_port, 
                           shiftLeftOnePos(0) => n_3172);
   shifter_2 : shifter_N64_29 port map( input(63) => plus2A_out_63_port, 
                           input(62) => plus2A_out_62_port, input(61) => 
                           plus2A_out_61_port, input(60) => plus2A_out_60_port,
                           input(59) => plus2A_out_59_port, input(58) => 
                           plus2A_out_58_port, input(57) => plus2A_out_57_port,
                           input(56) => plus2A_out_56_port, input(55) => 
                           plus2A_out_55_port, input(54) => plus2A_out_54_port,
                           input(53) => plus2A_out_53_port, input(52) => 
                           plus2A_out_52_port, input(51) => plus2A_out_51_port,
                           input(50) => plus2A_out_50_port, input(49) => 
                           plus2A_out_49_port, input(48) => plus2A_out_48_port,
                           input(47) => plus2A_out_47_port, input(46) => 
                           plus2A_out_46_port, input(45) => plus2A_out_45_port,
                           input(44) => plus2A_out_44_port, input(43) => 
                           plus2A_out_43_port, input(42) => plus2A_out_42_port,
                           input(41) => plus2A_out_41_port, input(40) => 
                           plus2A_out_40_port, input(39) => plus2A_out_39_port,
                           input(38) => plus2A_out_38_port, input(37) => 
                           plus2A_out_37_port, input(36) => plus2A_out_36_port,
                           input(35) => plus2A_out_35_port, input(34) => 
                           plus2A_out_34_port, input(33) => plus2A_out_33_port,
                           input(32) => plus2A_out_32_port, input(31) => 
                           plus2A_out_31_port, input(30) => plus2A_out_30_port,
                           input(29) => plus2A_out_29_port, input(28) => 
                           plus2A_out_28_port, input(27) => plus2A_out_27_port,
                           input(26) => plus2A_out_26_port, input(25) => 
                           plus2A_out_25_port, input(24) => plus2A_out_24_port,
                           input(23) => plus2A_out_23_port, input(22) => 
                           plus2A_out_22_port, input(21) => plus2A_out_21_port,
                           input(20) => plus2A_out_20_port, input(19) => 
                           plus2A_out_19_port, input(18) => plus2A_out_18_port,
                           input(17) => plus2A_out_17_port, input(16) => 
                           plus2A_out_16_port, input(15) => plus2A_out_15_port,
                           input(14) => plus2A_out_14_port, input(13) => 
                           plus2A_out_13_port, input(12) => plus2A_out_12_port,
                           input(11) => plus2A_out_11_port, input(10) => 
                           plus2A_out_10_port, input(9) => plus2A_out_9_port, 
                           input(8) => plus2A_out_8_port, input(7) => 
                           plus2A_out_7_port, input(6) => plus2A_out_6_port, 
                           input(5) => plus2A_out_5_port, input(4) => 
                           plus2A_out_4_port, input(3) => plus2A_out_3_port, 
                           input(2) => plus2A_out_2_port, input(1) => 
                           plus2A_out_1_port, input(0) => plus2A_out_0_port, 
                           shiftLeftOnePos(63) => plus4A_out_63_port, 
                           shiftLeftOnePos(62) => plus4A_out_62_port, 
                           shiftLeftOnePos(61) => plus4A_out_61_port, 
                           shiftLeftOnePos(60) => plus4A_out_60_port, 
                           shiftLeftOnePos(59) => plus4A_out_59_port, 
                           shiftLeftOnePos(58) => plus4A_out_58_port, 
                           shiftLeftOnePos(57) => plus4A_out_57_port, 
                           shiftLeftOnePos(56) => plus4A_out_56_port, 
                           shiftLeftOnePos(55) => plus4A_out_55_port, 
                           shiftLeftOnePos(54) => plus4A_out_54_port, 
                           shiftLeftOnePos(53) => n75, shiftLeftOnePos(52) => 
                           n76, shiftLeftOnePos(51) => plus4A_out_51_port, 
                           shiftLeftOnePos(50) => plus4A_out_50_port, 
                           shiftLeftOnePos(49) => plus4A_out_49_port, 
                           shiftLeftOnePos(48) => plus4A_out_48_port, 
                           shiftLeftOnePos(47) => plus4A_out_47_port, 
                           shiftLeftOnePos(46) => plus4A_out_46_port, 
                           shiftLeftOnePos(45) => plus4A_out_45_port, 
                           shiftLeftOnePos(44) => plus4A_out_44_port, 
                           shiftLeftOnePos(43) => n77, shiftLeftOnePos(42) => 
                           n78, shiftLeftOnePos(41) => plus4A_out_41_port, 
                           shiftLeftOnePos(40) => plus4A_out_40_port, 
                           shiftLeftOnePos(39) => plus4A_out_39_port, 
                           shiftLeftOnePos(38) => plus4A_out_38_port, 
                           shiftLeftOnePos(37) => plus4A_out_37_port, 
                           shiftLeftOnePos(36) => plus4A_out_36_port, 
                           shiftLeftOnePos(35) => plus4A_out_35_port, 
                           shiftLeftOnePos(34) => plus4A_out_34_port, 
                           shiftLeftOnePos(33) => plus4A_out_33_port, 
                           shiftLeftOnePos(32) => plus4A_out_32_port, 
                           shiftLeftOnePos(31) => plus4A_out_31_port, 
                           shiftLeftOnePos(30) => plus4A_out_30_port, 
                           shiftLeftOnePos(29) => plus4A_out_29_port, 
                           shiftLeftOnePos(28) => plus4A_out_28_port, 
                           shiftLeftOnePos(27) => plus4A_out_27_port, 
                           shiftLeftOnePos(26) => plus4A_out_26_port, 
                           shiftLeftOnePos(25) => plus4A_out_25_port, 
                           shiftLeftOnePos(24) => plus4A_out_24_port, 
                           shiftLeftOnePos(23) => plus4A_out_23_port, 
                           shiftLeftOnePos(22) => plus4A_out_22_port, 
                           shiftLeftOnePos(21) => plus4A_out_21_port, 
                           shiftLeftOnePos(20) => plus4A_out_20_port, 
                           shiftLeftOnePos(19) => plus4A_out_19_port, 
                           shiftLeftOnePos(18) => plus4A_out_18_port, 
                           shiftLeftOnePos(17) => plus4A_out_17_port, 
                           shiftLeftOnePos(16) => plus4A_out_16_port, 
                           shiftLeftOnePos(15) => plus4A_out_15_port, 
                           shiftLeftOnePos(14) => plus4A_out_14_port, 
                           shiftLeftOnePos(13) => plus4A_out_13_port, 
                           shiftLeftOnePos(12) => plus4A_out_12_port, 
                           shiftLeftOnePos(11) => plus4A_out_11_port, 
                           shiftLeftOnePos(10) => plus4A_out_10_port, 
                           shiftLeftOnePos(9) => plus4A_out_9_port, 
                           shiftLeftOnePos(8) => plus4A_out_8_port, 
                           shiftLeftOnePos(7) => plus4A_out_7_port, 
                           shiftLeftOnePos(6) => plus4A_out_6_port, 
                           shiftLeftOnePos(5) => plus4A_out_5_port, 
                           shiftLeftOnePos(4) => plus4A_out_4_port, 
                           shiftLeftOnePos(3) => plus4A_out_3_port, 
                           shiftLeftOnePos(2) => plus4A_out_2_port, 
                           shiftLeftOnePos(1) => plus4A_out_1_port, 
                           shiftLeftOnePos(0) => n_3173);
   complementer_1 : complementer_N64_30 port map( input(63) => 
                           plus2A_out_63_port, input(62) => plus2A_out_62_port,
                           input(61) => plus2A_out_61_port, input(60) => 
                           plus2A_out_60_port, input(59) => plus2A_out_59_port,
                           input(58) => plus2A_out_58_port, input(57) => 
                           plus2A_out_57_port, input(56) => plus2A_out_56_port,
                           input(55) => plus2A_out_55_port, input(54) => 
                           plus2A_out_54_port, input(53) => plus2A_out_53_port,
                           input(52) => plus2A_out_52_port, input(51) => 
                           plus2A_out_51_port, input(50) => plus2A_out_50_port,
                           input(49) => plus2A_out_49_port, input(48) => 
                           plus2A_out_48_port, input(47) => plus2A_out_47_port,
                           input(46) => plus2A_out_46_port, input(45) => 
                           plus2A_out_45_port, input(44) => plus2A_out_44_port,
                           input(43) => plus2A_out_43_port, input(42) => 
                           plus2A_out_42_port, input(41) => plus2A_out_41_port,
                           input(40) => plus2A_out_40_port, input(39) => 
                           plus2A_out_39_port, input(38) => plus2A_out_38_port,
                           input(37) => plus2A_out_37_port, input(36) => 
                           plus2A_out_36_port, input(35) => plus2A_out_35_port,
                           input(34) => plus2A_out_34_port, input(33) => 
                           plus2A_out_33_port, input(32) => plus2A_out_32_port,
                           input(31) => plus2A_out_31_port, input(30) => 
                           plus2A_out_30_port, input(29) => plus2A_out_29_port,
                           input(28) => plus2A_out_28_port, input(27) => 
                           plus2A_out_27_port, input(26) => plus2A_out_26_port,
                           input(25) => plus2A_out_25_port, input(24) => 
                           plus2A_out_24_port, input(23) => plus2A_out_23_port,
                           input(22) => plus2A_out_22_port, input(21) => 
                           plus2A_out_21_port, input(20) => plus2A_out_20_port,
                           input(19) => plus2A_out_19_port, input(18) => 
                           plus2A_out_18_port, input(17) => plus2A_out_17_port,
                           input(16) => plus2A_out_16_port, input(15) => 
                           plus2A_out_15_port, input(14) => plus2A_out_14_port,
                           input(13) => plus2A_out_13_port, input(12) => 
                           plus2A_out_12_port, input(11) => plus2A_out_11_port,
                           input(10) => plus2A_out_10_port, input(9) => 
                           plus2A_out_9_port, input(8) => plus2A_out_8_port, 
                           input(7) => plus2A_out_7_port, input(6) => 
                           plus2A_out_6_port, input(5) => plus2A_out_5_port, 
                           input(4) => plus2A_out_4_port, input(3) => 
                           plus2A_out_3_port, input(2) => plus2A_out_2_port, 
                           input(1) => plus2A_out_1_port, input(0) => 
                           plus2A_out_0_port, complement2(63) => 
                           minus2A_out(63), complement2(62) => minus2A_out(62),
                           complement2(61) => minus2A_out(61), complement2(60) 
                           => minus2A_out(60), complement2(59) => 
                           minus2A_out(59), complement2(58) => minus2A_out(58),
                           complement2(57) => minus2A_out(57), complement2(56) 
                           => minus2A_out(56), complement2(55) => 
                           minus2A_out(55), complement2(54) => minus2A_out(54),
                           complement2(53) => minus2A_out(53), complement2(52) 
                           => minus2A_out(52), complement2(51) => 
                           minus2A_out(51), complement2(50) => minus2A_out(50),
                           complement2(49) => minus2A_out(49), complement2(48) 
                           => minus2A_out(48), complement2(47) => 
                           minus2A_out(47), complement2(46) => minus2A_out(46),
                           complement2(45) => minus2A_out(45), complement2(44) 
                           => minus2A_out(44), complement2(43) => 
                           minus2A_out(43), complement2(42) => minus2A_out(42),
                           complement2(41) => minus2A_out(41), complement2(40) 
                           => minus2A_out(40), complement2(39) => 
                           minus2A_out(39), complement2(38) => minus2A_out(38),
                           complement2(37) => minus2A_out(37), complement2(36) 
                           => minus2A_out(36), complement2(35) => 
                           minus2A_out(35), complement2(34) => minus2A_out(34),
                           complement2(33) => minus2A_out(33), complement2(32) 
                           => minus2A_out(32), complement2(31) => 
                           minus2A_out(31), complement2(30) => minus2A_out(30),
                           complement2(29) => minus2A_out(29), complement2(28) 
                           => minus2A_out(28), complement2(27) => 
                           minus2A_out(27), complement2(26) => minus2A_out(26),
                           complement2(25) => minus2A_out(25), complement2(24) 
                           => minus2A_out(24), complement2(23) => 
                           minus2A_out(23), complement2(22) => minus2A_out(22),
                           complement2(21) => minus2A_out(21), complement2(20) 
                           => minus2A_out(20), complement2(19) => 
                           minus2A_out(19), complement2(18) => minus2A_out(18),
                           complement2(17) => minus2A_out(17), complement2(16) 
                           => minus2A_out(16), complement2(15) => 
                           minus2A_out(15), complement2(14) => minus2A_out(14),
                           complement2(13) => minus2A_out(13), complement2(12) 
                           => minus2A_out(12), complement2(11) => 
                           minus2A_out(11), complement2(10) => minus2A_out(10),
                           complement2(9) => minus2A_out(9), complement2(8) => 
                           minus2A_out(8), complement2(7) => minus2A_out(7), 
                           complement2(6) => minus2A_out(6), complement2(5) => 
                           minus2A_out(5), complement2(4) => minus2A_out(4), 
                           complement2(3) => minus2A_out(3), complement2(2) => 
                           minus2A_out(2), complement2(1) => minus2A_out(1), 
                           complement2(0) => minus2A_out(0));
   complementer_2 : complementer_N64_29 port map( input(63) => 
                           plus4A_out_63_port, input(62) => plus4A_out_62_port,
                           input(61) => plus4A_out_61_port, input(60) => 
                           plus4A_out_60_port, input(59) => plus4A_out_59_port,
                           input(58) => plus4A_out_58_port, input(57) => 
                           plus4A_out_57_port, input(56) => plus4A_out_56_port,
                           input(55) => plus4A_out_55_port, input(54) => 
                           plus4A_out_54_port, input(53) => plus4A_out_53_port,
                           input(52) => plus4A_out_52_port, input(51) => 
                           plus4A_out_51_port, input(50) => plus4A_out_50_port,
                           input(49) => plus4A_out_49_port, input(48) => 
                           plus4A_out_48_port, input(47) => plus4A_out_47_port,
                           input(46) => plus4A_out_46_port, input(45) => 
                           plus4A_out_45_port, input(44) => plus4A_out_44_port,
                           input(43) => plus4A_out_43_port, input(42) => 
                           plus4A_out_42_port, input(41) => plus4A_out_41_port,
                           input(40) => plus4A_out_40_port, input(39) => 
                           plus4A_out_39_port, input(38) => plus4A_out_38_port,
                           input(37) => plus4A_out_37_port, input(36) => 
                           plus4A_out_36_port, input(35) => plus4A_out_35_port,
                           input(34) => plus4A_out_34_port, input(33) => 
                           plus4A_out_33_port, input(32) => plus4A_out_32_port,
                           input(31) => plus4A_out_31_port, input(30) => 
                           plus4A_out_30_port, input(29) => plus4A_out_29_port,
                           input(28) => plus4A_out_28_port, input(27) => 
                           plus4A_out_27_port, input(26) => plus4A_out_26_port,
                           input(25) => plus4A_out_25_port, input(24) => 
                           plus4A_out_24_port, input(23) => plus4A_out_23_port,
                           input(22) => plus4A_out_22_port, input(21) => 
                           plus4A_out_21_port, input(20) => plus4A_out_20_port,
                           input(19) => plus4A_out_19_port, input(18) => 
                           plus4A_out_18_port, input(17) => plus4A_out_17_port,
                           input(16) => plus4A_out_16_port, input(15) => 
                           plus4A_out_15_port, input(14) => plus4A_out_14_port,
                           input(13) => plus4A_out_13_port, input(12) => 
                           plus4A_out_12_port, input(11) => plus4A_out_11_port,
                           input(10) => plus4A_out_10_port, input(9) => 
                           plus4A_out_9_port, input(8) => plus4A_out_8_port, 
                           input(7) => plus4A_out_7_port, input(6) => 
                           plus4A_out_6_port, input(5) => plus4A_out_5_port, 
                           input(4) => plus4A_out_4_port, input(3) => 
                           plus4A_out_3_port, input(2) => plus4A_out_2_port, 
                           input(1) => plus4A_out_1_port, input(0) => 
                           plus4A_out_0_port, complement2(63) => 
                           minus4A_out(63), complement2(62) => minus4A_out(62),
                           complement2(61) => minus4A_out(61), complement2(60) 
                           => minus4A_out(60), complement2(59) => 
                           minus4A_out(59), complement2(58) => minus4A_out(58),
                           complement2(57) => minus4A_out(57), complement2(56) 
                           => minus4A_out(56), complement2(55) => 
                           minus4A_out(55), complement2(54) => minus4A_out(54),
                           complement2(53) => minus4A_out(53), complement2(52) 
                           => minus4A_out(52), complement2(51) => 
                           minus4A_out(51), complement2(50) => minus4A_out(50),
                           complement2(49) => minus4A_out(49), complement2(48) 
                           => minus4A_out(48), complement2(47) => 
                           minus4A_out(47), complement2(46) => minus4A_out(46),
                           complement2(45) => minus4A_out(45), complement2(44) 
                           => minus4A_out(44), complement2(43) => 
                           minus4A_out(43), complement2(42) => minus4A_out(42),
                           complement2(41) => minus4A_out(41), complement2(40) 
                           => minus4A_out(40), complement2(39) => 
                           minus4A_out(39), complement2(38) => minus4A_out(38),
                           complement2(37) => minus4A_out(37), complement2(36) 
                           => minus4A_out(36), complement2(35) => 
                           minus4A_out(35), complement2(34) => minus4A_out(34),
                           complement2(33) => minus4A_out(33), complement2(32) 
                           => minus4A_out(32), complement2(31) => 
                           minus4A_out(31), complement2(30) => minus4A_out(30),
                           complement2(29) => minus4A_out(29), complement2(28) 
                           => minus4A_out(28), complement2(27) => 
                           minus4A_out(27), complement2(26) => minus4A_out(26),
                           complement2(25) => minus4A_out(25), complement2(24) 
                           => minus4A_out(24), complement2(23) => 
                           minus4A_out(23), complement2(22) => minus4A_out(22),
                           complement2(21) => minus4A_out(21), complement2(20) 
                           => minus4A_out(20), complement2(19) => 
                           minus4A_out(19), complement2(18) => minus4A_out(18),
                           complement2(17) => minus4A_out(17), complement2(16) 
                           => minus4A_out(16), complement2(15) => 
                           minus4A_out(15), complement2(14) => minus4A_out(14),
                           complement2(13) => minus4A_out(13), complement2(12) 
                           => minus4A_out(12), complement2(11) => 
                           minus4A_out(11), complement2(10) => minus4A_out(10),
                           complement2(9) => minus4A_out(9), complement2(8) => 
                           minus4A_out(8), complement2(7) => minus4A_out(7), 
                           complement2(6) => minus4A_out(6), complement2(5) => 
                           minus4A_out(5), complement2(4) => minus4A_out(4), 
                           complement2(3) => minus4A_out(3), complement2(2) => 
                           minus4A_out(2), complement2(1) => minus4A_out(1), 
                           complement2(0) => minus4A_out(0));
   U3 : BUF_X2 port map( A => n74, Z => plus2A_out_2_port);
   U4 : BUF_X1 port map( A => n72, Z => plus2A_out_4_port);
   U5 : BUF_X1 port map( A => n57, Z => plus2A_out_19_port);
   U6 : BUF_X1 port map( A => n61, Z => plus2A_out_15_port);
   U7 : BUF_X1 port map( A => n49, Z => plus2A_out_27_port);
   U8 : BUF_X1 port map( A => n53, Z => plus2A_out_23_port);
   U9 : BUF_X1 port map( A => n55, Z => plus2A_out_21_port);
   U10 : BUF_X1 port map( A => n59, Z => plus2A_out_17_port);
   U11 : BUF_X1 port map( A => n67, Z => plus2A_out_9_port);
   U12 : BUF_X1 port map( A => n63, Z => plus2A_out_13_port);
   U13 : BUF_X1 port map( A => n51, Z => plus2A_out_25_port);
   U14 : BUF_X1 port map( A => n54, Z => plus2A_out_22_port);
   U15 : BUF_X1 port map( A => n70, Z => plus2A_out_6_port);
   U16 : BUF_X1 port map( A => n58, Z => plus2A_out_18_port);
   U17 : BUF_X1 port map( A => n62, Z => plus2A_out_14_port);
   U18 : BUF_X1 port map( A => n50, Z => plus2A_out_26_port);
   U19 : BUF_X1 port map( A => n56, Z => plus2A_out_20_port);
   U20 : BUF_X1 port map( A => n68, Z => plus2A_out_8_port);
   U21 : BUF_X1 port map( A => n60, Z => plus2A_out_16_port);
   U22 : BUF_X1 port map( A => n64, Z => plus2A_out_12_port);
   U23 : BUF_X1 port map( A => n52, Z => plus2A_out_24_port);
   U24 : BUF_X1 port map( A => n45, Z => plus2A_out_31_port);
   U25 : BUF_X1 port map( A => n47, Z => plus2A_out_29_port);
   U26 : BUF_X1 port map( A => n44, Z => plus2A_out_37_port);
   U27 : BUF_X1 port map( A => n46, Z => plus2A_out_30_port);
   U28 : BUF_X1 port map( A => n43, Z => plus2A_out_38_port);
   U29 : BUF_X1 port map( A => n48, Z => plus2A_out_28_port);
   U30 : BUF_X1 port map( A => n42, Z => plus2A_out_47_port);
   U31 : BUF_X1 port map( A => n77, Z => plus4A_out_43_port);
   U32 : BUF_X1 port map( A => n78, Z => plus4A_out_42_port);
   U33 : BUF_X1 port map( A => n41, Z => plus2A_out_48_port);
   U34 : BUF_X1 port map( A => n40, Z => plus2A_out_57_port);
   U35 : BUF_X1 port map( A => n76, Z => plus4A_out_52_port);
   U36 : BUF_X1 port map( A => n75, Z => plus4A_out_53_port);
   U37 : BUF_X2 port map( A => n73, Z => plus2A_out_3_port);
   U38 : BUF_X2 port map( A => n71, Z => plus2A_out_5_port);
   U39 : BUF_X2 port map( A => n69, Z => plus2A_out_7_port);
   U40 : BUF_X2 port map( A => n65, Z => plus2A_out_11_port);
   U41 : BUF_X2 port map( A => n66, Z => plus2A_out_10_port);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity MUX_GENERIC_N64_RADIX3_0 is

   port( plusA, minusA, plus2A, minus2A : in std_logic_vector (63 downto 0);  
         SEL : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (63 
         downto 0));

end MUX_GENERIC_N64_RADIX3_0;

architecture SYN_beh of MUX_GENERIC_N64_RADIX3_0 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X8
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component TBUF_X2
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   component TBUF_X1
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   signal n207, n208, n209, n210, n211, n212, n213, n214, n215, n217, n218, 
      n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, 
      n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, 
      n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, 
      n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, 
      n267, n268, n269, n270, n271, n4, n5, n6, n8, n10, n11, n12, n13, n14, 
      n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29
      , n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, 
      n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58
      , n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, 
      n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87
      , n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
      n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, 
      n114, n115, n116, n117, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n134, net86764, net86762, net86760, 
      net86778, net86774, net86770, net86798, net86796, net86794, net89127, 
      net89124, net89171, net89170, net89204, net94788, n133, net119074, 
      net119196, net119210, net119299, net119289, net119279, net119278, 
      net119275, net119414, net119324, net119316, net119302, net119273, 
      net119270, net119268, net124921, net125048, net125043, net119320, n272, 
      n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, 
      n285 : std_logic;

begin
   
   Y_tri_3_inst : TBUF_X1 port map( A => n210, EN => net119196, Z => Y(3));
   Y_tri_4_inst : TBUF_X1 port map( A => n211, EN => net86762, Z => Y(4));
   Y_tri_5_inst : TBUF_X1 port map( A => n212, EN => net119196, Z => Y(5));
   Y_tri_6_inst : TBUF_X1 port map( A => n213, EN => net119196, Z => Y(6));
   Y_tri_7_inst : TBUF_X1 port map( A => n214, EN => net86762, Z => Y(7));
   Y_tri_8_inst : TBUF_X1 port map( A => n215, EN => net86760, Z => Y(8));
   Y_tri_9_inst : TBUF_X1 port map( A => n217, EN => net86760, Z => Y(9));
   Y_tri_10_inst : TBUF_X1 port map( A => n218, EN => net86764, Z => Y(10));
   Y_tri_11_inst : TBUF_X1 port map( A => n219, EN => net86764, Z => Y(11));
   Y_tri_60_inst : TBUF_X1 port map( A => n268, EN => net86764, Z => Y(60));
   Y_tri_61_inst : TBUF_X1 port map( A => n269, EN => net86764, Z => Y(61));
   Y_tri_62_inst : TBUF_X1 port map( A => n270, EN => net86764, Z => Y(62));
   Y_tri_63_inst : TBUF_X1 port map( A => n271, EN => net86764, Z => Y(63));
   Y_tri_42_inst : TBUF_X1 port map( A => n250, EN => net86764, Z => Y(42));
   Y_tri_43_inst : TBUF_X1 port map( A => n251, EN => net86764, Z => Y(43));
   Y_tri_44_inst : TBUF_X1 port map( A => n252, EN => net86764, Z => Y(44));
   Y_tri_45_inst : TBUF_X1 port map( A => n253, EN => net86764, Z => Y(45));
   Y_tri_46_inst : TBUF_X1 port map( A => n254, EN => net86764, Z => Y(46));
   Y_tri_47_inst : TBUF_X1 port map( A => n255, EN => net86764, Z => Y(47));
   Y_tri_48_inst : TBUF_X1 port map( A => n256, EN => net86764, Z => Y(48));
   Y_tri_49_inst : TBUF_X1 port map( A => n257, EN => net86764, Z => Y(49));
   Y_tri_50_inst : TBUF_X1 port map( A => n258, EN => net86764, Z => Y(50));
   Y_tri_51_inst : TBUF_X1 port map( A => n259, EN => net86764, Z => Y(51));
   Y_tri_52_inst : TBUF_X1 port map( A => n260, EN => net86764, Z => Y(52));
   Y_tri_53_inst : TBUF_X1 port map( A => n261, EN => net86764, Z => Y(53));
   Y_tri_54_inst : TBUF_X1 port map( A => n262, EN => net86764, Z => Y(54));
   Y_tri_55_inst : TBUF_X1 port map( A => n263, EN => net86764, Z => Y(55));
   Y_tri_56_inst : TBUF_X1 port map( A => n264, EN => net86764, Z => Y(56));
   Y_tri_57_inst : TBUF_X1 port map( A => n265, EN => net86764, Z => Y(57));
   Y_tri_58_inst : TBUF_X1 port map( A => n266, EN => net86764, Z => Y(58));
   Y_tri_59_inst : TBUF_X1 port map( A => n267, EN => net86764, Z => Y(59));
   Y_tri_36_inst : TBUF_X1 port map( A => n244, EN => net86764, Z => Y(36));
   Y_tri_31_inst : TBUF_X1 port map( A => n239, EN => net86764, Z => Y(31));
   Y_tri_14_inst : TBUF_X1 port map( A => n222, EN => net86764, Z => Y(14));
   Y_tri_13_inst : TBUF_X1 port map( A => n221, EN => net86764, Z => Y(13));
   Y_tri_15_inst : TBUF_X1 port map( A => n223, EN => net86764, Z => Y(15));
   Y_tri_16_inst : TBUF_X1 port map( A => n224, EN => net86764, Z => Y(16));
   Y_tri_12_inst : TBUF_X1 port map( A => n220, EN => net86764, Z => Y(12));
   Y_tri_17_inst : TBUF_X1 port map( A => n225, EN => net86764, Z => Y(17));
   Y_tri_18_inst : TBUF_X1 port map( A => n226, EN => net86764, Z => Y(18));
   Y_tri_19_inst : TBUF_X1 port map( A => n227, EN => net86764, Z => Y(19));
   Y_tri_20_inst : TBUF_X1 port map( A => n228, EN => net86764, Z => Y(20));
   Y_tri_21_inst : TBUF_X1 port map( A => n229, EN => net86764, Z => Y(21));
   Y_tri_22_inst : TBUF_X1 port map( A => n230, EN => net86764, Z => Y(22));
   Y_tri_23_inst : TBUF_X1 port map( A => n231, EN => net86764, Z => Y(23));
   Y_tri_24_inst : TBUF_X1 port map( A => n232, EN => net86764, Z => Y(24));
   Y_tri_25_inst : TBUF_X1 port map( A => n233, EN => net86764, Z => Y(25));
   Y_tri_26_inst : TBUF_X1 port map( A => n234, EN => net86764, Z => Y(26));
   Y_tri_27_inst : TBUF_X1 port map( A => n235, EN => net86764, Z => Y(27));
   Y_tri_32_inst : TBUF_X1 port map( A => n240, EN => net86764, Z => Y(32));
   Y_tri_28_inst : TBUF_X1 port map( A => n236, EN => net86764, Z => Y(28));
   Y_tri_33_inst : TBUF_X1 port map( A => n241, EN => net86764, Z => Y(33));
   Y_tri_34_inst : TBUF_X1 port map( A => n242, EN => net86764, Z => Y(34));
   Y_tri_29_inst : TBUF_X1 port map( A => n237, EN => net86764, Z => Y(29));
   Y_tri_37_inst : TBUF_X1 port map( A => n245, EN => net86764, Z => Y(37));
   Y_tri_38_inst : TBUF_X1 port map( A => n246, EN => net86764, Z => Y(38));
   Y_tri_39_inst : TBUF_X1 port map( A => n247, EN => net86764, Z => Y(39));
   Y_tri_30_inst : TBUF_X1 port map( A => n238, EN => net86764, Z => Y(30));
   Y_tri_35_inst : TBUF_X1 port map( A => n243, EN => net86764, Z => Y(35));
   Y_tri_40_inst : TBUF_X1 port map( A => n248, EN => net86764, Z => Y(40));
   Y_tri_41_inst : TBUF_X1 port map( A => n249, EN => net86764, Z => Y(41));
   Y_tri_1_inst : TBUF_X1 port map( A => n208, EN => net94788, Z => Y(1));
   Y_tri_2_inst : TBUF_X1 port map( A => n209, EN => net89204, Z => Y(2));
   Y_tri_0_inst : TBUF_X2 port map( A => n207, EN => net119210, Z => Y(0));
   U2 : AND2_X1 port map( A1 => net125043, A2 => net119320, ZN => n8);
   U3 : CLKBUF_X3 port map( A => net89127, Z => net119074);
   U4 : BUF_X4 port map( A => net89124, Z => net89127);
   U5 : BUF_X4 port map( A => net124921, Z => net86798);
   U6 : INV_X2 port map( A => n282, ZN => n6);
   U7 : BUF_X4 port map( A => n6, Z => net86778);
   U8 : AND2_X1 port map( A1 => n277, A2 => net119324, ZN => n272);
   U9 : AND2_X1 port map( A1 => net125048, A2 => net119273, ZN => n273);
   U10 : AND2_X1 port map( A1 => n273, A2 => minusA(1), ZN => n274);
   U11 : NOR2_X1 port map( A1 => n274, A2 => n276, ZN => n134);
   U12 : OAI21_X1 port map( B1 => net119320, B2 => net119299, A => SEL(2), ZN 
                           => n275);
   U13 : INV_X1 port map( A => n275, ZN => net94788);
   U14 : INV_X1 port map( A => n275, ZN => net119210);
   U15 : BUF_X2 port map( A => SEL(1), Z => net119299);
   U16 : BUF_X1 port map( A => SEL(0), Z => net119320);
   U17 : NOR2_X1 port map( A1 => net119299, A2 => net119320, ZN => net119275);
   U18 : BUF_X1 port map( A => SEL(1), Z => net125048);
   U19 : CLKBUF_X1 port map( A => SEL(0), Z => net119302);
   U20 : NOR2_X1 port map( A1 => SEL(0), A2 => SEL(2), ZN => net119273);
   U21 : NOR2_X1 port map( A1 => net125048, A2 => SEL(2), ZN => net125043);
   U22 : CLKBUF_X1 port map( A => n8, Z => net124921);
   U23 : NAND4_X1 port map( A1 => n278, A2 => n279, A3 => n280, A4 => n281, ZN 
                           => n207);
   U24 : NAND2_X1 port map( A1 => n273, A2 => minusA(0), ZN => n281);
   U25 : NAND2_X1 port map( A1 => net86770, A2 => minus2A(0), ZN => n280);
   U26 : INV_X1 port map( A => n282, ZN => net86770);
   U27 : NAND2_X1 port map( A1 => plus2A(0), A2 => n272, ZN => n279);
   U28 : AOI22_X1 port map( A1 => n272, A2 => plus2A(2), B1 => net124921, B2 =>
                           plusA(2), ZN => n131);
   U29 : CLKBUF_X1 port map( A => net119299, Z => net119324);
   U30 : AND2_X1 port map( A1 => n283, A2 => net119324, ZN => net89170);
   U31 : AND2_X4 port map( A1 => n283, A2 => net119324, ZN => net89171);
   U32 : NOR2_X1 port map( A1 => net119316, A2 => net119268, ZN => n277);
   U33 : INV_X1 port map( A => net119302, ZN => net119268);
   U34 : NOR2_X1 port map( A1 => net119316, A2 => net119268, ZN => n283);
   U35 : NAND2_X1 port map( A1 => net119270, A2 => net119302, ZN => net119279);
   U36 : NOR3_X1 port map( A1 => net119278, A2 => net119414, A3 => net119302, 
                           ZN => n276);
   U37 : INV_X1 port map( A => net119270, ZN => net119316);
   U38 : INV_X1 port map( A => SEL(2), ZN => net119270);
   U39 : NAND2_X1 port map( A1 => n8, A2 => plusA(0), ZN => n278);
   U40 : NAND2_X1 port map( A1 => net119273, A2 => net119299, ZN => net119289);
   U41 : NAND2_X1 port map( A1 => net119275, A2 => net119316, ZN => n282);
   U42 : CLKBUF_X1 port map( A => net119299, Z => net119414);
   U43 : BUF_X1 port map( A => net94788, Z => net89204);
   U44 : INV_X2 port map( A => net119289, ZN => net89124);
   U45 : NAND2_X1 port map( A1 => plus2A(1), A2 => net119299, ZN => n285);
   U46 : NAND2_X1 port map( A1 => minus2A(1), A2 => SEL(2), ZN => net119278);
   U47 : AOI21_X1 port map( B1 => n8, B2 => plusA(1), A => n284, ZN => n133);
   U48 : CLKBUF_X3 port map( A => net89204, Z => net119196);
   U49 : NOR2_X1 port map( A1 => net119279, A2 => n285, ZN => n284);
   U50 : BUF_X4 port map( A => n6, Z => net86774);
   U51 : NAND2_X1 port map( A1 => n134, A2 => n133, ZN => n208);
   U52 : BUF_X8 port map( A => net119196, Z => net86764);
   U53 : CLKBUF_X1 port map( A => net119196, Z => net86762);
   U54 : CLKBUF_X1 port map( A => net119196, Z => net86760);
   U55 : BUF_X1 port map( A => n8, Z => net86796);
   U56 : NAND2_X1 port map( A1 => n58, A2 => n59, ZN => n246);
   U57 : AOI22_X1 port map( A1 => plusA(38), A2 => net86798, B1 => plus2A(38), 
                           B2 => net89171, ZN => n58);
   U58 : AOI22_X1 port map( A1 => minus2A(38), A2 => net86778, B1 => minusA(38)
                           , B2 => net119074, ZN => n59);
   U59 : NAND2_X1 port map( A1 => n38, A2 => n39, ZN => n256);
   U60 : AOI22_X1 port map( A1 => plusA(48), A2 => net86798, B1 => plus2A(48), 
                           B2 => net89171, ZN => n38);
   U61 : AOI22_X1 port map( A1 => minus2A(48), A2 => net86778, B1 => minusA(48)
                           , B2 => net119074, ZN => n39);
   U62 : NAND2_X1 port map( A1 => n127, A2 => n128, ZN => n211);
   U63 : NAND2_X1 port map( A1 => n129, A2 => n130, ZN => n210);
   U64 : NAND2_X1 port map( A1 => n116, A2 => n117, ZN => n217);
   U65 : NAND2_X1 port map( A1 => n132, A2 => n131, ZN => n209);
   U66 : NAND2_X1 port map( A1 => n119, A2 => n120, ZN => n215);
   U67 : NAND2_X1 port map( A1 => n121, A2 => n122, ZN => n214);
   U68 : NAND2_X1 port map( A1 => n123, A2 => n124, ZN => n213);
   U69 : NAND2_X1 port map( A1 => n125, A2 => n126, ZN => n212);
   U70 : NAND2_X1 port map( A1 => n12, A2 => n13, ZN => n269);
   U71 : AOI22_X1 port map( A1 => plusA(61), A2 => net86796, B1 => plus2A(61), 
                           B2 => net89171, ZN => n12);
   U72 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => n271);
   U73 : AOI22_X1 port map( A1 => plusA(63), A2 => net86796, B1 => plus2A(63), 
                           B2 => net89171, ZN => n4);
   U74 : AOI22_X1 port map( A1 => minus2A(63), A2 => net86774, B1 => minusA(63)
                           , B2 => net119074, ZN => n5);
   U75 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => n268);
   U76 : AOI22_X1 port map( A1 => plusA(60), A2 => net86798, B1 => plus2A(60), 
                           B2 => net89171, ZN => n14);
   U77 : AOI22_X1 port map( A1 => minus2A(60), A2 => net86774, B1 => minusA(60)
                           , B2 => net89127, ZN => n15);
   U78 : NAND2_X1 port map( A1 => n110, A2 => n111, ZN => n220);
   U79 : AOI22_X1 port map( A1 => plusA(12), A2 => net86798, B1 => plus2A(12), 
                           B2 => net89171, ZN => n110);
   U80 : AOI22_X1 port map( A1 => minus2A(12), A2 => net86778, B1 => minusA(12)
                           , B2 => net89124, ZN => n111);
   U81 : NAND2_X1 port map( A1 => n104, A2 => n105, ZN => n223);
   U82 : AOI22_X1 port map( A1 => plusA(15), A2 => net86798, B1 => plus2A(15), 
                           B2 => net89171, ZN => n104);
   U83 : AOI22_X1 port map( A1 => minus2A(15), A2 => net86774, B1 => minusA(15)
                           , B2 => net119074, ZN => n105);
   U84 : NAND2_X1 port map( A1 => n108, A2 => n109, ZN => n221);
   U85 : AOI22_X1 port map( A1 => plusA(13), A2 => net86798, B1 => plus2A(13), 
                           B2 => net89171, ZN => n108);
   U86 : NAND2_X1 port map( A1 => n106, A2 => n107, ZN => n222);
   U87 : AOI22_X1 port map( A1 => plusA(14), A2 => net86798, B1 => plus2A(14), 
                           B2 => net89171, ZN => n106);
   U88 : AOI22_X1 port map( A1 => minus2A(14), A2 => net86774, B1 => minusA(14)
                           , B2 => net89127, ZN => n107);
   U89 : NAND2_X1 port map( A1 => n74, A2 => n75, ZN => n238);
   U90 : AOI22_X1 port map( A1 => plusA(30), A2 => net86796, B1 => plus2A(30), 
                           B2 => net89171, ZN => n74);
   U91 : NAND2_X1 port map( A1 => n102, A2 => n103, ZN => n224);
   U92 : AOI22_X1 port map( A1 => plusA(16), A2 => net86798, B1 => plus2A(16), 
                           B2 => net89171, ZN => n102);
   U93 : AOI22_X1 port map( A1 => minus2A(16), A2 => net86778, B1 => minusA(16)
                           , B2 => net119074, ZN => n103);
   U94 : NAND2_X1 port map( A1 => n100, A2 => n101, ZN => n225);
   U95 : AOI22_X1 port map( A1 => plusA(17), A2 => net86798, B1 => plus2A(17), 
                           B2 => net89171, ZN => n100);
   U96 : AOI22_X1 port map( A1 => minus2A(17), A2 => net86778, B1 => minusA(17)
                           , B2 => net89127, ZN => n101);
   U97 : NAND2_X1 port map( A1 => n98, A2 => n99, ZN => n226);
   U98 : AOI22_X1 port map( A1 => plusA(18), A2 => net86798, B1 => plus2A(18), 
                           B2 => net89171, ZN => n98);
   U99 : AOI22_X1 port map( A1 => minus2A(18), A2 => net86770, B1 => minusA(18)
                           , B2 => net89124, ZN => n99);
   U100 : NAND2_X1 port map( A1 => n96, A2 => n97, ZN => n227);
   U101 : AOI22_X1 port map( A1 => plusA(19), A2 => net86798, B1 => plus2A(19),
                           B2 => net89171, ZN => n96);
   U102 : NAND2_X1 port map( A1 => n94, A2 => n95, ZN => n228);
   U103 : AOI22_X1 port map( A1 => plusA(20), A2 => net86798, B1 => plus2A(20),
                           B2 => net89171, ZN => n94);
   U104 : AOI22_X1 port map( A1 => minus2A(20), A2 => net86778, B1 => 
                           minusA(20), B2 => net89127, ZN => n95);
   U105 : NAND2_X1 port map( A1 => n64, A2 => n65, ZN => n243);
   U106 : AOI22_X1 port map( A1 => plusA(35), A2 => net86796, B1 => plus2A(35),
                           B2 => net89171, ZN => n64);
   U107 : NAND2_X1 port map( A1 => n92, A2 => n93, ZN => n229);
   U108 : AOI22_X1 port map( A1 => plusA(21), A2 => net86798, B1 => plus2A(21),
                           B2 => net89171, ZN => n92);
   U109 : AOI22_X1 port map( A1 => minus2A(21), A2 => net86778, B1 => 
                           minusA(21), B2 => net119074, ZN => n93);
   U110 : NAND2_X1 port map( A1 => n90, A2 => n91, ZN => n230);
   U111 : AOI22_X1 port map( A1 => plusA(22), A2 => net86798, B1 => plus2A(22),
                           B2 => net89171, ZN => n90);
   U112 : AOI22_X1 port map( A1 => minus2A(22), A2 => net86770, B1 => 
                           minusA(22), B2 => net119074, ZN => n91);
   U113 : NAND2_X1 port map( A1 => n88, A2 => n89, ZN => n231);
   U114 : AOI22_X1 port map( A1 => plusA(23), A2 => net86798, B1 => plus2A(23),
                           B2 => net89171, ZN => n88);
   U115 : AOI22_X1 port map( A1 => minus2A(23), A2 => net86770, B1 => 
                           minusA(23), B2 => net89127, ZN => n89);
   U116 : NAND2_X1 port map( A1 => n86, A2 => n87, ZN => n232);
   U117 : AOI22_X1 port map( A1 => plusA(24), A2 => net86796, B1 => plus2A(24),
                           B2 => net89171, ZN => n86);
   U118 : AOI22_X1 port map( A1 => minus2A(24), A2 => net86778, B1 => 
                           minusA(24), B2 => net89124, ZN => n87);
   U119 : NAND2_X1 port map( A1 => n84, A2 => n85, ZN => n233);
   U120 : AOI22_X1 port map( A1 => plusA(25), A2 => net86796, B1 => plus2A(25),
                           B2 => net89171, ZN => n84);
   U121 : AOI22_X1 port map( A1 => minus2A(25), A2 => net86770, B1 => 
                           minusA(25), B2 => net89127, ZN => n85);
   U122 : NAND2_X1 port map( A1 => n82, A2 => n83, ZN => n234);
   U123 : AOI22_X1 port map( A1 => plusA(26), A2 => net86796, B1 => plus2A(26),
                           B2 => net89171, ZN => n82);
   U124 : AOI22_X1 port map( A1 => minus2A(26), A2 => net86774, B1 => 
                           minusA(26), B2 => net119074, ZN => n83);
   U125 : NAND2_X1 port map( A1 => n80, A2 => n81, ZN => n235);
   U126 : AOI22_X1 port map( A1 => plusA(27), A2 => net86796, B1 => plus2A(27),
                           B2 => net89171, ZN => n80);
   U127 : AOI22_X1 port map( A1 => minus2A(27), A2 => net86778, B1 => 
                           minusA(27), B2 => net119074, ZN => n81);
   U128 : NAND2_X1 port map( A1 => n78, A2 => n79, ZN => n236);
   U129 : AOI22_X1 port map( A1 => plusA(28), A2 => net86796, B1 => plus2A(28),
                           B2 => net89171, ZN => n78);
   U130 : AOI22_X1 port map( A1 => minus2A(28), A2 => net86778, B1 => 
                           minusA(28), B2 => net89127, ZN => n79);
   U131 : NAND2_X1 port map( A1 => n52, A2 => n53, ZN => n249);
   U132 : AOI22_X1 port map( A1 => plusA(41), A2 => net86798, B1 => plus2A(41),
                           B2 => net89171, ZN => n52);
   U133 : AOI22_X1 port map( A1 => minus2A(41), A2 => net86774, B1 => 
                           minusA(41), B2 => net89127, ZN => n53);
   U134 : NAND2_X1 port map( A1 => n54, A2 => n55, ZN => n248);
   U135 : AOI22_X1 port map( A1 => plusA(40), A2 => net86798, B1 => plus2A(40),
                           B2 => net89171, ZN => n54);
   U136 : AOI22_X1 port map( A1 => minus2A(40), A2 => net86774, B1 => 
                           minusA(40), B2 => net119074, ZN => n55);
   U137 : NAND2_X1 port map( A1 => n56, A2 => n57, ZN => n247);
   U138 : AOI22_X1 port map( A1 => plusA(39), A2 => net86798, B1 => plus2A(39),
                           B2 => net89171, ZN => n56);
   U139 : AOI22_X1 port map( A1 => minus2A(39), A2 => net86770, B1 => 
                           minusA(39), B2 => net119074, ZN => n57);
   U140 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => n245);
   U141 : AOI22_X1 port map( A1 => plusA(37), A2 => net86798, B1 => plus2A(37),
                           B2 => net89171, ZN => n60);
   U142 : NAND2_X1 port map( A1 => n76, A2 => n77, ZN => n237);
   U143 : AOI22_X1 port map( A1 => plusA(29), A2 => net86796, B1 => plus2A(29),
                           B2 => net89171, ZN => n76);
   U144 : AOI22_X1 port map( A1 => minus2A(29), A2 => net86770, B1 => 
                           minusA(29), B2 => net119074, ZN => n77);
   U145 : NAND2_X1 port map( A1 => n72, A2 => n73, ZN => n239);
   U146 : AOI22_X1 port map( A1 => plusA(31), A2 => net86796, B1 => plus2A(31),
                           B2 => net89171, ZN => n72);
   U147 : AOI22_X1 port map( A1 => minus2A(31), A2 => net86774, B1 => 
                           minusA(31), B2 => net89127, ZN => n73);
   U148 : NAND2_X1 port map( A1 => n70, A2 => n71, ZN => n240);
   U149 : AOI22_X1 port map( A1 => plusA(32), A2 => net86796, B1 => plus2A(32),
                           B2 => net89171, ZN => n70);
   U150 : AOI22_X1 port map( A1 => minus2A(32), A2 => net86770, B1 => 
                           minusA(32), B2 => net119074, ZN => n71);
   U151 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => n241);
   U152 : AOI22_X1 port map( A1 => plusA(33), A2 => net86796, B1 => plus2A(33),
                           B2 => net89171, ZN => n68);
   U153 : AOI22_X1 port map( A1 => minus2A(33), A2 => net86778, B1 => 
                           minusA(33), B2 => net119074, ZN => n69);
   U154 : NAND2_X1 port map( A1 => n66, A2 => n67, ZN => n242);
   U155 : AOI22_X1 port map( A1 => plusA(34), A2 => net86796, B1 => plus2A(34),
                           B2 => net89171, ZN => n66);
   U156 : AOI22_X1 port map( A1 => minus2A(34), A2 => net86770, B1 => 
                           minusA(34), B2 => net89127, ZN => n67);
   U157 : NAND2_X1 port map( A1 => n62, A2 => n63, ZN => n244);
   U158 : AOI22_X1 port map( A1 => plusA(36), A2 => net86798, B1 => plus2A(36),
                           B2 => net89171, ZN => n62);
   U159 : AOI22_X1 port map( A1 => minus2A(36), A2 => net86774, B1 => 
                           minusA(36), B2 => net89127, ZN => n63);
   U160 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => n267);
   U161 : AOI22_X1 port map( A1 => plusA(59), A2 => net86798, B1 => plus2A(59),
                           B2 => net89171, ZN => n16);
   U162 : AOI22_X1 port map( A1 => minus2A(59), A2 => net86770, B1 => 
                           minusA(59), B2 => net89127, ZN => n17);
   U163 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => n266);
   U164 : AOI22_X1 port map( A1 => plusA(58), A2 => net86798, B1 => plus2A(58),
                           B2 => net89171, ZN => n18);
   U165 : AOI22_X1 port map( A1 => minus2A(58), A2 => net86778, B1 => 
                           minusA(58), B2 => net119074, ZN => n19);
   U166 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => n265);
   U167 : AOI22_X1 port map( A1 => plusA(57), A2 => net86798, B1 => plus2A(57),
                           B2 => net89171, ZN => n20);
   U168 : AOI22_X1 port map( A1 => minus2A(57), A2 => net86778, B1 => 
                           minusA(57), B2 => net119074, ZN => n21);
   U169 : NAND2_X1 port map( A1 => n22, A2 => n23, ZN => n264);
   U170 : AOI22_X1 port map( A1 => plusA(56), A2 => net86798, B1 => plus2A(56),
                           B2 => net89171, ZN => n22);
   U171 : AOI22_X1 port map( A1 => minus2A(56), A2 => net86774, B1 => 
                           minusA(56), B2 => net119074, ZN => n23);
   U172 : NAND2_X1 port map( A1 => n24, A2 => n25, ZN => n263);
   U173 : AOI22_X1 port map( A1 => plusA(55), A2 => net86798, B1 => plus2A(55),
                           B2 => net89171, ZN => n24);
   U174 : NAND2_X1 port map( A1 => n26, A2 => n27, ZN => n262);
   U175 : AOI22_X1 port map( A1 => plusA(54), A2 => net86798, B1 => plus2A(54),
                           B2 => net89171, ZN => n26);
   U176 : AOI22_X1 port map( A1 => minus2A(54), A2 => net86770, B1 => 
                           minusA(54), B2 => net89124, ZN => n27);
   U177 : NAND2_X1 port map( A1 => n28, A2 => n29, ZN => n261);
   U178 : AOI22_X1 port map( A1 => plusA(53), A2 => net86798, B1 => plus2A(53),
                           B2 => net89171, ZN => n28);
   U179 : AOI22_X1 port map( A1 => minus2A(53), A2 => net86778, B1 => 
                           minusA(53), B2 => net89127, ZN => n29);
   U180 : NAND2_X1 port map( A1 => n30, A2 => n31, ZN => n260);
   U181 : AOI22_X1 port map( A1 => plusA(52), A2 => net86798, B1 => plus2A(52),
                           B2 => net89171, ZN => n30);
   U182 : AOI22_X1 port map( A1 => minus2A(52), A2 => net86770, B1 => 
                           minusA(52), B2 => net119074, ZN => n31);
   U183 : NAND2_X1 port map( A1 => n32, A2 => n33, ZN => n259);
   U184 : AOI22_X1 port map( A1 => plusA(51), A2 => net86798, B1 => plus2A(51),
                           B2 => net89171, ZN => n32);
   U185 : AOI22_X1 port map( A1 => minus2A(51), A2 => net86774, B1 => 
                           minusA(51), B2 => net119074, ZN => n33);
   U186 : NAND2_X1 port map( A1 => n34, A2 => n35, ZN => n258);
   U187 : AOI22_X1 port map( A1 => plusA(50), A2 => net86798, B1 => plus2A(50),
                           B2 => net89171, ZN => n34);
   U188 : AOI22_X1 port map( A1 => minus2A(50), A2 => net86770, B1 => 
                           minusA(50), B2 => net89127, ZN => n35);
   U189 : NAND2_X1 port map( A1 => n36, A2 => n37, ZN => n257);
   U190 : AOI22_X1 port map( A1 => plusA(49), A2 => net86798, B1 => plus2A(49),
                           B2 => net89171, ZN => n36);
   U191 : NAND2_X1 port map( A1 => n40, A2 => n41, ZN => n255);
   U192 : AOI22_X1 port map( A1 => plusA(47), A2 => net86798, B1 => plus2A(47),
                           B2 => net89171, ZN => n40);
   U193 : AOI22_X1 port map( A1 => minus2A(47), A2 => net86774, B1 => 
                           minusA(47), B2 => net89127, ZN => n41);
   U194 : NAND2_X1 port map( A1 => n42, A2 => n43, ZN => n254);
   U195 : AOI22_X1 port map( A1 => plusA(46), A2 => net86798, B1 => plus2A(46),
                           B2 => net89171, ZN => n42);
   U196 : AOI22_X1 port map( A1 => minus2A(46), A2 => net86774, B1 => 
                           minusA(46), B2 => net119074, ZN => n43);
   U197 : NAND2_X1 port map( A1 => n44, A2 => n45, ZN => n253);
   U198 : AOI22_X1 port map( A1 => plusA(45), A2 => net86798, B1 => plus2A(45),
                           B2 => net89171, ZN => n44);
   U199 : AOI22_X1 port map( A1 => minus2A(45), A2 => net86770, B1 => 
                           minusA(45), B2 => net119074, ZN => n45);
   U200 : NAND2_X1 port map( A1 => n46, A2 => n47, ZN => n252);
   U201 : AOI22_X1 port map( A1 => plusA(44), A2 => net86798, B1 => plus2A(44),
                           B2 => net89171, ZN => n46);
   U202 : AOI22_X1 port map( A1 => minus2A(44), A2 => net86778, B1 => 
                           minusA(44), B2 => net89127, ZN => n47);
   U203 : NAND2_X1 port map( A1 => n48, A2 => n49, ZN => n251);
   U204 : AOI22_X1 port map( A1 => plusA(43), A2 => net86798, B1 => plus2A(43),
                           B2 => net89171, ZN => n48);
   U205 : NAND2_X1 port map( A1 => n50, A2 => n51, ZN => n250);
   U206 : AOI22_X1 port map( A1 => plusA(42), A2 => net86798, B1 => plus2A(42),
                           B2 => net89171, ZN => n50);
   U207 : AOI22_X1 port map( A1 => minus2A(42), A2 => net86774, B1 => 
                           minusA(42), B2 => net89124, ZN => n51);
   U208 : NAND2_X1 port map( A1 => n10, A2 => n11, ZN => n270);
   U209 : AOI22_X1 port map( A1 => plusA(62), A2 => net86796, B1 => plus2A(62),
                           B2 => net89171, ZN => n10);
   U210 : AOI22_X1 port map( A1 => minus2A(62), A2 => net86778, B1 => 
                           minusA(62), B2 => net89127, ZN => n11);
   U211 : NAND2_X1 port map( A1 => n114, A2 => n115, ZN => n218);
   U212 : NAND2_X1 port map( A1 => n112, A2 => n113, ZN => n219);
   U213 : AOI22_X1 port map( A1 => minus2A(61), A2 => net86770, B1 => 
                           minusA(61), B2 => net119074, ZN => n13);
   U214 : AOI22_X1 port map( A1 => minus2A(55), A2 => net86774, B1 => 
                           minusA(55), B2 => net119074, ZN => n25);
   U215 : AOI22_X1 port map( A1 => minus2A(49), A2 => net86778, B1 => 
                           minusA(49), B2 => net119074, ZN => n37);
   U216 : AOI22_X1 port map( A1 => minus2A(43), A2 => net86770, B1 => 
                           minusA(43), B2 => net119074, ZN => n49);
   U217 : AOI22_X1 port map( A1 => minus2A(37), A2 => net86778, B1 => 
                           minusA(37), B2 => net89124, ZN => n61);
   U218 : AOI22_X1 port map( A1 => minus2A(35), A2 => net86774, B1 => 
                           minusA(35), B2 => net89127, ZN => n65);
   U219 : AOI22_X1 port map( A1 => minus2A(30), A2 => net86774, B1 => 
                           minusA(30), B2 => net89124, ZN => n75);
   U220 : AOI22_X1 port map( A1 => minus2A(19), A2 => net86774, B1 => 
                           minusA(19), B2 => net89124, ZN => n97);
   U221 : AOI22_X1 port map( A1 => minus2A(13), A2 => n6, B1 => minusA(13), B2 
                           => net89127, ZN => n109);
   U222 : CLKBUF_X1 port map( A => net124921, Z => net86794);
   U223 : AOI22_X1 port map( A1 => minus2A(11), A2 => net86778, B1 => 
                           minusA(11), B2 => net89127, ZN => n113);
   U224 : AOI22_X1 port map( A1 => minus2A(10), A2 => net86774, B1 => 
                           minusA(10), B2 => net119074, ZN => n115);
   U225 : AOI22_X1 port map( A1 => minus2A(9), A2 => net86774, B1 => minusA(9),
                           B2 => net119074, ZN => n117);
   U226 : AOI22_X1 port map( A1 => minus2A(8), A2 => n6, B1 => minusA(8), B2 =>
                           net89124, ZN => n120);
   U227 : AOI22_X1 port map( A1 => minus2A(7), A2 => net86778, B1 => minusA(7),
                           B2 => net89124, ZN => n122);
   U228 : AOI22_X1 port map( A1 => minus2A(6), A2 => net86770, B1 => minusA(6),
                           B2 => net89127, ZN => n124);
   U229 : AOI22_X1 port map( A1 => minus2A(5), A2 => net86774, B1 => minusA(5),
                           B2 => net89127, ZN => n126);
   U230 : AOI22_X1 port map( A1 => minus2A(4), A2 => net86774, B1 => minusA(4),
                           B2 => net89127, ZN => n128);
   U231 : AOI22_X1 port map( A1 => minus2A(3), A2 => n6, B1 => minusA(3), B2 =>
                           net89124, ZN => n130);
   U232 : AOI22_X1 port map( A1 => minus2A(2), A2 => n6, B1 => minusA(2), B2 =>
                           net89124, ZN => n132);
   U233 : AOI22_X1 port map( A1 => plusA(11), A2 => net86796, B1 => plus2A(11),
                           B2 => net89171, ZN => n112);
   U234 : AOI22_X1 port map( A1 => plusA(10), A2 => net86796, B1 => plus2A(10),
                           B2 => net89171, ZN => n114);
   U235 : AOI22_X1 port map( A1 => plusA(9), A2 => net86796, B1 => plus2A(9), 
                           B2 => net89171, ZN => n116);
   U236 : AOI22_X1 port map( A1 => plusA(8), A2 => net86796, B1 => plus2A(8), 
                           B2 => net89171, ZN => n119);
   U237 : AOI22_X1 port map( A1 => plusA(7), A2 => net86796, B1 => plus2A(7), 
                           B2 => net89171, ZN => n121);
   U238 : AOI22_X1 port map( A1 => plusA(6), A2 => net86796, B1 => plus2A(6), 
                           B2 => net89171, ZN => n123);
   U239 : AOI22_X1 port map( A1 => plusA(5), A2 => net86796, B1 => plus2A(5), 
                           B2 => net89171, ZN => n125);
   U240 : AOI22_X1 port map( A1 => plusA(4), A2 => net86796, B1 => plus2A(4), 
                           B2 => net89170, ZN => n127);
   U241 : AOI22_X1 port map( A1 => plusA(3), A2 => net86794, B1 => plus2A(3), 
                           B2 => net89170, ZN => n129);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity ShiftnCompl_special_N64 is

   port( plusA : in std_logic_vector (63 downto 0);  plusA_out, minusA_out, 
         plus2A_out, minus2A_out : out std_logic_vector (63 downto 0));

end ShiftnCompl_special_N64;

architecture SYN_struct of ShiftnCompl_special_N64 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component complementer_N64_31
      port( input : in std_logic_vector (63 downto 0);  complement2 : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component complementer_N64_0
      port( input : in std_logic_vector (63 downto 0);  complement2 : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component shifter_N64_0
      port( input : in std_logic_vector (63 downto 0);  shiftLeftOnePos : out 
            std_logic_vector (63 downto 0));
   end component;
   
   signal plus2A_out_63_port, plus2A_out_62_port, plus2A_out_61_port, 
      plus2A_out_60_port, plus2A_out_59_port, plus2A_out_58_port, 
      plus2A_out_57_port, plus2A_out_56_port, plus2A_out_55_port, 
      plus2A_out_54_port, n13, n14, plus2A_out_51_port, plus2A_out_50_port, 
      plus2A_out_49_port, plus2A_out_48_port, plus2A_out_47_port, 
      plus2A_out_46_port, plus2A_out_45_port, plus2A_out_44_port, n15, n16, 
      plus2A_out_41_port, plus2A_out_40_port, plus2A_out_39_port, 
      plus2A_out_38_port, plus2A_out_37_port, plus2A_out_36_port, 
      plus2A_out_35_port, plus2A_out_34_port, n17, n18, n19, plus2A_out_30_port
      , plus2A_out_29_port, plus2A_out_28_port, plus2A_out_27_port, 
      plus2A_out_26_port, plus2A_out_25_port, plus2A_out_24_port, 
      plus2A_out_23_port, plus2A_out_22_port, plus2A_out_21_port, 
      plus2A_out_20_port, plus2A_out_19_port, plus2A_out_18_port, 
      plus2A_out_17_port, plus2A_out_16_port, plus2A_out_15_port, 
      plus2A_out_14_port, plus2A_out_13_port, plus2A_out_12_port, 
      plus2A_out_11_port, plus2A_out_10_port, plus2A_out_9_port, 
      plus2A_out_8_port, plus2A_out_7_port, plus2A_out_6_port, 
      plus2A_out_5_port, plus2A_out_4_port, plus2A_out_3_port, 
      plus2A_out_2_port, plus2A_out_1_port, plus2A_out_0_port, 
      plus2A_out_31_port, plus2A_out_32_port, plus2A_out_33_port, 
      plusA_out_37_port, plusA_out_38_port, plus2A_out_42_port, 
      plus2A_out_43_port, plusA_out_47_port, plusA_out_48_port, 
      plus2A_out_52_port, plus2A_out_53_port, plusA_out_57_port, n_3174 : 
      std_logic;

begin
   plusA_out <= ( plusA(63), plusA(62), plusA(61), plusA(60), plusA(59), 
      plusA(58), plusA_out_57_port, plusA(56), plusA(55), plusA(54), plusA(53),
      plusA(52), plusA(51), plusA(50), plusA(49), plusA_out_48_port, 
      plusA_out_47_port, plusA(46), plusA(45), plusA(44), plusA(43), plusA(42),
      plusA(41), plusA(40), plusA(39), plusA_out_38_port, plusA_out_37_port, 
      plusA(36), plusA(35), plusA(34), plusA(33), plusA(32), plusA(31), 
      plusA(30), plusA(29), plusA(28), plusA(27), plusA(26), plusA(25), 
      plusA(24), plusA(23), plusA(22), plusA(21), plusA(20), plusA(19), 
      plusA(18), plusA(17), plusA(16), plusA(15), plusA(14), plusA(13), 
      plusA(12), plusA(11), plusA(10), plusA(9), plusA(8), plusA(7), plusA(6), 
      plusA(5), plusA(4), plusA(3), plusA(2), plusA(1), plusA(0) );
   plus2A_out <= ( plus2A_out_63_port, plus2A_out_62_port, plus2A_out_61_port, 
      plus2A_out_60_port, plus2A_out_59_port, plus2A_out_58_port, 
      plus2A_out_57_port, plus2A_out_56_port, plus2A_out_55_port, 
      plus2A_out_54_port, plus2A_out_53_port, plus2A_out_52_port, 
      plus2A_out_51_port, plus2A_out_50_port, plus2A_out_49_port, 
      plus2A_out_48_port, plus2A_out_47_port, plus2A_out_46_port, 
      plus2A_out_45_port, plus2A_out_44_port, plus2A_out_43_port, 
      plus2A_out_42_port, plus2A_out_41_port, plus2A_out_40_port, 
      plus2A_out_39_port, plus2A_out_38_port, plus2A_out_37_port, 
      plus2A_out_36_port, plus2A_out_35_port, plus2A_out_34_port, 
      plus2A_out_33_port, plus2A_out_32_port, plus2A_out_31_port, 
      plus2A_out_30_port, plus2A_out_29_port, plus2A_out_28_port, 
      plus2A_out_27_port, plus2A_out_26_port, plus2A_out_25_port, 
      plus2A_out_24_port, plus2A_out_23_port, plus2A_out_22_port, 
      plus2A_out_21_port, plus2A_out_20_port, plus2A_out_19_port, 
      plus2A_out_18_port, plus2A_out_17_port, plus2A_out_16_port, 
      plus2A_out_15_port, plus2A_out_14_port, plus2A_out_13_port, 
      plus2A_out_12_port, plus2A_out_11_port, plus2A_out_10_port, 
      plus2A_out_9_port, plus2A_out_8_port, plus2A_out_7_port, 
      plus2A_out_6_port, plus2A_out_5_port, plus2A_out_4_port, 
      plus2A_out_3_port, plus2A_out_2_port, plus2A_out_1_port, 
      plus2A_out_0_port );
   
   plus2A_out_0_port <= '0';
   shifter_1 : shifter_N64_0 port map( input(63) => plusA(63), input(62) => 
                           plusA(62), input(61) => plusA(61), input(60) => 
                           plusA(60), input(59) => plusA(59), input(58) => 
                           plusA(58), input(57) => plusA_out_57_port, input(56)
                           => plusA(56), input(55) => plusA(55), input(54) => 
                           plusA(54), input(53) => plusA(53), input(52) => 
                           plusA(52), input(51) => plusA(51), input(50) => 
                           plusA(50), input(49) => plusA(49), input(48) => 
                           plusA_out_48_port, input(47) => plusA_out_47_port, 
                           input(46) => plusA(46), input(45) => plusA(45), 
                           input(44) => plusA(44), input(43) => plusA(43), 
                           input(42) => plusA(42), input(41) => plusA(41), 
                           input(40) => plusA(40), input(39) => plusA(39), 
                           input(38) => plusA_out_38_port, input(37) => 
                           plusA_out_37_port, input(36) => plusA(36), input(35)
                           => plusA(35), input(34) => plusA(34), input(33) => 
                           plusA(33), input(32) => plusA(32), input(31) => 
                           plusA(31), input(30) => plusA(30), input(29) => 
                           plusA(29), input(28) => plusA(28), input(27) => 
                           plusA(27), input(26) => plusA(26), input(25) => 
                           plusA(25), input(24) => plusA(24), input(23) => 
                           plusA(23), input(22) => plusA(22), input(21) => 
                           plusA(21), input(20) => plusA(20), input(19) => 
                           plusA(19), input(18) => plusA(18), input(17) => 
                           plusA(17), input(16) => plusA(16), input(15) => 
                           plusA(15), input(14) => plusA(14), input(13) => 
                           plusA(13), input(12) => plusA(12), input(11) => 
                           plusA(11), input(10) => plusA(10), input(9) => 
                           plusA(9), input(8) => plusA(8), input(7) => plusA(7)
                           , input(6) => plusA(6), input(5) => plusA(5), 
                           input(4) => plusA(4), input(3) => plusA(3), input(2)
                           => plusA(2), input(1) => plusA(1), input(0) => 
                           plusA(0), shiftLeftOnePos(63) => plus2A_out_63_port,
                           shiftLeftOnePos(62) => plus2A_out_62_port, 
                           shiftLeftOnePos(61) => plus2A_out_61_port, 
                           shiftLeftOnePos(60) => plus2A_out_60_port, 
                           shiftLeftOnePos(59) => plus2A_out_59_port, 
                           shiftLeftOnePos(58) => plus2A_out_58_port, 
                           shiftLeftOnePos(57) => plus2A_out_57_port, 
                           shiftLeftOnePos(56) => plus2A_out_56_port, 
                           shiftLeftOnePos(55) => plus2A_out_55_port, 
                           shiftLeftOnePos(54) => plus2A_out_54_port, 
                           shiftLeftOnePos(53) => n13, shiftLeftOnePos(52) => 
                           n14, shiftLeftOnePos(51) => plus2A_out_51_port, 
                           shiftLeftOnePos(50) => plus2A_out_50_port, 
                           shiftLeftOnePos(49) => plus2A_out_49_port, 
                           shiftLeftOnePos(48) => plus2A_out_48_port, 
                           shiftLeftOnePos(47) => plus2A_out_47_port, 
                           shiftLeftOnePos(46) => plus2A_out_46_port, 
                           shiftLeftOnePos(45) => plus2A_out_45_port, 
                           shiftLeftOnePos(44) => plus2A_out_44_port, 
                           shiftLeftOnePos(43) => n15, shiftLeftOnePos(42) => 
                           n16, shiftLeftOnePos(41) => plus2A_out_41_port, 
                           shiftLeftOnePos(40) => plus2A_out_40_port, 
                           shiftLeftOnePos(39) => plus2A_out_39_port, 
                           shiftLeftOnePos(38) => plus2A_out_38_port, 
                           shiftLeftOnePos(37) => plus2A_out_37_port, 
                           shiftLeftOnePos(36) => plus2A_out_36_port, 
                           shiftLeftOnePos(35) => plus2A_out_35_port, 
                           shiftLeftOnePos(34) => plus2A_out_34_port, 
                           shiftLeftOnePos(33) => n17, shiftLeftOnePos(32) => 
                           n18, shiftLeftOnePos(31) => n19, shiftLeftOnePos(30)
                           => plus2A_out_30_port, shiftLeftOnePos(29) => 
                           plus2A_out_29_port, shiftLeftOnePos(28) => 
                           plus2A_out_28_port, shiftLeftOnePos(27) => 
                           plus2A_out_27_port, shiftLeftOnePos(26) => 
                           plus2A_out_26_port, shiftLeftOnePos(25) => 
                           plus2A_out_25_port, shiftLeftOnePos(24) => 
                           plus2A_out_24_port, shiftLeftOnePos(23) => 
                           plus2A_out_23_port, shiftLeftOnePos(22) => 
                           plus2A_out_22_port, shiftLeftOnePos(21) => 
                           plus2A_out_21_port, shiftLeftOnePos(20) => 
                           plus2A_out_20_port, shiftLeftOnePos(19) => 
                           plus2A_out_19_port, shiftLeftOnePos(18) => 
                           plus2A_out_18_port, shiftLeftOnePos(17) => 
                           plus2A_out_17_port, shiftLeftOnePos(16) => 
                           plus2A_out_16_port, shiftLeftOnePos(15) => 
                           plus2A_out_15_port, shiftLeftOnePos(14) => 
                           plus2A_out_14_port, shiftLeftOnePos(13) => 
                           plus2A_out_13_port, shiftLeftOnePos(12) => 
                           plus2A_out_12_port, shiftLeftOnePos(11) => 
                           plus2A_out_11_port, shiftLeftOnePos(10) => 
                           plus2A_out_10_port, shiftLeftOnePos(9) => 
                           plus2A_out_9_port, shiftLeftOnePos(8) => 
                           plus2A_out_8_port, shiftLeftOnePos(7) => 
                           plus2A_out_7_port, shiftLeftOnePos(6) => 
                           plus2A_out_6_port, shiftLeftOnePos(5) => 
                           plus2A_out_5_port, shiftLeftOnePos(4) => 
                           plus2A_out_4_port, shiftLeftOnePos(3) => 
                           plus2A_out_3_port, shiftLeftOnePos(2) => 
                           plus2A_out_2_port, shiftLeftOnePos(1) => 
                           plus2A_out_1_port, shiftLeftOnePos(0) => n_3174);
   complementer_1 : complementer_N64_0 port map( input(63) => plusA(63), 
                           input(62) => plusA(62), input(61) => plusA(61), 
                           input(60) => plusA(60), input(59) => plusA(59), 
                           input(58) => plusA(58), input(57) => 
                           plusA_out_57_port, input(56) => plusA(56), input(55)
                           => plusA(55), input(54) => plusA(54), input(53) => 
                           plusA(53), input(52) => plusA(52), input(51) => 
                           plusA(51), input(50) => plusA(50), input(49) => 
                           plusA(49), input(48) => plusA_out_48_port, input(47)
                           => plusA_out_47_port, input(46) => plusA(46), 
                           input(45) => plusA(45), input(44) => plusA(44), 
                           input(43) => plusA(43), input(42) => plusA(42), 
                           input(41) => plusA(41), input(40) => plusA(40), 
                           input(39) => plusA(39), input(38) => 
                           plusA_out_38_port, input(37) => plusA_out_37_port, 
                           input(36) => plusA(36), input(35) => plusA(35), 
                           input(34) => plusA(34), input(33) => plusA(33), 
                           input(32) => plusA(32), input(31) => plusA(31), 
                           input(30) => plusA(30), input(29) => plusA(29), 
                           input(28) => plusA(28), input(27) => plusA(27), 
                           input(26) => plusA(26), input(25) => plusA(25), 
                           input(24) => plusA(24), input(23) => plusA(23), 
                           input(22) => plusA(22), input(21) => plusA(21), 
                           input(20) => plusA(20), input(19) => plusA(19), 
                           input(18) => plusA(18), input(17) => plusA(17), 
                           input(16) => plusA(16), input(15) => plusA(15), 
                           input(14) => plusA(14), input(13) => plusA(13), 
                           input(12) => plusA(12), input(11) => plusA(11), 
                           input(10) => plusA(10), input(9) => plusA(9), 
                           input(8) => plusA(8), input(7) => plusA(7), input(6)
                           => plusA(6), input(5) => plusA(5), input(4) => 
                           plusA(4), input(3) => plusA(3), input(2) => plusA(2)
                           , input(1) => plusA(1), input(0) => plusA(0), 
                           complement2(63) => minusA_out(63), complement2(62) 
                           => minusA_out(62), complement2(61) => minusA_out(61)
                           , complement2(60) => minusA_out(60), complement2(59)
                           => minusA_out(59), complement2(58) => minusA_out(58)
                           , complement2(57) => minusA_out(57), complement2(56)
                           => minusA_out(56), complement2(55) => minusA_out(55)
                           , complement2(54) => minusA_out(54), complement2(53)
                           => minusA_out(53), complement2(52) => minusA_out(52)
                           , complement2(51) => minusA_out(51), complement2(50)
                           => minusA_out(50), complement2(49) => minusA_out(49)
                           , complement2(48) => minusA_out(48), complement2(47)
                           => minusA_out(47), complement2(46) => minusA_out(46)
                           , complement2(45) => minusA_out(45), complement2(44)
                           => minusA_out(44), complement2(43) => minusA_out(43)
                           , complement2(42) => minusA_out(42), complement2(41)
                           => minusA_out(41), complement2(40) => minusA_out(40)
                           , complement2(39) => minusA_out(39), complement2(38)
                           => minusA_out(38), complement2(37) => minusA_out(37)
                           , complement2(36) => minusA_out(36), complement2(35)
                           => minusA_out(35), complement2(34) => minusA_out(34)
                           , complement2(33) => minusA_out(33), complement2(32)
                           => minusA_out(32), complement2(31) => minusA_out(31)
                           , complement2(30) => minusA_out(30), complement2(29)
                           => minusA_out(29), complement2(28) => minusA_out(28)
                           , complement2(27) => minusA_out(27), complement2(26)
                           => minusA_out(26), complement2(25) => minusA_out(25)
                           , complement2(24) => minusA_out(24), complement2(23)
                           => minusA_out(23), complement2(22) => minusA_out(22)
                           , complement2(21) => minusA_out(21), complement2(20)
                           => minusA_out(20), complement2(19) => minusA_out(19)
                           , complement2(18) => minusA_out(18), complement2(17)
                           => minusA_out(17), complement2(16) => minusA_out(16)
                           , complement2(15) => minusA_out(15), complement2(14)
                           => minusA_out(14), complement2(13) => minusA_out(13)
                           , complement2(12) => minusA_out(12), complement2(11)
                           => minusA_out(11), complement2(10) => minusA_out(10)
                           , complement2(9) => minusA_out(9), complement2(8) =>
                           minusA_out(8), complement2(7) => minusA_out(7), 
                           complement2(6) => minusA_out(6), complement2(5) => 
                           minusA_out(5), complement2(4) => minusA_out(4), 
                           complement2(3) => minusA_out(3), complement2(2) => 
                           minusA_out(2), complement2(1) => minusA_out(1), 
                           complement2(0) => minusA_out(0));
   complementer_2 : complementer_N64_31 port map( input(63) => 
                           plus2A_out_63_port, input(62) => plus2A_out_62_port,
                           input(61) => plus2A_out_61_port, input(60) => 
                           plus2A_out_60_port, input(59) => plus2A_out_59_port,
                           input(58) => plus2A_out_58_port, input(57) => 
                           plus2A_out_57_port, input(56) => plus2A_out_56_port,
                           input(55) => plus2A_out_55_port, input(54) => 
                           plus2A_out_54_port, input(53) => plus2A_out_53_port,
                           input(52) => plus2A_out_52_port, input(51) => 
                           plus2A_out_51_port, input(50) => plus2A_out_50_port,
                           input(49) => plus2A_out_49_port, input(48) => 
                           plus2A_out_48_port, input(47) => plus2A_out_47_port,
                           input(46) => plus2A_out_46_port, input(45) => 
                           plus2A_out_45_port, input(44) => plus2A_out_44_port,
                           input(43) => plus2A_out_43_port, input(42) => 
                           plus2A_out_42_port, input(41) => plus2A_out_41_port,
                           input(40) => plus2A_out_40_port, input(39) => 
                           plus2A_out_39_port, input(38) => plus2A_out_38_port,
                           input(37) => plus2A_out_37_port, input(36) => 
                           plus2A_out_36_port, input(35) => plus2A_out_35_port,
                           input(34) => plus2A_out_34_port, input(33) => 
                           plus2A_out_33_port, input(32) => plus2A_out_32_port,
                           input(31) => plus2A_out_31_port, input(30) => 
                           plus2A_out_30_port, input(29) => plus2A_out_29_port,
                           input(28) => plus2A_out_28_port, input(27) => 
                           plus2A_out_27_port, input(26) => plus2A_out_26_port,
                           input(25) => plus2A_out_25_port, input(24) => 
                           plus2A_out_24_port, input(23) => plus2A_out_23_port,
                           input(22) => plus2A_out_22_port, input(21) => 
                           plus2A_out_21_port, input(20) => plus2A_out_20_port,
                           input(19) => plus2A_out_19_port, input(18) => 
                           plus2A_out_18_port, input(17) => plus2A_out_17_port,
                           input(16) => plus2A_out_16_port, input(15) => 
                           plus2A_out_15_port, input(14) => plus2A_out_14_port,
                           input(13) => plus2A_out_13_port, input(12) => 
                           plus2A_out_12_port, input(11) => plus2A_out_11_port,
                           input(10) => plus2A_out_10_port, input(9) => 
                           plus2A_out_9_port, input(8) => plus2A_out_8_port, 
                           input(7) => plus2A_out_7_port, input(6) => 
                           plus2A_out_6_port, input(5) => plus2A_out_5_port, 
                           input(4) => plus2A_out_4_port, input(3) => 
                           plus2A_out_3_port, input(2) => plus2A_out_2_port, 
                           input(1) => plus2A_out_1_port, input(0) => 
                           plus2A_out_0_port, complement2(63) => 
                           minus2A_out(63), complement2(62) => minus2A_out(62),
                           complement2(61) => minus2A_out(61), complement2(60) 
                           => minus2A_out(60), complement2(59) => 
                           minus2A_out(59), complement2(58) => minus2A_out(58),
                           complement2(57) => minus2A_out(57), complement2(56) 
                           => minus2A_out(56), complement2(55) => 
                           minus2A_out(55), complement2(54) => minus2A_out(54),
                           complement2(53) => minus2A_out(53), complement2(52) 
                           => minus2A_out(52), complement2(51) => 
                           minus2A_out(51), complement2(50) => minus2A_out(50),
                           complement2(49) => minus2A_out(49), complement2(48) 
                           => minus2A_out(48), complement2(47) => 
                           minus2A_out(47), complement2(46) => minus2A_out(46),
                           complement2(45) => minus2A_out(45), complement2(44) 
                           => minus2A_out(44), complement2(43) => 
                           minus2A_out(43), complement2(42) => minus2A_out(42),
                           complement2(41) => minus2A_out(41), complement2(40) 
                           => minus2A_out(40), complement2(39) => 
                           minus2A_out(39), complement2(38) => minus2A_out(38),
                           complement2(37) => minus2A_out(37), complement2(36) 
                           => minus2A_out(36), complement2(35) => 
                           minus2A_out(35), complement2(34) => minus2A_out(34),
                           complement2(33) => minus2A_out(33), complement2(32) 
                           => minus2A_out(32), complement2(31) => 
                           minus2A_out(31), complement2(30) => minus2A_out(30),
                           complement2(29) => minus2A_out(29), complement2(28) 
                           => minus2A_out(28), complement2(27) => 
                           minus2A_out(27), complement2(26) => minus2A_out(26),
                           complement2(25) => minus2A_out(25), complement2(24) 
                           => minus2A_out(24), complement2(23) => 
                           minus2A_out(23), complement2(22) => minus2A_out(22),
                           complement2(21) => minus2A_out(21), complement2(20) 
                           => minus2A_out(20), complement2(19) => 
                           minus2A_out(19), complement2(18) => minus2A_out(18),
                           complement2(17) => minus2A_out(17), complement2(16) 
                           => minus2A_out(16), complement2(15) => 
                           minus2A_out(15), complement2(14) => minus2A_out(14),
                           complement2(13) => minus2A_out(13), complement2(12) 
                           => minus2A_out(12), complement2(11) => 
                           minus2A_out(11), complement2(10) => minus2A_out(10),
                           complement2(9) => minus2A_out(9), complement2(8) => 
                           minus2A_out(8), complement2(7) => minus2A_out(7), 
                           complement2(6) => minus2A_out(6), complement2(5) => 
                           minus2A_out(5), complement2(4) => minus2A_out(4), 
                           complement2(3) => minus2A_out(3), complement2(2) => 
                           minus2A_out(2), complement2(1) => minus2A_out(1), 
                           complement2(0) => minus2A_out(0));
   U2 : BUF_X1 port map( A => plusA(37), Z => plusA_out_37_port);
   U3 : BUF_X1 port map( A => n19, Z => plus2A_out_31_port);
   U4 : BUF_X1 port map( A => n18, Z => plus2A_out_32_port);
   U5 : BUF_X1 port map( A => plusA(38), Z => plusA_out_38_port);
   U6 : BUF_X1 port map( A => plusA(47), Z => plusA_out_47_port);
   U7 : BUF_X1 port map( A => n15, Z => plus2A_out_43_port);
   U8 : BUF_X1 port map( A => n16, Z => plus2A_out_42_port);
   U9 : BUF_X1 port map( A => plusA(48), Z => plusA_out_48_port);
   U10 : BUF_X1 port map( A => plusA(57), Z => plusA_out_57_port);
   U11 : BUF_X1 port map( A => n14, Z => plus2A_out_52_port);
   U12 : BUF_X1 port map( A => n13, Z => plus2A_out_53_port);
   U13 : BUF_X1 port map( A => n17, Z => plus2A_out_33_port);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity encoder_N64_RADIX3_0 is

   port( X : in std_logic_vector (2 downto 0);  Z : out std_logic_vector (2 
         downto 0));

end encoder_N64_RADIX3_0;

architecture SYN_beh of encoder_N64_RADIX3_0 is

   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, net92849, net85021, n3, n5 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => X(1), A2 => X(0), ZN => n3);
   U2 : OAI21_X1 port map( B1 => X(1), B2 => X(0), A => n3, ZN => n5);
   U3 : AOI21_X1 port map( B1 => n5, B2 => n3, A => X(2), ZN => Z(0));
   U4 : OAI22_X1 port map( A1 => n5, A2 => net85021, B1 => X(2), B2 => n3, ZN 
                           => Z(1));
   U5 : OAI21_X1 port map( B1 => X(1), B2 => X(0), A => n3, ZN => n2);
   U6 : INV_X1 port map( A => X(2), ZN => net85021);
   U7 : AND2_X1 port map( A1 => n3, A2 => X(2), ZN => net92849);
   U8 : AND2_X2 port map( A1 => n2, A2 => net92849, ZN => Z(2));

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity booth_mul_row_N64_RADIX3_1 is

   port( prevA, prevSum : in std_logic_vector (63 downto 0);  encoderIn : in 
         std_logic_vector (2 downto 0);  nextA, nextSum : out std_logic_vector 
         (63 downto 0));

end booth_mul_row_N64_RADIX3_1;

architecture SYN_struct of booth_mul_row_N64_RADIX3_1 is

   component RCA_N64_1
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component MUX_GENERIC_N64_RADIX3_1
      port( plusA, minusA, plus2A, minus2A : in std_logic_vector (63 downto 0);
            SEL : in std_logic_vector (2 downto 0);  Y : out std_logic_vector 
            (63 downto 0));
   end component;
   
   component ShiftnCompl_N64_1
      port( plusA : in std_logic_vector (63 downto 0);  plus2A_out, minus2A_out
            , plus4A_out, minus4A_out : out std_logic_vector (63 downto 0));
   end component;
   
   component encoder_N64_RADIX3_1
      port( X : in std_logic_vector (2 downto 0);  Z : out std_logic_vector (2 
            downto 0));
   end component;
   
   signal X_Logic0_port, nextA_63_port, nextA_62_port, nextA_61_port, 
      nextA_60_port, nextA_59_port, nextA_58_port, nextA_57_port, nextA_56_port
      , nextA_55_port, nextA_54_port, nextA_53_port, nextA_52_port, 
      nextA_51_port, nextA_50_port, nextA_49_port, nextA_48_port, nextA_47_port
      , nextA_46_port, nextA_45_port, nextA_44_port, nextA_43_port, 
      nextA_42_port, nextA_41_port, nextA_40_port, nextA_39_port, nextA_38_port
      , nextA_37_port, nextA_36_port, nextA_35_port, nextA_34_port, 
      nextA_33_port, nextA_32_port, nextA_31_port, nextA_30_port, nextA_29_port
      , nextA_28_port, nextA_27_port, nextA_26_port, nextA_25_port, 
      nextA_24_port, nextA_23_port, nextA_22_port, nextA_21_port, nextA_20_port
      , nextA_19_port, nextA_18_port, nextA_17_port, nextA_16_port, 
      nextA_15_port, nextA_14_port, nextA_13_port, nextA_12_port, nextA_11_port
      , nextA_10_port, nextA_9_port, nextA_8_port, nextA_7_port, nextA_6_port, 
      nextA_5_port, nextA_4_port, nextA_3_port, nextA_2_port, nextA_1_port, 
      encoder_to_mux_2_port, encoder_to_mux_1_port, encoder_to_mux_0_port, 
      plus2A_s_63_port, plus2A_s_62_port, plus2A_s_61_port, plus2A_s_60_port, 
      plus2A_s_59_port, plus2A_s_58_port, plus2A_s_57_port, plus2A_s_56_port, 
      plus2A_s_55_port, plus2A_s_54_port, plus2A_s_53_port, plus2A_s_52_port, 
      plus2A_s_51_port, plus2A_s_50_port, plus2A_s_49_port, plus2A_s_48_port, 
      plus2A_s_47_port, plus2A_s_46_port, plus2A_s_45_port, plus2A_s_44_port, 
      plus2A_s_43_port, plus2A_s_42_port, plus2A_s_41_port, plus2A_s_40_port, 
      plus2A_s_39_port, plus2A_s_38_port, plus2A_s_37_port, plus2A_s_36_port, 
      plus2A_s_35_port, plus2A_s_34_port, plus2A_s_33_port, plus2A_s_32_port, 
      plus2A_s_31_port, plus2A_s_30_port, plus2A_s_29_port, plus2A_s_28_port, 
      plus2A_s_27_port, plus2A_s_26_port, plus2A_s_25_port, plus2A_s_24_port, 
      plus2A_s_23_port, plus2A_s_22_port, plus2A_s_21_port, plus2A_s_20_port, 
      plus2A_s_19_port, plus2A_s_18_port, plus2A_s_17_port, plus2A_s_16_port, 
      plus2A_s_15_port, plus2A_s_14_port, plus2A_s_13_port, plus2A_s_12_port, 
      plus2A_s_11_port, plus2A_s_10_port, plus2A_s_9_port, plus2A_s_8_port, 
      plus2A_s_7_port, plus2A_s_6_port, plus2A_s_5_port, plus2A_s_4_port, 
      plus2A_s_3_port, plus2A_s_2_port, plus2A_s_1_port, minus2A_s_63_port, 
      minus2A_s_62_port, minus2A_s_61_port, minus2A_s_60_port, 
      minus2A_s_59_port, minus2A_s_58_port, minus2A_s_57_port, 
      minus2A_s_56_port, minus2A_s_55_port, minus2A_s_54_port, 
      minus2A_s_53_port, minus2A_s_52_port, minus2A_s_51_port, 
      minus2A_s_50_port, minus2A_s_49_port, minus2A_s_48_port, 
      minus2A_s_47_port, minus2A_s_46_port, minus2A_s_45_port, 
      minus2A_s_44_port, minus2A_s_43_port, minus2A_s_42_port, 
      minus2A_s_41_port, minus2A_s_40_port, minus2A_s_39_port, 
      minus2A_s_38_port, minus2A_s_37_port, minus2A_s_36_port, 
      minus2A_s_35_port, minus2A_s_34_port, minus2A_s_33_port, 
      minus2A_s_32_port, minus2A_s_31_port, minus2A_s_30_port, 
      minus2A_s_29_port, minus2A_s_28_port, minus2A_s_27_port, 
      minus2A_s_26_port, minus2A_s_25_port, minus2A_s_24_port, 
      minus2A_s_23_port, minus2A_s_22_port, minus2A_s_21_port, 
      minus2A_s_20_port, minus2A_s_19_port, minus2A_s_18_port, 
      minus2A_s_17_port, minus2A_s_16_port, minus2A_s_15_port, 
      minus2A_s_14_port, minus2A_s_13_port, minus2A_s_12_port, 
      minus2A_s_11_port, minus2A_s_10_port, minus2A_s_9_port, minus2A_s_8_port,
      minus2A_s_7_port, minus2A_s_6_port, minus2A_s_5_port, minus2A_s_4_port, 
      minus2A_s_3_port, minus2A_s_2_port, minus2A_s_1_port, minus2A_s_0_port, 
      minus4A_s_63_port, minus4A_s_62_port, minus4A_s_61_port, 
      minus4A_s_60_port, minus4A_s_59_port, minus4A_s_58_port, 
      minus4A_s_57_port, minus4A_s_56_port, minus4A_s_55_port, 
      minus4A_s_54_port, minus4A_s_53_port, minus4A_s_52_port, 
      minus4A_s_51_port, minus4A_s_50_port, minus4A_s_49_port, 
      minus4A_s_48_port, minus4A_s_47_port, minus4A_s_46_port, 
      minus4A_s_45_port, minus4A_s_44_port, minus4A_s_43_port, 
      minus4A_s_42_port, minus4A_s_41_port, minus4A_s_40_port, 
      minus4A_s_39_port, minus4A_s_38_port, minus4A_s_37_port, 
      minus4A_s_36_port, minus4A_s_35_port, minus4A_s_34_port, 
      minus4A_s_33_port, minus4A_s_32_port, minus4A_s_31_port, 
      minus4A_s_30_port, minus4A_s_29_port, minus4A_s_28_port, 
      minus4A_s_27_port, minus4A_s_26_port, minus4A_s_25_port, 
      minus4A_s_24_port, minus4A_s_23_port, minus4A_s_22_port, 
      minus4A_s_21_port, minus4A_s_20_port, minus4A_s_19_port, 
      minus4A_s_18_port, minus4A_s_17_port, minus4A_s_16_port, 
      minus4A_s_15_port, minus4A_s_14_port, minus4A_s_13_port, 
      minus4A_s_12_port, minus4A_s_11_port, minus4A_s_10_port, minus4A_s_9_port
      , minus4A_s_8_port, minus4A_s_7_port, minus4A_s_6_port, minus4A_s_5_port,
      minus4A_s_4_port, minus4A_s_3_port, minus4A_s_2_port, minus4A_s_1_port, 
      minus4A_s_0_port, mux_to_adder_63_port, mux_to_adder_62_port, 
      mux_to_adder_61_port, mux_to_adder_60_port, mux_to_adder_59_port, 
      mux_to_adder_58_port, mux_to_adder_57_port, mux_to_adder_56_port, 
      mux_to_adder_55_port, mux_to_adder_54_port, mux_to_adder_53_port, 
      mux_to_adder_52_port, mux_to_adder_51_port, mux_to_adder_50_port, 
      mux_to_adder_49_port, mux_to_adder_48_port, mux_to_adder_47_port, 
      mux_to_adder_46_port, mux_to_adder_45_port, mux_to_adder_44_port, 
      mux_to_adder_43_port, mux_to_adder_42_port, mux_to_adder_41_port, 
      mux_to_adder_40_port, mux_to_adder_39_port, mux_to_adder_38_port, 
      mux_to_adder_37_port, mux_to_adder_36_port, mux_to_adder_35_port, 
      mux_to_adder_34_port, mux_to_adder_33_port, mux_to_adder_32_port, 
      mux_to_adder_31_port, mux_to_adder_30_port, mux_to_adder_29_port, 
      mux_to_adder_28_port, mux_to_adder_27_port, mux_to_adder_26_port, 
      mux_to_adder_25_port, mux_to_adder_24_port, mux_to_adder_23_port, 
      mux_to_adder_22_port, mux_to_adder_21_port, mux_to_adder_20_port, 
      mux_to_adder_19_port, mux_to_adder_18_port, mux_to_adder_17_port, 
      mux_to_adder_16_port, mux_to_adder_15_port, mux_to_adder_14_port, 
      mux_to_adder_13_port, mux_to_adder_12_port, mux_to_adder_11_port, 
      mux_to_adder_10_port, mux_to_adder_9_port, mux_to_adder_8_port, 
      mux_to_adder_7_port, mux_to_adder_6_port, mux_to_adder_5_port, 
      mux_to_adder_4_port, mux_to_adder_3_port, mux_to_adder_2_port, 
      mux_to_adder_1_port, mux_to_adder_0_port, nextA_0_port, n_3175, n_3176, 
      n_3177 : std_logic;

begin
   nextA <= ( nextA_63_port, nextA_62_port, nextA_61_port, nextA_60_port, 
      nextA_59_port, nextA_58_port, nextA_57_port, nextA_56_port, nextA_55_port
      , nextA_54_port, nextA_53_port, nextA_52_port, nextA_51_port, 
      nextA_50_port, nextA_49_port, nextA_48_port, nextA_47_port, nextA_46_port
      , nextA_45_port, nextA_44_port, nextA_43_port, nextA_42_port, 
      nextA_41_port, nextA_40_port, nextA_39_port, nextA_38_port, nextA_37_port
      , nextA_36_port, nextA_35_port, nextA_34_port, nextA_33_port, 
      nextA_32_port, nextA_31_port, nextA_30_port, nextA_29_port, nextA_28_port
      , nextA_27_port, nextA_26_port, nextA_25_port, nextA_24_port, 
      nextA_23_port, nextA_22_port, nextA_21_port, nextA_20_port, nextA_19_port
      , nextA_18_port, nextA_17_port, nextA_16_port, nextA_15_port, 
      nextA_14_port, nextA_13_port, nextA_12_port, nextA_11_port, nextA_10_port
      , nextA_9_port, nextA_8_port, nextA_7_port, nextA_6_port, nextA_5_port, 
      nextA_4_port, nextA_3_port, nextA_2_port, nextA_1_port, nextA_0_port );
   
   X_Logic0_port <= '0';
   nextA_0_port <= '0';
   encoder_1 : encoder_N64_RADIX3_1 port map( X(2) => encoderIn(2), X(1) => 
                           encoderIn(1), X(0) => encoderIn(0), Z(2) => 
                           encoder_to_mux_2_port, Z(1) => encoder_to_mux_1_port
                           , Z(0) => encoder_to_mux_0_port);
   ShiftnCompl_1 : ShiftnCompl_N64_1 port map( plusA(63) => prevA(63), 
                           plusA(62) => prevA(62), plusA(61) => prevA(61), 
                           plusA(60) => prevA(60), plusA(59) => prevA(59), 
                           plusA(58) => prevA(58), plusA(57) => prevA(57), 
                           plusA(56) => prevA(56), plusA(55) => prevA(55), 
                           plusA(54) => prevA(54), plusA(53) => prevA(53), 
                           plusA(52) => prevA(52), plusA(51) => prevA(51), 
                           plusA(50) => prevA(50), plusA(49) => prevA(49), 
                           plusA(48) => prevA(48), plusA(47) => prevA(47), 
                           plusA(46) => prevA(46), plusA(45) => prevA(45), 
                           plusA(44) => prevA(44), plusA(43) => prevA(43), 
                           plusA(42) => prevA(42), plusA(41) => prevA(41), 
                           plusA(40) => prevA(40), plusA(39) => prevA(39), 
                           plusA(38) => prevA(38), plusA(37) => prevA(37), 
                           plusA(36) => prevA(36), plusA(35) => prevA(35), 
                           plusA(34) => prevA(34), plusA(33) => prevA(33), 
                           plusA(32) => prevA(32), plusA(31) => prevA(31), 
                           plusA(30) => prevA(30), plusA(29) => prevA(29), 
                           plusA(28) => prevA(28), plusA(27) => prevA(27), 
                           plusA(26) => prevA(26), plusA(25) => prevA(25), 
                           plusA(24) => prevA(24), plusA(23) => prevA(23), 
                           plusA(22) => prevA(22), plusA(21) => prevA(21), 
                           plusA(20) => prevA(20), plusA(19) => prevA(19), 
                           plusA(18) => prevA(18), plusA(17) => prevA(17), 
                           plusA(16) => prevA(16), plusA(15) => prevA(15), 
                           plusA(14) => prevA(14), plusA(13) => prevA(13), 
                           plusA(12) => prevA(12), plusA(11) => prevA(11), 
                           plusA(10) => prevA(10), plusA(9) => prevA(9), 
                           plusA(8) => prevA(8), plusA(7) => prevA(7), plusA(6)
                           => prevA(6), plusA(5) => prevA(5), plusA(4) => 
                           prevA(4), plusA(3) => prevA(3), plusA(2) => prevA(2)
                           , plusA(1) => prevA(1), plusA(0) => prevA(0), 
                           plus2A_out(63) => plus2A_s_63_port, plus2A_out(62) 
                           => plus2A_s_62_port, plus2A_out(61) => 
                           plus2A_s_61_port, plus2A_out(60) => plus2A_s_60_port
                           , plus2A_out(59) => plus2A_s_59_port, plus2A_out(58)
                           => plus2A_s_58_port, plus2A_out(57) => 
                           plus2A_s_57_port, plus2A_out(56) => plus2A_s_56_port
                           , plus2A_out(55) => plus2A_s_55_port, plus2A_out(54)
                           => plus2A_s_54_port, plus2A_out(53) => 
                           plus2A_s_53_port, plus2A_out(52) => plus2A_s_52_port
                           , plus2A_out(51) => plus2A_s_51_port, plus2A_out(50)
                           => plus2A_s_50_port, plus2A_out(49) => 
                           plus2A_s_49_port, plus2A_out(48) => plus2A_s_48_port
                           , plus2A_out(47) => plus2A_s_47_port, plus2A_out(46)
                           => plus2A_s_46_port, plus2A_out(45) => 
                           plus2A_s_45_port, plus2A_out(44) => plus2A_s_44_port
                           , plus2A_out(43) => plus2A_s_43_port, plus2A_out(42)
                           => plus2A_s_42_port, plus2A_out(41) => 
                           plus2A_s_41_port, plus2A_out(40) => plus2A_s_40_port
                           , plus2A_out(39) => plus2A_s_39_port, plus2A_out(38)
                           => plus2A_s_38_port, plus2A_out(37) => 
                           plus2A_s_37_port, plus2A_out(36) => plus2A_s_36_port
                           , plus2A_out(35) => plus2A_s_35_port, plus2A_out(34)
                           => plus2A_s_34_port, plus2A_out(33) => 
                           plus2A_s_33_port, plus2A_out(32) => plus2A_s_32_port
                           , plus2A_out(31) => plus2A_s_31_port, plus2A_out(30)
                           => plus2A_s_30_port, plus2A_out(29) => 
                           plus2A_s_29_port, plus2A_out(28) => plus2A_s_28_port
                           , plus2A_out(27) => plus2A_s_27_port, plus2A_out(26)
                           => plus2A_s_26_port, plus2A_out(25) => 
                           plus2A_s_25_port, plus2A_out(24) => plus2A_s_24_port
                           , plus2A_out(23) => plus2A_s_23_port, plus2A_out(22)
                           => plus2A_s_22_port, plus2A_out(21) => 
                           plus2A_s_21_port, plus2A_out(20) => plus2A_s_20_port
                           , plus2A_out(19) => plus2A_s_19_port, plus2A_out(18)
                           => plus2A_s_18_port, plus2A_out(17) => 
                           plus2A_s_17_port, plus2A_out(16) => plus2A_s_16_port
                           , plus2A_out(15) => plus2A_s_15_port, plus2A_out(14)
                           => plus2A_s_14_port, plus2A_out(13) => 
                           plus2A_s_13_port, plus2A_out(12) => plus2A_s_12_port
                           , plus2A_out(11) => plus2A_s_11_port, plus2A_out(10)
                           => plus2A_s_10_port, plus2A_out(9) => 
                           plus2A_s_9_port, plus2A_out(8) => plus2A_s_8_port, 
                           plus2A_out(7) => plus2A_s_7_port, plus2A_out(6) => 
                           plus2A_s_6_port, plus2A_out(5) => plus2A_s_5_port, 
                           plus2A_out(4) => plus2A_s_4_port, plus2A_out(3) => 
                           plus2A_s_3_port, plus2A_out(2) => plus2A_s_2_port, 
                           plus2A_out(1) => plus2A_s_1_port, plus2A_out(0) => 
                           n_3175, minus2A_out(63) => minus2A_s_63_port, 
                           minus2A_out(62) => minus2A_s_62_port, 
                           minus2A_out(61) => minus2A_s_61_port, 
                           minus2A_out(60) => minus2A_s_60_port, 
                           minus2A_out(59) => minus2A_s_59_port, 
                           minus2A_out(58) => minus2A_s_58_port, 
                           minus2A_out(57) => minus2A_s_57_port, 
                           minus2A_out(56) => minus2A_s_56_port, 
                           minus2A_out(55) => minus2A_s_55_port, 
                           minus2A_out(54) => minus2A_s_54_port, 
                           minus2A_out(53) => minus2A_s_53_port, 
                           minus2A_out(52) => minus2A_s_52_port, 
                           minus2A_out(51) => minus2A_s_51_port, 
                           minus2A_out(50) => minus2A_s_50_port, 
                           minus2A_out(49) => minus2A_s_49_port, 
                           minus2A_out(48) => minus2A_s_48_port, 
                           minus2A_out(47) => minus2A_s_47_port, 
                           minus2A_out(46) => minus2A_s_46_port, 
                           minus2A_out(45) => minus2A_s_45_port, 
                           minus2A_out(44) => minus2A_s_44_port, 
                           minus2A_out(43) => minus2A_s_43_port, 
                           minus2A_out(42) => minus2A_s_42_port, 
                           minus2A_out(41) => minus2A_s_41_port, 
                           minus2A_out(40) => minus2A_s_40_port, 
                           minus2A_out(39) => minus2A_s_39_port, 
                           minus2A_out(38) => minus2A_s_38_port, 
                           minus2A_out(37) => minus2A_s_37_port, 
                           minus2A_out(36) => minus2A_s_36_port, 
                           minus2A_out(35) => minus2A_s_35_port, 
                           minus2A_out(34) => minus2A_s_34_port, 
                           minus2A_out(33) => minus2A_s_33_port, 
                           minus2A_out(32) => minus2A_s_32_port, 
                           minus2A_out(31) => minus2A_s_31_port, 
                           minus2A_out(30) => minus2A_s_30_port, 
                           minus2A_out(29) => minus2A_s_29_port, 
                           minus2A_out(28) => minus2A_s_28_port, 
                           minus2A_out(27) => minus2A_s_27_port, 
                           minus2A_out(26) => minus2A_s_26_port, 
                           minus2A_out(25) => minus2A_s_25_port, 
                           minus2A_out(24) => minus2A_s_24_port, 
                           minus2A_out(23) => minus2A_s_23_port, 
                           minus2A_out(22) => minus2A_s_22_port, 
                           minus2A_out(21) => minus2A_s_21_port, 
                           minus2A_out(20) => minus2A_s_20_port, 
                           minus2A_out(19) => minus2A_s_19_port, 
                           minus2A_out(18) => minus2A_s_18_port, 
                           minus2A_out(17) => minus2A_s_17_port, 
                           minus2A_out(16) => minus2A_s_16_port, 
                           minus2A_out(15) => minus2A_s_15_port, 
                           minus2A_out(14) => minus2A_s_14_port, 
                           minus2A_out(13) => minus2A_s_13_port, 
                           minus2A_out(12) => minus2A_s_12_port, 
                           minus2A_out(11) => minus2A_s_11_port, 
                           minus2A_out(10) => minus2A_s_10_port, minus2A_out(9)
                           => minus2A_s_9_port, minus2A_out(8) => 
                           minus2A_s_8_port, minus2A_out(7) => minus2A_s_7_port
                           , minus2A_out(6) => minus2A_s_6_port, minus2A_out(5)
                           => minus2A_s_5_port, minus2A_out(4) => 
                           minus2A_s_4_port, minus2A_out(3) => minus2A_s_3_port
                           , minus2A_out(2) => minus2A_s_2_port, minus2A_out(1)
                           => minus2A_s_1_port, minus2A_out(0) => 
                           minus2A_s_0_port, plus4A_out(63) => nextA_63_port, 
                           plus4A_out(62) => nextA_62_port, plus4A_out(61) => 
                           nextA_61_port, plus4A_out(60) => nextA_60_port, 
                           plus4A_out(59) => nextA_59_port, plus4A_out(58) => 
                           nextA_58_port, plus4A_out(57) => nextA_57_port, 
                           plus4A_out(56) => nextA_56_port, plus4A_out(55) => 
                           nextA_55_port, plus4A_out(54) => nextA_54_port, 
                           plus4A_out(53) => nextA_53_port, plus4A_out(52) => 
                           nextA_52_port, plus4A_out(51) => nextA_51_port, 
                           plus4A_out(50) => nextA_50_port, plus4A_out(49) => 
                           nextA_49_port, plus4A_out(48) => nextA_48_port, 
                           plus4A_out(47) => nextA_47_port, plus4A_out(46) => 
                           nextA_46_port, plus4A_out(45) => nextA_45_port, 
                           plus4A_out(44) => nextA_44_port, plus4A_out(43) => 
                           nextA_43_port, plus4A_out(42) => nextA_42_port, 
                           plus4A_out(41) => nextA_41_port, plus4A_out(40) => 
                           nextA_40_port, plus4A_out(39) => nextA_39_port, 
                           plus4A_out(38) => nextA_38_port, plus4A_out(37) => 
                           nextA_37_port, plus4A_out(36) => nextA_36_port, 
                           plus4A_out(35) => nextA_35_port, plus4A_out(34) => 
                           nextA_34_port, plus4A_out(33) => nextA_33_port, 
                           plus4A_out(32) => nextA_32_port, plus4A_out(31) => 
                           nextA_31_port, plus4A_out(30) => nextA_30_port, 
                           plus4A_out(29) => nextA_29_port, plus4A_out(28) => 
                           nextA_28_port, plus4A_out(27) => nextA_27_port, 
                           plus4A_out(26) => nextA_26_port, plus4A_out(25) => 
                           nextA_25_port, plus4A_out(24) => nextA_24_port, 
                           plus4A_out(23) => nextA_23_port, plus4A_out(22) => 
                           nextA_22_port, plus4A_out(21) => nextA_21_port, 
                           plus4A_out(20) => nextA_20_port, plus4A_out(19) => 
                           nextA_19_port, plus4A_out(18) => nextA_18_port, 
                           plus4A_out(17) => nextA_17_port, plus4A_out(16) => 
                           nextA_16_port, plus4A_out(15) => nextA_15_port, 
                           plus4A_out(14) => nextA_14_port, plus4A_out(13) => 
                           nextA_13_port, plus4A_out(12) => nextA_12_port, 
                           plus4A_out(11) => nextA_11_port, plus4A_out(10) => 
                           nextA_10_port, plus4A_out(9) => nextA_9_port, 
                           plus4A_out(8) => nextA_8_port, plus4A_out(7) => 
                           nextA_7_port, plus4A_out(6) => nextA_6_port, 
                           plus4A_out(5) => nextA_5_port, plus4A_out(4) => 
                           nextA_4_port, plus4A_out(3) => nextA_3_port, 
                           plus4A_out(2) => nextA_2_port, plus4A_out(1) => 
                           nextA_1_port, plus4A_out(0) => n_3176, 
                           minus4A_out(63) => minus4A_s_63_port, 
                           minus4A_out(62) => minus4A_s_62_port, 
                           minus4A_out(61) => minus4A_s_61_port, 
                           minus4A_out(60) => minus4A_s_60_port, 
                           minus4A_out(59) => minus4A_s_59_port, 
                           minus4A_out(58) => minus4A_s_58_port, 
                           minus4A_out(57) => minus4A_s_57_port, 
                           minus4A_out(56) => minus4A_s_56_port, 
                           minus4A_out(55) => minus4A_s_55_port, 
                           minus4A_out(54) => minus4A_s_54_port, 
                           minus4A_out(53) => minus4A_s_53_port, 
                           minus4A_out(52) => minus4A_s_52_port, 
                           minus4A_out(51) => minus4A_s_51_port, 
                           minus4A_out(50) => minus4A_s_50_port, 
                           minus4A_out(49) => minus4A_s_49_port, 
                           minus4A_out(48) => minus4A_s_48_port, 
                           minus4A_out(47) => minus4A_s_47_port, 
                           minus4A_out(46) => minus4A_s_46_port, 
                           minus4A_out(45) => minus4A_s_45_port, 
                           minus4A_out(44) => minus4A_s_44_port, 
                           minus4A_out(43) => minus4A_s_43_port, 
                           minus4A_out(42) => minus4A_s_42_port, 
                           minus4A_out(41) => minus4A_s_41_port, 
                           minus4A_out(40) => minus4A_s_40_port, 
                           minus4A_out(39) => minus4A_s_39_port, 
                           minus4A_out(38) => minus4A_s_38_port, 
                           minus4A_out(37) => minus4A_s_37_port, 
                           minus4A_out(36) => minus4A_s_36_port, 
                           minus4A_out(35) => minus4A_s_35_port, 
                           minus4A_out(34) => minus4A_s_34_port, 
                           minus4A_out(33) => minus4A_s_33_port, 
                           minus4A_out(32) => minus4A_s_32_port, 
                           minus4A_out(31) => minus4A_s_31_port, 
                           minus4A_out(30) => minus4A_s_30_port, 
                           minus4A_out(29) => minus4A_s_29_port, 
                           minus4A_out(28) => minus4A_s_28_port, 
                           minus4A_out(27) => minus4A_s_27_port, 
                           minus4A_out(26) => minus4A_s_26_port, 
                           minus4A_out(25) => minus4A_s_25_port, 
                           minus4A_out(24) => minus4A_s_24_port, 
                           minus4A_out(23) => minus4A_s_23_port, 
                           minus4A_out(22) => minus4A_s_22_port, 
                           minus4A_out(21) => minus4A_s_21_port, 
                           minus4A_out(20) => minus4A_s_20_port, 
                           minus4A_out(19) => minus4A_s_19_port, 
                           minus4A_out(18) => minus4A_s_18_port, 
                           minus4A_out(17) => minus4A_s_17_port, 
                           minus4A_out(16) => minus4A_s_16_port, 
                           minus4A_out(15) => minus4A_s_15_port, 
                           minus4A_out(14) => minus4A_s_14_port, 
                           minus4A_out(13) => minus4A_s_13_port, 
                           minus4A_out(12) => minus4A_s_12_port, 
                           minus4A_out(11) => minus4A_s_11_port, 
                           minus4A_out(10) => minus4A_s_10_port, minus4A_out(9)
                           => minus4A_s_9_port, minus4A_out(8) => 
                           minus4A_s_8_port, minus4A_out(7) => minus4A_s_7_port
                           , minus4A_out(6) => minus4A_s_6_port, minus4A_out(5)
                           => minus4A_s_5_port, minus4A_out(4) => 
                           minus4A_s_4_port, minus4A_out(3) => minus4A_s_3_port
                           , minus4A_out(2) => minus4A_s_2_port, minus4A_out(1)
                           => minus4A_s_1_port, minus4A_out(0) => 
                           minus4A_s_0_port);
   mux_1 : MUX_GENERIC_N64_RADIX3_1 port map( plusA(63) => plus2A_s_63_port, 
                           plusA(62) => plus2A_s_62_port, plusA(61) => 
                           plus2A_s_61_port, plusA(60) => plus2A_s_60_port, 
                           plusA(59) => plus2A_s_59_port, plusA(58) => 
                           plus2A_s_58_port, plusA(57) => plus2A_s_57_port, 
                           plusA(56) => plus2A_s_56_port, plusA(55) => 
                           plus2A_s_55_port, plusA(54) => plus2A_s_54_port, 
                           plusA(53) => plus2A_s_53_port, plusA(52) => 
                           plus2A_s_52_port, plusA(51) => plus2A_s_51_port, 
                           plusA(50) => plus2A_s_50_port, plusA(49) => 
                           plus2A_s_49_port, plusA(48) => plus2A_s_48_port, 
                           plusA(47) => plus2A_s_47_port, plusA(46) => 
                           plus2A_s_46_port, plusA(45) => plus2A_s_45_port, 
                           plusA(44) => plus2A_s_44_port, plusA(43) => 
                           plus2A_s_43_port, plusA(42) => plus2A_s_42_port, 
                           plusA(41) => plus2A_s_41_port, plusA(40) => 
                           plus2A_s_40_port, plusA(39) => plus2A_s_39_port, 
                           plusA(38) => plus2A_s_38_port, plusA(37) => 
                           plus2A_s_37_port, plusA(36) => plus2A_s_36_port, 
                           plusA(35) => plus2A_s_35_port, plusA(34) => 
                           plus2A_s_34_port, plusA(33) => plus2A_s_33_port, 
                           plusA(32) => plus2A_s_32_port, plusA(31) => 
                           plus2A_s_31_port, plusA(30) => plus2A_s_30_port, 
                           plusA(29) => plus2A_s_29_port, plusA(28) => 
                           plus2A_s_28_port, plusA(27) => plus2A_s_27_port, 
                           plusA(26) => plus2A_s_26_port, plusA(25) => 
                           plus2A_s_25_port, plusA(24) => plus2A_s_24_port, 
                           plusA(23) => plus2A_s_23_port, plusA(22) => 
                           plus2A_s_22_port, plusA(21) => plus2A_s_21_port, 
                           plusA(20) => plus2A_s_20_port, plusA(19) => 
                           plus2A_s_19_port, plusA(18) => plus2A_s_18_port, 
                           plusA(17) => plus2A_s_17_port, plusA(16) => 
                           plus2A_s_16_port, plusA(15) => plus2A_s_15_port, 
                           plusA(14) => plus2A_s_14_port, plusA(13) => 
                           plus2A_s_13_port, plusA(12) => plus2A_s_12_port, 
                           plusA(11) => plus2A_s_11_port, plusA(10) => 
                           plus2A_s_10_port, plusA(9) => plus2A_s_9_port, 
                           plusA(8) => plus2A_s_8_port, plusA(7) => 
                           plus2A_s_7_port, plusA(6) => plus2A_s_6_port, 
                           plusA(5) => plus2A_s_5_port, plusA(4) => 
                           plus2A_s_4_port, plusA(3) => plus2A_s_3_port, 
                           plusA(2) => plus2A_s_2_port, plusA(1) => 
                           plus2A_s_1_port, plusA(0) => nextA_0_port, 
                           minusA(63) => minus2A_s_63_port, minusA(62) => 
                           minus2A_s_62_port, minusA(61) => minus2A_s_61_port, 
                           minusA(60) => minus2A_s_60_port, minusA(59) => 
                           minus2A_s_59_port, minusA(58) => minus2A_s_58_port, 
                           minusA(57) => minus2A_s_57_port, minusA(56) => 
                           minus2A_s_56_port, minusA(55) => minus2A_s_55_port, 
                           minusA(54) => minus2A_s_54_port, minusA(53) => 
                           minus2A_s_53_port, minusA(52) => minus2A_s_52_port, 
                           minusA(51) => minus2A_s_51_port, minusA(50) => 
                           minus2A_s_50_port, minusA(49) => minus2A_s_49_port, 
                           minusA(48) => minus2A_s_48_port, minusA(47) => 
                           minus2A_s_47_port, minusA(46) => minus2A_s_46_port, 
                           minusA(45) => minus2A_s_45_port, minusA(44) => 
                           minus2A_s_44_port, minusA(43) => minus2A_s_43_port, 
                           minusA(42) => minus2A_s_42_port, minusA(41) => 
                           minus2A_s_41_port, minusA(40) => minus2A_s_40_port, 
                           minusA(39) => minus2A_s_39_port, minusA(38) => 
                           minus2A_s_38_port, minusA(37) => minus2A_s_37_port, 
                           minusA(36) => minus2A_s_36_port, minusA(35) => 
                           minus2A_s_35_port, minusA(34) => minus2A_s_34_port, 
                           minusA(33) => minus2A_s_33_port, minusA(32) => 
                           minus2A_s_32_port, minusA(31) => minus2A_s_31_port, 
                           minusA(30) => minus2A_s_30_port, minusA(29) => 
                           minus2A_s_29_port, minusA(28) => minus2A_s_28_port, 
                           minusA(27) => minus2A_s_27_port, minusA(26) => 
                           minus2A_s_26_port, minusA(25) => minus2A_s_25_port, 
                           minusA(24) => minus2A_s_24_port, minusA(23) => 
                           minus2A_s_23_port, minusA(22) => minus2A_s_22_port, 
                           minusA(21) => minus2A_s_21_port, minusA(20) => 
                           minus2A_s_20_port, minusA(19) => minus2A_s_19_port, 
                           minusA(18) => minus2A_s_18_port, minusA(17) => 
                           minus2A_s_17_port, minusA(16) => minus2A_s_16_port, 
                           minusA(15) => minus2A_s_15_port, minusA(14) => 
                           minus2A_s_14_port, minusA(13) => minus2A_s_13_port, 
                           minusA(12) => minus2A_s_12_port, minusA(11) => 
                           minus2A_s_11_port, minusA(10) => minus2A_s_10_port, 
                           minusA(9) => minus2A_s_9_port, minusA(8) => 
                           minus2A_s_8_port, minusA(7) => minus2A_s_7_port, 
                           minusA(6) => minus2A_s_6_port, minusA(5) => 
                           minus2A_s_5_port, minusA(4) => minus2A_s_4_port, 
                           minusA(3) => minus2A_s_3_port, minusA(2) => 
                           minus2A_s_2_port, minusA(1) => minus2A_s_1_port, 
                           minusA(0) => minus2A_s_0_port, plus2A(63) => 
                           nextA_63_port, plus2A(62) => nextA_62_port, 
                           plus2A(61) => nextA_61_port, plus2A(60) => 
                           nextA_60_port, plus2A(59) => nextA_59_port, 
                           plus2A(58) => nextA_58_port, plus2A(57) => 
                           nextA_57_port, plus2A(56) => nextA_56_port, 
                           plus2A(55) => nextA_55_port, plus2A(54) => 
                           nextA_54_port, plus2A(53) => nextA_53_port, 
                           plus2A(52) => nextA_52_port, plus2A(51) => 
                           nextA_51_port, plus2A(50) => nextA_50_port, 
                           plus2A(49) => nextA_49_port, plus2A(48) => 
                           nextA_48_port, plus2A(47) => nextA_47_port, 
                           plus2A(46) => nextA_46_port, plus2A(45) => 
                           nextA_45_port, plus2A(44) => nextA_44_port, 
                           plus2A(43) => nextA_43_port, plus2A(42) => 
                           nextA_42_port, plus2A(41) => nextA_41_port, 
                           plus2A(40) => nextA_40_port, plus2A(39) => 
                           nextA_39_port, plus2A(38) => nextA_38_port, 
                           plus2A(37) => nextA_37_port, plus2A(36) => 
                           nextA_36_port, plus2A(35) => nextA_35_port, 
                           plus2A(34) => nextA_34_port, plus2A(33) => 
                           nextA_33_port, plus2A(32) => nextA_32_port, 
                           plus2A(31) => nextA_31_port, plus2A(30) => 
                           nextA_30_port, plus2A(29) => nextA_29_port, 
                           plus2A(28) => nextA_28_port, plus2A(27) => 
                           nextA_27_port, plus2A(26) => nextA_26_port, 
                           plus2A(25) => nextA_25_port, plus2A(24) => 
                           nextA_24_port, plus2A(23) => nextA_23_port, 
                           plus2A(22) => nextA_22_port, plus2A(21) => 
                           nextA_21_port, plus2A(20) => nextA_20_port, 
                           plus2A(19) => nextA_19_port, plus2A(18) => 
                           nextA_18_port, plus2A(17) => nextA_17_port, 
                           plus2A(16) => nextA_16_port, plus2A(15) => 
                           nextA_15_port, plus2A(14) => nextA_14_port, 
                           plus2A(13) => nextA_13_port, plus2A(12) => 
                           nextA_12_port, plus2A(11) => nextA_11_port, 
                           plus2A(10) => nextA_10_port, plus2A(9) => 
                           nextA_9_port, plus2A(8) => nextA_8_port, plus2A(7) 
                           => nextA_7_port, plus2A(6) => nextA_6_port, 
                           plus2A(5) => nextA_5_port, plus2A(4) => nextA_4_port
                           , plus2A(3) => nextA_3_port, plus2A(2) => 
                           nextA_2_port, plus2A(1) => nextA_1_port, plus2A(0) 
                           => nextA_0_port, minus2A(63) => minus4A_s_63_port, 
                           minus2A(62) => minus4A_s_62_port, minus2A(61) => 
                           minus4A_s_61_port, minus2A(60) => minus4A_s_60_port,
                           minus2A(59) => minus4A_s_59_port, minus2A(58) => 
                           minus4A_s_58_port, minus2A(57) => minus4A_s_57_port,
                           minus2A(56) => minus4A_s_56_port, minus2A(55) => 
                           minus4A_s_55_port, minus2A(54) => minus4A_s_54_port,
                           minus2A(53) => minus4A_s_53_port, minus2A(52) => 
                           minus4A_s_52_port, minus2A(51) => minus4A_s_51_port,
                           minus2A(50) => minus4A_s_50_port, minus2A(49) => 
                           minus4A_s_49_port, minus2A(48) => minus4A_s_48_port,
                           minus2A(47) => minus4A_s_47_port, minus2A(46) => 
                           minus4A_s_46_port, minus2A(45) => minus4A_s_45_port,
                           minus2A(44) => minus4A_s_44_port, minus2A(43) => 
                           minus4A_s_43_port, minus2A(42) => minus4A_s_42_port,
                           minus2A(41) => minus4A_s_41_port, minus2A(40) => 
                           minus4A_s_40_port, minus2A(39) => minus4A_s_39_port,
                           minus2A(38) => minus4A_s_38_port, minus2A(37) => 
                           minus4A_s_37_port, minus2A(36) => minus4A_s_36_port,
                           minus2A(35) => minus4A_s_35_port, minus2A(34) => 
                           minus4A_s_34_port, minus2A(33) => minus4A_s_33_port,
                           minus2A(32) => minus4A_s_32_port, minus2A(31) => 
                           minus4A_s_31_port, minus2A(30) => minus4A_s_30_port,
                           minus2A(29) => minus4A_s_29_port, minus2A(28) => 
                           minus4A_s_28_port, minus2A(27) => minus4A_s_27_port,
                           minus2A(26) => minus4A_s_26_port, minus2A(25) => 
                           minus4A_s_25_port, minus2A(24) => minus4A_s_24_port,
                           minus2A(23) => minus4A_s_23_port, minus2A(22) => 
                           minus4A_s_22_port, minus2A(21) => minus4A_s_21_port,
                           minus2A(20) => minus4A_s_20_port, minus2A(19) => 
                           minus4A_s_19_port, minus2A(18) => minus4A_s_18_port,
                           minus2A(17) => minus4A_s_17_port, minus2A(16) => 
                           minus4A_s_16_port, minus2A(15) => minus4A_s_15_port,
                           minus2A(14) => minus4A_s_14_port, minus2A(13) => 
                           minus4A_s_13_port, minus2A(12) => minus4A_s_12_port,
                           minus2A(11) => minus4A_s_11_port, minus2A(10) => 
                           minus4A_s_10_port, minus2A(9) => minus4A_s_9_port, 
                           minus2A(8) => minus4A_s_8_port, minus2A(7) => 
                           minus4A_s_7_port, minus2A(6) => minus4A_s_6_port, 
                           minus2A(5) => minus4A_s_5_port, minus2A(4) => 
                           minus4A_s_4_port, minus2A(3) => minus4A_s_3_port, 
                           minus2A(2) => minus4A_s_2_port, minus2A(1) => 
                           minus4A_s_1_port, minus2A(0) => minus4A_s_0_port, 
                           SEL(2) => encoder_to_mux_2_port, SEL(1) => 
                           encoder_to_mux_1_port, SEL(0) => 
                           encoder_to_mux_0_port, Y(63) => mux_to_adder_63_port
                           , Y(62) => mux_to_adder_62_port, Y(61) => 
                           mux_to_adder_61_port, Y(60) => mux_to_adder_60_port,
                           Y(59) => mux_to_adder_59_port, Y(58) => 
                           mux_to_adder_58_port, Y(57) => mux_to_adder_57_port,
                           Y(56) => mux_to_adder_56_port, Y(55) => 
                           mux_to_adder_55_port, Y(54) => mux_to_adder_54_port,
                           Y(53) => mux_to_adder_53_port, Y(52) => 
                           mux_to_adder_52_port, Y(51) => mux_to_adder_51_port,
                           Y(50) => mux_to_adder_50_port, Y(49) => 
                           mux_to_adder_49_port, Y(48) => mux_to_adder_48_port,
                           Y(47) => mux_to_adder_47_port, Y(46) => 
                           mux_to_adder_46_port, Y(45) => mux_to_adder_45_port,
                           Y(44) => mux_to_adder_44_port, Y(43) => 
                           mux_to_adder_43_port, Y(42) => mux_to_adder_42_port,
                           Y(41) => mux_to_adder_41_port, Y(40) => 
                           mux_to_adder_40_port, Y(39) => mux_to_adder_39_port,
                           Y(38) => mux_to_adder_38_port, Y(37) => 
                           mux_to_adder_37_port, Y(36) => mux_to_adder_36_port,
                           Y(35) => mux_to_adder_35_port, Y(34) => 
                           mux_to_adder_34_port, Y(33) => mux_to_adder_33_port,
                           Y(32) => mux_to_adder_32_port, Y(31) => 
                           mux_to_adder_31_port, Y(30) => mux_to_adder_30_port,
                           Y(29) => mux_to_adder_29_port, Y(28) => 
                           mux_to_adder_28_port, Y(27) => mux_to_adder_27_port,
                           Y(26) => mux_to_adder_26_port, Y(25) => 
                           mux_to_adder_25_port, Y(24) => mux_to_adder_24_port,
                           Y(23) => mux_to_adder_23_port, Y(22) => 
                           mux_to_adder_22_port, Y(21) => mux_to_adder_21_port,
                           Y(20) => mux_to_adder_20_port, Y(19) => 
                           mux_to_adder_19_port, Y(18) => mux_to_adder_18_port,
                           Y(17) => mux_to_adder_17_port, Y(16) => 
                           mux_to_adder_16_port, Y(15) => mux_to_adder_15_port,
                           Y(14) => mux_to_adder_14_port, Y(13) => 
                           mux_to_adder_13_port, Y(12) => mux_to_adder_12_port,
                           Y(11) => mux_to_adder_11_port, Y(10) => 
                           mux_to_adder_10_port, Y(9) => mux_to_adder_9_port, 
                           Y(8) => mux_to_adder_8_port, Y(7) => 
                           mux_to_adder_7_port, Y(6) => mux_to_adder_6_port, 
                           Y(5) => mux_to_adder_5_port, Y(4) => 
                           mux_to_adder_4_port, Y(3) => mux_to_adder_3_port, 
                           Y(2) => mux_to_adder_2_port, Y(1) => 
                           mux_to_adder_1_port, Y(0) => mux_to_adder_0_port);
   rca_1 : RCA_N64_1 port map( A(63) => mux_to_adder_63_port, A(62) => 
                           mux_to_adder_62_port, A(61) => mux_to_adder_61_port,
                           A(60) => mux_to_adder_60_port, A(59) => 
                           mux_to_adder_59_port, A(58) => mux_to_adder_58_port,
                           A(57) => mux_to_adder_57_port, A(56) => 
                           mux_to_adder_56_port, A(55) => mux_to_adder_55_port,
                           A(54) => mux_to_adder_54_port, A(53) => 
                           mux_to_adder_53_port, A(52) => mux_to_adder_52_port,
                           A(51) => mux_to_adder_51_port, A(50) => 
                           mux_to_adder_50_port, A(49) => mux_to_adder_49_port,
                           A(48) => mux_to_adder_48_port, A(47) => 
                           mux_to_adder_47_port, A(46) => mux_to_adder_46_port,
                           A(45) => mux_to_adder_45_port, A(44) => 
                           mux_to_adder_44_port, A(43) => mux_to_adder_43_port,
                           A(42) => mux_to_adder_42_port, A(41) => 
                           mux_to_adder_41_port, A(40) => mux_to_adder_40_port,
                           A(39) => mux_to_adder_39_port, A(38) => 
                           mux_to_adder_38_port, A(37) => mux_to_adder_37_port,
                           A(36) => mux_to_adder_36_port, A(35) => 
                           mux_to_adder_35_port, A(34) => mux_to_adder_34_port,
                           A(33) => mux_to_adder_33_port, A(32) => 
                           mux_to_adder_32_port, A(31) => mux_to_adder_31_port,
                           A(30) => mux_to_adder_30_port, A(29) => 
                           mux_to_adder_29_port, A(28) => mux_to_adder_28_port,
                           A(27) => mux_to_adder_27_port, A(26) => 
                           mux_to_adder_26_port, A(25) => mux_to_adder_25_port,
                           A(24) => mux_to_adder_24_port, A(23) => 
                           mux_to_adder_23_port, A(22) => mux_to_adder_22_port,
                           A(21) => mux_to_adder_21_port, A(20) => 
                           mux_to_adder_20_port, A(19) => mux_to_adder_19_port,
                           A(18) => mux_to_adder_18_port, A(17) => 
                           mux_to_adder_17_port, A(16) => mux_to_adder_16_port,
                           A(15) => mux_to_adder_15_port, A(14) => 
                           mux_to_adder_14_port, A(13) => mux_to_adder_13_port,
                           A(12) => mux_to_adder_12_port, A(11) => 
                           mux_to_adder_11_port, A(10) => mux_to_adder_10_port,
                           A(9) => mux_to_adder_9_port, A(8) => 
                           mux_to_adder_8_port, A(7) => mux_to_adder_7_port, 
                           A(6) => mux_to_adder_6_port, A(5) => 
                           mux_to_adder_5_port, A(4) => mux_to_adder_4_port, 
                           A(3) => mux_to_adder_3_port, A(2) => 
                           mux_to_adder_2_port, A(1) => mux_to_adder_1_port, 
                           A(0) => mux_to_adder_0_port, B(63) => prevSum(63), 
                           B(62) => prevSum(62), B(61) => prevSum(61), B(60) =>
                           prevSum(60), B(59) => prevSum(59), B(58) => 
                           prevSum(58), B(57) => prevSum(57), B(56) => 
                           prevSum(56), B(55) => prevSum(55), B(54) => 
                           prevSum(54), B(53) => prevSum(53), B(52) => 
                           prevSum(52), B(51) => prevSum(51), B(50) => 
                           prevSum(50), B(49) => prevSum(49), B(48) => 
                           prevSum(48), B(47) => prevSum(47), B(46) => 
                           prevSum(46), B(45) => prevSum(45), B(44) => 
                           prevSum(44), B(43) => prevSum(43), B(42) => 
                           prevSum(42), B(41) => prevSum(41), B(40) => 
                           prevSum(40), B(39) => prevSum(39), B(38) => 
                           prevSum(38), B(37) => prevSum(37), B(36) => 
                           prevSum(36), B(35) => prevSum(35), B(34) => 
                           prevSum(34), B(33) => prevSum(33), B(32) => 
                           prevSum(32), B(31) => prevSum(31), B(30) => 
                           prevSum(30), B(29) => prevSum(29), B(28) => 
                           prevSum(28), B(27) => prevSum(27), B(26) => 
                           prevSum(26), B(25) => prevSum(25), B(24) => 
                           prevSum(24), B(23) => prevSum(23), B(22) => 
                           prevSum(22), B(21) => prevSum(21), B(20) => 
                           prevSum(20), B(19) => prevSum(19), B(18) => 
                           prevSum(18), B(17) => prevSum(17), B(16) => 
                           prevSum(16), B(15) => prevSum(15), B(14) => 
                           prevSum(14), B(13) => prevSum(13), B(12) => 
                           prevSum(12), B(11) => prevSum(11), B(10) => 
                           prevSum(10), B(9) => prevSum(9), B(8) => prevSum(8),
                           B(7) => prevSum(7), B(6) => prevSum(6), B(5) => 
                           prevSum(5), B(4) => prevSum(4), B(3) => prevSum(3), 
                           B(2) => prevSum(2), B(1) => prevSum(1), B(0) => 
                           prevSum(0), Ci => X_Logic0_port, S(63) => 
                           nextSum(63), S(62) => nextSum(62), S(61) => 
                           nextSum(61), S(60) => nextSum(60), S(59) => 
                           nextSum(59), S(58) => nextSum(58), S(57) => 
                           nextSum(57), S(56) => nextSum(56), S(55) => 
                           nextSum(55), S(54) => nextSum(54), S(53) => 
                           nextSum(53), S(52) => nextSum(52), S(51) => 
                           nextSum(51), S(50) => nextSum(50), S(49) => 
                           nextSum(49), S(48) => nextSum(48), S(47) => 
                           nextSum(47), S(46) => nextSum(46), S(45) => 
                           nextSum(45), S(44) => nextSum(44), S(43) => 
                           nextSum(43), S(42) => nextSum(42), S(41) => 
                           nextSum(41), S(40) => nextSum(40), S(39) => 
                           nextSum(39), S(38) => nextSum(38), S(37) => 
                           nextSum(37), S(36) => nextSum(36), S(35) => 
                           nextSum(35), S(34) => nextSum(34), S(33) => 
                           nextSum(33), S(32) => nextSum(32), S(31) => 
                           nextSum(31), S(30) => nextSum(30), S(29) => 
                           nextSum(29), S(28) => nextSum(28), S(27) => 
                           nextSum(27), S(26) => nextSum(26), S(25) => 
                           nextSum(25), S(24) => nextSum(24), S(23) => 
                           nextSum(23), S(22) => nextSum(22), S(21) => 
                           nextSum(21), S(20) => nextSum(20), S(19) => 
                           nextSum(19), S(18) => nextSum(18), S(17) => 
                           nextSum(17), S(16) => nextSum(16), S(15) => 
                           nextSum(15), S(14) => nextSum(14), S(13) => 
                           nextSum(13), S(12) => nextSum(12), S(11) => 
                           nextSum(11), S(10) => nextSum(10), S(9) => 
                           nextSum(9), S(8) => nextSum(8), S(7) => nextSum(7), 
                           S(6) => nextSum(6), S(5) => nextSum(5), S(4) => 
                           nextSum(4), S(3) => nextSum(3), S(2) => nextSum(2), 
                           S(1) => nextSum(1), S(0) => nextSum(0), Co => n_3177
                           );

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity booth_mul_row_N64_RADIX3_2 is

   port( prevA, prevSum : in std_logic_vector (63 downto 0);  encoderIn : in 
         std_logic_vector (2 downto 0);  nextA, nextSum : out std_logic_vector 
         (63 downto 0));

end booth_mul_row_N64_RADIX3_2;

architecture SYN_struct of booth_mul_row_N64_RADIX3_2 is

   component RCA_N64_2
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component MUX_GENERIC_N64_RADIX3_2
      port( plusA, minusA, plus2A, minus2A : in std_logic_vector (63 downto 0);
            SEL : in std_logic_vector (2 downto 0);  Y : out std_logic_vector 
            (63 downto 0));
   end component;
   
   component ShiftnCompl_N64_2
      port( plusA : in std_logic_vector (63 downto 0);  plus2A_out, minus2A_out
            , plus4A_out, minus4A_out : out std_logic_vector (63 downto 0));
   end component;
   
   component encoder_N64_RADIX3_2
      port( X : in std_logic_vector (2 downto 0);  Z : out std_logic_vector (2 
            downto 0));
   end component;
   
   signal X_Logic0_port, nextA_63_port, nextA_62_port, nextA_61_port, 
      nextA_60_port, nextA_59_port, nextA_58_port, nextA_57_port, nextA_56_port
      , nextA_55_port, nextA_54_port, nextA_53_port, nextA_52_port, 
      nextA_51_port, nextA_50_port, nextA_49_port, nextA_48_port, nextA_47_port
      , nextA_46_port, nextA_45_port, nextA_44_port, nextA_43_port, 
      nextA_42_port, nextA_41_port, nextA_40_port, nextA_39_port, nextA_38_port
      , nextA_37_port, nextA_36_port, nextA_35_port, nextA_34_port, 
      nextA_33_port, nextA_32_port, nextA_31_port, nextA_30_port, nextA_29_port
      , nextA_28_port, nextA_27_port, nextA_26_port, nextA_25_port, 
      nextA_24_port, nextA_23_port, nextA_22_port, nextA_21_port, nextA_20_port
      , nextA_19_port, nextA_18_port, nextA_17_port, nextA_16_port, 
      nextA_15_port, nextA_14_port, nextA_13_port, nextA_12_port, nextA_11_port
      , nextA_10_port, nextA_9_port, nextA_8_port, nextA_7_port, nextA_6_port, 
      nextA_5_port, nextA_4_port, nextA_3_port, nextA_2_port, nextA_1_port, 
      encoder_to_mux_2_port, encoder_to_mux_1_port, encoder_to_mux_0_port, 
      plus2A_s_63_port, plus2A_s_62_port, plus2A_s_61_port, plus2A_s_60_port, 
      plus2A_s_59_port, plus2A_s_58_port, plus2A_s_57_port, plus2A_s_56_port, 
      plus2A_s_55_port, plus2A_s_54_port, plus2A_s_53_port, plus2A_s_52_port, 
      plus2A_s_51_port, plus2A_s_50_port, plus2A_s_49_port, plus2A_s_48_port, 
      plus2A_s_47_port, plus2A_s_46_port, plus2A_s_45_port, plus2A_s_44_port, 
      plus2A_s_43_port, plus2A_s_42_port, plus2A_s_41_port, plus2A_s_40_port, 
      plus2A_s_39_port, plus2A_s_38_port, plus2A_s_37_port, plus2A_s_36_port, 
      plus2A_s_35_port, plus2A_s_34_port, plus2A_s_33_port, plus2A_s_32_port, 
      plus2A_s_31_port, plus2A_s_30_port, plus2A_s_29_port, plus2A_s_28_port, 
      plus2A_s_27_port, plus2A_s_26_port, plus2A_s_25_port, plus2A_s_24_port, 
      plus2A_s_23_port, plus2A_s_22_port, plus2A_s_21_port, plus2A_s_20_port, 
      plus2A_s_19_port, plus2A_s_18_port, plus2A_s_17_port, plus2A_s_16_port, 
      plus2A_s_15_port, plus2A_s_14_port, plus2A_s_13_port, plus2A_s_12_port, 
      plus2A_s_11_port, plus2A_s_10_port, plus2A_s_9_port, plus2A_s_8_port, 
      plus2A_s_7_port, plus2A_s_6_port, plus2A_s_5_port, plus2A_s_4_port, 
      plus2A_s_3_port, plus2A_s_2_port, plus2A_s_1_port, minus2A_s_63_port, 
      minus2A_s_62_port, minus2A_s_61_port, minus2A_s_60_port, 
      minus2A_s_59_port, minus2A_s_58_port, minus2A_s_57_port, 
      minus2A_s_56_port, minus2A_s_55_port, minus2A_s_54_port, 
      minus2A_s_53_port, minus2A_s_52_port, minus2A_s_51_port, 
      minus2A_s_50_port, minus2A_s_49_port, minus2A_s_48_port, 
      minus2A_s_47_port, minus2A_s_46_port, minus2A_s_45_port, 
      minus2A_s_44_port, minus2A_s_43_port, minus2A_s_42_port, 
      minus2A_s_41_port, minus2A_s_40_port, minus2A_s_39_port, 
      minus2A_s_38_port, minus2A_s_37_port, minus2A_s_36_port, 
      minus2A_s_35_port, minus2A_s_34_port, minus2A_s_33_port, 
      minus2A_s_32_port, minus2A_s_31_port, minus2A_s_30_port, 
      minus2A_s_29_port, minus2A_s_28_port, minus2A_s_27_port, 
      minus2A_s_26_port, minus2A_s_25_port, minus2A_s_24_port, 
      minus2A_s_23_port, minus2A_s_22_port, minus2A_s_21_port, 
      minus2A_s_20_port, minus2A_s_19_port, minus2A_s_18_port, 
      minus2A_s_17_port, minus2A_s_16_port, minus2A_s_15_port, 
      minus2A_s_14_port, minus2A_s_13_port, minus2A_s_12_port, 
      minus2A_s_11_port, minus2A_s_10_port, minus2A_s_9_port, minus2A_s_8_port,
      minus2A_s_7_port, minus2A_s_6_port, minus2A_s_5_port, minus2A_s_4_port, 
      minus2A_s_3_port, minus2A_s_2_port, minus2A_s_1_port, minus2A_s_0_port, 
      minus4A_s_63_port, minus4A_s_62_port, minus4A_s_61_port, 
      minus4A_s_60_port, minus4A_s_59_port, minus4A_s_58_port, 
      minus4A_s_57_port, minus4A_s_56_port, minus4A_s_55_port, 
      minus4A_s_54_port, minus4A_s_53_port, minus4A_s_52_port, 
      minus4A_s_51_port, minus4A_s_50_port, minus4A_s_49_port, 
      minus4A_s_48_port, minus4A_s_47_port, minus4A_s_46_port, 
      minus4A_s_45_port, minus4A_s_44_port, minus4A_s_43_port, 
      minus4A_s_42_port, minus4A_s_41_port, minus4A_s_40_port, 
      minus4A_s_39_port, minus4A_s_38_port, minus4A_s_37_port, 
      minus4A_s_36_port, minus4A_s_35_port, minus4A_s_34_port, 
      minus4A_s_33_port, minus4A_s_32_port, minus4A_s_31_port, 
      minus4A_s_30_port, minus4A_s_29_port, minus4A_s_28_port, 
      minus4A_s_27_port, minus4A_s_26_port, minus4A_s_25_port, 
      minus4A_s_24_port, minus4A_s_23_port, minus4A_s_22_port, 
      minus4A_s_21_port, minus4A_s_20_port, minus4A_s_19_port, 
      minus4A_s_18_port, minus4A_s_17_port, minus4A_s_16_port, 
      minus4A_s_15_port, minus4A_s_14_port, minus4A_s_13_port, 
      minus4A_s_12_port, minus4A_s_11_port, minus4A_s_10_port, minus4A_s_9_port
      , minus4A_s_8_port, minus4A_s_7_port, minus4A_s_6_port, minus4A_s_5_port,
      minus4A_s_4_port, minus4A_s_3_port, minus4A_s_2_port, minus4A_s_1_port, 
      minus4A_s_0_port, mux_to_adder_63_port, mux_to_adder_62_port, 
      mux_to_adder_61_port, mux_to_adder_60_port, mux_to_adder_59_port, 
      mux_to_adder_58_port, mux_to_adder_57_port, mux_to_adder_56_port, 
      mux_to_adder_55_port, mux_to_adder_54_port, mux_to_adder_53_port, 
      mux_to_adder_52_port, mux_to_adder_51_port, mux_to_adder_50_port, 
      mux_to_adder_49_port, mux_to_adder_48_port, mux_to_adder_47_port, 
      mux_to_adder_46_port, mux_to_adder_45_port, mux_to_adder_44_port, 
      mux_to_adder_43_port, mux_to_adder_42_port, mux_to_adder_41_port, 
      mux_to_adder_40_port, mux_to_adder_39_port, mux_to_adder_38_port, 
      mux_to_adder_37_port, mux_to_adder_36_port, mux_to_adder_35_port, 
      mux_to_adder_34_port, mux_to_adder_33_port, mux_to_adder_32_port, 
      mux_to_adder_31_port, mux_to_adder_30_port, mux_to_adder_29_port, 
      mux_to_adder_28_port, mux_to_adder_27_port, mux_to_adder_26_port, 
      mux_to_adder_25_port, mux_to_adder_24_port, mux_to_adder_23_port, 
      mux_to_adder_22_port, mux_to_adder_21_port, mux_to_adder_20_port, 
      mux_to_adder_19_port, mux_to_adder_18_port, mux_to_adder_17_port, 
      mux_to_adder_16_port, mux_to_adder_15_port, mux_to_adder_14_port, 
      mux_to_adder_13_port, mux_to_adder_12_port, mux_to_adder_11_port, 
      mux_to_adder_10_port, mux_to_adder_9_port, mux_to_adder_8_port, 
      mux_to_adder_7_port, mux_to_adder_6_port, mux_to_adder_5_port, 
      mux_to_adder_4_port, mux_to_adder_3_port, mux_to_adder_2_port, 
      mux_to_adder_1_port, mux_to_adder_0_port, nextA_0_port, n_3178, n_3179, 
      n_3180 : std_logic;

begin
   nextA <= ( nextA_63_port, nextA_62_port, nextA_61_port, nextA_60_port, 
      nextA_59_port, nextA_58_port, nextA_57_port, nextA_56_port, nextA_55_port
      , nextA_54_port, nextA_53_port, nextA_52_port, nextA_51_port, 
      nextA_50_port, nextA_49_port, nextA_48_port, nextA_47_port, nextA_46_port
      , nextA_45_port, nextA_44_port, nextA_43_port, nextA_42_port, 
      nextA_41_port, nextA_40_port, nextA_39_port, nextA_38_port, nextA_37_port
      , nextA_36_port, nextA_35_port, nextA_34_port, nextA_33_port, 
      nextA_32_port, nextA_31_port, nextA_30_port, nextA_29_port, nextA_28_port
      , nextA_27_port, nextA_26_port, nextA_25_port, nextA_24_port, 
      nextA_23_port, nextA_22_port, nextA_21_port, nextA_20_port, nextA_19_port
      , nextA_18_port, nextA_17_port, nextA_16_port, nextA_15_port, 
      nextA_14_port, nextA_13_port, nextA_12_port, nextA_11_port, nextA_10_port
      , nextA_9_port, nextA_8_port, nextA_7_port, nextA_6_port, nextA_5_port, 
      nextA_4_port, nextA_3_port, nextA_2_port, nextA_1_port, nextA_0_port );
   
   X_Logic0_port <= '0';
   nextA_0_port <= '0';
   encoder_1 : encoder_N64_RADIX3_2 port map( X(2) => encoderIn(2), X(1) => 
                           encoderIn(1), X(0) => encoderIn(0), Z(2) => 
                           encoder_to_mux_2_port, Z(1) => encoder_to_mux_1_port
                           , Z(0) => encoder_to_mux_0_port);
   ShiftnCompl_1 : ShiftnCompl_N64_2 port map( plusA(63) => prevA(63), 
                           plusA(62) => prevA(62), plusA(61) => prevA(61), 
                           plusA(60) => prevA(60), plusA(59) => prevA(59), 
                           plusA(58) => prevA(58), plusA(57) => prevA(57), 
                           plusA(56) => prevA(56), plusA(55) => prevA(55), 
                           plusA(54) => prevA(54), plusA(53) => prevA(53), 
                           plusA(52) => prevA(52), plusA(51) => prevA(51), 
                           plusA(50) => prevA(50), plusA(49) => prevA(49), 
                           plusA(48) => prevA(48), plusA(47) => prevA(47), 
                           plusA(46) => prevA(46), plusA(45) => prevA(45), 
                           plusA(44) => prevA(44), plusA(43) => prevA(43), 
                           plusA(42) => prevA(42), plusA(41) => prevA(41), 
                           plusA(40) => prevA(40), plusA(39) => prevA(39), 
                           plusA(38) => prevA(38), plusA(37) => prevA(37), 
                           plusA(36) => prevA(36), plusA(35) => prevA(35), 
                           plusA(34) => prevA(34), plusA(33) => prevA(33), 
                           plusA(32) => prevA(32), plusA(31) => prevA(31), 
                           plusA(30) => prevA(30), plusA(29) => prevA(29), 
                           plusA(28) => prevA(28), plusA(27) => prevA(27), 
                           plusA(26) => prevA(26), plusA(25) => prevA(25), 
                           plusA(24) => prevA(24), plusA(23) => prevA(23), 
                           plusA(22) => prevA(22), plusA(21) => prevA(21), 
                           plusA(20) => prevA(20), plusA(19) => prevA(19), 
                           plusA(18) => prevA(18), plusA(17) => prevA(17), 
                           plusA(16) => prevA(16), plusA(15) => prevA(15), 
                           plusA(14) => prevA(14), plusA(13) => prevA(13), 
                           plusA(12) => prevA(12), plusA(11) => prevA(11), 
                           plusA(10) => prevA(10), plusA(9) => prevA(9), 
                           plusA(8) => prevA(8), plusA(7) => prevA(7), plusA(6)
                           => prevA(6), plusA(5) => prevA(5), plusA(4) => 
                           prevA(4), plusA(3) => prevA(3), plusA(2) => prevA(2)
                           , plusA(1) => prevA(1), plusA(0) => prevA(0), 
                           plus2A_out(63) => plus2A_s_63_port, plus2A_out(62) 
                           => plus2A_s_62_port, plus2A_out(61) => 
                           plus2A_s_61_port, plus2A_out(60) => plus2A_s_60_port
                           , plus2A_out(59) => plus2A_s_59_port, plus2A_out(58)
                           => plus2A_s_58_port, plus2A_out(57) => 
                           plus2A_s_57_port, plus2A_out(56) => plus2A_s_56_port
                           , plus2A_out(55) => plus2A_s_55_port, plus2A_out(54)
                           => plus2A_s_54_port, plus2A_out(53) => 
                           plus2A_s_53_port, plus2A_out(52) => plus2A_s_52_port
                           , plus2A_out(51) => plus2A_s_51_port, plus2A_out(50)
                           => plus2A_s_50_port, plus2A_out(49) => 
                           plus2A_s_49_port, plus2A_out(48) => plus2A_s_48_port
                           , plus2A_out(47) => plus2A_s_47_port, plus2A_out(46)
                           => plus2A_s_46_port, plus2A_out(45) => 
                           plus2A_s_45_port, plus2A_out(44) => plus2A_s_44_port
                           , plus2A_out(43) => plus2A_s_43_port, plus2A_out(42)
                           => plus2A_s_42_port, plus2A_out(41) => 
                           plus2A_s_41_port, plus2A_out(40) => plus2A_s_40_port
                           , plus2A_out(39) => plus2A_s_39_port, plus2A_out(38)
                           => plus2A_s_38_port, plus2A_out(37) => 
                           plus2A_s_37_port, plus2A_out(36) => plus2A_s_36_port
                           , plus2A_out(35) => plus2A_s_35_port, plus2A_out(34)
                           => plus2A_s_34_port, plus2A_out(33) => 
                           plus2A_s_33_port, plus2A_out(32) => plus2A_s_32_port
                           , plus2A_out(31) => plus2A_s_31_port, plus2A_out(30)
                           => plus2A_s_30_port, plus2A_out(29) => 
                           plus2A_s_29_port, plus2A_out(28) => plus2A_s_28_port
                           , plus2A_out(27) => plus2A_s_27_port, plus2A_out(26)
                           => plus2A_s_26_port, plus2A_out(25) => 
                           plus2A_s_25_port, plus2A_out(24) => plus2A_s_24_port
                           , plus2A_out(23) => plus2A_s_23_port, plus2A_out(22)
                           => plus2A_s_22_port, plus2A_out(21) => 
                           plus2A_s_21_port, plus2A_out(20) => plus2A_s_20_port
                           , plus2A_out(19) => plus2A_s_19_port, plus2A_out(18)
                           => plus2A_s_18_port, plus2A_out(17) => 
                           plus2A_s_17_port, plus2A_out(16) => plus2A_s_16_port
                           , plus2A_out(15) => plus2A_s_15_port, plus2A_out(14)
                           => plus2A_s_14_port, plus2A_out(13) => 
                           plus2A_s_13_port, plus2A_out(12) => plus2A_s_12_port
                           , plus2A_out(11) => plus2A_s_11_port, plus2A_out(10)
                           => plus2A_s_10_port, plus2A_out(9) => 
                           plus2A_s_9_port, plus2A_out(8) => plus2A_s_8_port, 
                           plus2A_out(7) => plus2A_s_7_port, plus2A_out(6) => 
                           plus2A_s_6_port, plus2A_out(5) => plus2A_s_5_port, 
                           plus2A_out(4) => plus2A_s_4_port, plus2A_out(3) => 
                           plus2A_s_3_port, plus2A_out(2) => plus2A_s_2_port, 
                           plus2A_out(1) => plus2A_s_1_port, plus2A_out(0) => 
                           n_3178, minus2A_out(63) => minus2A_s_63_port, 
                           minus2A_out(62) => minus2A_s_62_port, 
                           minus2A_out(61) => minus2A_s_61_port, 
                           minus2A_out(60) => minus2A_s_60_port, 
                           minus2A_out(59) => minus2A_s_59_port, 
                           minus2A_out(58) => minus2A_s_58_port, 
                           minus2A_out(57) => minus2A_s_57_port, 
                           minus2A_out(56) => minus2A_s_56_port, 
                           minus2A_out(55) => minus2A_s_55_port, 
                           minus2A_out(54) => minus2A_s_54_port, 
                           minus2A_out(53) => minus2A_s_53_port, 
                           minus2A_out(52) => minus2A_s_52_port, 
                           minus2A_out(51) => minus2A_s_51_port, 
                           minus2A_out(50) => minus2A_s_50_port, 
                           minus2A_out(49) => minus2A_s_49_port, 
                           minus2A_out(48) => minus2A_s_48_port, 
                           minus2A_out(47) => minus2A_s_47_port, 
                           minus2A_out(46) => minus2A_s_46_port, 
                           minus2A_out(45) => minus2A_s_45_port, 
                           minus2A_out(44) => minus2A_s_44_port, 
                           minus2A_out(43) => minus2A_s_43_port, 
                           minus2A_out(42) => minus2A_s_42_port, 
                           minus2A_out(41) => minus2A_s_41_port, 
                           minus2A_out(40) => minus2A_s_40_port, 
                           minus2A_out(39) => minus2A_s_39_port, 
                           minus2A_out(38) => minus2A_s_38_port, 
                           minus2A_out(37) => minus2A_s_37_port, 
                           minus2A_out(36) => minus2A_s_36_port, 
                           minus2A_out(35) => minus2A_s_35_port, 
                           minus2A_out(34) => minus2A_s_34_port, 
                           minus2A_out(33) => minus2A_s_33_port, 
                           minus2A_out(32) => minus2A_s_32_port, 
                           minus2A_out(31) => minus2A_s_31_port, 
                           minus2A_out(30) => minus2A_s_30_port, 
                           minus2A_out(29) => minus2A_s_29_port, 
                           minus2A_out(28) => minus2A_s_28_port, 
                           minus2A_out(27) => minus2A_s_27_port, 
                           minus2A_out(26) => minus2A_s_26_port, 
                           minus2A_out(25) => minus2A_s_25_port, 
                           minus2A_out(24) => minus2A_s_24_port, 
                           minus2A_out(23) => minus2A_s_23_port, 
                           minus2A_out(22) => minus2A_s_22_port, 
                           minus2A_out(21) => minus2A_s_21_port, 
                           minus2A_out(20) => minus2A_s_20_port, 
                           minus2A_out(19) => minus2A_s_19_port, 
                           minus2A_out(18) => minus2A_s_18_port, 
                           minus2A_out(17) => minus2A_s_17_port, 
                           minus2A_out(16) => minus2A_s_16_port, 
                           minus2A_out(15) => minus2A_s_15_port, 
                           minus2A_out(14) => minus2A_s_14_port, 
                           minus2A_out(13) => minus2A_s_13_port, 
                           minus2A_out(12) => minus2A_s_12_port, 
                           minus2A_out(11) => minus2A_s_11_port, 
                           minus2A_out(10) => minus2A_s_10_port, minus2A_out(9)
                           => minus2A_s_9_port, minus2A_out(8) => 
                           minus2A_s_8_port, minus2A_out(7) => minus2A_s_7_port
                           , minus2A_out(6) => minus2A_s_6_port, minus2A_out(5)
                           => minus2A_s_5_port, minus2A_out(4) => 
                           minus2A_s_4_port, minus2A_out(3) => minus2A_s_3_port
                           , minus2A_out(2) => minus2A_s_2_port, minus2A_out(1)
                           => minus2A_s_1_port, minus2A_out(0) => 
                           minus2A_s_0_port, plus4A_out(63) => nextA_63_port, 
                           plus4A_out(62) => nextA_62_port, plus4A_out(61) => 
                           nextA_61_port, plus4A_out(60) => nextA_60_port, 
                           plus4A_out(59) => nextA_59_port, plus4A_out(58) => 
                           nextA_58_port, plus4A_out(57) => nextA_57_port, 
                           plus4A_out(56) => nextA_56_port, plus4A_out(55) => 
                           nextA_55_port, plus4A_out(54) => nextA_54_port, 
                           plus4A_out(53) => nextA_53_port, plus4A_out(52) => 
                           nextA_52_port, plus4A_out(51) => nextA_51_port, 
                           plus4A_out(50) => nextA_50_port, plus4A_out(49) => 
                           nextA_49_port, plus4A_out(48) => nextA_48_port, 
                           plus4A_out(47) => nextA_47_port, plus4A_out(46) => 
                           nextA_46_port, plus4A_out(45) => nextA_45_port, 
                           plus4A_out(44) => nextA_44_port, plus4A_out(43) => 
                           nextA_43_port, plus4A_out(42) => nextA_42_port, 
                           plus4A_out(41) => nextA_41_port, plus4A_out(40) => 
                           nextA_40_port, plus4A_out(39) => nextA_39_port, 
                           plus4A_out(38) => nextA_38_port, plus4A_out(37) => 
                           nextA_37_port, plus4A_out(36) => nextA_36_port, 
                           plus4A_out(35) => nextA_35_port, plus4A_out(34) => 
                           nextA_34_port, plus4A_out(33) => nextA_33_port, 
                           plus4A_out(32) => nextA_32_port, plus4A_out(31) => 
                           nextA_31_port, plus4A_out(30) => nextA_30_port, 
                           plus4A_out(29) => nextA_29_port, plus4A_out(28) => 
                           nextA_28_port, plus4A_out(27) => nextA_27_port, 
                           plus4A_out(26) => nextA_26_port, plus4A_out(25) => 
                           nextA_25_port, plus4A_out(24) => nextA_24_port, 
                           plus4A_out(23) => nextA_23_port, plus4A_out(22) => 
                           nextA_22_port, plus4A_out(21) => nextA_21_port, 
                           plus4A_out(20) => nextA_20_port, plus4A_out(19) => 
                           nextA_19_port, plus4A_out(18) => nextA_18_port, 
                           plus4A_out(17) => nextA_17_port, plus4A_out(16) => 
                           nextA_16_port, plus4A_out(15) => nextA_15_port, 
                           plus4A_out(14) => nextA_14_port, plus4A_out(13) => 
                           nextA_13_port, plus4A_out(12) => nextA_12_port, 
                           plus4A_out(11) => nextA_11_port, plus4A_out(10) => 
                           nextA_10_port, plus4A_out(9) => nextA_9_port, 
                           plus4A_out(8) => nextA_8_port, plus4A_out(7) => 
                           nextA_7_port, plus4A_out(6) => nextA_6_port, 
                           plus4A_out(5) => nextA_5_port, plus4A_out(4) => 
                           nextA_4_port, plus4A_out(3) => nextA_3_port, 
                           plus4A_out(2) => nextA_2_port, plus4A_out(1) => 
                           nextA_1_port, plus4A_out(0) => n_3179, 
                           minus4A_out(63) => minus4A_s_63_port, 
                           minus4A_out(62) => minus4A_s_62_port, 
                           minus4A_out(61) => minus4A_s_61_port, 
                           minus4A_out(60) => minus4A_s_60_port, 
                           minus4A_out(59) => minus4A_s_59_port, 
                           minus4A_out(58) => minus4A_s_58_port, 
                           minus4A_out(57) => minus4A_s_57_port, 
                           minus4A_out(56) => minus4A_s_56_port, 
                           minus4A_out(55) => minus4A_s_55_port, 
                           minus4A_out(54) => minus4A_s_54_port, 
                           minus4A_out(53) => minus4A_s_53_port, 
                           minus4A_out(52) => minus4A_s_52_port, 
                           minus4A_out(51) => minus4A_s_51_port, 
                           minus4A_out(50) => minus4A_s_50_port, 
                           minus4A_out(49) => minus4A_s_49_port, 
                           minus4A_out(48) => minus4A_s_48_port, 
                           minus4A_out(47) => minus4A_s_47_port, 
                           minus4A_out(46) => minus4A_s_46_port, 
                           minus4A_out(45) => minus4A_s_45_port, 
                           minus4A_out(44) => minus4A_s_44_port, 
                           minus4A_out(43) => minus4A_s_43_port, 
                           minus4A_out(42) => minus4A_s_42_port, 
                           minus4A_out(41) => minus4A_s_41_port, 
                           minus4A_out(40) => minus4A_s_40_port, 
                           minus4A_out(39) => minus4A_s_39_port, 
                           minus4A_out(38) => minus4A_s_38_port, 
                           minus4A_out(37) => minus4A_s_37_port, 
                           minus4A_out(36) => minus4A_s_36_port, 
                           minus4A_out(35) => minus4A_s_35_port, 
                           minus4A_out(34) => minus4A_s_34_port, 
                           minus4A_out(33) => minus4A_s_33_port, 
                           minus4A_out(32) => minus4A_s_32_port, 
                           minus4A_out(31) => minus4A_s_31_port, 
                           minus4A_out(30) => minus4A_s_30_port, 
                           minus4A_out(29) => minus4A_s_29_port, 
                           minus4A_out(28) => minus4A_s_28_port, 
                           minus4A_out(27) => minus4A_s_27_port, 
                           minus4A_out(26) => minus4A_s_26_port, 
                           minus4A_out(25) => minus4A_s_25_port, 
                           minus4A_out(24) => minus4A_s_24_port, 
                           minus4A_out(23) => minus4A_s_23_port, 
                           minus4A_out(22) => minus4A_s_22_port, 
                           minus4A_out(21) => minus4A_s_21_port, 
                           minus4A_out(20) => minus4A_s_20_port, 
                           minus4A_out(19) => minus4A_s_19_port, 
                           minus4A_out(18) => minus4A_s_18_port, 
                           minus4A_out(17) => minus4A_s_17_port, 
                           minus4A_out(16) => minus4A_s_16_port, 
                           minus4A_out(15) => minus4A_s_15_port, 
                           minus4A_out(14) => minus4A_s_14_port, 
                           minus4A_out(13) => minus4A_s_13_port, 
                           minus4A_out(12) => minus4A_s_12_port, 
                           minus4A_out(11) => minus4A_s_11_port, 
                           minus4A_out(10) => minus4A_s_10_port, minus4A_out(9)
                           => minus4A_s_9_port, minus4A_out(8) => 
                           minus4A_s_8_port, minus4A_out(7) => minus4A_s_7_port
                           , minus4A_out(6) => minus4A_s_6_port, minus4A_out(5)
                           => minus4A_s_5_port, minus4A_out(4) => 
                           minus4A_s_4_port, minus4A_out(3) => minus4A_s_3_port
                           , minus4A_out(2) => minus4A_s_2_port, minus4A_out(1)
                           => minus4A_s_1_port, minus4A_out(0) => 
                           minus4A_s_0_port);
   mux_1 : MUX_GENERIC_N64_RADIX3_2 port map( plusA(63) => plus2A_s_63_port, 
                           plusA(62) => plus2A_s_62_port, plusA(61) => 
                           plus2A_s_61_port, plusA(60) => plus2A_s_60_port, 
                           plusA(59) => plus2A_s_59_port, plusA(58) => 
                           plus2A_s_58_port, plusA(57) => plus2A_s_57_port, 
                           plusA(56) => plus2A_s_56_port, plusA(55) => 
                           plus2A_s_55_port, plusA(54) => plus2A_s_54_port, 
                           plusA(53) => plus2A_s_53_port, plusA(52) => 
                           plus2A_s_52_port, plusA(51) => plus2A_s_51_port, 
                           plusA(50) => plus2A_s_50_port, plusA(49) => 
                           plus2A_s_49_port, plusA(48) => plus2A_s_48_port, 
                           plusA(47) => plus2A_s_47_port, plusA(46) => 
                           plus2A_s_46_port, plusA(45) => plus2A_s_45_port, 
                           plusA(44) => plus2A_s_44_port, plusA(43) => 
                           plus2A_s_43_port, plusA(42) => plus2A_s_42_port, 
                           plusA(41) => plus2A_s_41_port, plusA(40) => 
                           plus2A_s_40_port, plusA(39) => plus2A_s_39_port, 
                           plusA(38) => plus2A_s_38_port, plusA(37) => 
                           plus2A_s_37_port, plusA(36) => plus2A_s_36_port, 
                           plusA(35) => plus2A_s_35_port, plusA(34) => 
                           plus2A_s_34_port, plusA(33) => plus2A_s_33_port, 
                           plusA(32) => plus2A_s_32_port, plusA(31) => 
                           plus2A_s_31_port, plusA(30) => plus2A_s_30_port, 
                           plusA(29) => plus2A_s_29_port, plusA(28) => 
                           plus2A_s_28_port, plusA(27) => plus2A_s_27_port, 
                           plusA(26) => plus2A_s_26_port, plusA(25) => 
                           plus2A_s_25_port, plusA(24) => plus2A_s_24_port, 
                           plusA(23) => plus2A_s_23_port, plusA(22) => 
                           plus2A_s_22_port, plusA(21) => plus2A_s_21_port, 
                           plusA(20) => plus2A_s_20_port, plusA(19) => 
                           plus2A_s_19_port, plusA(18) => plus2A_s_18_port, 
                           plusA(17) => plus2A_s_17_port, plusA(16) => 
                           plus2A_s_16_port, plusA(15) => plus2A_s_15_port, 
                           plusA(14) => plus2A_s_14_port, plusA(13) => 
                           plus2A_s_13_port, plusA(12) => plus2A_s_12_port, 
                           plusA(11) => plus2A_s_11_port, plusA(10) => 
                           plus2A_s_10_port, plusA(9) => plus2A_s_9_port, 
                           plusA(8) => plus2A_s_8_port, plusA(7) => 
                           plus2A_s_7_port, plusA(6) => plus2A_s_6_port, 
                           plusA(5) => plus2A_s_5_port, plusA(4) => 
                           plus2A_s_4_port, plusA(3) => plus2A_s_3_port, 
                           plusA(2) => plus2A_s_2_port, plusA(1) => 
                           plus2A_s_1_port, plusA(0) => nextA_0_port, 
                           minusA(63) => minus2A_s_63_port, minusA(62) => 
                           minus2A_s_62_port, minusA(61) => minus2A_s_61_port, 
                           minusA(60) => minus2A_s_60_port, minusA(59) => 
                           minus2A_s_59_port, minusA(58) => minus2A_s_58_port, 
                           minusA(57) => minus2A_s_57_port, minusA(56) => 
                           minus2A_s_56_port, minusA(55) => minus2A_s_55_port, 
                           minusA(54) => minus2A_s_54_port, minusA(53) => 
                           minus2A_s_53_port, minusA(52) => minus2A_s_52_port, 
                           minusA(51) => minus2A_s_51_port, minusA(50) => 
                           minus2A_s_50_port, minusA(49) => minus2A_s_49_port, 
                           minusA(48) => minus2A_s_48_port, minusA(47) => 
                           minus2A_s_47_port, minusA(46) => minus2A_s_46_port, 
                           minusA(45) => minus2A_s_45_port, minusA(44) => 
                           minus2A_s_44_port, minusA(43) => minus2A_s_43_port, 
                           minusA(42) => minus2A_s_42_port, minusA(41) => 
                           minus2A_s_41_port, minusA(40) => minus2A_s_40_port, 
                           minusA(39) => minus2A_s_39_port, minusA(38) => 
                           minus2A_s_38_port, minusA(37) => minus2A_s_37_port, 
                           minusA(36) => minus2A_s_36_port, minusA(35) => 
                           minus2A_s_35_port, minusA(34) => minus2A_s_34_port, 
                           minusA(33) => minus2A_s_33_port, minusA(32) => 
                           minus2A_s_32_port, minusA(31) => minus2A_s_31_port, 
                           minusA(30) => minus2A_s_30_port, minusA(29) => 
                           minus2A_s_29_port, minusA(28) => minus2A_s_28_port, 
                           minusA(27) => minus2A_s_27_port, minusA(26) => 
                           minus2A_s_26_port, minusA(25) => minus2A_s_25_port, 
                           minusA(24) => minus2A_s_24_port, minusA(23) => 
                           minus2A_s_23_port, minusA(22) => minus2A_s_22_port, 
                           minusA(21) => minus2A_s_21_port, minusA(20) => 
                           minus2A_s_20_port, minusA(19) => minus2A_s_19_port, 
                           minusA(18) => minus2A_s_18_port, minusA(17) => 
                           minus2A_s_17_port, minusA(16) => minus2A_s_16_port, 
                           minusA(15) => minus2A_s_15_port, minusA(14) => 
                           minus2A_s_14_port, minusA(13) => minus2A_s_13_port, 
                           minusA(12) => minus2A_s_12_port, minusA(11) => 
                           minus2A_s_11_port, minusA(10) => minus2A_s_10_port, 
                           minusA(9) => minus2A_s_9_port, minusA(8) => 
                           minus2A_s_8_port, minusA(7) => minus2A_s_7_port, 
                           minusA(6) => minus2A_s_6_port, minusA(5) => 
                           minus2A_s_5_port, minusA(4) => minus2A_s_4_port, 
                           minusA(3) => minus2A_s_3_port, minusA(2) => 
                           minus2A_s_2_port, minusA(1) => minus2A_s_1_port, 
                           minusA(0) => minus2A_s_0_port, plus2A(63) => 
                           nextA_63_port, plus2A(62) => nextA_62_port, 
                           plus2A(61) => nextA_61_port, plus2A(60) => 
                           nextA_60_port, plus2A(59) => nextA_59_port, 
                           plus2A(58) => nextA_58_port, plus2A(57) => 
                           nextA_57_port, plus2A(56) => nextA_56_port, 
                           plus2A(55) => nextA_55_port, plus2A(54) => 
                           nextA_54_port, plus2A(53) => nextA_53_port, 
                           plus2A(52) => nextA_52_port, plus2A(51) => 
                           nextA_51_port, plus2A(50) => nextA_50_port, 
                           plus2A(49) => nextA_49_port, plus2A(48) => 
                           nextA_48_port, plus2A(47) => nextA_47_port, 
                           plus2A(46) => nextA_46_port, plus2A(45) => 
                           nextA_45_port, plus2A(44) => nextA_44_port, 
                           plus2A(43) => nextA_43_port, plus2A(42) => 
                           nextA_42_port, plus2A(41) => nextA_41_port, 
                           plus2A(40) => nextA_40_port, plus2A(39) => 
                           nextA_39_port, plus2A(38) => nextA_38_port, 
                           plus2A(37) => nextA_37_port, plus2A(36) => 
                           nextA_36_port, plus2A(35) => nextA_35_port, 
                           plus2A(34) => nextA_34_port, plus2A(33) => 
                           nextA_33_port, plus2A(32) => nextA_32_port, 
                           plus2A(31) => nextA_31_port, plus2A(30) => 
                           nextA_30_port, plus2A(29) => nextA_29_port, 
                           plus2A(28) => nextA_28_port, plus2A(27) => 
                           nextA_27_port, plus2A(26) => nextA_26_port, 
                           plus2A(25) => nextA_25_port, plus2A(24) => 
                           nextA_24_port, plus2A(23) => nextA_23_port, 
                           plus2A(22) => nextA_22_port, plus2A(21) => 
                           nextA_21_port, plus2A(20) => nextA_20_port, 
                           plus2A(19) => nextA_19_port, plus2A(18) => 
                           nextA_18_port, plus2A(17) => nextA_17_port, 
                           plus2A(16) => nextA_16_port, plus2A(15) => 
                           nextA_15_port, plus2A(14) => nextA_14_port, 
                           plus2A(13) => nextA_13_port, plus2A(12) => 
                           nextA_12_port, plus2A(11) => nextA_11_port, 
                           plus2A(10) => nextA_10_port, plus2A(9) => 
                           nextA_9_port, plus2A(8) => nextA_8_port, plus2A(7) 
                           => nextA_7_port, plus2A(6) => nextA_6_port, 
                           plus2A(5) => nextA_5_port, plus2A(4) => nextA_4_port
                           , plus2A(3) => nextA_3_port, plus2A(2) => 
                           nextA_2_port, plus2A(1) => nextA_1_port, plus2A(0) 
                           => nextA_0_port, minus2A(63) => minus4A_s_63_port, 
                           minus2A(62) => minus4A_s_62_port, minus2A(61) => 
                           minus4A_s_61_port, minus2A(60) => minus4A_s_60_port,
                           minus2A(59) => minus4A_s_59_port, minus2A(58) => 
                           minus4A_s_58_port, minus2A(57) => minus4A_s_57_port,
                           minus2A(56) => minus4A_s_56_port, minus2A(55) => 
                           minus4A_s_55_port, minus2A(54) => minus4A_s_54_port,
                           minus2A(53) => minus4A_s_53_port, minus2A(52) => 
                           minus4A_s_52_port, minus2A(51) => minus4A_s_51_port,
                           minus2A(50) => minus4A_s_50_port, minus2A(49) => 
                           minus4A_s_49_port, minus2A(48) => minus4A_s_48_port,
                           minus2A(47) => minus4A_s_47_port, minus2A(46) => 
                           minus4A_s_46_port, minus2A(45) => minus4A_s_45_port,
                           minus2A(44) => minus4A_s_44_port, minus2A(43) => 
                           minus4A_s_43_port, minus2A(42) => minus4A_s_42_port,
                           minus2A(41) => minus4A_s_41_port, minus2A(40) => 
                           minus4A_s_40_port, minus2A(39) => minus4A_s_39_port,
                           minus2A(38) => minus4A_s_38_port, minus2A(37) => 
                           minus4A_s_37_port, minus2A(36) => minus4A_s_36_port,
                           minus2A(35) => minus4A_s_35_port, minus2A(34) => 
                           minus4A_s_34_port, minus2A(33) => minus4A_s_33_port,
                           minus2A(32) => minus4A_s_32_port, minus2A(31) => 
                           minus4A_s_31_port, minus2A(30) => minus4A_s_30_port,
                           minus2A(29) => minus4A_s_29_port, minus2A(28) => 
                           minus4A_s_28_port, minus2A(27) => minus4A_s_27_port,
                           minus2A(26) => minus4A_s_26_port, minus2A(25) => 
                           minus4A_s_25_port, minus2A(24) => minus4A_s_24_port,
                           minus2A(23) => minus4A_s_23_port, minus2A(22) => 
                           minus4A_s_22_port, minus2A(21) => minus4A_s_21_port,
                           minus2A(20) => minus4A_s_20_port, minus2A(19) => 
                           minus4A_s_19_port, minus2A(18) => minus4A_s_18_port,
                           minus2A(17) => minus4A_s_17_port, minus2A(16) => 
                           minus4A_s_16_port, minus2A(15) => minus4A_s_15_port,
                           minus2A(14) => minus4A_s_14_port, minus2A(13) => 
                           minus4A_s_13_port, minus2A(12) => minus4A_s_12_port,
                           minus2A(11) => minus4A_s_11_port, minus2A(10) => 
                           minus4A_s_10_port, minus2A(9) => minus4A_s_9_port, 
                           minus2A(8) => minus4A_s_8_port, minus2A(7) => 
                           minus4A_s_7_port, minus2A(6) => minus4A_s_6_port, 
                           minus2A(5) => minus4A_s_5_port, minus2A(4) => 
                           minus4A_s_4_port, minus2A(3) => minus4A_s_3_port, 
                           minus2A(2) => minus4A_s_2_port, minus2A(1) => 
                           minus4A_s_1_port, minus2A(0) => minus4A_s_0_port, 
                           SEL(2) => encoder_to_mux_2_port, SEL(1) => 
                           encoder_to_mux_1_port, SEL(0) => 
                           encoder_to_mux_0_port, Y(63) => mux_to_adder_63_port
                           , Y(62) => mux_to_adder_62_port, Y(61) => 
                           mux_to_adder_61_port, Y(60) => mux_to_adder_60_port,
                           Y(59) => mux_to_adder_59_port, Y(58) => 
                           mux_to_adder_58_port, Y(57) => mux_to_adder_57_port,
                           Y(56) => mux_to_adder_56_port, Y(55) => 
                           mux_to_adder_55_port, Y(54) => mux_to_adder_54_port,
                           Y(53) => mux_to_adder_53_port, Y(52) => 
                           mux_to_adder_52_port, Y(51) => mux_to_adder_51_port,
                           Y(50) => mux_to_adder_50_port, Y(49) => 
                           mux_to_adder_49_port, Y(48) => mux_to_adder_48_port,
                           Y(47) => mux_to_adder_47_port, Y(46) => 
                           mux_to_adder_46_port, Y(45) => mux_to_adder_45_port,
                           Y(44) => mux_to_adder_44_port, Y(43) => 
                           mux_to_adder_43_port, Y(42) => mux_to_adder_42_port,
                           Y(41) => mux_to_adder_41_port, Y(40) => 
                           mux_to_adder_40_port, Y(39) => mux_to_adder_39_port,
                           Y(38) => mux_to_adder_38_port, Y(37) => 
                           mux_to_adder_37_port, Y(36) => mux_to_adder_36_port,
                           Y(35) => mux_to_adder_35_port, Y(34) => 
                           mux_to_adder_34_port, Y(33) => mux_to_adder_33_port,
                           Y(32) => mux_to_adder_32_port, Y(31) => 
                           mux_to_adder_31_port, Y(30) => mux_to_adder_30_port,
                           Y(29) => mux_to_adder_29_port, Y(28) => 
                           mux_to_adder_28_port, Y(27) => mux_to_adder_27_port,
                           Y(26) => mux_to_adder_26_port, Y(25) => 
                           mux_to_adder_25_port, Y(24) => mux_to_adder_24_port,
                           Y(23) => mux_to_adder_23_port, Y(22) => 
                           mux_to_adder_22_port, Y(21) => mux_to_adder_21_port,
                           Y(20) => mux_to_adder_20_port, Y(19) => 
                           mux_to_adder_19_port, Y(18) => mux_to_adder_18_port,
                           Y(17) => mux_to_adder_17_port, Y(16) => 
                           mux_to_adder_16_port, Y(15) => mux_to_adder_15_port,
                           Y(14) => mux_to_adder_14_port, Y(13) => 
                           mux_to_adder_13_port, Y(12) => mux_to_adder_12_port,
                           Y(11) => mux_to_adder_11_port, Y(10) => 
                           mux_to_adder_10_port, Y(9) => mux_to_adder_9_port, 
                           Y(8) => mux_to_adder_8_port, Y(7) => 
                           mux_to_adder_7_port, Y(6) => mux_to_adder_6_port, 
                           Y(5) => mux_to_adder_5_port, Y(4) => 
                           mux_to_adder_4_port, Y(3) => mux_to_adder_3_port, 
                           Y(2) => mux_to_adder_2_port, Y(1) => 
                           mux_to_adder_1_port, Y(0) => mux_to_adder_0_port);
   rca_1 : RCA_N64_2 port map( A(63) => mux_to_adder_63_port, A(62) => 
                           mux_to_adder_62_port, A(61) => mux_to_adder_61_port,
                           A(60) => mux_to_adder_60_port, A(59) => 
                           mux_to_adder_59_port, A(58) => mux_to_adder_58_port,
                           A(57) => mux_to_adder_57_port, A(56) => 
                           mux_to_adder_56_port, A(55) => mux_to_adder_55_port,
                           A(54) => mux_to_adder_54_port, A(53) => 
                           mux_to_adder_53_port, A(52) => mux_to_adder_52_port,
                           A(51) => mux_to_adder_51_port, A(50) => 
                           mux_to_adder_50_port, A(49) => mux_to_adder_49_port,
                           A(48) => mux_to_adder_48_port, A(47) => 
                           mux_to_adder_47_port, A(46) => mux_to_adder_46_port,
                           A(45) => mux_to_adder_45_port, A(44) => 
                           mux_to_adder_44_port, A(43) => mux_to_adder_43_port,
                           A(42) => mux_to_adder_42_port, A(41) => 
                           mux_to_adder_41_port, A(40) => mux_to_adder_40_port,
                           A(39) => mux_to_adder_39_port, A(38) => 
                           mux_to_adder_38_port, A(37) => mux_to_adder_37_port,
                           A(36) => mux_to_adder_36_port, A(35) => 
                           mux_to_adder_35_port, A(34) => mux_to_adder_34_port,
                           A(33) => mux_to_adder_33_port, A(32) => 
                           mux_to_adder_32_port, A(31) => mux_to_adder_31_port,
                           A(30) => mux_to_adder_30_port, A(29) => 
                           mux_to_adder_29_port, A(28) => mux_to_adder_28_port,
                           A(27) => mux_to_adder_27_port, A(26) => 
                           mux_to_adder_26_port, A(25) => mux_to_adder_25_port,
                           A(24) => mux_to_adder_24_port, A(23) => 
                           mux_to_adder_23_port, A(22) => mux_to_adder_22_port,
                           A(21) => mux_to_adder_21_port, A(20) => 
                           mux_to_adder_20_port, A(19) => mux_to_adder_19_port,
                           A(18) => mux_to_adder_18_port, A(17) => 
                           mux_to_adder_17_port, A(16) => mux_to_adder_16_port,
                           A(15) => mux_to_adder_15_port, A(14) => 
                           mux_to_adder_14_port, A(13) => mux_to_adder_13_port,
                           A(12) => mux_to_adder_12_port, A(11) => 
                           mux_to_adder_11_port, A(10) => mux_to_adder_10_port,
                           A(9) => mux_to_adder_9_port, A(8) => 
                           mux_to_adder_8_port, A(7) => mux_to_adder_7_port, 
                           A(6) => mux_to_adder_6_port, A(5) => 
                           mux_to_adder_5_port, A(4) => mux_to_adder_4_port, 
                           A(3) => mux_to_adder_3_port, A(2) => 
                           mux_to_adder_2_port, A(1) => mux_to_adder_1_port, 
                           A(0) => mux_to_adder_0_port, B(63) => prevSum(63), 
                           B(62) => prevSum(62), B(61) => prevSum(61), B(60) =>
                           prevSum(60), B(59) => prevSum(59), B(58) => 
                           prevSum(58), B(57) => prevSum(57), B(56) => 
                           prevSum(56), B(55) => prevSum(55), B(54) => 
                           prevSum(54), B(53) => prevSum(53), B(52) => 
                           prevSum(52), B(51) => prevSum(51), B(50) => 
                           prevSum(50), B(49) => prevSum(49), B(48) => 
                           prevSum(48), B(47) => prevSum(47), B(46) => 
                           prevSum(46), B(45) => prevSum(45), B(44) => 
                           prevSum(44), B(43) => prevSum(43), B(42) => 
                           prevSum(42), B(41) => prevSum(41), B(40) => 
                           prevSum(40), B(39) => prevSum(39), B(38) => 
                           prevSum(38), B(37) => prevSum(37), B(36) => 
                           prevSum(36), B(35) => prevSum(35), B(34) => 
                           prevSum(34), B(33) => prevSum(33), B(32) => 
                           prevSum(32), B(31) => prevSum(31), B(30) => 
                           prevSum(30), B(29) => prevSum(29), B(28) => 
                           prevSum(28), B(27) => prevSum(27), B(26) => 
                           prevSum(26), B(25) => prevSum(25), B(24) => 
                           prevSum(24), B(23) => prevSum(23), B(22) => 
                           prevSum(22), B(21) => prevSum(21), B(20) => 
                           prevSum(20), B(19) => prevSum(19), B(18) => 
                           prevSum(18), B(17) => prevSum(17), B(16) => 
                           prevSum(16), B(15) => prevSum(15), B(14) => 
                           prevSum(14), B(13) => prevSum(13), B(12) => 
                           prevSum(12), B(11) => prevSum(11), B(10) => 
                           prevSum(10), B(9) => prevSum(9), B(8) => prevSum(8),
                           B(7) => prevSum(7), B(6) => prevSum(6), B(5) => 
                           prevSum(5), B(4) => prevSum(4), B(3) => prevSum(3), 
                           B(2) => prevSum(2), B(1) => prevSum(1), B(0) => 
                           prevSum(0), Ci => X_Logic0_port, S(63) => 
                           nextSum(63), S(62) => nextSum(62), S(61) => 
                           nextSum(61), S(60) => nextSum(60), S(59) => 
                           nextSum(59), S(58) => nextSum(58), S(57) => 
                           nextSum(57), S(56) => nextSum(56), S(55) => 
                           nextSum(55), S(54) => nextSum(54), S(53) => 
                           nextSum(53), S(52) => nextSum(52), S(51) => 
                           nextSum(51), S(50) => nextSum(50), S(49) => 
                           nextSum(49), S(48) => nextSum(48), S(47) => 
                           nextSum(47), S(46) => nextSum(46), S(45) => 
                           nextSum(45), S(44) => nextSum(44), S(43) => 
                           nextSum(43), S(42) => nextSum(42), S(41) => 
                           nextSum(41), S(40) => nextSum(40), S(39) => 
                           nextSum(39), S(38) => nextSum(38), S(37) => 
                           nextSum(37), S(36) => nextSum(36), S(35) => 
                           nextSum(35), S(34) => nextSum(34), S(33) => 
                           nextSum(33), S(32) => nextSum(32), S(31) => 
                           nextSum(31), S(30) => nextSum(30), S(29) => 
                           nextSum(29), S(28) => nextSum(28), S(27) => 
                           nextSum(27), S(26) => nextSum(26), S(25) => 
                           nextSum(25), S(24) => nextSum(24), S(23) => 
                           nextSum(23), S(22) => nextSum(22), S(21) => 
                           nextSum(21), S(20) => nextSum(20), S(19) => 
                           nextSum(19), S(18) => nextSum(18), S(17) => 
                           nextSum(17), S(16) => nextSum(16), S(15) => 
                           nextSum(15), S(14) => nextSum(14), S(13) => 
                           nextSum(13), S(12) => nextSum(12), S(11) => 
                           nextSum(11), S(10) => nextSum(10), S(9) => 
                           nextSum(9), S(8) => nextSum(8), S(7) => nextSum(7), 
                           S(6) => nextSum(6), S(5) => nextSum(5), S(4) => 
                           nextSum(4), S(3) => nextSum(3), S(2) => nextSum(2), 
                           S(1) => nextSum(1), S(0) => nextSum(0), Co => n_3180
                           );

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity booth_mul_row_N64_RADIX3_3 is

   port( prevA, prevSum : in std_logic_vector (63 downto 0);  encoderIn : in 
         std_logic_vector (2 downto 0);  nextA, nextSum : out std_logic_vector 
         (63 downto 0));

end booth_mul_row_N64_RADIX3_3;

architecture SYN_struct of booth_mul_row_N64_RADIX3_3 is

   component RCA_N64_3
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component MUX_GENERIC_N64_RADIX3_3
      port( plusA, minusA, plus2A, minus2A : in std_logic_vector (63 downto 0);
            SEL : in std_logic_vector (2 downto 0);  Y : out std_logic_vector 
            (63 downto 0));
   end component;
   
   component ShiftnCompl_N64_3
      port( plusA : in std_logic_vector (63 downto 0);  plus2A_out, minus2A_out
            , plus4A_out, minus4A_out : out std_logic_vector (63 downto 0));
   end component;
   
   component encoder_N64_RADIX3_3
      port( X : in std_logic_vector (2 downto 0);  Z : out std_logic_vector (2 
            downto 0));
   end component;
   
   signal X_Logic0_port, nextA_63_port, nextA_62_port, nextA_61_port, 
      nextA_60_port, nextA_59_port, nextA_58_port, nextA_57_port, nextA_56_port
      , nextA_55_port, nextA_54_port, nextA_53_port, nextA_52_port, 
      nextA_51_port, nextA_50_port, nextA_49_port, nextA_48_port, nextA_47_port
      , nextA_46_port, nextA_45_port, nextA_44_port, nextA_43_port, 
      nextA_42_port, nextA_41_port, nextA_40_port, nextA_39_port, nextA_38_port
      , nextA_37_port, nextA_36_port, nextA_35_port, nextA_34_port, 
      nextA_33_port, nextA_32_port, nextA_31_port, nextA_30_port, nextA_29_port
      , nextA_28_port, nextA_27_port, nextA_26_port, nextA_25_port, 
      nextA_24_port, nextA_23_port, nextA_22_port, nextA_21_port, nextA_20_port
      , nextA_19_port, nextA_18_port, nextA_17_port, nextA_16_port, 
      nextA_15_port, nextA_14_port, nextA_13_port, nextA_12_port, nextA_11_port
      , nextA_10_port, nextA_9_port, nextA_8_port, nextA_7_port, nextA_6_port, 
      nextA_5_port, nextA_4_port, nextA_3_port, nextA_2_port, nextA_1_port, 
      encoder_to_mux_2_port, encoder_to_mux_1_port, encoder_to_mux_0_port, 
      plus2A_s_63_port, plus2A_s_62_port, plus2A_s_61_port, plus2A_s_60_port, 
      plus2A_s_59_port, plus2A_s_58_port, plus2A_s_57_port, plus2A_s_56_port, 
      plus2A_s_55_port, plus2A_s_54_port, plus2A_s_53_port, plus2A_s_52_port, 
      plus2A_s_51_port, plus2A_s_50_port, plus2A_s_49_port, plus2A_s_48_port, 
      plus2A_s_47_port, plus2A_s_46_port, plus2A_s_45_port, plus2A_s_44_port, 
      plus2A_s_43_port, plus2A_s_42_port, plus2A_s_41_port, plus2A_s_40_port, 
      plus2A_s_39_port, plus2A_s_38_port, plus2A_s_37_port, plus2A_s_36_port, 
      plus2A_s_35_port, plus2A_s_34_port, plus2A_s_33_port, plus2A_s_32_port, 
      plus2A_s_31_port, plus2A_s_30_port, plus2A_s_29_port, plus2A_s_28_port, 
      plus2A_s_27_port, plus2A_s_26_port, plus2A_s_25_port, plus2A_s_24_port, 
      plus2A_s_23_port, plus2A_s_22_port, plus2A_s_21_port, plus2A_s_20_port, 
      plus2A_s_19_port, plus2A_s_18_port, plus2A_s_17_port, plus2A_s_16_port, 
      plus2A_s_15_port, plus2A_s_14_port, plus2A_s_13_port, plus2A_s_12_port, 
      plus2A_s_11_port, plus2A_s_10_port, plus2A_s_9_port, plus2A_s_8_port, 
      plus2A_s_7_port, plus2A_s_6_port, plus2A_s_5_port, plus2A_s_4_port, 
      plus2A_s_3_port, plus2A_s_2_port, plus2A_s_1_port, minus2A_s_63_port, 
      minus2A_s_62_port, minus2A_s_61_port, minus2A_s_60_port, 
      minus2A_s_59_port, minus2A_s_58_port, minus2A_s_57_port, 
      minus2A_s_56_port, minus2A_s_55_port, minus2A_s_54_port, 
      minus2A_s_53_port, minus2A_s_52_port, minus2A_s_51_port, 
      minus2A_s_50_port, minus2A_s_49_port, minus2A_s_48_port, 
      minus2A_s_47_port, minus2A_s_46_port, minus2A_s_45_port, 
      minus2A_s_44_port, minus2A_s_43_port, minus2A_s_42_port, 
      minus2A_s_41_port, minus2A_s_40_port, minus2A_s_39_port, 
      minus2A_s_38_port, minus2A_s_37_port, minus2A_s_36_port, 
      minus2A_s_35_port, minus2A_s_34_port, minus2A_s_33_port, 
      minus2A_s_32_port, minus2A_s_31_port, minus2A_s_30_port, 
      minus2A_s_29_port, minus2A_s_28_port, minus2A_s_27_port, 
      minus2A_s_26_port, minus2A_s_25_port, minus2A_s_24_port, 
      minus2A_s_23_port, minus2A_s_22_port, minus2A_s_21_port, 
      minus2A_s_20_port, minus2A_s_19_port, minus2A_s_18_port, 
      minus2A_s_17_port, minus2A_s_16_port, minus2A_s_15_port, 
      minus2A_s_14_port, minus2A_s_13_port, minus2A_s_12_port, 
      minus2A_s_11_port, minus2A_s_10_port, minus2A_s_9_port, minus2A_s_8_port,
      minus2A_s_7_port, minus2A_s_6_port, minus2A_s_5_port, minus2A_s_4_port, 
      minus2A_s_3_port, minus2A_s_2_port, minus2A_s_1_port, minus2A_s_0_port, 
      minus4A_s_63_port, minus4A_s_62_port, minus4A_s_61_port, 
      minus4A_s_60_port, minus4A_s_59_port, minus4A_s_58_port, 
      minus4A_s_57_port, minus4A_s_56_port, minus4A_s_55_port, 
      minus4A_s_54_port, minus4A_s_53_port, minus4A_s_52_port, 
      minus4A_s_51_port, minus4A_s_50_port, minus4A_s_49_port, 
      minus4A_s_48_port, minus4A_s_47_port, minus4A_s_46_port, 
      minus4A_s_45_port, minus4A_s_44_port, minus4A_s_43_port, 
      minus4A_s_42_port, minus4A_s_41_port, minus4A_s_40_port, 
      minus4A_s_39_port, minus4A_s_38_port, minus4A_s_37_port, 
      minus4A_s_36_port, minus4A_s_35_port, minus4A_s_34_port, 
      minus4A_s_33_port, minus4A_s_32_port, minus4A_s_31_port, 
      minus4A_s_30_port, minus4A_s_29_port, minus4A_s_28_port, 
      minus4A_s_27_port, minus4A_s_26_port, minus4A_s_25_port, 
      minus4A_s_24_port, minus4A_s_23_port, minus4A_s_22_port, 
      minus4A_s_21_port, minus4A_s_20_port, minus4A_s_19_port, 
      minus4A_s_18_port, minus4A_s_17_port, minus4A_s_16_port, 
      minus4A_s_15_port, minus4A_s_14_port, minus4A_s_13_port, 
      minus4A_s_12_port, minus4A_s_11_port, minus4A_s_10_port, minus4A_s_9_port
      , minus4A_s_8_port, minus4A_s_7_port, minus4A_s_6_port, minus4A_s_5_port,
      minus4A_s_4_port, minus4A_s_3_port, minus4A_s_2_port, minus4A_s_1_port, 
      minus4A_s_0_port, mux_to_adder_63_port, mux_to_adder_62_port, 
      mux_to_adder_61_port, mux_to_adder_60_port, mux_to_adder_59_port, 
      mux_to_adder_58_port, mux_to_adder_57_port, mux_to_adder_56_port, 
      mux_to_adder_55_port, mux_to_adder_54_port, mux_to_adder_53_port, 
      mux_to_adder_52_port, mux_to_adder_51_port, mux_to_adder_50_port, 
      mux_to_adder_49_port, mux_to_adder_48_port, mux_to_adder_47_port, 
      mux_to_adder_46_port, mux_to_adder_45_port, mux_to_adder_44_port, 
      mux_to_adder_43_port, mux_to_adder_42_port, mux_to_adder_41_port, 
      mux_to_adder_40_port, mux_to_adder_39_port, mux_to_adder_38_port, 
      mux_to_adder_37_port, mux_to_adder_36_port, mux_to_adder_35_port, 
      mux_to_adder_34_port, mux_to_adder_33_port, mux_to_adder_32_port, 
      mux_to_adder_31_port, mux_to_adder_30_port, mux_to_adder_29_port, 
      mux_to_adder_28_port, mux_to_adder_27_port, mux_to_adder_26_port, 
      mux_to_adder_25_port, mux_to_adder_24_port, mux_to_adder_23_port, 
      mux_to_adder_22_port, mux_to_adder_21_port, mux_to_adder_20_port, 
      mux_to_adder_19_port, mux_to_adder_18_port, mux_to_adder_17_port, 
      mux_to_adder_16_port, mux_to_adder_15_port, mux_to_adder_14_port, 
      mux_to_adder_13_port, mux_to_adder_12_port, mux_to_adder_11_port, 
      mux_to_adder_10_port, mux_to_adder_9_port, mux_to_adder_8_port, 
      mux_to_adder_7_port, mux_to_adder_6_port, mux_to_adder_5_port, 
      mux_to_adder_4_port, mux_to_adder_3_port, mux_to_adder_2_port, 
      mux_to_adder_1_port, mux_to_adder_0_port, nextA_0_port, n_3181, n_3182, 
      n_3183 : std_logic;

begin
   nextA <= ( nextA_63_port, nextA_62_port, nextA_61_port, nextA_60_port, 
      nextA_59_port, nextA_58_port, nextA_57_port, nextA_56_port, nextA_55_port
      , nextA_54_port, nextA_53_port, nextA_52_port, nextA_51_port, 
      nextA_50_port, nextA_49_port, nextA_48_port, nextA_47_port, nextA_46_port
      , nextA_45_port, nextA_44_port, nextA_43_port, nextA_42_port, 
      nextA_41_port, nextA_40_port, nextA_39_port, nextA_38_port, nextA_37_port
      , nextA_36_port, nextA_35_port, nextA_34_port, nextA_33_port, 
      nextA_32_port, nextA_31_port, nextA_30_port, nextA_29_port, nextA_28_port
      , nextA_27_port, nextA_26_port, nextA_25_port, nextA_24_port, 
      nextA_23_port, nextA_22_port, nextA_21_port, nextA_20_port, nextA_19_port
      , nextA_18_port, nextA_17_port, nextA_16_port, nextA_15_port, 
      nextA_14_port, nextA_13_port, nextA_12_port, nextA_11_port, nextA_10_port
      , nextA_9_port, nextA_8_port, nextA_7_port, nextA_6_port, nextA_5_port, 
      nextA_4_port, nextA_3_port, nextA_2_port, nextA_1_port, nextA_0_port );
   
   X_Logic0_port <= '0';
   nextA_0_port <= '0';
   encoder_1 : encoder_N64_RADIX3_3 port map( X(2) => encoderIn(2), X(1) => 
                           encoderIn(1), X(0) => encoderIn(0), Z(2) => 
                           encoder_to_mux_2_port, Z(1) => encoder_to_mux_1_port
                           , Z(0) => encoder_to_mux_0_port);
   ShiftnCompl_1 : ShiftnCompl_N64_3 port map( plusA(63) => prevA(63), 
                           plusA(62) => prevA(62), plusA(61) => prevA(61), 
                           plusA(60) => prevA(60), plusA(59) => prevA(59), 
                           plusA(58) => prevA(58), plusA(57) => prevA(57), 
                           plusA(56) => prevA(56), plusA(55) => prevA(55), 
                           plusA(54) => prevA(54), plusA(53) => prevA(53), 
                           plusA(52) => prevA(52), plusA(51) => prevA(51), 
                           plusA(50) => prevA(50), plusA(49) => prevA(49), 
                           plusA(48) => prevA(48), plusA(47) => prevA(47), 
                           plusA(46) => prevA(46), plusA(45) => prevA(45), 
                           plusA(44) => prevA(44), plusA(43) => prevA(43), 
                           plusA(42) => prevA(42), plusA(41) => prevA(41), 
                           plusA(40) => prevA(40), plusA(39) => prevA(39), 
                           plusA(38) => prevA(38), plusA(37) => prevA(37), 
                           plusA(36) => prevA(36), plusA(35) => prevA(35), 
                           plusA(34) => prevA(34), plusA(33) => prevA(33), 
                           plusA(32) => prevA(32), plusA(31) => prevA(31), 
                           plusA(30) => prevA(30), plusA(29) => prevA(29), 
                           plusA(28) => prevA(28), plusA(27) => prevA(27), 
                           plusA(26) => prevA(26), plusA(25) => prevA(25), 
                           plusA(24) => prevA(24), plusA(23) => prevA(23), 
                           plusA(22) => prevA(22), plusA(21) => prevA(21), 
                           plusA(20) => prevA(20), plusA(19) => prevA(19), 
                           plusA(18) => prevA(18), plusA(17) => prevA(17), 
                           plusA(16) => prevA(16), plusA(15) => prevA(15), 
                           plusA(14) => prevA(14), plusA(13) => prevA(13), 
                           plusA(12) => prevA(12), plusA(11) => prevA(11), 
                           plusA(10) => prevA(10), plusA(9) => prevA(9), 
                           plusA(8) => prevA(8), plusA(7) => prevA(7), plusA(6)
                           => prevA(6), plusA(5) => prevA(5), plusA(4) => 
                           prevA(4), plusA(3) => prevA(3), plusA(2) => prevA(2)
                           , plusA(1) => prevA(1), plusA(0) => prevA(0), 
                           plus2A_out(63) => plus2A_s_63_port, plus2A_out(62) 
                           => plus2A_s_62_port, plus2A_out(61) => 
                           plus2A_s_61_port, plus2A_out(60) => plus2A_s_60_port
                           , plus2A_out(59) => plus2A_s_59_port, plus2A_out(58)
                           => plus2A_s_58_port, plus2A_out(57) => 
                           plus2A_s_57_port, plus2A_out(56) => plus2A_s_56_port
                           , plus2A_out(55) => plus2A_s_55_port, plus2A_out(54)
                           => plus2A_s_54_port, plus2A_out(53) => 
                           plus2A_s_53_port, plus2A_out(52) => plus2A_s_52_port
                           , plus2A_out(51) => plus2A_s_51_port, plus2A_out(50)
                           => plus2A_s_50_port, plus2A_out(49) => 
                           plus2A_s_49_port, plus2A_out(48) => plus2A_s_48_port
                           , plus2A_out(47) => plus2A_s_47_port, plus2A_out(46)
                           => plus2A_s_46_port, plus2A_out(45) => 
                           plus2A_s_45_port, plus2A_out(44) => plus2A_s_44_port
                           , plus2A_out(43) => plus2A_s_43_port, plus2A_out(42)
                           => plus2A_s_42_port, plus2A_out(41) => 
                           plus2A_s_41_port, plus2A_out(40) => plus2A_s_40_port
                           , plus2A_out(39) => plus2A_s_39_port, plus2A_out(38)
                           => plus2A_s_38_port, plus2A_out(37) => 
                           plus2A_s_37_port, plus2A_out(36) => plus2A_s_36_port
                           , plus2A_out(35) => plus2A_s_35_port, plus2A_out(34)
                           => plus2A_s_34_port, plus2A_out(33) => 
                           plus2A_s_33_port, plus2A_out(32) => plus2A_s_32_port
                           , plus2A_out(31) => plus2A_s_31_port, plus2A_out(30)
                           => plus2A_s_30_port, plus2A_out(29) => 
                           plus2A_s_29_port, plus2A_out(28) => plus2A_s_28_port
                           , plus2A_out(27) => plus2A_s_27_port, plus2A_out(26)
                           => plus2A_s_26_port, plus2A_out(25) => 
                           plus2A_s_25_port, plus2A_out(24) => plus2A_s_24_port
                           , plus2A_out(23) => plus2A_s_23_port, plus2A_out(22)
                           => plus2A_s_22_port, plus2A_out(21) => 
                           plus2A_s_21_port, plus2A_out(20) => plus2A_s_20_port
                           , plus2A_out(19) => plus2A_s_19_port, plus2A_out(18)
                           => plus2A_s_18_port, plus2A_out(17) => 
                           plus2A_s_17_port, plus2A_out(16) => plus2A_s_16_port
                           , plus2A_out(15) => plus2A_s_15_port, plus2A_out(14)
                           => plus2A_s_14_port, plus2A_out(13) => 
                           plus2A_s_13_port, plus2A_out(12) => plus2A_s_12_port
                           , plus2A_out(11) => plus2A_s_11_port, plus2A_out(10)
                           => plus2A_s_10_port, plus2A_out(9) => 
                           plus2A_s_9_port, plus2A_out(8) => plus2A_s_8_port, 
                           plus2A_out(7) => plus2A_s_7_port, plus2A_out(6) => 
                           plus2A_s_6_port, plus2A_out(5) => plus2A_s_5_port, 
                           plus2A_out(4) => plus2A_s_4_port, plus2A_out(3) => 
                           plus2A_s_3_port, plus2A_out(2) => plus2A_s_2_port, 
                           plus2A_out(1) => plus2A_s_1_port, plus2A_out(0) => 
                           n_3181, minus2A_out(63) => minus2A_s_63_port, 
                           minus2A_out(62) => minus2A_s_62_port, 
                           minus2A_out(61) => minus2A_s_61_port, 
                           minus2A_out(60) => minus2A_s_60_port, 
                           minus2A_out(59) => minus2A_s_59_port, 
                           minus2A_out(58) => minus2A_s_58_port, 
                           minus2A_out(57) => minus2A_s_57_port, 
                           minus2A_out(56) => minus2A_s_56_port, 
                           minus2A_out(55) => minus2A_s_55_port, 
                           minus2A_out(54) => minus2A_s_54_port, 
                           minus2A_out(53) => minus2A_s_53_port, 
                           minus2A_out(52) => minus2A_s_52_port, 
                           minus2A_out(51) => minus2A_s_51_port, 
                           minus2A_out(50) => minus2A_s_50_port, 
                           minus2A_out(49) => minus2A_s_49_port, 
                           minus2A_out(48) => minus2A_s_48_port, 
                           minus2A_out(47) => minus2A_s_47_port, 
                           minus2A_out(46) => minus2A_s_46_port, 
                           minus2A_out(45) => minus2A_s_45_port, 
                           minus2A_out(44) => minus2A_s_44_port, 
                           minus2A_out(43) => minus2A_s_43_port, 
                           minus2A_out(42) => minus2A_s_42_port, 
                           minus2A_out(41) => minus2A_s_41_port, 
                           minus2A_out(40) => minus2A_s_40_port, 
                           minus2A_out(39) => minus2A_s_39_port, 
                           minus2A_out(38) => minus2A_s_38_port, 
                           minus2A_out(37) => minus2A_s_37_port, 
                           minus2A_out(36) => minus2A_s_36_port, 
                           minus2A_out(35) => minus2A_s_35_port, 
                           minus2A_out(34) => minus2A_s_34_port, 
                           minus2A_out(33) => minus2A_s_33_port, 
                           minus2A_out(32) => minus2A_s_32_port, 
                           minus2A_out(31) => minus2A_s_31_port, 
                           minus2A_out(30) => minus2A_s_30_port, 
                           minus2A_out(29) => minus2A_s_29_port, 
                           minus2A_out(28) => minus2A_s_28_port, 
                           minus2A_out(27) => minus2A_s_27_port, 
                           minus2A_out(26) => minus2A_s_26_port, 
                           minus2A_out(25) => minus2A_s_25_port, 
                           minus2A_out(24) => minus2A_s_24_port, 
                           minus2A_out(23) => minus2A_s_23_port, 
                           minus2A_out(22) => minus2A_s_22_port, 
                           minus2A_out(21) => minus2A_s_21_port, 
                           minus2A_out(20) => minus2A_s_20_port, 
                           minus2A_out(19) => minus2A_s_19_port, 
                           minus2A_out(18) => minus2A_s_18_port, 
                           minus2A_out(17) => minus2A_s_17_port, 
                           minus2A_out(16) => minus2A_s_16_port, 
                           minus2A_out(15) => minus2A_s_15_port, 
                           minus2A_out(14) => minus2A_s_14_port, 
                           minus2A_out(13) => minus2A_s_13_port, 
                           minus2A_out(12) => minus2A_s_12_port, 
                           minus2A_out(11) => minus2A_s_11_port, 
                           minus2A_out(10) => minus2A_s_10_port, minus2A_out(9)
                           => minus2A_s_9_port, minus2A_out(8) => 
                           minus2A_s_8_port, minus2A_out(7) => minus2A_s_7_port
                           , minus2A_out(6) => minus2A_s_6_port, minus2A_out(5)
                           => minus2A_s_5_port, minus2A_out(4) => 
                           minus2A_s_4_port, minus2A_out(3) => minus2A_s_3_port
                           , minus2A_out(2) => minus2A_s_2_port, minus2A_out(1)
                           => minus2A_s_1_port, minus2A_out(0) => 
                           minus2A_s_0_port, plus4A_out(63) => nextA_63_port, 
                           plus4A_out(62) => nextA_62_port, plus4A_out(61) => 
                           nextA_61_port, plus4A_out(60) => nextA_60_port, 
                           plus4A_out(59) => nextA_59_port, plus4A_out(58) => 
                           nextA_58_port, plus4A_out(57) => nextA_57_port, 
                           plus4A_out(56) => nextA_56_port, plus4A_out(55) => 
                           nextA_55_port, plus4A_out(54) => nextA_54_port, 
                           plus4A_out(53) => nextA_53_port, plus4A_out(52) => 
                           nextA_52_port, plus4A_out(51) => nextA_51_port, 
                           plus4A_out(50) => nextA_50_port, plus4A_out(49) => 
                           nextA_49_port, plus4A_out(48) => nextA_48_port, 
                           plus4A_out(47) => nextA_47_port, plus4A_out(46) => 
                           nextA_46_port, plus4A_out(45) => nextA_45_port, 
                           plus4A_out(44) => nextA_44_port, plus4A_out(43) => 
                           nextA_43_port, plus4A_out(42) => nextA_42_port, 
                           plus4A_out(41) => nextA_41_port, plus4A_out(40) => 
                           nextA_40_port, plus4A_out(39) => nextA_39_port, 
                           plus4A_out(38) => nextA_38_port, plus4A_out(37) => 
                           nextA_37_port, plus4A_out(36) => nextA_36_port, 
                           plus4A_out(35) => nextA_35_port, plus4A_out(34) => 
                           nextA_34_port, plus4A_out(33) => nextA_33_port, 
                           plus4A_out(32) => nextA_32_port, plus4A_out(31) => 
                           nextA_31_port, plus4A_out(30) => nextA_30_port, 
                           plus4A_out(29) => nextA_29_port, plus4A_out(28) => 
                           nextA_28_port, plus4A_out(27) => nextA_27_port, 
                           plus4A_out(26) => nextA_26_port, plus4A_out(25) => 
                           nextA_25_port, plus4A_out(24) => nextA_24_port, 
                           plus4A_out(23) => nextA_23_port, plus4A_out(22) => 
                           nextA_22_port, plus4A_out(21) => nextA_21_port, 
                           plus4A_out(20) => nextA_20_port, plus4A_out(19) => 
                           nextA_19_port, plus4A_out(18) => nextA_18_port, 
                           plus4A_out(17) => nextA_17_port, plus4A_out(16) => 
                           nextA_16_port, plus4A_out(15) => nextA_15_port, 
                           plus4A_out(14) => nextA_14_port, plus4A_out(13) => 
                           nextA_13_port, plus4A_out(12) => nextA_12_port, 
                           plus4A_out(11) => nextA_11_port, plus4A_out(10) => 
                           nextA_10_port, plus4A_out(9) => nextA_9_port, 
                           plus4A_out(8) => nextA_8_port, plus4A_out(7) => 
                           nextA_7_port, plus4A_out(6) => nextA_6_port, 
                           plus4A_out(5) => nextA_5_port, plus4A_out(4) => 
                           nextA_4_port, plus4A_out(3) => nextA_3_port, 
                           plus4A_out(2) => nextA_2_port, plus4A_out(1) => 
                           nextA_1_port, plus4A_out(0) => n_3182, 
                           minus4A_out(63) => minus4A_s_63_port, 
                           minus4A_out(62) => minus4A_s_62_port, 
                           minus4A_out(61) => minus4A_s_61_port, 
                           minus4A_out(60) => minus4A_s_60_port, 
                           minus4A_out(59) => minus4A_s_59_port, 
                           minus4A_out(58) => minus4A_s_58_port, 
                           minus4A_out(57) => minus4A_s_57_port, 
                           minus4A_out(56) => minus4A_s_56_port, 
                           minus4A_out(55) => minus4A_s_55_port, 
                           minus4A_out(54) => minus4A_s_54_port, 
                           minus4A_out(53) => minus4A_s_53_port, 
                           minus4A_out(52) => minus4A_s_52_port, 
                           minus4A_out(51) => minus4A_s_51_port, 
                           minus4A_out(50) => minus4A_s_50_port, 
                           minus4A_out(49) => minus4A_s_49_port, 
                           minus4A_out(48) => minus4A_s_48_port, 
                           minus4A_out(47) => minus4A_s_47_port, 
                           minus4A_out(46) => minus4A_s_46_port, 
                           minus4A_out(45) => minus4A_s_45_port, 
                           minus4A_out(44) => minus4A_s_44_port, 
                           minus4A_out(43) => minus4A_s_43_port, 
                           minus4A_out(42) => minus4A_s_42_port, 
                           minus4A_out(41) => minus4A_s_41_port, 
                           minus4A_out(40) => minus4A_s_40_port, 
                           minus4A_out(39) => minus4A_s_39_port, 
                           minus4A_out(38) => minus4A_s_38_port, 
                           minus4A_out(37) => minus4A_s_37_port, 
                           minus4A_out(36) => minus4A_s_36_port, 
                           minus4A_out(35) => minus4A_s_35_port, 
                           minus4A_out(34) => minus4A_s_34_port, 
                           minus4A_out(33) => minus4A_s_33_port, 
                           minus4A_out(32) => minus4A_s_32_port, 
                           minus4A_out(31) => minus4A_s_31_port, 
                           minus4A_out(30) => minus4A_s_30_port, 
                           minus4A_out(29) => minus4A_s_29_port, 
                           minus4A_out(28) => minus4A_s_28_port, 
                           minus4A_out(27) => minus4A_s_27_port, 
                           minus4A_out(26) => minus4A_s_26_port, 
                           minus4A_out(25) => minus4A_s_25_port, 
                           minus4A_out(24) => minus4A_s_24_port, 
                           minus4A_out(23) => minus4A_s_23_port, 
                           minus4A_out(22) => minus4A_s_22_port, 
                           minus4A_out(21) => minus4A_s_21_port, 
                           minus4A_out(20) => minus4A_s_20_port, 
                           minus4A_out(19) => minus4A_s_19_port, 
                           minus4A_out(18) => minus4A_s_18_port, 
                           minus4A_out(17) => minus4A_s_17_port, 
                           minus4A_out(16) => minus4A_s_16_port, 
                           minus4A_out(15) => minus4A_s_15_port, 
                           minus4A_out(14) => minus4A_s_14_port, 
                           minus4A_out(13) => minus4A_s_13_port, 
                           minus4A_out(12) => minus4A_s_12_port, 
                           minus4A_out(11) => minus4A_s_11_port, 
                           minus4A_out(10) => minus4A_s_10_port, minus4A_out(9)
                           => minus4A_s_9_port, minus4A_out(8) => 
                           minus4A_s_8_port, minus4A_out(7) => minus4A_s_7_port
                           , minus4A_out(6) => minus4A_s_6_port, minus4A_out(5)
                           => minus4A_s_5_port, minus4A_out(4) => 
                           minus4A_s_4_port, minus4A_out(3) => minus4A_s_3_port
                           , minus4A_out(2) => minus4A_s_2_port, minus4A_out(1)
                           => minus4A_s_1_port, minus4A_out(0) => 
                           minus4A_s_0_port);
   mux_1 : MUX_GENERIC_N64_RADIX3_3 port map( plusA(63) => plus2A_s_63_port, 
                           plusA(62) => plus2A_s_62_port, plusA(61) => 
                           plus2A_s_61_port, plusA(60) => plus2A_s_60_port, 
                           plusA(59) => plus2A_s_59_port, plusA(58) => 
                           plus2A_s_58_port, plusA(57) => plus2A_s_57_port, 
                           plusA(56) => plus2A_s_56_port, plusA(55) => 
                           plus2A_s_55_port, plusA(54) => plus2A_s_54_port, 
                           plusA(53) => plus2A_s_53_port, plusA(52) => 
                           plus2A_s_52_port, plusA(51) => plus2A_s_51_port, 
                           plusA(50) => plus2A_s_50_port, plusA(49) => 
                           plus2A_s_49_port, plusA(48) => plus2A_s_48_port, 
                           plusA(47) => plus2A_s_47_port, plusA(46) => 
                           plus2A_s_46_port, plusA(45) => plus2A_s_45_port, 
                           plusA(44) => plus2A_s_44_port, plusA(43) => 
                           plus2A_s_43_port, plusA(42) => plus2A_s_42_port, 
                           plusA(41) => plus2A_s_41_port, plusA(40) => 
                           plus2A_s_40_port, plusA(39) => plus2A_s_39_port, 
                           plusA(38) => plus2A_s_38_port, plusA(37) => 
                           plus2A_s_37_port, plusA(36) => plus2A_s_36_port, 
                           plusA(35) => plus2A_s_35_port, plusA(34) => 
                           plus2A_s_34_port, plusA(33) => plus2A_s_33_port, 
                           plusA(32) => plus2A_s_32_port, plusA(31) => 
                           plus2A_s_31_port, plusA(30) => plus2A_s_30_port, 
                           plusA(29) => plus2A_s_29_port, plusA(28) => 
                           plus2A_s_28_port, plusA(27) => plus2A_s_27_port, 
                           plusA(26) => plus2A_s_26_port, plusA(25) => 
                           plus2A_s_25_port, plusA(24) => plus2A_s_24_port, 
                           plusA(23) => plus2A_s_23_port, plusA(22) => 
                           plus2A_s_22_port, plusA(21) => plus2A_s_21_port, 
                           plusA(20) => plus2A_s_20_port, plusA(19) => 
                           plus2A_s_19_port, plusA(18) => plus2A_s_18_port, 
                           plusA(17) => plus2A_s_17_port, plusA(16) => 
                           plus2A_s_16_port, plusA(15) => plus2A_s_15_port, 
                           plusA(14) => plus2A_s_14_port, plusA(13) => 
                           plus2A_s_13_port, plusA(12) => plus2A_s_12_port, 
                           plusA(11) => plus2A_s_11_port, plusA(10) => 
                           plus2A_s_10_port, plusA(9) => plus2A_s_9_port, 
                           plusA(8) => plus2A_s_8_port, plusA(7) => 
                           plus2A_s_7_port, plusA(6) => plus2A_s_6_port, 
                           plusA(5) => plus2A_s_5_port, plusA(4) => 
                           plus2A_s_4_port, plusA(3) => plus2A_s_3_port, 
                           plusA(2) => plus2A_s_2_port, plusA(1) => 
                           plus2A_s_1_port, plusA(0) => nextA_0_port, 
                           minusA(63) => minus2A_s_63_port, minusA(62) => 
                           minus2A_s_62_port, minusA(61) => minus2A_s_61_port, 
                           minusA(60) => minus2A_s_60_port, minusA(59) => 
                           minus2A_s_59_port, minusA(58) => minus2A_s_58_port, 
                           minusA(57) => minus2A_s_57_port, minusA(56) => 
                           minus2A_s_56_port, minusA(55) => minus2A_s_55_port, 
                           minusA(54) => minus2A_s_54_port, minusA(53) => 
                           minus2A_s_53_port, minusA(52) => minus2A_s_52_port, 
                           minusA(51) => minus2A_s_51_port, minusA(50) => 
                           minus2A_s_50_port, minusA(49) => minus2A_s_49_port, 
                           minusA(48) => minus2A_s_48_port, minusA(47) => 
                           minus2A_s_47_port, minusA(46) => minus2A_s_46_port, 
                           minusA(45) => minus2A_s_45_port, minusA(44) => 
                           minus2A_s_44_port, minusA(43) => minus2A_s_43_port, 
                           minusA(42) => minus2A_s_42_port, minusA(41) => 
                           minus2A_s_41_port, minusA(40) => minus2A_s_40_port, 
                           minusA(39) => minus2A_s_39_port, minusA(38) => 
                           minus2A_s_38_port, minusA(37) => minus2A_s_37_port, 
                           minusA(36) => minus2A_s_36_port, minusA(35) => 
                           minus2A_s_35_port, minusA(34) => minus2A_s_34_port, 
                           minusA(33) => minus2A_s_33_port, minusA(32) => 
                           minus2A_s_32_port, minusA(31) => minus2A_s_31_port, 
                           minusA(30) => minus2A_s_30_port, minusA(29) => 
                           minus2A_s_29_port, minusA(28) => minus2A_s_28_port, 
                           minusA(27) => minus2A_s_27_port, minusA(26) => 
                           minus2A_s_26_port, minusA(25) => minus2A_s_25_port, 
                           minusA(24) => minus2A_s_24_port, minusA(23) => 
                           minus2A_s_23_port, minusA(22) => minus2A_s_22_port, 
                           minusA(21) => minus2A_s_21_port, minusA(20) => 
                           minus2A_s_20_port, minusA(19) => minus2A_s_19_port, 
                           minusA(18) => minus2A_s_18_port, minusA(17) => 
                           minus2A_s_17_port, minusA(16) => minus2A_s_16_port, 
                           minusA(15) => minus2A_s_15_port, minusA(14) => 
                           minus2A_s_14_port, minusA(13) => minus2A_s_13_port, 
                           minusA(12) => minus2A_s_12_port, minusA(11) => 
                           minus2A_s_11_port, minusA(10) => minus2A_s_10_port, 
                           minusA(9) => minus2A_s_9_port, minusA(8) => 
                           minus2A_s_8_port, minusA(7) => minus2A_s_7_port, 
                           minusA(6) => minus2A_s_6_port, minusA(5) => 
                           minus2A_s_5_port, minusA(4) => minus2A_s_4_port, 
                           minusA(3) => minus2A_s_3_port, minusA(2) => 
                           minus2A_s_2_port, minusA(1) => minus2A_s_1_port, 
                           minusA(0) => minus2A_s_0_port, plus2A(63) => 
                           nextA_63_port, plus2A(62) => nextA_62_port, 
                           plus2A(61) => nextA_61_port, plus2A(60) => 
                           nextA_60_port, plus2A(59) => nextA_59_port, 
                           plus2A(58) => nextA_58_port, plus2A(57) => 
                           nextA_57_port, plus2A(56) => nextA_56_port, 
                           plus2A(55) => nextA_55_port, plus2A(54) => 
                           nextA_54_port, plus2A(53) => nextA_53_port, 
                           plus2A(52) => nextA_52_port, plus2A(51) => 
                           nextA_51_port, plus2A(50) => nextA_50_port, 
                           plus2A(49) => nextA_49_port, plus2A(48) => 
                           nextA_48_port, plus2A(47) => nextA_47_port, 
                           plus2A(46) => nextA_46_port, plus2A(45) => 
                           nextA_45_port, plus2A(44) => nextA_44_port, 
                           plus2A(43) => nextA_43_port, plus2A(42) => 
                           nextA_42_port, plus2A(41) => nextA_41_port, 
                           plus2A(40) => nextA_40_port, plus2A(39) => 
                           nextA_39_port, plus2A(38) => nextA_38_port, 
                           plus2A(37) => nextA_37_port, plus2A(36) => 
                           nextA_36_port, plus2A(35) => nextA_35_port, 
                           plus2A(34) => nextA_34_port, plus2A(33) => 
                           nextA_33_port, plus2A(32) => nextA_32_port, 
                           plus2A(31) => nextA_31_port, plus2A(30) => 
                           nextA_30_port, plus2A(29) => nextA_29_port, 
                           plus2A(28) => nextA_28_port, plus2A(27) => 
                           nextA_27_port, plus2A(26) => nextA_26_port, 
                           plus2A(25) => nextA_25_port, plus2A(24) => 
                           nextA_24_port, plus2A(23) => nextA_23_port, 
                           plus2A(22) => nextA_22_port, plus2A(21) => 
                           nextA_21_port, plus2A(20) => nextA_20_port, 
                           plus2A(19) => nextA_19_port, plus2A(18) => 
                           nextA_18_port, plus2A(17) => nextA_17_port, 
                           plus2A(16) => nextA_16_port, plus2A(15) => 
                           nextA_15_port, plus2A(14) => nextA_14_port, 
                           plus2A(13) => nextA_13_port, plus2A(12) => 
                           nextA_12_port, plus2A(11) => nextA_11_port, 
                           plus2A(10) => nextA_10_port, plus2A(9) => 
                           nextA_9_port, plus2A(8) => nextA_8_port, plus2A(7) 
                           => nextA_7_port, plus2A(6) => nextA_6_port, 
                           plus2A(5) => nextA_5_port, plus2A(4) => nextA_4_port
                           , plus2A(3) => nextA_3_port, plus2A(2) => 
                           nextA_2_port, plus2A(1) => nextA_1_port, plus2A(0) 
                           => nextA_0_port, minus2A(63) => minus4A_s_63_port, 
                           minus2A(62) => minus4A_s_62_port, minus2A(61) => 
                           minus4A_s_61_port, minus2A(60) => minus4A_s_60_port,
                           minus2A(59) => minus4A_s_59_port, minus2A(58) => 
                           minus4A_s_58_port, minus2A(57) => minus4A_s_57_port,
                           minus2A(56) => minus4A_s_56_port, minus2A(55) => 
                           minus4A_s_55_port, minus2A(54) => minus4A_s_54_port,
                           minus2A(53) => minus4A_s_53_port, minus2A(52) => 
                           minus4A_s_52_port, minus2A(51) => minus4A_s_51_port,
                           minus2A(50) => minus4A_s_50_port, minus2A(49) => 
                           minus4A_s_49_port, minus2A(48) => minus4A_s_48_port,
                           minus2A(47) => minus4A_s_47_port, minus2A(46) => 
                           minus4A_s_46_port, minus2A(45) => minus4A_s_45_port,
                           minus2A(44) => minus4A_s_44_port, minus2A(43) => 
                           minus4A_s_43_port, minus2A(42) => minus4A_s_42_port,
                           minus2A(41) => minus4A_s_41_port, minus2A(40) => 
                           minus4A_s_40_port, minus2A(39) => minus4A_s_39_port,
                           minus2A(38) => minus4A_s_38_port, minus2A(37) => 
                           minus4A_s_37_port, minus2A(36) => minus4A_s_36_port,
                           minus2A(35) => minus4A_s_35_port, minus2A(34) => 
                           minus4A_s_34_port, minus2A(33) => minus4A_s_33_port,
                           minus2A(32) => minus4A_s_32_port, minus2A(31) => 
                           minus4A_s_31_port, minus2A(30) => minus4A_s_30_port,
                           minus2A(29) => minus4A_s_29_port, minus2A(28) => 
                           minus4A_s_28_port, minus2A(27) => minus4A_s_27_port,
                           minus2A(26) => minus4A_s_26_port, minus2A(25) => 
                           minus4A_s_25_port, minus2A(24) => minus4A_s_24_port,
                           minus2A(23) => minus4A_s_23_port, minus2A(22) => 
                           minus4A_s_22_port, minus2A(21) => minus4A_s_21_port,
                           minus2A(20) => minus4A_s_20_port, minus2A(19) => 
                           minus4A_s_19_port, minus2A(18) => minus4A_s_18_port,
                           minus2A(17) => minus4A_s_17_port, minus2A(16) => 
                           minus4A_s_16_port, minus2A(15) => minus4A_s_15_port,
                           minus2A(14) => minus4A_s_14_port, minus2A(13) => 
                           minus4A_s_13_port, minus2A(12) => minus4A_s_12_port,
                           minus2A(11) => minus4A_s_11_port, minus2A(10) => 
                           minus4A_s_10_port, minus2A(9) => minus4A_s_9_port, 
                           minus2A(8) => minus4A_s_8_port, minus2A(7) => 
                           minus4A_s_7_port, minus2A(6) => minus4A_s_6_port, 
                           minus2A(5) => minus4A_s_5_port, minus2A(4) => 
                           minus4A_s_4_port, minus2A(3) => minus4A_s_3_port, 
                           minus2A(2) => minus4A_s_2_port, minus2A(1) => 
                           minus4A_s_1_port, minus2A(0) => minus4A_s_0_port, 
                           SEL(2) => encoder_to_mux_2_port, SEL(1) => 
                           encoder_to_mux_1_port, SEL(0) => 
                           encoder_to_mux_0_port, Y(63) => mux_to_adder_63_port
                           , Y(62) => mux_to_adder_62_port, Y(61) => 
                           mux_to_adder_61_port, Y(60) => mux_to_adder_60_port,
                           Y(59) => mux_to_adder_59_port, Y(58) => 
                           mux_to_adder_58_port, Y(57) => mux_to_adder_57_port,
                           Y(56) => mux_to_adder_56_port, Y(55) => 
                           mux_to_adder_55_port, Y(54) => mux_to_adder_54_port,
                           Y(53) => mux_to_adder_53_port, Y(52) => 
                           mux_to_adder_52_port, Y(51) => mux_to_adder_51_port,
                           Y(50) => mux_to_adder_50_port, Y(49) => 
                           mux_to_adder_49_port, Y(48) => mux_to_adder_48_port,
                           Y(47) => mux_to_adder_47_port, Y(46) => 
                           mux_to_adder_46_port, Y(45) => mux_to_adder_45_port,
                           Y(44) => mux_to_adder_44_port, Y(43) => 
                           mux_to_adder_43_port, Y(42) => mux_to_adder_42_port,
                           Y(41) => mux_to_adder_41_port, Y(40) => 
                           mux_to_adder_40_port, Y(39) => mux_to_adder_39_port,
                           Y(38) => mux_to_adder_38_port, Y(37) => 
                           mux_to_adder_37_port, Y(36) => mux_to_adder_36_port,
                           Y(35) => mux_to_adder_35_port, Y(34) => 
                           mux_to_adder_34_port, Y(33) => mux_to_adder_33_port,
                           Y(32) => mux_to_adder_32_port, Y(31) => 
                           mux_to_adder_31_port, Y(30) => mux_to_adder_30_port,
                           Y(29) => mux_to_adder_29_port, Y(28) => 
                           mux_to_adder_28_port, Y(27) => mux_to_adder_27_port,
                           Y(26) => mux_to_adder_26_port, Y(25) => 
                           mux_to_adder_25_port, Y(24) => mux_to_adder_24_port,
                           Y(23) => mux_to_adder_23_port, Y(22) => 
                           mux_to_adder_22_port, Y(21) => mux_to_adder_21_port,
                           Y(20) => mux_to_adder_20_port, Y(19) => 
                           mux_to_adder_19_port, Y(18) => mux_to_adder_18_port,
                           Y(17) => mux_to_adder_17_port, Y(16) => 
                           mux_to_adder_16_port, Y(15) => mux_to_adder_15_port,
                           Y(14) => mux_to_adder_14_port, Y(13) => 
                           mux_to_adder_13_port, Y(12) => mux_to_adder_12_port,
                           Y(11) => mux_to_adder_11_port, Y(10) => 
                           mux_to_adder_10_port, Y(9) => mux_to_adder_9_port, 
                           Y(8) => mux_to_adder_8_port, Y(7) => 
                           mux_to_adder_7_port, Y(6) => mux_to_adder_6_port, 
                           Y(5) => mux_to_adder_5_port, Y(4) => 
                           mux_to_adder_4_port, Y(3) => mux_to_adder_3_port, 
                           Y(2) => mux_to_adder_2_port, Y(1) => 
                           mux_to_adder_1_port, Y(0) => mux_to_adder_0_port);
   rca_1 : RCA_N64_3 port map( A(63) => mux_to_adder_63_port, A(62) => 
                           mux_to_adder_62_port, A(61) => mux_to_adder_61_port,
                           A(60) => mux_to_adder_60_port, A(59) => 
                           mux_to_adder_59_port, A(58) => mux_to_adder_58_port,
                           A(57) => mux_to_adder_57_port, A(56) => 
                           mux_to_adder_56_port, A(55) => mux_to_adder_55_port,
                           A(54) => mux_to_adder_54_port, A(53) => 
                           mux_to_adder_53_port, A(52) => mux_to_adder_52_port,
                           A(51) => mux_to_adder_51_port, A(50) => 
                           mux_to_adder_50_port, A(49) => mux_to_adder_49_port,
                           A(48) => mux_to_adder_48_port, A(47) => 
                           mux_to_adder_47_port, A(46) => mux_to_adder_46_port,
                           A(45) => mux_to_adder_45_port, A(44) => 
                           mux_to_adder_44_port, A(43) => mux_to_adder_43_port,
                           A(42) => mux_to_adder_42_port, A(41) => 
                           mux_to_adder_41_port, A(40) => mux_to_adder_40_port,
                           A(39) => mux_to_adder_39_port, A(38) => 
                           mux_to_adder_38_port, A(37) => mux_to_adder_37_port,
                           A(36) => mux_to_adder_36_port, A(35) => 
                           mux_to_adder_35_port, A(34) => mux_to_adder_34_port,
                           A(33) => mux_to_adder_33_port, A(32) => 
                           mux_to_adder_32_port, A(31) => mux_to_adder_31_port,
                           A(30) => mux_to_adder_30_port, A(29) => 
                           mux_to_adder_29_port, A(28) => mux_to_adder_28_port,
                           A(27) => mux_to_adder_27_port, A(26) => 
                           mux_to_adder_26_port, A(25) => mux_to_adder_25_port,
                           A(24) => mux_to_adder_24_port, A(23) => 
                           mux_to_adder_23_port, A(22) => mux_to_adder_22_port,
                           A(21) => mux_to_adder_21_port, A(20) => 
                           mux_to_adder_20_port, A(19) => mux_to_adder_19_port,
                           A(18) => mux_to_adder_18_port, A(17) => 
                           mux_to_adder_17_port, A(16) => mux_to_adder_16_port,
                           A(15) => mux_to_adder_15_port, A(14) => 
                           mux_to_adder_14_port, A(13) => mux_to_adder_13_port,
                           A(12) => mux_to_adder_12_port, A(11) => 
                           mux_to_adder_11_port, A(10) => mux_to_adder_10_port,
                           A(9) => mux_to_adder_9_port, A(8) => 
                           mux_to_adder_8_port, A(7) => mux_to_adder_7_port, 
                           A(6) => mux_to_adder_6_port, A(5) => 
                           mux_to_adder_5_port, A(4) => mux_to_adder_4_port, 
                           A(3) => mux_to_adder_3_port, A(2) => 
                           mux_to_adder_2_port, A(1) => mux_to_adder_1_port, 
                           A(0) => mux_to_adder_0_port, B(63) => prevSum(63), 
                           B(62) => prevSum(62), B(61) => prevSum(61), B(60) =>
                           prevSum(60), B(59) => prevSum(59), B(58) => 
                           prevSum(58), B(57) => prevSum(57), B(56) => 
                           prevSum(56), B(55) => prevSum(55), B(54) => 
                           prevSum(54), B(53) => prevSum(53), B(52) => 
                           prevSum(52), B(51) => prevSum(51), B(50) => 
                           prevSum(50), B(49) => prevSum(49), B(48) => 
                           prevSum(48), B(47) => prevSum(47), B(46) => 
                           prevSum(46), B(45) => prevSum(45), B(44) => 
                           prevSum(44), B(43) => prevSum(43), B(42) => 
                           prevSum(42), B(41) => prevSum(41), B(40) => 
                           prevSum(40), B(39) => prevSum(39), B(38) => 
                           prevSum(38), B(37) => prevSum(37), B(36) => 
                           prevSum(36), B(35) => prevSum(35), B(34) => 
                           prevSum(34), B(33) => prevSum(33), B(32) => 
                           prevSum(32), B(31) => prevSum(31), B(30) => 
                           prevSum(30), B(29) => prevSum(29), B(28) => 
                           prevSum(28), B(27) => prevSum(27), B(26) => 
                           prevSum(26), B(25) => prevSum(25), B(24) => 
                           prevSum(24), B(23) => prevSum(23), B(22) => 
                           prevSum(22), B(21) => prevSum(21), B(20) => 
                           prevSum(20), B(19) => prevSum(19), B(18) => 
                           prevSum(18), B(17) => prevSum(17), B(16) => 
                           prevSum(16), B(15) => prevSum(15), B(14) => 
                           prevSum(14), B(13) => prevSum(13), B(12) => 
                           prevSum(12), B(11) => prevSum(11), B(10) => 
                           prevSum(10), B(9) => prevSum(9), B(8) => prevSum(8),
                           B(7) => prevSum(7), B(6) => prevSum(6), B(5) => 
                           prevSum(5), B(4) => prevSum(4), B(3) => prevSum(3), 
                           B(2) => prevSum(2), B(1) => prevSum(1), B(0) => 
                           prevSum(0), Ci => X_Logic0_port, S(63) => 
                           nextSum(63), S(62) => nextSum(62), S(61) => 
                           nextSum(61), S(60) => nextSum(60), S(59) => 
                           nextSum(59), S(58) => nextSum(58), S(57) => 
                           nextSum(57), S(56) => nextSum(56), S(55) => 
                           nextSum(55), S(54) => nextSum(54), S(53) => 
                           nextSum(53), S(52) => nextSum(52), S(51) => 
                           nextSum(51), S(50) => nextSum(50), S(49) => 
                           nextSum(49), S(48) => nextSum(48), S(47) => 
                           nextSum(47), S(46) => nextSum(46), S(45) => 
                           nextSum(45), S(44) => nextSum(44), S(43) => 
                           nextSum(43), S(42) => nextSum(42), S(41) => 
                           nextSum(41), S(40) => nextSum(40), S(39) => 
                           nextSum(39), S(38) => nextSum(38), S(37) => 
                           nextSum(37), S(36) => nextSum(36), S(35) => 
                           nextSum(35), S(34) => nextSum(34), S(33) => 
                           nextSum(33), S(32) => nextSum(32), S(31) => 
                           nextSum(31), S(30) => nextSum(30), S(29) => 
                           nextSum(29), S(28) => nextSum(28), S(27) => 
                           nextSum(27), S(26) => nextSum(26), S(25) => 
                           nextSum(25), S(24) => nextSum(24), S(23) => 
                           nextSum(23), S(22) => nextSum(22), S(21) => 
                           nextSum(21), S(20) => nextSum(20), S(19) => 
                           nextSum(19), S(18) => nextSum(18), S(17) => 
                           nextSum(17), S(16) => nextSum(16), S(15) => 
                           nextSum(15), S(14) => nextSum(14), S(13) => 
                           nextSum(13), S(12) => nextSum(12), S(11) => 
                           nextSum(11), S(10) => nextSum(10), S(9) => 
                           nextSum(9), S(8) => nextSum(8), S(7) => nextSum(7), 
                           S(6) => nextSum(6), S(5) => nextSum(5), S(4) => 
                           nextSum(4), S(3) => nextSum(3), S(2) => nextSum(2), 
                           S(1) => nextSum(1), S(0) => nextSum(0), Co => n_3183
                           );

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity booth_mul_row_N64_RADIX3_4 is

   port( prevA, prevSum : in std_logic_vector (63 downto 0);  encoderIn : in 
         std_logic_vector (2 downto 0);  nextA, nextSum : out std_logic_vector 
         (63 downto 0));

end booth_mul_row_N64_RADIX3_4;

architecture SYN_struct of booth_mul_row_N64_RADIX3_4 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component RCA_N64_4
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component MUX_GENERIC_N64_RADIX3_4
      port( plusA, minusA, plus2A, minus2A : in std_logic_vector (63 downto 0);
            SEL : in std_logic_vector (2 downto 0);  Y : out std_logic_vector 
            (63 downto 0));
   end component;
   
   component ShiftnCompl_N64_4
      port( plusA : in std_logic_vector (63 downto 0);  plus2A_out, minus2A_out
            , plus4A_out, minus4A_out : out std_logic_vector (63 downto 0));
   end component;
   
   component encoder_N64_RADIX3_4
      port( X : in std_logic_vector (2 downto 0);  Z : out std_logic_vector (2 
            downto 0));
   end component;
   
   signal X_Logic0_port, nextA_63_port, nextA_62_port, nextA_61_port, 
      nextA_60_port, nextA_59_port, nextA_58_port, n3, nextA_56_port, 
      nextA_55_port, nextA_54_port, nextA_53_port, nextA_52_port, nextA_51_port
      , nextA_50_port, nextA_49_port, nextA_48_port, nextA_47_port, 
      nextA_46_port, nextA_45_port, nextA_44_port, nextA_43_port, nextA_42_port
      , nextA_41_port, nextA_40_port, nextA_39_port, nextA_38_port, 
      nextA_37_port, nextA_36_port, nextA_35_port, nextA_34_port, nextA_33_port
      , nextA_32_port, nextA_31_port, nextA_30_port, nextA_29_port, 
      nextA_28_port, nextA_27_port, nextA_26_port, nextA_25_port, nextA_24_port
      , nextA_23_port, nextA_22_port, nextA_21_port, nextA_20_port, 
      nextA_19_port, nextA_18_port, nextA_17_port, nextA_16_port, nextA_15_port
      , nextA_14_port, nextA_13_port, nextA_12_port, nextA_11_port, 
      nextA_10_port, nextA_9_port, nextA_8_port, nextA_7_port, nextA_6_port, 
      nextA_5_port, nextA_4_port, nextA_3_port, nextA_2_port, nextA_1_port, 
      encoder_to_mux_2_port, encoder_to_mux_1_port, encoder_to_mux_0_port, 
      plus2A_s_63_port, plus2A_s_62_port, plus2A_s_61_port, plus2A_s_60_port, 
      plus2A_s_59_port, plus2A_s_58_port, plus2A_s_57_port, plus2A_s_56_port, 
      plus2A_s_55_port, plus2A_s_54_port, plus2A_s_53_port, plus2A_s_52_port, 
      plus2A_s_51_port, plus2A_s_50_port, plus2A_s_49_port, plus2A_s_48_port, 
      plus2A_s_47_port, plus2A_s_46_port, plus2A_s_45_port, plus2A_s_44_port, 
      plus2A_s_43_port, plus2A_s_42_port, plus2A_s_41_port, plus2A_s_40_port, 
      plus2A_s_39_port, plus2A_s_38_port, plus2A_s_37_port, plus2A_s_36_port, 
      plus2A_s_35_port, plus2A_s_34_port, plus2A_s_33_port, plus2A_s_32_port, 
      plus2A_s_31_port, plus2A_s_30_port, plus2A_s_29_port, plus2A_s_28_port, 
      plus2A_s_27_port, plus2A_s_26_port, plus2A_s_25_port, plus2A_s_24_port, 
      plus2A_s_23_port, plus2A_s_22_port, plus2A_s_21_port, plus2A_s_20_port, 
      plus2A_s_19_port, plus2A_s_18_port, plus2A_s_17_port, plus2A_s_16_port, 
      plus2A_s_15_port, plus2A_s_14_port, plus2A_s_13_port, plus2A_s_12_port, 
      plus2A_s_11_port, plus2A_s_10_port, plus2A_s_9_port, plus2A_s_8_port, 
      plus2A_s_7_port, plus2A_s_6_port, plus2A_s_5_port, plus2A_s_4_port, 
      plus2A_s_3_port, plus2A_s_2_port, plus2A_s_1_port, minus2A_s_63_port, 
      minus2A_s_62_port, minus2A_s_61_port, minus2A_s_60_port, 
      minus2A_s_59_port, minus2A_s_58_port, minus2A_s_57_port, 
      minus2A_s_56_port, minus2A_s_55_port, minus2A_s_54_port, 
      minus2A_s_53_port, minus2A_s_52_port, minus2A_s_51_port, 
      minus2A_s_50_port, minus2A_s_49_port, minus2A_s_48_port, 
      minus2A_s_47_port, minus2A_s_46_port, minus2A_s_45_port, 
      minus2A_s_44_port, minus2A_s_43_port, minus2A_s_42_port, 
      minus2A_s_41_port, minus2A_s_40_port, minus2A_s_39_port, 
      minus2A_s_38_port, minus2A_s_37_port, minus2A_s_36_port, 
      minus2A_s_35_port, minus2A_s_34_port, minus2A_s_33_port, 
      minus2A_s_32_port, minus2A_s_31_port, minus2A_s_30_port, 
      minus2A_s_29_port, minus2A_s_28_port, minus2A_s_27_port, 
      minus2A_s_26_port, minus2A_s_25_port, minus2A_s_24_port, 
      minus2A_s_23_port, minus2A_s_22_port, minus2A_s_21_port, 
      minus2A_s_20_port, minus2A_s_19_port, minus2A_s_18_port, 
      minus2A_s_17_port, minus2A_s_16_port, minus2A_s_15_port, 
      minus2A_s_14_port, minus2A_s_13_port, minus2A_s_12_port, 
      minus2A_s_11_port, minus2A_s_10_port, minus2A_s_9_port, minus2A_s_8_port,
      minus2A_s_7_port, minus2A_s_6_port, minus2A_s_5_port, minus2A_s_4_port, 
      minus2A_s_3_port, minus2A_s_2_port, minus2A_s_1_port, minus2A_s_0_port, 
      minus4A_s_63_port, minus4A_s_62_port, minus4A_s_61_port, 
      minus4A_s_60_port, minus4A_s_59_port, minus4A_s_58_port, 
      minus4A_s_57_port, minus4A_s_56_port, minus4A_s_55_port, 
      minus4A_s_54_port, minus4A_s_53_port, minus4A_s_52_port, 
      minus4A_s_51_port, minus4A_s_50_port, minus4A_s_49_port, 
      minus4A_s_48_port, minus4A_s_47_port, minus4A_s_46_port, 
      minus4A_s_45_port, minus4A_s_44_port, minus4A_s_43_port, 
      minus4A_s_42_port, minus4A_s_41_port, minus4A_s_40_port, 
      minus4A_s_39_port, minus4A_s_38_port, minus4A_s_37_port, 
      minus4A_s_36_port, minus4A_s_35_port, minus4A_s_34_port, 
      minus4A_s_33_port, minus4A_s_32_port, minus4A_s_31_port, 
      minus4A_s_30_port, minus4A_s_29_port, minus4A_s_28_port, 
      minus4A_s_27_port, minus4A_s_26_port, minus4A_s_25_port, 
      minus4A_s_24_port, minus4A_s_23_port, minus4A_s_22_port, 
      minus4A_s_21_port, minus4A_s_20_port, minus4A_s_19_port, 
      minus4A_s_18_port, minus4A_s_17_port, minus4A_s_16_port, 
      minus4A_s_15_port, minus4A_s_14_port, minus4A_s_13_port, 
      minus4A_s_12_port, minus4A_s_11_port, minus4A_s_10_port, minus4A_s_9_port
      , minus4A_s_8_port, minus4A_s_7_port, minus4A_s_6_port, minus4A_s_5_port,
      minus4A_s_4_port, minus4A_s_3_port, minus4A_s_2_port, minus4A_s_1_port, 
      minus4A_s_0_port, mux_to_adder_63_port, mux_to_adder_62_port, 
      mux_to_adder_61_port, mux_to_adder_60_port, mux_to_adder_59_port, 
      mux_to_adder_58_port, mux_to_adder_57_port, mux_to_adder_56_port, 
      mux_to_adder_55_port, mux_to_adder_54_port, mux_to_adder_53_port, 
      mux_to_adder_52_port, mux_to_adder_51_port, mux_to_adder_50_port, 
      mux_to_adder_49_port, mux_to_adder_48_port, mux_to_adder_47_port, 
      mux_to_adder_46_port, mux_to_adder_45_port, mux_to_adder_44_port, 
      mux_to_adder_43_port, mux_to_adder_42_port, mux_to_adder_41_port, 
      mux_to_adder_40_port, mux_to_adder_39_port, mux_to_adder_38_port, 
      mux_to_adder_37_port, mux_to_adder_36_port, mux_to_adder_35_port, 
      mux_to_adder_34_port, mux_to_adder_33_port, mux_to_adder_32_port, 
      mux_to_adder_31_port, mux_to_adder_30_port, mux_to_adder_29_port, 
      mux_to_adder_28_port, mux_to_adder_27_port, mux_to_adder_26_port, 
      mux_to_adder_25_port, mux_to_adder_24_port, mux_to_adder_23_port, 
      mux_to_adder_22_port, mux_to_adder_21_port, mux_to_adder_20_port, 
      mux_to_adder_19_port, mux_to_adder_18_port, mux_to_adder_17_port, 
      mux_to_adder_16_port, mux_to_adder_15_port, mux_to_adder_14_port, 
      mux_to_adder_13_port, mux_to_adder_12_port, mux_to_adder_11_port, 
      mux_to_adder_10_port, mux_to_adder_9_port, mux_to_adder_8_port, 
      mux_to_adder_7_port, mux_to_adder_6_port, mux_to_adder_5_port, 
      mux_to_adder_4_port, mux_to_adder_3_port, mux_to_adder_2_port, 
      mux_to_adder_1_port, mux_to_adder_0_port, nextA_0_port, nextA_57_port, 
      n_3184, n_3185, n_3186 : std_logic;

begin
   nextA <= ( nextA_63_port, nextA_62_port, nextA_61_port, nextA_60_port, 
      nextA_59_port, nextA_58_port, nextA_57_port, nextA_56_port, nextA_55_port
      , nextA_54_port, nextA_53_port, nextA_52_port, nextA_51_port, 
      nextA_50_port, nextA_49_port, nextA_48_port, nextA_47_port, nextA_46_port
      , nextA_45_port, nextA_44_port, nextA_43_port, nextA_42_port, 
      nextA_41_port, nextA_40_port, nextA_39_port, nextA_38_port, nextA_37_port
      , nextA_36_port, nextA_35_port, nextA_34_port, nextA_33_port, 
      nextA_32_port, nextA_31_port, nextA_30_port, nextA_29_port, nextA_28_port
      , nextA_27_port, nextA_26_port, nextA_25_port, nextA_24_port, 
      nextA_23_port, nextA_22_port, nextA_21_port, nextA_20_port, nextA_19_port
      , nextA_18_port, nextA_17_port, nextA_16_port, nextA_15_port, 
      nextA_14_port, nextA_13_port, nextA_12_port, nextA_11_port, nextA_10_port
      , nextA_9_port, nextA_8_port, nextA_7_port, nextA_6_port, nextA_5_port, 
      nextA_4_port, nextA_3_port, nextA_2_port, nextA_1_port, nextA_0_port );
   
   X_Logic0_port <= '0';
   nextA_0_port <= '0';
   encoder_1 : encoder_N64_RADIX3_4 port map( X(2) => encoderIn(2), X(1) => 
                           encoderIn(1), X(0) => encoderIn(0), Z(2) => 
                           encoder_to_mux_2_port, Z(1) => encoder_to_mux_1_port
                           , Z(0) => encoder_to_mux_0_port);
   ShiftnCompl_1 : ShiftnCompl_N64_4 port map( plusA(63) => prevA(63), 
                           plusA(62) => prevA(62), plusA(61) => prevA(61), 
                           plusA(60) => prevA(60), plusA(59) => prevA(59), 
                           plusA(58) => prevA(58), plusA(57) => prevA(57), 
                           plusA(56) => prevA(56), plusA(55) => prevA(55), 
                           plusA(54) => prevA(54), plusA(53) => prevA(53), 
                           plusA(52) => prevA(52), plusA(51) => prevA(51), 
                           plusA(50) => prevA(50), plusA(49) => prevA(49), 
                           plusA(48) => prevA(48), plusA(47) => prevA(47), 
                           plusA(46) => prevA(46), plusA(45) => prevA(45), 
                           plusA(44) => prevA(44), plusA(43) => prevA(43), 
                           plusA(42) => prevA(42), plusA(41) => prevA(41), 
                           plusA(40) => prevA(40), plusA(39) => prevA(39), 
                           plusA(38) => prevA(38), plusA(37) => prevA(37), 
                           plusA(36) => prevA(36), plusA(35) => prevA(35), 
                           plusA(34) => prevA(34), plusA(33) => prevA(33), 
                           plusA(32) => prevA(32), plusA(31) => prevA(31), 
                           plusA(30) => prevA(30), plusA(29) => prevA(29), 
                           plusA(28) => prevA(28), plusA(27) => prevA(27), 
                           plusA(26) => prevA(26), plusA(25) => prevA(25), 
                           plusA(24) => prevA(24), plusA(23) => prevA(23), 
                           plusA(22) => prevA(22), plusA(21) => prevA(21), 
                           plusA(20) => prevA(20), plusA(19) => prevA(19), 
                           plusA(18) => prevA(18), plusA(17) => prevA(17), 
                           plusA(16) => prevA(16), plusA(15) => prevA(15), 
                           plusA(14) => prevA(14), plusA(13) => prevA(13), 
                           plusA(12) => prevA(12), plusA(11) => prevA(11), 
                           plusA(10) => prevA(10), plusA(9) => prevA(9), 
                           plusA(8) => prevA(8), plusA(7) => prevA(7), plusA(6)
                           => prevA(6), plusA(5) => prevA(5), plusA(4) => 
                           prevA(4), plusA(3) => prevA(3), plusA(2) => prevA(2)
                           , plusA(1) => prevA(1), plusA(0) => prevA(0), 
                           plus2A_out(63) => plus2A_s_63_port, plus2A_out(62) 
                           => plus2A_s_62_port, plus2A_out(61) => 
                           plus2A_s_61_port, plus2A_out(60) => plus2A_s_60_port
                           , plus2A_out(59) => plus2A_s_59_port, plus2A_out(58)
                           => plus2A_s_58_port, plus2A_out(57) => 
                           plus2A_s_57_port, plus2A_out(56) => plus2A_s_56_port
                           , plus2A_out(55) => plus2A_s_55_port, plus2A_out(54)
                           => plus2A_s_54_port, plus2A_out(53) => 
                           plus2A_s_53_port, plus2A_out(52) => plus2A_s_52_port
                           , plus2A_out(51) => plus2A_s_51_port, plus2A_out(50)
                           => plus2A_s_50_port, plus2A_out(49) => 
                           plus2A_s_49_port, plus2A_out(48) => plus2A_s_48_port
                           , plus2A_out(47) => plus2A_s_47_port, plus2A_out(46)
                           => plus2A_s_46_port, plus2A_out(45) => 
                           plus2A_s_45_port, plus2A_out(44) => plus2A_s_44_port
                           , plus2A_out(43) => plus2A_s_43_port, plus2A_out(42)
                           => plus2A_s_42_port, plus2A_out(41) => 
                           plus2A_s_41_port, plus2A_out(40) => plus2A_s_40_port
                           , plus2A_out(39) => plus2A_s_39_port, plus2A_out(38)
                           => plus2A_s_38_port, plus2A_out(37) => 
                           plus2A_s_37_port, plus2A_out(36) => plus2A_s_36_port
                           , plus2A_out(35) => plus2A_s_35_port, plus2A_out(34)
                           => plus2A_s_34_port, plus2A_out(33) => 
                           plus2A_s_33_port, plus2A_out(32) => plus2A_s_32_port
                           , plus2A_out(31) => plus2A_s_31_port, plus2A_out(30)
                           => plus2A_s_30_port, plus2A_out(29) => 
                           plus2A_s_29_port, plus2A_out(28) => plus2A_s_28_port
                           , plus2A_out(27) => plus2A_s_27_port, plus2A_out(26)
                           => plus2A_s_26_port, plus2A_out(25) => 
                           plus2A_s_25_port, plus2A_out(24) => plus2A_s_24_port
                           , plus2A_out(23) => plus2A_s_23_port, plus2A_out(22)
                           => plus2A_s_22_port, plus2A_out(21) => 
                           plus2A_s_21_port, plus2A_out(20) => plus2A_s_20_port
                           , plus2A_out(19) => plus2A_s_19_port, plus2A_out(18)
                           => plus2A_s_18_port, plus2A_out(17) => 
                           plus2A_s_17_port, plus2A_out(16) => plus2A_s_16_port
                           , plus2A_out(15) => plus2A_s_15_port, plus2A_out(14)
                           => plus2A_s_14_port, plus2A_out(13) => 
                           plus2A_s_13_port, plus2A_out(12) => plus2A_s_12_port
                           , plus2A_out(11) => plus2A_s_11_port, plus2A_out(10)
                           => plus2A_s_10_port, plus2A_out(9) => 
                           plus2A_s_9_port, plus2A_out(8) => plus2A_s_8_port, 
                           plus2A_out(7) => plus2A_s_7_port, plus2A_out(6) => 
                           plus2A_s_6_port, plus2A_out(5) => plus2A_s_5_port, 
                           plus2A_out(4) => plus2A_s_4_port, plus2A_out(3) => 
                           plus2A_s_3_port, plus2A_out(2) => plus2A_s_2_port, 
                           plus2A_out(1) => plus2A_s_1_port, plus2A_out(0) => 
                           n_3184, minus2A_out(63) => minus2A_s_63_port, 
                           minus2A_out(62) => minus2A_s_62_port, 
                           minus2A_out(61) => minus2A_s_61_port, 
                           minus2A_out(60) => minus2A_s_60_port, 
                           minus2A_out(59) => minus2A_s_59_port, 
                           minus2A_out(58) => minus2A_s_58_port, 
                           minus2A_out(57) => minus2A_s_57_port, 
                           minus2A_out(56) => minus2A_s_56_port, 
                           minus2A_out(55) => minus2A_s_55_port, 
                           minus2A_out(54) => minus2A_s_54_port, 
                           minus2A_out(53) => minus2A_s_53_port, 
                           minus2A_out(52) => minus2A_s_52_port, 
                           minus2A_out(51) => minus2A_s_51_port, 
                           minus2A_out(50) => minus2A_s_50_port, 
                           minus2A_out(49) => minus2A_s_49_port, 
                           minus2A_out(48) => minus2A_s_48_port, 
                           minus2A_out(47) => minus2A_s_47_port, 
                           minus2A_out(46) => minus2A_s_46_port, 
                           minus2A_out(45) => minus2A_s_45_port, 
                           minus2A_out(44) => minus2A_s_44_port, 
                           minus2A_out(43) => minus2A_s_43_port, 
                           minus2A_out(42) => minus2A_s_42_port, 
                           minus2A_out(41) => minus2A_s_41_port, 
                           minus2A_out(40) => minus2A_s_40_port, 
                           minus2A_out(39) => minus2A_s_39_port, 
                           minus2A_out(38) => minus2A_s_38_port, 
                           minus2A_out(37) => minus2A_s_37_port, 
                           minus2A_out(36) => minus2A_s_36_port, 
                           minus2A_out(35) => minus2A_s_35_port, 
                           minus2A_out(34) => minus2A_s_34_port, 
                           minus2A_out(33) => minus2A_s_33_port, 
                           minus2A_out(32) => minus2A_s_32_port, 
                           minus2A_out(31) => minus2A_s_31_port, 
                           minus2A_out(30) => minus2A_s_30_port, 
                           minus2A_out(29) => minus2A_s_29_port, 
                           minus2A_out(28) => minus2A_s_28_port, 
                           minus2A_out(27) => minus2A_s_27_port, 
                           minus2A_out(26) => minus2A_s_26_port, 
                           minus2A_out(25) => minus2A_s_25_port, 
                           minus2A_out(24) => minus2A_s_24_port, 
                           minus2A_out(23) => minus2A_s_23_port, 
                           minus2A_out(22) => minus2A_s_22_port, 
                           minus2A_out(21) => minus2A_s_21_port, 
                           minus2A_out(20) => minus2A_s_20_port, 
                           minus2A_out(19) => minus2A_s_19_port, 
                           minus2A_out(18) => minus2A_s_18_port, 
                           minus2A_out(17) => minus2A_s_17_port, 
                           minus2A_out(16) => minus2A_s_16_port, 
                           minus2A_out(15) => minus2A_s_15_port, 
                           minus2A_out(14) => minus2A_s_14_port, 
                           minus2A_out(13) => minus2A_s_13_port, 
                           minus2A_out(12) => minus2A_s_12_port, 
                           minus2A_out(11) => minus2A_s_11_port, 
                           minus2A_out(10) => minus2A_s_10_port, minus2A_out(9)
                           => minus2A_s_9_port, minus2A_out(8) => 
                           minus2A_s_8_port, minus2A_out(7) => minus2A_s_7_port
                           , minus2A_out(6) => minus2A_s_6_port, minus2A_out(5)
                           => minus2A_s_5_port, minus2A_out(4) => 
                           minus2A_s_4_port, minus2A_out(3) => minus2A_s_3_port
                           , minus2A_out(2) => minus2A_s_2_port, minus2A_out(1)
                           => minus2A_s_1_port, minus2A_out(0) => 
                           minus2A_s_0_port, plus4A_out(63) => nextA_63_port, 
                           plus4A_out(62) => nextA_62_port, plus4A_out(61) => 
                           nextA_61_port, plus4A_out(60) => nextA_60_port, 
                           plus4A_out(59) => nextA_59_port, plus4A_out(58) => 
                           nextA_58_port, plus4A_out(57) => n3, plus4A_out(56) 
                           => nextA_56_port, plus4A_out(55) => nextA_55_port, 
                           plus4A_out(54) => nextA_54_port, plus4A_out(53) => 
                           nextA_53_port, plus4A_out(52) => nextA_52_port, 
                           plus4A_out(51) => nextA_51_port, plus4A_out(50) => 
                           nextA_50_port, plus4A_out(49) => nextA_49_port, 
                           plus4A_out(48) => nextA_48_port, plus4A_out(47) => 
                           nextA_47_port, plus4A_out(46) => nextA_46_port, 
                           plus4A_out(45) => nextA_45_port, plus4A_out(44) => 
                           nextA_44_port, plus4A_out(43) => nextA_43_port, 
                           plus4A_out(42) => nextA_42_port, plus4A_out(41) => 
                           nextA_41_port, plus4A_out(40) => nextA_40_port, 
                           plus4A_out(39) => nextA_39_port, plus4A_out(38) => 
                           nextA_38_port, plus4A_out(37) => nextA_37_port, 
                           plus4A_out(36) => nextA_36_port, plus4A_out(35) => 
                           nextA_35_port, plus4A_out(34) => nextA_34_port, 
                           plus4A_out(33) => nextA_33_port, plus4A_out(32) => 
                           nextA_32_port, plus4A_out(31) => nextA_31_port, 
                           plus4A_out(30) => nextA_30_port, plus4A_out(29) => 
                           nextA_29_port, plus4A_out(28) => nextA_28_port, 
                           plus4A_out(27) => nextA_27_port, plus4A_out(26) => 
                           nextA_26_port, plus4A_out(25) => nextA_25_port, 
                           plus4A_out(24) => nextA_24_port, plus4A_out(23) => 
                           nextA_23_port, plus4A_out(22) => nextA_22_port, 
                           plus4A_out(21) => nextA_21_port, plus4A_out(20) => 
                           nextA_20_port, plus4A_out(19) => nextA_19_port, 
                           plus4A_out(18) => nextA_18_port, plus4A_out(17) => 
                           nextA_17_port, plus4A_out(16) => nextA_16_port, 
                           plus4A_out(15) => nextA_15_port, plus4A_out(14) => 
                           nextA_14_port, plus4A_out(13) => nextA_13_port, 
                           plus4A_out(12) => nextA_12_port, plus4A_out(11) => 
                           nextA_11_port, plus4A_out(10) => nextA_10_port, 
                           plus4A_out(9) => nextA_9_port, plus4A_out(8) => 
                           nextA_8_port, plus4A_out(7) => nextA_7_port, 
                           plus4A_out(6) => nextA_6_port, plus4A_out(5) => 
                           nextA_5_port, plus4A_out(4) => nextA_4_port, 
                           plus4A_out(3) => nextA_3_port, plus4A_out(2) => 
                           nextA_2_port, plus4A_out(1) => nextA_1_port, 
                           plus4A_out(0) => n_3185, minus4A_out(63) => 
                           minus4A_s_63_port, minus4A_out(62) => 
                           minus4A_s_62_port, minus4A_out(61) => 
                           minus4A_s_61_port, minus4A_out(60) => 
                           minus4A_s_60_port, minus4A_out(59) => 
                           minus4A_s_59_port, minus4A_out(58) => 
                           minus4A_s_58_port, minus4A_out(57) => 
                           minus4A_s_57_port, minus4A_out(56) => 
                           minus4A_s_56_port, minus4A_out(55) => 
                           minus4A_s_55_port, minus4A_out(54) => 
                           minus4A_s_54_port, minus4A_out(53) => 
                           minus4A_s_53_port, minus4A_out(52) => 
                           minus4A_s_52_port, minus4A_out(51) => 
                           minus4A_s_51_port, minus4A_out(50) => 
                           minus4A_s_50_port, minus4A_out(49) => 
                           minus4A_s_49_port, minus4A_out(48) => 
                           minus4A_s_48_port, minus4A_out(47) => 
                           minus4A_s_47_port, minus4A_out(46) => 
                           minus4A_s_46_port, minus4A_out(45) => 
                           minus4A_s_45_port, minus4A_out(44) => 
                           minus4A_s_44_port, minus4A_out(43) => 
                           minus4A_s_43_port, minus4A_out(42) => 
                           minus4A_s_42_port, minus4A_out(41) => 
                           minus4A_s_41_port, minus4A_out(40) => 
                           minus4A_s_40_port, minus4A_out(39) => 
                           minus4A_s_39_port, minus4A_out(38) => 
                           minus4A_s_38_port, minus4A_out(37) => 
                           minus4A_s_37_port, minus4A_out(36) => 
                           minus4A_s_36_port, minus4A_out(35) => 
                           minus4A_s_35_port, minus4A_out(34) => 
                           minus4A_s_34_port, minus4A_out(33) => 
                           minus4A_s_33_port, minus4A_out(32) => 
                           minus4A_s_32_port, minus4A_out(31) => 
                           minus4A_s_31_port, minus4A_out(30) => 
                           minus4A_s_30_port, minus4A_out(29) => 
                           minus4A_s_29_port, minus4A_out(28) => 
                           minus4A_s_28_port, minus4A_out(27) => 
                           minus4A_s_27_port, minus4A_out(26) => 
                           minus4A_s_26_port, minus4A_out(25) => 
                           minus4A_s_25_port, minus4A_out(24) => 
                           minus4A_s_24_port, minus4A_out(23) => 
                           minus4A_s_23_port, minus4A_out(22) => 
                           minus4A_s_22_port, minus4A_out(21) => 
                           minus4A_s_21_port, minus4A_out(20) => 
                           minus4A_s_20_port, minus4A_out(19) => 
                           minus4A_s_19_port, minus4A_out(18) => 
                           minus4A_s_18_port, minus4A_out(17) => 
                           minus4A_s_17_port, minus4A_out(16) => 
                           minus4A_s_16_port, minus4A_out(15) => 
                           minus4A_s_15_port, minus4A_out(14) => 
                           minus4A_s_14_port, minus4A_out(13) => 
                           minus4A_s_13_port, minus4A_out(12) => 
                           minus4A_s_12_port, minus4A_out(11) => 
                           minus4A_s_11_port, minus4A_out(10) => 
                           minus4A_s_10_port, minus4A_out(9) => 
                           minus4A_s_9_port, minus4A_out(8) => minus4A_s_8_port
                           , minus4A_out(7) => minus4A_s_7_port, minus4A_out(6)
                           => minus4A_s_6_port, minus4A_out(5) => 
                           minus4A_s_5_port, minus4A_out(4) => minus4A_s_4_port
                           , minus4A_out(3) => minus4A_s_3_port, minus4A_out(2)
                           => minus4A_s_2_port, minus4A_out(1) => 
                           minus4A_s_1_port, minus4A_out(0) => minus4A_s_0_port
                           );
   mux_1 : MUX_GENERIC_N64_RADIX3_4 port map( plusA(63) => plus2A_s_63_port, 
                           plusA(62) => plus2A_s_62_port, plusA(61) => 
                           plus2A_s_61_port, plusA(60) => plus2A_s_60_port, 
                           plusA(59) => plus2A_s_59_port, plusA(58) => 
                           plus2A_s_58_port, plusA(57) => plus2A_s_57_port, 
                           plusA(56) => plus2A_s_56_port, plusA(55) => 
                           plus2A_s_55_port, plusA(54) => plus2A_s_54_port, 
                           plusA(53) => plus2A_s_53_port, plusA(52) => 
                           plus2A_s_52_port, plusA(51) => plus2A_s_51_port, 
                           plusA(50) => plus2A_s_50_port, plusA(49) => 
                           plus2A_s_49_port, plusA(48) => plus2A_s_48_port, 
                           plusA(47) => plus2A_s_47_port, plusA(46) => 
                           plus2A_s_46_port, plusA(45) => plus2A_s_45_port, 
                           plusA(44) => plus2A_s_44_port, plusA(43) => 
                           plus2A_s_43_port, plusA(42) => plus2A_s_42_port, 
                           plusA(41) => plus2A_s_41_port, plusA(40) => 
                           plus2A_s_40_port, plusA(39) => plus2A_s_39_port, 
                           plusA(38) => plus2A_s_38_port, plusA(37) => 
                           plus2A_s_37_port, plusA(36) => plus2A_s_36_port, 
                           plusA(35) => plus2A_s_35_port, plusA(34) => 
                           plus2A_s_34_port, plusA(33) => plus2A_s_33_port, 
                           plusA(32) => plus2A_s_32_port, plusA(31) => 
                           plus2A_s_31_port, plusA(30) => plus2A_s_30_port, 
                           plusA(29) => plus2A_s_29_port, plusA(28) => 
                           plus2A_s_28_port, plusA(27) => plus2A_s_27_port, 
                           plusA(26) => plus2A_s_26_port, plusA(25) => 
                           plus2A_s_25_port, plusA(24) => plus2A_s_24_port, 
                           plusA(23) => plus2A_s_23_port, plusA(22) => 
                           plus2A_s_22_port, plusA(21) => plus2A_s_21_port, 
                           plusA(20) => plus2A_s_20_port, plusA(19) => 
                           plus2A_s_19_port, plusA(18) => plus2A_s_18_port, 
                           plusA(17) => plus2A_s_17_port, plusA(16) => 
                           plus2A_s_16_port, plusA(15) => plus2A_s_15_port, 
                           plusA(14) => plus2A_s_14_port, plusA(13) => 
                           plus2A_s_13_port, plusA(12) => plus2A_s_12_port, 
                           plusA(11) => plus2A_s_11_port, plusA(10) => 
                           plus2A_s_10_port, plusA(9) => plus2A_s_9_port, 
                           plusA(8) => plus2A_s_8_port, plusA(7) => 
                           plus2A_s_7_port, plusA(6) => plus2A_s_6_port, 
                           plusA(5) => plus2A_s_5_port, plusA(4) => 
                           plus2A_s_4_port, plusA(3) => plus2A_s_3_port, 
                           plusA(2) => plus2A_s_2_port, plusA(1) => 
                           plus2A_s_1_port, plusA(0) => nextA_0_port, 
                           minusA(63) => minus2A_s_63_port, minusA(62) => 
                           minus2A_s_62_port, minusA(61) => minus2A_s_61_port, 
                           minusA(60) => minus2A_s_60_port, minusA(59) => 
                           minus2A_s_59_port, minusA(58) => minus2A_s_58_port, 
                           minusA(57) => minus2A_s_57_port, minusA(56) => 
                           minus2A_s_56_port, minusA(55) => minus2A_s_55_port, 
                           minusA(54) => minus2A_s_54_port, minusA(53) => 
                           minus2A_s_53_port, minusA(52) => minus2A_s_52_port, 
                           minusA(51) => minus2A_s_51_port, minusA(50) => 
                           minus2A_s_50_port, minusA(49) => minus2A_s_49_port, 
                           minusA(48) => minus2A_s_48_port, minusA(47) => 
                           minus2A_s_47_port, minusA(46) => minus2A_s_46_port, 
                           minusA(45) => minus2A_s_45_port, minusA(44) => 
                           minus2A_s_44_port, minusA(43) => minus2A_s_43_port, 
                           minusA(42) => minus2A_s_42_port, minusA(41) => 
                           minus2A_s_41_port, minusA(40) => minus2A_s_40_port, 
                           minusA(39) => minus2A_s_39_port, minusA(38) => 
                           minus2A_s_38_port, minusA(37) => minus2A_s_37_port, 
                           minusA(36) => minus2A_s_36_port, minusA(35) => 
                           minus2A_s_35_port, minusA(34) => minus2A_s_34_port, 
                           minusA(33) => minus2A_s_33_port, minusA(32) => 
                           minus2A_s_32_port, minusA(31) => minus2A_s_31_port, 
                           minusA(30) => minus2A_s_30_port, minusA(29) => 
                           minus2A_s_29_port, minusA(28) => minus2A_s_28_port, 
                           minusA(27) => minus2A_s_27_port, minusA(26) => 
                           minus2A_s_26_port, minusA(25) => minus2A_s_25_port, 
                           minusA(24) => minus2A_s_24_port, minusA(23) => 
                           minus2A_s_23_port, minusA(22) => minus2A_s_22_port, 
                           minusA(21) => minus2A_s_21_port, minusA(20) => 
                           minus2A_s_20_port, minusA(19) => minus2A_s_19_port, 
                           minusA(18) => minus2A_s_18_port, minusA(17) => 
                           minus2A_s_17_port, minusA(16) => minus2A_s_16_port, 
                           minusA(15) => minus2A_s_15_port, minusA(14) => 
                           minus2A_s_14_port, minusA(13) => minus2A_s_13_port, 
                           minusA(12) => minus2A_s_12_port, minusA(11) => 
                           minus2A_s_11_port, minusA(10) => minus2A_s_10_port, 
                           minusA(9) => minus2A_s_9_port, minusA(8) => 
                           minus2A_s_8_port, minusA(7) => minus2A_s_7_port, 
                           minusA(6) => minus2A_s_6_port, minusA(5) => 
                           minus2A_s_5_port, minusA(4) => minus2A_s_4_port, 
                           minusA(3) => minus2A_s_3_port, minusA(2) => 
                           minus2A_s_2_port, minusA(1) => minus2A_s_1_port, 
                           minusA(0) => minus2A_s_0_port, plus2A(63) => 
                           nextA_63_port, plus2A(62) => nextA_62_port, 
                           plus2A(61) => nextA_61_port, plus2A(60) => 
                           nextA_60_port, plus2A(59) => nextA_59_port, 
                           plus2A(58) => nextA_58_port, plus2A(57) => 
                           nextA_57_port, plus2A(56) => nextA_56_port, 
                           plus2A(55) => nextA_55_port, plus2A(54) => 
                           nextA_54_port, plus2A(53) => nextA_53_port, 
                           plus2A(52) => nextA_52_port, plus2A(51) => 
                           nextA_51_port, plus2A(50) => nextA_50_port, 
                           plus2A(49) => nextA_49_port, plus2A(48) => 
                           nextA_48_port, plus2A(47) => nextA_47_port, 
                           plus2A(46) => nextA_46_port, plus2A(45) => 
                           nextA_45_port, plus2A(44) => nextA_44_port, 
                           plus2A(43) => nextA_43_port, plus2A(42) => 
                           nextA_42_port, plus2A(41) => nextA_41_port, 
                           plus2A(40) => nextA_40_port, plus2A(39) => 
                           nextA_39_port, plus2A(38) => nextA_38_port, 
                           plus2A(37) => nextA_37_port, plus2A(36) => 
                           nextA_36_port, plus2A(35) => nextA_35_port, 
                           plus2A(34) => nextA_34_port, plus2A(33) => 
                           nextA_33_port, plus2A(32) => nextA_32_port, 
                           plus2A(31) => nextA_31_port, plus2A(30) => 
                           nextA_30_port, plus2A(29) => nextA_29_port, 
                           plus2A(28) => nextA_28_port, plus2A(27) => 
                           nextA_27_port, plus2A(26) => nextA_26_port, 
                           plus2A(25) => nextA_25_port, plus2A(24) => 
                           nextA_24_port, plus2A(23) => nextA_23_port, 
                           plus2A(22) => nextA_22_port, plus2A(21) => 
                           nextA_21_port, plus2A(20) => nextA_20_port, 
                           plus2A(19) => nextA_19_port, plus2A(18) => 
                           nextA_18_port, plus2A(17) => nextA_17_port, 
                           plus2A(16) => nextA_16_port, plus2A(15) => 
                           nextA_15_port, plus2A(14) => nextA_14_port, 
                           plus2A(13) => nextA_13_port, plus2A(12) => 
                           nextA_12_port, plus2A(11) => nextA_11_port, 
                           plus2A(10) => nextA_10_port, plus2A(9) => 
                           nextA_9_port, plus2A(8) => nextA_8_port, plus2A(7) 
                           => nextA_7_port, plus2A(6) => nextA_6_port, 
                           plus2A(5) => nextA_5_port, plus2A(4) => nextA_4_port
                           , plus2A(3) => nextA_3_port, plus2A(2) => 
                           nextA_2_port, plus2A(1) => nextA_1_port, plus2A(0) 
                           => nextA_0_port, minus2A(63) => minus4A_s_63_port, 
                           minus2A(62) => minus4A_s_62_port, minus2A(61) => 
                           minus4A_s_61_port, minus2A(60) => minus4A_s_60_port,
                           minus2A(59) => minus4A_s_59_port, minus2A(58) => 
                           minus4A_s_58_port, minus2A(57) => minus4A_s_57_port,
                           minus2A(56) => minus4A_s_56_port, minus2A(55) => 
                           minus4A_s_55_port, minus2A(54) => minus4A_s_54_port,
                           minus2A(53) => minus4A_s_53_port, minus2A(52) => 
                           minus4A_s_52_port, minus2A(51) => minus4A_s_51_port,
                           minus2A(50) => minus4A_s_50_port, minus2A(49) => 
                           minus4A_s_49_port, minus2A(48) => minus4A_s_48_port,
                           minus2A(47) => minus4A_s_47_port, minus2A(46) => 
                           minus4A_s_46_port, minus2A(45) => minus4A_s_45_port,
                           minus2A(44) => minus4A_s_44_port, minus2A(43) => 
                           minus4A_s_43_port, minus2A(42) => minus4A_s_42_port,
                           minus2A(41) => minus4A_s_41_port, minus2A(40) => 
                           minus4A_s_40_port, minus2A(39) => minus4A_s_39_port,
                           minus2A(38) => minus4A_s_38_port, minus2A(37) => 
                           minus4A_s_37_port, minus2A(36) => minus4A_s_36_port,
                           minus2A(35) => minus4A_s_35_port, minus2A(34) => 
                           minus4A_s_34_port, minus2A(33) => minus4A_s_33_port,
                           minus2A(32) => minus4A_s_32_port, minus2A(31) => 
                           minus4A_s_31_port, minus2A(30) => minus4A_s_30_port,
                           minus2A(29) => minus4A_s_29_port, minus2A(28) => 
                           minus4A_s_28_port, minus2A(27) => minus4A_s_27_port,
                           minus2A(26) => minus4A_s_26_port, minus2A(25) => 
                           minus4A_s_25_port, minus2A(24) => minus4A_s_24_port,
                           minus2A(23) => minus4A_s_23_port, minus2A(22) => 
                           minus4A_s_22_port, minus2A(21) => minus4A_s_21_port,
                           minus2A(20) => minus4A_s_20_port, minus2A(19) => 
                           minus4A_s_19_port, minus2A(18) => minus4A_s_18_port,
                           minus2A(17) => minus4A_s_17_port, minus2A(16) => 
                           minus4A_s_16_port, minus2A(15) => minus4A_s_15_port,
                           minus2A(14) => minus4A_s_14_port, minus2A(13) => 
                           minus4A_s_13_port, minus2A(12) => minus4A_s_12_port,
                           minus2A(11) => minus4A_s_11_port, minus2A(10) => 
                           minus4A_s_10_port, minus2A(9) => minus4A_s_9_port, 
                           minus2A(8) => minus4A_s_8_port, minus2A(7) => 
                           minus4A_s_7_port, minus2A(6) => minus4A_s_6_port, 
                           minus2A(5) => minus4A_s_5_port, minus2A(4) => 
                           minus4A_s_4_port, minus2A(3) => minus4A_s_3_port, 
                           minus2A(2) => minus4A_s_2_port, minus2A(1) => 
                           minus4A_s_1_port, minus2A(0) => minus4A_s_0_port, 
                           SEL(2) => encoder_to_mux_2_port, SEL(1) => 
                           encoder_to_mux_1_port, SEL(0) => 
                           encoder_to_mux_0_port, Y(63) => mux_to_adder_63_port
                           , Y(62) => mux_to_adder_62_port, Y(61) => 
                           mux_to_adder_61_port, Y(60) => mux_to_adder_60_port,
                           Y(59) => mux_to_adder_59_port, Y(58) => 
                           mux_to_adder_58_port, Y(57) => mux_to_adder_57_port,
                           Y(56) => mux_to_adder_56_port, Y(55) => 
                           mux_to_adder_55_port, Y(54) => mux_to_adder_54_port,
                           Y(53) => mux_to_adder_53_port, Y(52) => 
                           mux_to_adder_52_port, Y(51) => mux_to_adder_51_port,
                           Y(50) => mux_to_adder_50_port, Y(49) => 
                           mux_to_adder_49_port, Y(48) => mux_to_adder_48_port,
                           Y(47) => mux_to_adder_47_port, Y(46) => 
                           mux_to_adder_46_port, Y(45) => mux_to_adder_45_port,
                           Y(44) => mux_to_adder_44_port, Y(43) => 
                           mux_to_adder_43_port, Y(42) => mux_to_adder_42_port,
                           Y(41) => mux_to_adder_41_port, Y(40) => 
                           mux_to_adder_40_port, Y(39) => mux_to_adder_39_port,
                           Y(38) => mux_to_adder_38_port, Y(37) => 
                           mux_to_adder_37_port, Y(36) => mux_to_adder_36_port,
                           Y(35) => mux_to_adder_35_port, Y(34) => 
                           mux_to_adder_34_port, Y(33) => mux_to_adder_33_port,
                           Y(32) => mux_to_adder_32_port, Y(31) => 
                           mux_to_adder_31_port, Y(30) => mux_to_adder_30_port,
                           Y(29) => mux_to_adder_29_port, Y(28) => 
                           mux_to_adder_28_port, Y(27) => mux_to_adder_27_port,
                           Y(26) => mux_to_adder_26_port, Y(25) => 
                           mux_to_adder_25_port, Y(24) => mux_to_adder_24_port,
                           Y(23) => mux_to_adder_23_port, Y(22) => 
                           mux_to_adder_22_port, Y(21) => mux_to_adder_21_port,
                           Y(20) => mux_to_adder_20_port, Y(19) => 
                           mux_to_adder_19_port, Y(18) => mux_to_adder_18_port,
                           Y(17) => mux_to_adder_17_port, Y(16) => 
                           mux_to_adder_16_port, Y(15) => mux_to_adder_15_port,
                           Y(14) => mux_to_adder_14_port, Y(13) => 
                           mux_to_adder_13_port, Y(12) => mux_to_adder_12_port,
                           Y(11) => mux_to_adder_11_port, Y(10) => 
                           mux_to_adder_10_port, Y(9) => mux_to_adder_9_port, 
                           Y(8) => mux_to_adder_8_port, Y(7) => 
                           mux_to_adder_7_port, Y(6) => mux_to_adder_6_port, 
                           Y(5) => mux_to_adder_5_port, Y(4) => 
                           mux_to_adder_4_port, Y(3) => mux_to_adder_3_port, 
                           Y(2) => mux_to_adder_2_port, Y(1) => 
                           mux_to_adder_1_port, Y(0) => mux_to_adder_0_port);
   rca_1 : RCA_N64_4 port map( A(63) => mux_to_adder_63_port, A(62) => 
                           mux_to_adder_62_port, A(61) => mux_to_adder_61_port,
                           A(60) => mux_to_adder_60_port, A(59) => 
                           mux_to_adder_59_port, A(58) => mux_to_adder_58_port,
                           A(57) => mux_to_adder_57_port, A(56) => 
                           mux_to_adder_56_port, A(55) => mux_to_adder_55_port,
                           A(54) => mux_to_adder_54_port, A(53) => 
                           mux_to_adder_53_port, A(52) => mux_to_adder_52_port,
                           A(51) => mux_to_adder_51_port, A(50) => 
                           mux_to_adder_50_port, A(49) => mux_to_adder_49_port,
                           A(48) => mux_to_adder_48_port, A(47) => 
                           mux_to_adder_47_port, A(46) => mux_to_adder_46_port,
                           A(45) => mux_to_adder_45_port, A(44) => 
                           mux_to_adder_44_port, A(43) => mux_to_adder_43_port,
                           A(42) => mux_to_adder_42_port, A(41) => 
                           mux_to_adder_41_port, A(40) => mux_to_adder_40_port,
                           A(39) => mux_to_adder_39_port, A(38) => 
                           mux_to_adder_38_port, A(37) => mux_to_adder_37_port,
                           A(36) => mux_to_adder_36_port, A(35) => 
                           mux_to_adder_35_port, A(34) => mux_to_adder_34_port,
                           A(33) => mux_to_adder_33_port, A(32) => 
                           mux_to_adder_32_port, A(31) => mux_to_adder_31_port,
                           A(30) => mux_to_adder_30_port, A(29) => 
                           mux_to_adder_29_port, A(28) => mux_to_adder_28_port,
                           A(27) => mux_to_adder_27_port, A(26) => 
                           mux_to_adder_26_port, A(25) => mux_to_adder_25_port,
                           A(24) => mux_to_adder_24_port, A(23) => 
                           mux_to_adder_23_port, A(22) => mux_to_adder_22_port,
                           A(21) => mux_to_adder_21_port, A(20) => 
                           mux_to_adder_20_port, A(19) => mux_to_adder_19_port,
                           A(18) => mux_to_adder_18_port, A(17) => 
                           mux_to_adder_17_port, A(16) => mux_to_adder_16_port,
                           A(15) => mux_to_adder_15_port, A(14) => 
                           mux_to_adder_14_port, A(13) => mux_to_adder_13_port,
                           A(12) => mux_to_adder_12_port, A(11) => 
                           mux_to_adder_11_port, A(10) => mux_to_adder_10_port,
                           A(9) => mux_to_adder_9_port, A(8) => 
                           mux_to_adder_8_port, A(7) => mux_to_adder_7_port, 
                           A(6) => mux_to_adder_6_port, A(5) => 
                           mux_to_adder_5_port, A(4) => mux_to_adder_4_port, 
                           A(3) => mux_to_adder_3_port, A(2) => 
                           mux_to_adder_2_port, A(1) => mux_to_adder_1_port, 
                           A(0) => mux_to_adder_0_port, B(63) => prevSum(63), 
                           B(62) => prevSum(62), B(61) => prevSum(61), B(60) =>
                           prevSum(60), B(59) => prevSum(59), B(58) => 
                           prevSum(58), B(57) => prevSum(57), B(56) => 
                           prevSum(56), B(55) => prevSum(55), B(54) => 
                           prevSum(54), B(53) => prevSum(53), B(52) => 
                           prevSum(52), B(51) => prevSum(51), B(50) => 
                           prevSum(50), B(49) => prevSum(49), B(48) => 
                           prevSum(48), B(47) => prevSum(47), B(46) => 
                           prevSum(46), B(45) => prevSum(45), B(44) => 
                           prevSum(44), B(43) => prevSum(43), B(42) => 
                           prevSum(42), B(41) => prevSum(41), B(40) => 
                           prevSum(40), B(39) => prevSum(39), B(38) => 
                           prevSum(38), B(37) => prevSum(37), B(36) => 
                           prevSum(36), B(35) => prevSum(35), B(34) => 
                           prevSum(34), B(33) => prevSum(33), B(32) => 
                           prevSum(32), B(31) => prevSum(31), B(30) => 
                           prevSum(30), B(29) => prevSum(29), B(28) => 
                           prevSum(28), B(27) => prevSum(27), B(26) => 
                           prevSum(26), B(25) => prevSum(25), B(24) => 
                           prevSum(24), B(23) => prevSum(23), B(22) => 
                           prevSum(22), B(21) => prevSum(21), B(20) => 
                           prevSum(20), B(19) => prevSum(19), B(18) => 
                           prevSum(18), B(17) => prevSum(17), B(16) => 
                           prevSum(16), B(15) => prevSum(15), B(14) => 
                           prevSum(14), B(13) => prevSum(13), B(12) => 
                           prevSum(12), B(11) => prevSum(11), B(10) => 
                           prevSum(10), B(9) => prevSum(9), B(8) => prevSum(8),
                           B(7) => prevSum(7), B(6) => prevSum(6), B(5) => 
                           prevSum(5), B(4) => prevSum(4), B(3) => prevSum(3), 
                           B(2) => prevSum(2), B(1) => prevSum(1), B(0) => 
                           prevSum(0), Ci => X_Logic0_port, S(63) => 
                           nextSum(63), S(62) => nextSum(62), S(61) => 
                           nextSum(61), S(60) => nextSum(60), S(59) => 
                           nextSum(59), S(58) => nextSum(58), S(57) => 
                           nextSum(57), S(56) => nextSum(56), S(55) => 
                           nextSum(55), S(54) => nextSum(54), S(53) => 
                           nextSum(53), S(52) => nextSum(52), S(51) => 
                           nextSum(51), S(50) => nextSum(50), S(49) => 
                           nextSum(49), S(48) => nextSum(48), S(47) => 
                           nextSum(47), S(46) => nextSum(46), S(45) => 
                           nextSum(45), S(44) => nextSum(44), S(43) => 
                           nextSum(43), S(42) => nextSum(42), S(41) => 
                           nextSum(41), S(40) => nextSum(40), S(39) => 
                           nextSum(39), S(38) => nextSum(38), S(37) => 
                           nextSum(37), S(36) => nextSum(36), S(35) => 
                           nextSum(35), S(34) => nextSum(34), S(33) => 
                           nextSum(33), S(32) => nextSum(32), S(31) => 
                           nextSum(31), S(30) => nextSum(30), S(29) => 
                           nextSum(29), S(28) => nextSum(28), S(27) => 
                           nextSum(27), S(26) => nextSum(26), S(25) => 
                           nextSum(25), S(24) => nextSum(24), S(23) => 
                           nextSum(23), S(22) => nextSum(22), S(21) => 
                           nextSum(21), S(20) => nextSum(20), S(19) => 
                           nextSum(19), S(18) => nextSum(18), S(17) => 
                           nextSum(17), S(16) => nextSum(16), S(15) => 
                           nextSum(15), S(14) => nextSum(14), S(13) => 
                           nextSum(13), S(12) => nextSum(12), S(11) => 
                           nextSum(11), S(10) => nextSum(10), S(9) => 
                           nextSum(9), S(8) => nextSum(8), S(7) => nextSum(7), 
                           S(6) => nextSum(6), S(5) => nextSum(5), S(4) => 
                           nextSum(4), S(3) => nextSum(3), S(2) => nextSum(2), 
                           S(1) => nextSum(1), S(0) => nextSum(0), Co => n_3186
                           );
   U3 : BUF_X1 port map( A => n3, Z => nextA_57_port);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity booth_mul_row_N64_RADIX3_5 is

   port( prevA, prevSum : in std_logic_vector (63 downto 0);  encoderIn : in 
         std_logic_vector (2 downto 0);  nextA, nextSum : out std_logic_vector 
         (63 downto 0));

end booth_mul_row_N64_RADIX3_5;

architecture SYN_struct of booth_mul_row_N64_RADIX3_5 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component RCA_N64_5
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component MUX_GENERIC_N64_RADIX3_5
      port( plusA, minusA, plus2A, minus2A : in std_logic_vector (63 downto 0);
            SEL : in std_logic_vector (2 downto 0);  Y : out std_logic_vector 
            (63 downto 0));
   end component;
   
   component ShiftnCompl_N64_5
      port( plusA : in std_logic_vector (63 downto 0);  plus2A_out, minus2A_out
            , plus4A_out, minus4A_out : out std_logic_vector (63 downto 0));
   end component;
   
   component encoder_N64_RADIX3_5
      port( X : in std_logic_vector (2 downto 0);  Z : out std_logic_vector (2 
            downto 0));
   end component;
   
   signal X_Logic0_port, nextA_63_port, nextA_62_port, nextA_61_port, 
      nextA_60_port, nextA_59_port, nextA_58_port, n3, nextA_56_port, 
      nextA_55_port, nextA_54_port, nextA_53_port, nextA_52_port, nextA_51_port
      , nextA_50_port, nextA_49_port, nextA_48_port, nextA_47_port, 
      nextA_46_port, nextA_45_port, nextA_44_port, nextA_43_port, nextA_42_port
      , nextA_41_port, nextA_40_port, nextA_39_port, nextA_38_port, 
      nextA_37_port, nextA_36_port, nextA_35_port, nextA_34_port, nextA_33_port
      , nextA_32_port, nextA_31_port, nextA_30_port, nextA_29_port, 
      nextA_28_port, nextA_27_port, nextA_26_port, nextA_25_port, nextA_24_port
      , nextA_23_port, nextA_22_port, nextA_21_port, nextA_20_port, 
      nextA_19_port, nextA_18_port, nextA_17_port, nextA_16_port, nextA_15_port
      , nextA_14_port, nextA_13_port, nextA_12_port, nextA_11_port, 
      nextA_10_port, nextA_9_port, nextA_8_port, nextA_7_port, nextA_6_port, 
      nextA_5_port, nextA_4_port, nextA_3_port, nextA_2_port, nextA_1_port, 
      encoder_to_mux_2_port, encoder_to_mux_1_port, encoder_to_mux_0_port, 
      plus2A_s_63_port, plus2A_s_62_port, plus2A_s_61_port, plus2A_s_60_port, 
      plus2A_s_59_port, plus2A_s_58_port, plus2A_s_57_port, plus2A_s_56_port, 
      plus2A_s_55_port, plus2A_s_54_port, plus2A_s_53_port, plus2A_s_52_port, 
      plus2A_s_51_port, plus2A_s_50_port, plus2A_s_49_port, plus2A_s_48_port, 
      plus2A_s_47_port, plus2A_s_46_port, plus2A_s_45_port, plus2A_s_44_port, 
      plus2A_s_43_port, plus2A_s_42_port, plus2A_s_41_port, plus2A_s_40_port, 
      plus2A_s_39_port, plus2A_s_38_port, plus2A_s_37_port, plus2A_s_36_port, 
      plus2A_s_35_port, plus2A_s_34_port, plus2A_s_33_port, plus2A_s_32_port, 
      plus2A_s_31_port, plus2A_s_30_port, plus2A_s_29_port, plus2A_s_28_port, 
      plus2A_s_27_port, plus2A_s_26_port, plus2A_s_25_port, plus2A_s_24_port, 
      plus2A_s_23_port, plus2A_s_22_port, plus2A_s_21_port, plus2A_s_20_port, 
      plus2A_s_19_port, plus2A_s_18_port, plus2A_s_17_port, plus2A_s_16_port, 
      plus2A_s_15_port, plus2A_s_14_port, plus2A_s_13_port, plus2A_s_12_port, 
      plus2A_s_11_port, plus2A_s_10_port, plus2A_s_9_port, plus2A_s_8_port, 
      plus2A_s_7_port, plus2A_s_6_port, plus2A_s_5_port, plus2A_s_4_port, 
      plus2A_s_3_port, plus2A_s_2_port, plus2A_s_1_port, minus2A_s_63_port, 
      minus2A_s_62_port, minus2A_s_61_port, minus2A_s_60_port, 
      minus2A_s_59_port, minus2A_s_58_port, minus2A_s_57_port, 
      minus2A_s_56_port, minus2A_s_55_port, minus2A_s_54_port, 
      minus2A_s_53_port, minus2A_s_52_port, minus2A_s_51_port, 
      minus2A_s_50_port, minus2A_s_49_port, minus2A_s_48_port, 
      minus2A_s_47_port, minus2A_s_46_port, minus2A_s_45_port, 
      minus2A_s_44_port, minus2A_s_43_port, minus2A_s_42_port, 
      minus2A_s_41_port, minus2A_s_40_port, minus2A_s_39_port, 
      minus2A_s_38_port, minus2A_s_37_port, minus2A_s_36_port, 
      minus2A_s_35_port, minus2A_s_34_port, minus2A_s_33_port, 
      minus2A_s_32_port, minus2A_s_31_port, minus2A_s_30_port, 
      minus2A_s_29_port, minus2A_s_28_port, minus2A_s_27_port, 
      minus2A_s_26_port, minus2A_s_25_port, minus2A_s_24_port, 
      minus2A_s_23_port, minus2A_s_22_port, minus2A_s_21_port, 
      minus2A_s_20_port, minus2A_s_19_port, minus2A_s_18_port, 
      minus2A_s_17_port, minus2A_s_16_port, minus2A_s_15_port, 
      minus2A_s_14_port, minus2A_s_13_port, minus2A_s_12_port, 
      minus2A_s_11_port, minus2A_s_10_port, minus2A_s_9_port, minus2A_s_8_port,
      minus2A_s_7_port, minus2A_s_6_port, minus2A_s_5_port, minus2A_s_4_port, 
      minus2A_s_3_port, minus2A_s_2_port, minus2A_s_1_port, minus2A_s_0_port, 
      minus4A_s_63_port, minus4A_s_62_port, minus4A_s_61_port, 
      minus4A_s_60_port, minus4A_s_59_port, minus4A_s_58_port, 
      minus4A_s_57_port, minus4A_s_56_port, minus4A_s_55_port, 
      minus4A_s_54_port, minus4A_s_53_port, minus4A_s_52_port, 
      minus4A_s_51_port, minus4A_s_50_port, minus4A_s_49_port, 
      minus4A_s_48_port, minus4A_s_47_port, minus4A_s_46_port, 
      minus4A_s_45_port, minus4A_s_44_port, minus4A_s_43_port, 
      minus4A_s_42_port, minus4A_s_41_port, minus4A_s_40_port, 
      minus4A_s_39_port, minus4A_s_38_port, minus4A_s_37_port, 
      minus4A_s_36_port, minus4A_s_35_port, minus4A_s_34_port, 
      minus4A_s_33_port, minus4A_s_32_port, minus4A_s_31_port, 
      minus4A_s_30_port, minus4A_s_29_port, minus4A_s_28_port, 
      minus4A_s_27_port, minus4A_s_26_port, minus4A_s_25_port, 
      minus4A_s_24_port, minus4A_s_23_port, minus4A_s_22_port, 
      minus4A_s_21_port, minus4A_s_20_port, minus4A_s_19_port, 
      minus4A_s_18_port, minus4A_s_17_port, minus4A_s_16_port, 
      minus4A_s_15_port, minus4A_s_14_port, minus4A_s_13_port, 
      minus4A_s_12_port, minus4A_s_11_port, minus4A_s_10_port, minus4A_s_9_port
      , minus4A_s_8_port, minus4A_s_7_port, minus4A_s_6_port, minus4A_s_5_port,
      minus4A_s_4_port, minus4A_s_3_port, minus4A_s_2_port, minus4A_s_1_port, 
      minus4A_s_0_port, mux_to_adder_63_port, mux_to_adder_62_port, 
      mux_to_adder_61_port, mux_to_adder_60_port, mux_to_adder_59_port, 
      mux_to_adder_58_port, mux_to_adder_57_port, mux_to_adder_56_port, 
      mux_to_adder_55_port, mux_to_adder_54_port, mux_to_adder_53_port, 
      mux_to_adder_52_port, mux_to_adder_51_port, mux_to_adder_50_port, 
      mux_to_adder_49_port, mux_to_adder_48_port, mux_to_adder_47_port, 
      mux_to_adder_46_port, mux_to_adder_45_port, mux_to_adder_44_port, 
      mux_to_adder_43_port, mux_to_adder_42_port, mux_to_adder_41_port, 
      mux_to_adder_40_port, mux_to_adder_39_port, mux_to_adder_38_port, 
      mux_to_adder_37_port, mux_to_adder_36_port, mux_to_adder_35_port, 
      mux_to_adder_34_port, mux_to_adder_33_port, mux_to_adder_32_port, 
      mux_to_adder_31_port, mux_to_adder_30_port, mux_to_adder_29_port, 
      mux_to_adder_28_port, mux_to_adder_27_port, mux_to_adder_26_port, 
      mux_to_adder_25_port, mux_to_adder_24_port, mux_to_adder_23_port, 
      mux_to_adder_22_port, mux_to_adder_21_port, mux_to_adder_20_port, 
      mux_to_adder_19_port, mux_to_adder_18_port, mux_to_adder_17_port, 
      mux_to_adder_16_port, mux_to_adder_15_port, mux_to_adder_14_port, 
      mux_to_adder_13_port, mux_to_adder_12_port, mux_to_adder_11_port, 
      mux_to_adder_10_port, mux_to_adder_9_port, mux_to_adder_8_port, 
      mux_to_adder_7_port, mux_to_adder_6_port, mux_to_adder_5_port, 
      mux_to_adder_4_port, mux_to_adder_3_port, mux_to_adder_2_port, 
      mux_to_adder_1_port, mux_to_adder_0_port, nextA_0_port, nextA_57_port, 
      n_3187, n_3188, n_3189 : std_logic;

begin
   nextA <= ( nextA_63_port, nextA_62_port, nextA_61_port, nextA_60_port, 
      nextA_59_port, nextA_58_port, nextA_57_port, nextA_56_port, nextA_55_port
      , nextA_54_port, nextA_53_port, nextA_52_port, nextA_51_port, 
      nextA_50_port, nextA_49_port, nextA_48_port, nextA_47_port, nextA_46_port
      , nextA_45_port, nextA_44_port, nextA_43_port, nextA_42_port, 
      nextA_41_port, nextA_40_port, nextA_39_port, nextA_38_port, nextA_37_port
      , nextA_36_port, nextA_35_port, nextA_34_port, nextA_33_port, 
      nextA_32_port, nextA_31_port, nextA_30_port, nextA_29_port, nextA_28_port
      , nextA_27_port, nextA_26_port, nextA_25_port, nextA_24_port, 
      nextA_23_port, nextA_22_port, nextA_21_port, nextA_20_port, nextA_19_port
      , nextA_18_port, nextA_17_port, nextA_16_port, nextA_15_port, 
      nextA_14_port, nextA_13_port, nextA_12_port, nextA_11_port, nextA_10_port
      , nextA_9_port, nextA_8_port, nextA_7_port, nextA_6_port, nextA_5_port, 
      nextA_4_port, nextA_3_port, nextA_2_port, nextA_1_port, nextA_0_port );
   
   X_Logic0_port <= '0';
   nextA_0_port <= '0';
   encoder_1 : encoder_N64_RADIX3_5 port map( X(2) => encoderIn(2), X(1) => 
                           encoderIn(1), X(0) => encoderIn(0), Z(2) => 
                           encoder_to_mux_2_port, Z(1) => encoder_to_mux_1_port
                           , Z(0) => encoder_to_mux_0_port);
   ShiftnCompl_1 : ShiftnCompl_N64_5 port map( plusA(63) => prevA(63), 
                           plusA(62) => prevA(62), plusA(61) => prevA(61), 
                           plusA(60) => prevA(60), plusA(59) => prevA(59), 
                           plusA(58) => prevA(58), plusA(57) => prevA(57), 
                           plusA(56) => prevA(56), plusA(55) => prevA(55), 
                           plusA(54) => prevA(54), plusA(53) => prevA(53), 
                           plusA(52) => prevA(52), plusA(51) => prevA(51), 
                           plusA(50) => prevA(50), plusA(49) => prevA(49), 
                           plusA(48) => prevA(48), plusA(47) => prevA(47), 
                           plusA(46) => prevA(46), plusA(45) => prevA(45), 
                           plusA(44) => prevA(44), plusA(43) => prevA(43), 
                           plusA(42) => prevA(42), plusA(41) => prevA(41), 
                           plusA(40) => prevA(40), plusA(39) => prevA(39), 
                           plusA(38) => prevA(38), plusA(37) => prevA(37), 
                           plusA(36) => prevA(36), plusA(35) => prevA(35), 
                           plusA(34) => prevA(34), plusA(33) => prevA(33), 
                           plusA(32) => prevA(32), plusA(31) => prevA(31), 
                           plusA(30) => prevA(30), plusA(29) => prevA(29), 
                           plusA(28) => prevA(28), plusA(27) => prevA(27), 
                           plusA(26) => prevA(26), plusA(25) => prevA(25), 
                           plusA(24) => prevA(24), plusA(23) => prevA(23), 
                           plusA(22) => prevA(22), plusA(21) => prevA(21), 
                           plusA(20) => prevA(20), plusA(19) => prevA(19), 
                           plusA(18) => prevA(18), plusA(17) => prevA(17), 
                           plusA(16) => prevA(16), plusA(15) => prevA(15), 
                           plusA(14) => prevA(14), plusA(13) => prevA(13), 
                           plusA(12) => prevA(12), plusA(11) => prevA(11), 
                           plusA(10) => prevA(10), plusA(9) => prevA(9), 
                           plusA(8) => prevA(8), plusA(7) => prevA(7), plusA(6)
                           => prevA(6), plusA(5) => prevA(5), plusA(4) => 
                           prevA(4), plusA(3) => prevA(3), plusA(2) => prevA(2)
                           , plusA(1) => prevA(1), plusA(0) => prevA(0), 
                           plus2A_out(63) => plus2A_s_63_port, plus2A_out(62) 
                           => plus2A_s_62_port, plus2A_out(61) => 
                           plus2A_s_61_port, plus2A_out(60) => plus2A_s_60_port
                           , plus2A_out(59) => plus2A_s_59_port, plus2A_out(58)
                           => plus2A_s_58_port, plus2A_out(57) => 
                           plus2A_s_57_port, plus2A_out(56) => plus2A_s_56_port
                           , plus2A_out(55) => plus2A_s_55_port, plus2A_out(54)
                           => plus2A_s_54_port, plus2A_out(53) => 
                           plus2A_s_53_port, plus2A_out(52) => plus2A_s_52_port
                           , plus2A_out(51) => plus2A_s_51_port, plus2A_out(50)
                           => plus2A_s_50_port, plus2A_out(49) => 
                           plus2A_s_49_port, plus2A_out(48) => plus2A_s_48_port
                           , plus2A_out(47) => plus2A_s_47_port, plus2A_out(46)
                           => plus2A_s_46_port, plus2A_out(45) => 
                           plus2A_s_45_port, plus2A_out(44) => plus2A_s_44_port
                           , plus2A_out(43) => plus2A_s_43_port, plus2A_out(42)
                           => plus2A_s_42_port, plus2A_out(41) => 
                           plus2A_s_41_port, plus2A_out(40) => plus2A_s_40_port
                           , plus2A_out(39) => plus2A_s_39_port, plus2A_out(38)
                           => plus2A_s_38_port, plus2A_out(37) => 
                           plus2A_s_37_port, plus2A_out(36) => plus2A_s_36_port
                           , plus2A_out(35) => plus2A_s_35_port, plus2A_out(34)
                           => plus2A_s_34_port, plus2A_out(33) => 
                           plus2A_s_33_port, plus2A_out(32) => plus2A_s_32_port
                           , plus2A_out(31) => plus2A_s_31_port, plus2A_out(30)
                           => plus2A_s_30_port, plus2A_out(29) => 
                           plus2A_s_29_port, plus2A_out(28) => plus2A_s_28_port
                           , plus2A_out(27) => plus2A_s_27_port, plus2A_out(26)
                           => plus2A_s_26_port, plus2A_out(25) => 
                           plus2A_s_25_port, plus2A_out(24) => plus2A_s_24_port
                           , plus2A_out(23) => plus2A_s_23_port, plus2A_out(22)
                           => plus2A_s_22_port, plus2A_out(21) => 
                           plus2A_s_21_port, plus2A_out(20) => plus2A_s_20_port
                           , plus2A_out(19) => plus2A_s_19_port, plus2A_out(18)
                           => plus2A_s_18_port, plus2A_out(17) => 
                           plus2A_s_17_port, plus2A_out(16) => plus2A_s_16_port
                           , plus2A_out(15) => plus2A_s_15_port, plus2A_out(14)
                           => plus2A_s_14_port, plus2A_out(13) => 
                           plus2A_s_13_port, plus2A_out(12) => plus2A_s_12_port
                           , plus2A_out(11) => plus2A_s_11_port, plus2A_out(10)
                           => plus2A_s_10_port, plus2A_out(9) => 
                           plus2A_s_9_port, plus2A_out(8) => plus2A_s_8_port, 
                           plus2A_out(7) => plus2A_s_7_port, plus2A_out(6) => 
                           plus2A_s_6_port, plus2A_out(5) => plus2A_s_5_port, 
                           plus2A_out(4) => plus2A_s_4_port, plus2A_out(3) => 
                           plus2A_s_3_port, plus2A_out(2) => plus2A_s_2_port, 
                           plus2A_out(1) => plus2A_s_1_port, plus2A_out(0) => 
                           n_3187, minus2A_out(63) => minus2A_s_63_port, 
                           minus2A_out(62) => minus2A_s_62_port, 
                           minus2A_out(61) => minus2A_s_61_port, 
                           minus2A_out(60) => minus2A_s_60_port, 
                           minus2A_out(59) => minus2A_s_59_port, 
                           minus2A_out(58) => minus2A_s_58_port, 
                           minus2A_out(57) => minus2A_s_57_port, 
                           minus2A_out(56) => minus2A_s_56_port, 
                           minus2A_out(55) => minus2A_s_55_port, 
                           minus2A_out(54) => minus2A_s_54_port, 
                           minus2A_out(53) => minus2A_s_53_port, 
                           minus2A_out(52) => minus2A_s_52_port, 
                           minus2A_out(51) => minus2A_s_51_port, 
                           minus2A_out(50) => minus2A_s_50_port, 
                           minus2A_out(49) => minus2A_s_49_port, 
                           minus2A_out(48) => minus2A_s_48_port, 
                           minus2A_out(47) => minus2A_s_47_port, 
                           minus2A_out(46) => minus2A_s_46_port, 
                           minus2A_out(45) => minus2A_s_45_port, 
                           minus2A_out(44) => minus2A_s_44_port, 
                           minus2A_out(43) => minus2A_s_43_port, 
                           minus2A_out(42) => minus2A_s_42_port, 
                           minus2A_out(41) => minus2A_s_41_port, 
                           minus2A_out(40) => minus2A_s_40_port, 
                           minus2A_out(39) => minus2A_s_39_port, 
                           minus2A_out(38) => minus2A_s_38_port, 
                           minus2A_out(37) => minus2A_s_37_port, 
                           minus2A_out(36) => minus2A_s_36_port, 
                           minus2A_out(35) => minus2A_s_35_port, 
                           minus2A_out(34) => minus2A_s_34_port, 
                           minus2A_out(33) => minus2A_s_33_port, 
                           minus2A_out(32) => minus2A_s_32_port, 
                           minus2A_out(31) => minus2A_s_31_port, 
                           minus2A_out(30) => minus2A_s_30_port, 
                           minus2A_out(29) => minus2A_s_29_port, 
                           minus2A_out(28) => minus2A_s_28_port, 
                           minus2A_out(27) => minus2A_s_27_port, 
                           minus2A_out(26) => minus2A_s_26_port, 
                           minus2A_out(25) => minus2A_s_25_port, 
                           minus2A_out(24) => minus2A_s_24_port, 
                           minus2A_out(23) => minus2A_s_23_port, 
                           minus2A_out(22) => minus2A_s_22_port, 
                           minus2A_out(21) => minus2A_s_21_port, 
                           minus2A_out(20) => minus2A_s_20_port, 
                           minus2A_out(19) => minus2A_s_19_port, 
                           minus2A_out(18) => minus2A_s_18_port, 
                           minus2A_out(17) => minus2A_s_17_port, 
                           minus2A_out(16) => minus2A_s_16_port, 
                           minus2A_out(15) => minus2A_s_15_port, 
                           minus2A_out(14) => minus2A_s_14_port, 
                           minus2A_out(13) => minus2A_s_13_port, 
                           minus2A_out(12) => minus2A_s_12_port, 
                           minus2A_out(11) => minus2A_s_11_port, 
                           minus2A_out(10) => minus2A_s_10_port, minus2A_out(9)
                           => minus2A_s_9_port, minus2A_out(8) => 
                           minus2A_s_8_port, minus2A_out(7) => minus2A_s_7_port
                           , minus2A_out(6) => minus2A_s_6_port, minus2A_out(5)
                           => minus2A_s_5_port, minus2A_out(4) => 
                           minus2A_s_4_port, minus2A_out(3) => minus2A_s_3_port
                           , minus2A_out(2) => minus2A_s_2_port, minus2A_out(1)
                           => minus2A_s_1_port, minus2A_out(0) => 
                           minus2A_s_0_port, plus4A_out(63) => nextA_63_port, 
                           plus4A_out(62) => nextA_62_port, plus4A_out(61) => 
                           nextA_61_port, plus4A_out(60) => nextA_60_port, 
                           plus4A_out(59) => nextA_59_port, plus4A_out(58) => 
                           nextA_58_port, plus4A_out(57) => n3, plus4A_out(56) 
                           => nextA_56_port, plus4A_out(55) => nextA_55_port, 
                           plus4A_out(54) => nextA_54_port, plus4A_out(53) => 
                           nextA_53_port, plus4A_out(52) => nextA_52_port, 
                           plus4A_out(51) => nextA_51_port, plus4A_out(50) => 
                           nextA_50_port, plus4A_out(49) => nextA_49_port, 
                           plus4A_out(48) => nextA_48_port, plus4A_out(47) => 
                           nextA_47_port, plus4A_out(46) => nextA_46_port, 
                           plus4A_out(45) => nextA_45_port, plus4A_out(44) => 
                           nextA_44_port, plus4A_out(43) => nextA_43_port, 
                           plus4A_out(42) => nextA_42_port, plus4A_out(41) => 
                           nextA_41_port, plus4A_out(40) => nextA_40_port, 
                           plus4A_out(39) => nextA_39_port, plus4A_out(38) => 
                           nextA_38_port, plus4A_out(37) => nextA_37_port, 
                           plus4A_out(36) => nextA_36_port, plus4A_out(35) => 
                           nextA_35_port, plus4A_out(34) => nextA_34_port, 
                           plus4A_out(33) => nextA_33_port, plus4A_out(32) => 
                           nextA_32_port, plus4A_out(31) => nextA_31_port, 
                           plus4A_out(30) => nextA_30_port, plus4A_out(29) => 
                           nextA_29_port, plus4A_out(28) => nextA_28_port, 
                           plus4A_out(27) => nextA_27_port, plus4A_out(26) => 
                           nextA_26_port, plus4A_out(25) => nextA_25_port, 
                           plus4A_out(24) => nextA_24_port, plus4A_out(23) => 
                           nextA_23_port, plus4A_out(22) => nextA_22_port, 
                           plus4A_out(21) => nextA_21_port, plus4A_out(20) => 
                           nextA_20_port, plus4A_out(19) => nextA_19_port, 
                           plus4A_out(18) => nextA_18_port, plus4A_out(17) => 
                           nextA_17_port, plus4A_out(16) => nextA_16_port, 
                           plus4A_out(15) => nextA_15_port, plus4A_out(14) => 
                           nextA_14_port, plus4A_out(13) => nextA_13_port, 
                           plus4A_out(12) => nextA_12_port, plus4A_out(11) => 
                           nextA_11_port, plus4A_out(10) => nextA_10_port, 
                           plus4A_out(9) => nextA_9_port, plus4A_out(8) => 
                           nextA_8_port, plus4A_out(7) => nextA_7_port, 
                           plus4A_out(6) => nextA_6_port, plus4A_out(5) => 
                           nextA_5_port, plus4A_out(4) => nextA_4_port, 
                           plus4A_out(3) => nextA_3_port, plus4A_out(2) => 
                           nextA_2_port, plus4A_out(1) => nextA_1_port, 
                           plus4A_out(0) => n_3188, minus4A_out(63) => 
                           minus4A_s_63_port, minus4A_out(62) => 
                           minus4A_s_62_port, minus4A_out(61) => 
                           minus4A_s_61_port, minus4A_out(60) => 
                           minus4A_s_60_port, minus4A_out(59) => 
                           minus4A_s_59_port, minus4A_out(58) => 
                           minus4A_s_58_port, minus4A_out(57) => 
                           minus4A_s_57_port, minus4A_out(56) => 
                           minus4A_s_56_port, minus4A_out(55) => 
                           minus4A_s_55_port, minus4A_out(54) => 
                           minus4A_s_54_port, minus4A_out(53) => 
                           minus4A_s_53_port, minus4A_out(52) => 
                           minus4A_s_52_port, minus4A_out(51) => 
                           minus4A_s_51_port, minus4A_out(50) => 
                           minus4A_s_50_port, minus4A_out(49) => 
                           minus4A_s_49_port, minus4A_out(48) => 
                           minus4A_s_48_port, minus4A_out(47) => 
                           minus4A_s_47_port, minus4A_out(46) => 
                           minus4A_s_46_port, minus4A_out(45) => 
                           minus4A_s_45_port, minus4A_out(44) => 
                           minus4A_s_44_port, minus4A_out(43) => 
                           minus4A_s_43_port, minus4A_out(42) => 
                           minus4A_s_42_port, minus4A_out(41) => 
                           minus4A_s_41_port, minus4A_out(40) => 
                           minus4A_s_40_port, minus4A_out(39) => 
                           minus4A_s_39_port, minus4A_out(38) => 
                           minus4A_s_38_port, minus4A_out(37) => 
                           minus4A_s_37_port, minus4A_out(36) => 
                           minus4A_s_36_port, minus4A_out(35) => 
                           minus4A_s_35_port, minus4A_out(34) => 
                           minus4A_s_34_port, minus4A_out(33) => 
                           minus4A_s_33_port, minus4A_out(32) => 
                           minus4A_s_32_port, minus4A_out(31) => 
                           minus4A_s_31_port, minus4A_out(30) => 
                           minus4A_s_30_port, minus4A_out(29) => 
                           minus4A_s_29_port, minus4A_out(28) => 
                           minus4A_s_28_port, minus4A_out(27) => 
                           minus4A_s_27_port, minus4A_out(26) => 
                           minus4A_s_26_port, minus4A_out(25) => 
                           minus4A_s_25_port, minus4A_out(24) => 
                           minus4A_s_24_port, minus4A_out(23) => 
                           minus4A_s_23_port, minus4A_out(22) => 
                           minus4A_s_22_port, minus4A_out(21) => 
                           minus4A_s_21_port, minus4A_out(20) => 
                           minus4A_s_20_port, minus4A_out(19) => 
                           minus4A_s_19_port, minus4A_out(18) => 
                           minus4A_s_18_port, minus4A_out(17) => 
                           minus4A_s_17_port, minus4A_out(16) => 
                           minus4A_s_16_port, minus4A_out(15) => 
                           minus4A_s_15_port, minus4A_out(14) => 
                           minus4A_s_14_port, minus4A_out(13) => 
                           minus4A_s_13_port, minus4A_out(12) => 
                           minus4A_s_12_port, minus4A_out(11) => 
                           minus4A_s_11_port, minus4A_out(10) => 
                           minus4A_s_10_port, minus4A_out(9) => 
                           minus4A_s_9_port, minus4A_out(8) => minus4A_s_8_port
                           , minus4A_out(7) => minus4A_s_7_port, minus4A_out(6)
                           => minus4A_s_6_port, minus4A_out(5) => 
                           minus4A_s_5_port, minus4A_out(4) => minus4A_s_4_port
                           , minus4A_out(3) => minus4A_s_3_port, minus4A_out(2)
                           => minus4A_s_2_port, minus4A_out(1) => 
                           minus4A_s_1_port, minus4A_out(0) => minus4A_s_0_port
                           );
   mux_1 : MUX_GENERIC_N64_RADIX3_5 port map( plusA(63) => plus2A_s_63_port, 
                           plusA(62) => plus2A_s_62_port, plusA(61) => 
                           plus2A_s_61_port, plusA(60) => plus2A_s_60_port, 
                           plusA(59) => plus2A_s_59_port, plusA(58) => 
                           plus2A_s_58_port, plusA(57) => plus2A_s_57_port, 
                           plusA(56) => plus2A_s_56_port, plusA(55) => 
                           plus2A_s_55_port, plusA(54) => plus2A_s_54_port, 
                           plusA(53) => plus2A_s_53_port, plusA(52) => 
                           plus2A_s_52_port, plusA(51) => plus2A_s_51_port, 
                           plusA(50) => plus2A_s_50_port, plusA(49) => 
                           plus2A_s_49_port, plusA(48) => plus2A_s_48_port, 
                           plusA(47) => plus2A_s_47_port, plusA(46) => 
                           plus2A_s_46_port, plusA(45) => plus2A_s_45_port, 
                           plusA(44) => plus2A_s_44_port, plusA(43) => 
                           plus2A_s_43_port, plusA(42) => plus2A_s_42_port, 
                           plusA(41) => plus2A_s_41_port, plusA(40) => 
                           plus2A_s_40_port, plusA(39) => plus2A_s_39_port, 
                           plusA(38) => plus2A_s_38_port, plusA(37) => 
                           plus2A_s_37_port, plusA(36) => plus2A_s_36_port, 
                           plusA(35) => plus2A_s_35_port, plusA(34) => 
                           plus2A_s_34_port, plusA(33) => plus2A_s_33_port, 
                           plusA(32) => plus2A_s_32_port, plusA(31) => 
                           plus2A_s_31_port, plusA(30) => plus2A_s_30_port, 
                           plusA(29) => plus2A_s_29_port, plusA(28) => 
                           plus2A_s_28_port, plusA(27) => plus2A_s_27_port, 
                           plusA(26) => plus2A_s_26_port, plusA(25) => 
                           plus2A_s_25_port, plusA(24) => plus2A_s_24_port, 
                           plusA(23) => plus2A_s_23_port, plusA(22) => 
                           plus2A_s_22_port, plusA(21) => plus2A_s_21_port, 
                           plusA(20) => plus2A_s_20_port, plusA(19) => 
                           plus2A_s_19_port, plusA(18) => plus2A_s_18_port, 
                           plusA(17) => plus2A_s_17_port, plusA(16) => 
                           plus2A_s_16_port, plusA(15) => plus2A_s_15_port, 
                           plusA(14) => plus2A_s_14_port, plusA(13) => 
                           plus2A_s_13_port, plusA(12) => plus2A_s_12_port, 
                           plusA(11) => plus2A_s_11_port, plusA(10) => 
                           plus2A_s_10_port, plusA(9) => plus2A_s_9_port, 
                           plusA(8) => plus2A_s_8_port, plusA(7) => 
                           plus2A_s_7_port, plusA(6) => plus2A_s_6_port, 
                           plusA(5) => plus2A_s_5_port, plusA(4) => 
                           plus2A_s_4_port, plusA(3) => plus2A_s_3_port, 
                           plusA(2) => plus2A_s_2_port, plusA(1) => 
                           plus2A_s_1_port, plusA(0) => nextA_0_port, 
                           minusA(63) => minus2A_s_63_port, minusA(62) => 
                           minus2A_s_62_port, minusA(61) => minus2A_s_61_port, 
                           minusA(60) => minus2A_s_60_port, minusA(59) => 
                           minus2A_s_59_port, minusA(58) => minus2A_s_58_port, 
                           minusA(57) => minus2A_s_57_port, minusA(56) => 
                           minus2A_s_56_port, minusA(55) => minus2A_s_55_port, 
                           minusA(54) => minus2A_s_54_port, minusA(53) => 
                           minus2A_s_53_port, minusA(52) => minus2A_s_52_port, 
                           minusA(51) => minus2A_s_51_port, minusA(50) => 
                           minus2A_s_50_port, minusA(49) => minus2A_s_49_port, 
                           minusA(48) => minus2A_s_48_port, minusA(47) => 
                           minus2A_s_47_port, minusA(46) => minus2A_s_46_port, 
                           minusA(45) => minus2A_s_45_port, minusA(44) => 
                           minus2A_s_44_port, minusA(43) => minus2A_s_43_port, 
                           minusA(42) => minus2A_s_42_port, minusA(41) => 
                           minus2A_s_41_port, minusA(40) => minus2A_s_40_port, 
                           minusA(39) => minus2A_s_39_port, minusA(38) => 
                           minus2A_s_38_port, minusA(37) => minus2A_s_37_port, 
                           minusA(36) => minus2A_s_36_port, minusA(35) => 
                           minus2A_s_35_port, minusA(34) => minus2A_s_34_port, 
                           minusA(33) => minus2A_s_33_port, minusA(32) => 
                           minus2A_s_32_port, minusA(31) => minus2A_s_31_port, 
                           minusA(30) => minus2A_s_30_port, minusA(29) => 
                           minus2A_s_29_port, minusA(28) => minus2A_s_28_port, 
                           minusA(27) => minus2A_s_27_port, minusA(26) => 
                           minus2A_s_26_port, minusA(25) => minus2A_s_25_port, 
                           minusA(24) => minus2A_s_24_port, minusA(23) => 
                           minus2A_s_23_port, minusA(22) => minus2A_s_22_port, 
                           minusA(21) => minus2A_s_21_port, minusA(20) => 
                           minus2A_s_20_port, minusA(19) => minus2A_s_19_port, 
                           minusA(18) => minus2A_s_18_port, minusA(17) => 
                           minus2A_s_17_port, minusA(16) => minus2A_s_16_port, 
                           minusA(15) => minus2A_s_15_port, minusA(14) => 
                           minus2A_s_14_port, minusA(13) => minus2A_s_13_port, 
                           minusA(12) => minus2A_s_12_port, minusA(11) => 
                           minus2A_s_11_port, minusA(10) => minus2A_s_10_port, 
                           minusA(9) => minus2A_s_9_port, minusA(8) => 
                           minus2A_s_8_port, minusA(7) => minus2A_s_7_port, 
                           minusA(6) => minus2A_s_6_port, minusA(5) => 
                           minus2A_s_5_port, minusA(4) => minus2A_s_4_port, 
                           minusA(3) => minus2A_s_3_port, minusA(2) => 
                           minus2A_s_2_port, minusA(1) => minus2A_s_1_port, 
                           minusA(0) => minus2A_s_0_port, plus2A(63) => 
                           nextA_63_port, plus2A(62) => nextA_62_port, 
                           plus2A(61) => nextA_61_port, plus2A(60) => 
                           nextA_60_port, plus2A(59) => nextA_59_port, 
                           plus2A(58) => nextA_58_port, plus2A(57) => 
                           nextA_57_port, plus2A(56) => nextA_56_port, 
                           plus2A(55) => nextA_55_port, plus2A(54) => 
                           nextA_54_port, plus2A(53) => nextA_53_port, 
                           plus2A(52) => nextA_52_port, plus2A(51) => 
                           nextA_51_port, plus2A(50) => nextA_50_port, 
                           plus2A(49) => nextA_49_port, plus2A(48) => 
                           nextA_48_port, plus2A(47) => nextA_47_port, 
                           plus2A(46) => nextA_46_port, plus2A(45) => 
                           nextA_45_port, plus2A(44) => nextA_44_port, 
                           plus2A(43) => nextA_43_port, plus2A(42) => 
                           nextA_42_port, plus2A(41) => nextA_41_port, 
                           plus2A(40) => nextA_40_port, plus2A(39) => 
                           nextA_39_port, plus2A(38) => nextA_38_port, 
                           plus2A(37) => nextA_37_port, plus2A(36) => 
                           nextA_36_port, plus2A(35) => nextA_35_port, 
                           plus2A(34) => nextA_34_port, plus2A(33) => 
                           nextA_33_port, plus2A(32) => nextA_32_port, 
                           plus2A(31) => nextA_31_port, plus2A(30) => 
                           nextA_30_port, plus2A(29) => nextA_29_port, 
                           plus2A(28) => nextA_28_port, plus2A(27) => 
                           nextA_27_port, plus2A(26) => nextA_26_port, 
                           plus2A(25) => nextA_25_port, plus2A(24) => 
                           nextA_24_port, plus2A(23) => nextA_23_port, 
                           plus2A(22) => nextA_22_port, plus2A(21) => 
                           nextA_21_port, plus2A(20) => nextA_20_port, 
                           plus2A(19) => nextA_19_port, plus2A(18) => 
                           nextA_18_port, plus2A(17) => nextA_17_port, 
                           plus2A(16) => nextA_16_port, plus2A(15) => 
                           nextA_15_port, plus2A(14) => nextA_14_port, 
                           plus2A(13) => nextA_13_port, plus2A(12) => 
                           nextA_12_port, plus2A(11) => nextA_11_port, 
                           plus2A(10) => nextA_10_port, plus2A(9) => 
                           nextA_9_port, plus2A(8) => nextA_8_port, plus2A(7) 
                           => nextA_7_port, plus2A(6) => nextA_6_port, 
                           plus2A(5) => nextA_5_port, plus2A(4) => nextA_4_port
                           , plus2A(3) => nextA_3_port, plus2A(2) => 
                           nextA_2_port, plus2A(1) => nextA_1_port, plus2A(0) 
                           => nextA_0_port, minus2A(63) => minus4A_s_63_port, 
                           minus2A(62) => minus4A_s_62_port, minus2A(61) => 
                           minus4A_s_61_port, minus2A(60) => minus4A_s_60_port,
                           minus2A(59) => minus4A_s_59_port, minus2A(58) => 
                           minus4A_s_58_port, minus2A(57) => minus4A_s_57_port,
                           minus2A(56) => minus4A_s_56_port, minus2A(55) => 
                           minus4A_s_55_port, minus2A(54) => minus4A_s_54_port,
                           minus2A(53) => minus4A_s_53_port, minus2A(52) => 
                           minus4A_s_52_port, minus2A(51) => minus4A_s_51_port,
                           minus2A(50) => minus4A_s_50_port, minus2A(49) => 
                           minus4A_s_49_port, minus2A(48) => minus4A_s_48_port,
                           minus2A(47) => minus4A_s_47_port, minus2A(46) => 
                           minus4A_s_46_port, minus2A(45) => minus4A_s_45_port,
                           minus2A(44) => minus4A_s_44_port, minus2A(43) => 
                           minus4A_s_43_port, minus2A(42) => minus4A_s_42_port,
                           minus2A(41) => minus4A_s_41_port, minus2A(40) => 
                           minus4A_s_40_port, minus2A(39) => minus4A_s_39_port,
                           minus2A(38) => minus4A_s_38_port, minus2A(37) => 
                           minus4A_s_37_port, minus2A(36) => minus4A_s_36_port,
                           minus2A(35) => minus4A_s_35_port, minus2A(34) => 
                           minus4A_s_34_port, minus2A(33) => minus4A_s_33_port,
                           minus2A(32) => minus4A_s_32_port, minus2A(31) => 
                           minus4A_s_31_port, minus2A(30) => minus4A_s_30_port,
                           minus2A(29) => minus4A_s_29_port, minus2A(28) => 
                           minus4A_s_28_port, minus2A(27) => minus4A_s_27_port,
                           minus2A(26) => minus4A_s_26_port, minus2A(25) => 
                           minus4A_s_25_port, minus2A(24) => minus4A_s_24_port,
                           minus2A(23) => minus4A_s_23_port, minus2A(22) => 
                           minus4A_s_22_port, minus2A(21) => minus4A_s_21_port,
                           minus2A(20) => minus4A_s_20_port, minus2A(19) => 
                           minus4A_s_19_port, minus2A(18) => minus4A_s_18_port,
                           minus2A(17) => minus4A_s_17_port, minus2A(16) => 
                           minus4A_s_16_port, minus2A(15) => minus4A_s_15_port,
                           minus2A(14) => minus4A_s_14_port, minus2A(13) => 
                           minus4A_s_13_port, minus2A(12) => minus4A_s_12_port,
                           minus2A(11) => minus4A_s_11_port, minus2A(10) => 
                           minus4A_s_10_port, minus2A(9) => minus4A_s_9_port, 
                           minus2A(8) => minus4A_s_8_port, minus2A(7) => 
                           minus4A_s_7_port, minus2A(6) => minus4A_s_6_port, 
                           minus2A(5) => minus4A_s_5_port, minus2A(4) => 
                           minus4A_s_4_port, minus2A(3) => minus4A_s_3_port, 
                           minus2A(2) => minus4A_s_2_port, minus2A(1) => 
                           minus4A_s_1_port, minus2A(0) => minus4A_s_0_port, 
                           SEL(2) => encoder_to_mux_2_port, SEL(1) => 
                           encoder_to_mux_1_port, SEL(0) => 
                           encoder_to_mux_0_port, Y(63) => mux_to_adder_63_port
                           , Y(62) => mux_to_adder_62_port, Y(61) => 
                           mux_to_adder_61_port, Y(60) => mux_to_adder_60_port,
                           Y(59) => mux_to_adder_59_port, Y(58) => 
                           mux_to_adder_58_port, Y(57) => mux_to_adder_57_port,
                           Y(56) => mux_to_adder_56_port, Y(55) => 
                           mux_to_adder_55_port, Y(54) => mux_to_adder_54_port,
                           Y(53) => mux_to_adder_53_port, Y(52) => 
                           mux_to_adder_52_port, Y(51) => mux_to_adder_51_port,
                           Y(50) => mux_to_adder_50_port, Y(49) => 
                           mux_to_adder_49_port, Y(48) => mux_to_adder_48_port,
                           Y(47) => mux_to_adder_47_port, Y(46) => 
                           mux_to_adder_46_port, Y(45) => mux_to_adder_45_port,
                           Y(44) => mux_to_adder_44_port, Y(43) => 
                           mux_to_adder_43_port, Y(42) => mux_to_adder_42_port,
                           Y(41) => mux_to_adder_41_port, Y(40) => 
                           mux_to_adder_40_port, Y(39) => mux_to_adder_39_port,
                           Y(38) => mux_to_adder_38_port, Y(37) => 
                           mux_to_adder_37_port, Y(36) => mux_to_adder_36_port,
                           Y(35) => mux_to_adder_35_port, Y(34) => 
                           mux_to_adder_34_port, Y(33) => mux_to_adder_33_port,
                           Y(32) => mux_to_adder_32_port, Y(31) => 
                           mux_to_adder_31_port, Y(30) => mux_to_adder_30_port,
                           Y(29) => mux_to_adder_29_port, Y(28) => 
                           mux_to_adder_28_port, Y(27) => mux_to_adder_27_port,
                           Y(26) => mux_to_adder_26_port, Y(25) => 
                           mux_to_adder_25_port, Y(24) => mux_to_adder_24_port,
                           Y(23) => mux_to_adder_23_port, Y(22) => 
                           mux_to_adder_22_port, Y(21) => mux_to_adder_21_port,
                           Y(20) => mux_to_adder_20_port, Y(19) => 
                           mux_to_adder_19_port, Y(18) => mux_to_adder_18_port,
                           Y(17) => mux_to_adder_17_port, Y(16) => 
                           mux_to_adder_16_port, Y(15) => mux_to_adder_15_port,
                           Y(14) => mux_to_adder_14_port, Y(13) => 
                           mux_to_adder_13_port, Y(12) => mux_to_adder_12_port,
                           Y(11) => mux_to_adder_11_port, Y(10) => 
                           mux_to_adder_10_port, Y(9) => mux_to_adder_9_port, 
                           Y(8) => mux_to_adder_8_port, Y(7) => 
                           mux_to_adder_7_port, Y(6) => mux_to_adder_6_port, 
                           Y(5) => mux_to_adder_5_port, Y(4) => 
                           mux_to_adder_4_port, Y(3) => mux_to_adder_3_port, 
                           Y(2) => mux_to_adder_2_port, Y(1) => 
                           mux_to_adder_1_port, Y(0) => mux_to_adder_0_port);
   rca_1 : RCA_N64_5 port map( A(63) => mux_to_adder_63_port, A(62) => 
                           mux_to_adder_62_port, A(61) => mux_to_adder_61_port,
                           A(60) => mux_to_adder_60_port, A(59) => 
                           mux_to_adder_59_port, A(58) => mux_to_adder_58_port,
                           A(57) => mux_to_adder_57_port, A(56) => 
                           mux_to_adder_56_port, A(55) => mux_to_adder_55_port,
                           A(54) => mux_to_adder_54_port, A(53) => 
                           mux_to_adder_53_port, A(52) => mux_to_adder_52_port,
                           A(51) => mux_to_adder_51_port, A(50) => 
                           mux_to_adder_50_port, A(49) => mux_to_adder_49_port,
                           A(48) => mux_to_adder_48_port, A(47) => 
                           mux_to_adder_47_port, A(46) => mux_to_adder_46_port,
                           A(45) => mux_to_adder_45_port, A(44) => 
                           mux_to_adder_44_port, A(43) => mux_to_adder_43_port,
                           A(42) => mux_to_adder_42_port, A(41) => 
                           mux_to_adder_41_port, A(40) => mux_to_adder_40_port,
                           A(39) => mux_to_adder_39_port, A(38) => 
                           mux_to_adder_38_port, A(37) => mux_to_adder_37_port,
                           A(36) => mux_to_adder_36_port, A(35) => 
                           mux_to_adder_35_port, A(34) => mux_to_adder_34_port,
                           A(33) => mux_to_adder_33_port, A(32) => 
                           mux_to_adder_32_port, A(31) => mux_to_adder_31_port,
                           A(30) => mux_to_adder_30_port, A(29) => 
                           mux_to_adder_29_port, A(28) => mux_to_adder_28_port,
                           A(27) => mux_to_adder_27_port, A(26) => 
                           mux_to_adder_26_port, A(25) => mux_to_adder_25_port,
                           A(24) => mux_to_adder_24_port, A(23) => 
                           mux_to_adder_23_port, A(22) => mux_to_adder_22_port,
                           A(21) => mux_to_adder_21_port, A(20) => 
                           mux_to_adder_20_port, A(19) => mux_to_adder_19_port,
                           A(18) => mux_to_adder_18_port, A(17) => 
                           mux_to_adder_17_port, A(16) => mux_to_adder_16_port,
                           A(15) => mux_to_adder_15_port, A(14) => 
                           mux_to_adder_14_port, A(13) => mux_to_adder_13_port,
                           A(12) => mux_to_adder_12_port, A(11) => 
                           mux_to_adder_11_port, A(10) => mux_to_adder_10_port,
                           A(9) => mux_to_adder_9_port, A(8) => 
                           mux_to_adder_8_port, A(7) => mux_to_adder_7_port, 
                           A(6) => mux_to_adder_6_port, A(5) => 
                           mux_to_adder_5_port, A(4) => mux_to_adder_4_port, 
                           A(3) => mux_to_adder_3_port, A(2) => 
                           mux_to_adder_2_port, A(1) => mux_to_adder_1_port, 
                           A(0) => mux_to_adder_0_port, B(63) => prevSum(63), 
                           B(62) => prevSum(62), B(61) => prevSum(61), B(60) =>
                           prevSum(60), B(59) => prevSum(59), B(58) => 
                           prevSum(58), B(57) => prevSum(57), B(56) => 
                           prevSum(56), B(55) => prevSum(55), B(54) => 
                           prevSum(54), B(53) => prevSum(53), B(52) => 
                           prevSum(52), B(51) => prevSum(51), B(50) => 
                           prevSum(50), B(49) => prevSum(49), B(48) => 
                           prevSum(48), B(47) => prevSum(47), B(46) => 
                           prevSum(46), B(45) => prevSum(45), B(44) => 
                           prevSum(44), B(43) => prevSum(43), B(42) => 
                           prevSum(42), B(41) => prevSum(41), B(40) => 
                           prevSum(40), B(39) => prevSum(39), B(38) => 
                           prevSum(38), B(37) => prevSum(37), B(36) => 
                           prevSum(36), B(35) => prevSum(35), B(34) => 
                           prevSum(34), B(33) => prevSum(33), B(32) => 
                           prevSum(32), B(31) => prevSum(31), B(30) => 
                           prevSum(30), B(29) => prevSum(29), B(28) => 
                           prevSum(28), B(27) => prevSum(27), B(26) => 
                           prevSum(26), B(25) => prevSum(25), B(24) => 
                           prevSum(24), B(23) => prevSum(23), B(22) => 
                           prevSum(22), B(21) => prevSum(21), B(20) => 
                           prevSum(20), B(19) => prevSum(19), B(18) => 
                           prevSum(18), B(17) => prevSum(17), B(16) => 
                           prevSum(16), B(15) => prevSum(15), B(14) => 
                           prevSum(14), B(13) => prevSum(13), B(12) => 
                           prevSum(12), B(11) => prevSum(11), B(10) => 
                           prevSum(10), B(9) => prevSum(9), B(8) => prevSum(8),
                           B(7) => prevSum(7), B(6) => prevSum(6), B(5) => 
                           prevSum(5), B(4) => prevSum(4), B(3) => prevSum(3), 
                           B(2) => prevSum(2), B(1) => prevSum(1), B(0) => 
                           prevSum(0), Ci => X_Logic0_port, S(63) => 
                           nextSum(63), S(62) => nextSum(62), S(61) => 
                           nextSum(61), S(60) => nextSum(60), S(59) => 
                           nextSum(59), S(58) => nextSum(58), S(57) => 
                           nextSum(57), S(56) => nextSum(56), S(55) => 
                           nextSum(55), S(54) => nextSum(54), S(53) => 
                           nextSum(53), S(52) => nextSum(52), S(51) => 
                           nextSum(51), S(50) => nextSum(50), S(49) => 
                           nextSum(49), S(48) => nextSum(48), S(47) => 
                           nextSum(47), S(46) => nextSum(46), S(45) => 
                           nextSum(45), S(44) => nextSum(44), S(43) => 
                           nextSum(43), S(42) => nextSum(42), S(41) => 
                           nextSum(41), S(40) => nextSum(40), S(39) => 
                           nextSum(39), S(38) => nextSum(38), S(37) => 
                           nextSum(37), S(36) => nextSum(36), S(35) => 
                           nextSum(35), S(34) => nextSum(34), S(33) => 
                           nextSum(33), S(32) => nextSum(32), S(31) => 
                           nextSum(31), S(30) => nextSum(30), S(29) => 
                           nextSum(29), S(28) => nextSum(28), S(27) => 
                           nextSum(27), S(26) => nextSum(26), S(25) => 
                           nextSum(25), S(24) => nextSum(24), S(23) => 
                           nextSum(23), S(22) => nextSum(22), S(21) => 
                           nextSum(21), S(20) => nextSum(20), S(19) => 
                           nextSum(19), S(18) => nextSum(18), S(17) => 
                           nextSum(17), S(16) => nextSum(16), S(15) => 
                           nextSum(15), S(14) => nextSum(14), S(13) => 
                           nextSum(13), S(12) => nextSum(12), S(11) => 
                           nextSum(11), S(10) => nextSum(10), S(9) => 
                           nextSum(9), S(8) => nextSum(8), S(7) => nextSum(7), 
                           S(6) => nextSum(6), S(5) => nextSum(5), S(4) => 
                           nextSum(4), S(3) => nextSum(3), S(2) => nextSum(2), 
                           S(1) => nextSum(1), S(0) => nextSum(0), Co => n_3189
                           );
   U3 : BUF_X1 port map( A => n3, Z => nextA_57_port);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity booth_mul_row_N64_RADIX3_6 is

   port( prevA, prevSum : in std_logic_vector (63 downto 0);  encoderIn : in 
         std_logic_vector (2 downto 0);  nextA, nextSum : out std_logic_vector 
         (63 downto 0));

end booth_mul_row_N64_RADIX3_6;

architecture SYN_struct of booth_mul_row_N64_RADIX3_6 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component RCA_N64_6
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component MUX_GENERIC_N64_RADIX3_6
      port( plusA, minusA, plus2A, minus2A : in std_logic_vector (63 downto 0);
            SEL : in std_logic_vector (2 downto 0);  Y : out std_logic_vector 
            (63 downto 0));
   end component;
   
   component ShiftnCompl_N64_6
      port( plusA : in std_logic_vector (63 downto 0);  plus2A_out, minus2A_out
            , plus4A_out, minus4A_out : out std_logic_vector (63 downto 0));
   end component;
   
   component encoder_N64_RADIX3_6
      port( X : in std_logic_vector (2 downto 0);  Z : out std_logic_vector (2 
            downto 0));
   end component;
   
   signal X_Logic0_port, nextA_63_port, nextA_62_port, nextA_61_port, 
      nextA_60_port, nextA_59_port, nextA_58_port, n3, nextA_56_port, 
      nextA_55_port, nextA_54_port, nextA_53_port, nextA_52_port, nextA_51_port
      , nextA_50_port, nextA_49_port, nextA_48_port, nextA_47_port, 
      nextA_46_port, nextA_45_port, nextA_44_port, nextA_43_port, nextA_42_port
      , nextA_41_port, nextA_40_port, nextA_39_port, nextA_38_port, 
      nextA_37_port, nextA_36_port, nextA_35_port, nextA_34_port, nextA_33_port
      , nextA_32_port, nextA_31_port, nextA_30_port, nextA_29_port, 
      nextA_28_port, nextA_27_port, nextA_26_port, nextA_25_port, nextA_24_port
      , nextA_23_port, nextA_22_port, nextA_21_port, nextA_20_port, 
      nextA_19_port, nextA_18_port, nextA_17_port, nextA_16_port, nextA_15_port
      , nextA_14_port, nextA_13_port, nextA_12_port, nextA_11_port, 
      nextA_10_port, nextA_9_port, nextA_8_port, nextA_7_port, nextA_6_port, 
      nextA_5_port, nextA_4_port, nextA_3_port, nextA_2_port, nextA_1_port, 
      encoder_to_mux_2_port, encoder_to_mux_1_port, encoder_to_mux_0_port, 
      plus2A_s_63_port, plus2A_s_62_port, plus2A_s_61_port, plus2A_s_60_port, 
      plus2A_s_59_port, plus2A_s_58_port, plus2A_s_57_port, plus2A_s_56_port, 
      plus2A_s_55_port, plus2A_s_54_port, plus2A_s_53_port, plus2A_s_52_port, 
      plus2A_s_51_port, plus2A_s_50_port, plus2A_s_49_port, plus2A_s_48_port, 
      plus2A_s_47_port, plus2A_s_46_port, plus2A_s_45_port, plus2A_s_44_port, 
      plus2A_s_43_port, plus2A_s_42_port, plus2A_s_41_port, plus2A_s_40_port, 
      plus2A_s_39_port, plus2A_s_38_port, plus2A_s_37_port, plus2A_s_36_port, 
      plus2A_s_35_port, plus2A_s_34_port, plus2A_s_33_port, plus2A_s_32_port, 
      plus2A_s_31_port, plus2A_s_30_port, plus2A_s_29_port, plus2A_s_28_port, 
      plus2A_s_27_port, plus2A_s_26_port, plus2A_s_25_port, plus2A_s_24_port, 
      plus2A_s_23_port, plus2A_s_22_port, plus2A_s_21_port, plus2A_s_20_port, 
      plus2A_s_19_port, plus2A_s_18_port, plus2A_s_17_port, plus2A_s_16_port, 
      plus2A_s_15_port, plus2A_s_14_port, plus2A_s_13_port, plus2A_s_12_port, 
      plus2A_s_11_port, plus2A_s_10_port, plus2A_s_9_port, plus2A_s_8_port, 
      plus2A_s_7_port, plus2A_s_6_port, plus2A_s_5_port, plus2A_s_4_port, 
      plus2A_s_3_port, plus2A_s_2_port, plus2A_s_1_port, minus2A_s_63_port, 
      minus2A_s_62_port, minus2A_s_61_port, minus2A_s_60_port, 
      minus2A_s_59_port, minus2A_s_58_port, minus2A_s_57_port, 
      minus2A_s_56_port, minus2A_s_55_port, minus2A_s_54_port, 
      minus2A_s_53_port, minus2A_s_52_port, minus2A_s_51_port, 
      minus2A_s_50_port, minus2A_s_49_port, minus2A_s_48_port, 
      minus2A_s_47_port, minus2A_s_46_port, minus2A_s_45_port, 
      minus2A_s_44_port, minus2A_s_43_port, minus2A_s_42_port, 
      minus2A_s_41_port, minus2A_s_40_port, minus2A_s_39_port, 
      minus2A_s_38_port, minus2A_s_37_port, minus2A_s_36_port, 
      minus2A_s_35_port, minus2A_s_34_port, minus2A_s_33_port, 
      minus2A_s_32_port, minus2A_s_31_port, minus2A_s_30_port, 
      minus2A_s_29_port, minus2A_s_28_port, minus2A_s_27_port, 
      minus2A_s_26_port, minus2A_s_25_port, minus2A_s_24_port, 
      minus2A_s_23_port, minus2A_s_22_port, minus2A_s_21_port, 
      minus2A_s_20_port, minus2A_s_19_port, minus2A_s_18_port, 
      minus2A_s_17_port, minus2A_s_16_port, minus2A_s_15_port, 
      minus2A_s_14_port, minus2A_s_13_port, minus2A_s_12_port, 
      minus2A_s_11_port, minus2A_s_10_port, minus2A_s_9_port, minus2A_s_8_port,
      minus2A_s_7_port, minus2A_s_6_port, minus2A_s_5_port, minus2A_s_4_port, 
      minus2A_s_3_port, minus2A_s_2_port, minus2A_s_1_port, minus2A_s_0_port, 
      minus4A_s_63_port, minus4A_s_62_port, minus4A_s_61_port, 
      minus4A_s_60_port, minus4A_s_59_port, minus4A_s_58_port, 
      minus4A_s_57_port, minus4A_s_56_port, minus4A_s_55_port, 
      minus4A_s_54_port, minus4A_s_53_port, minus4A_s_52_port, 
      minus4A_s_51_port, minus4A_s_50_port, minus4A_s_49_port, 
      minus4A_s_48_port, minus4A_s_47_port, minus4A_s_46_port, 
      minus4A_s_45_port, minus4A_s_44_port, minus4A_s_43_port, 
      minus4A_s_42_port, minus4A_s_41_port, minus4A_s_40_port, 
      minus4A_s_39_port, minus4A_s_38_port, minus4A_s_37_port, 
      minus4A_s_36_port, minus4A_s_35_port, minus4A_s_34_port, 
      minus4A_s_33_port, minus4A_s_32_port, minus4A_s_31_port, 
      minus4A_s_30_port, minus4A_s_29_port, minus4A_s_28_port, 
      minus4A_s_27_port, minus4A_s_26_port, minus4A_s_25_port, 
      minus4A_s_24_port, minus4A_s_23_port, minus4A_s_22_port, 
      minus4A_s_21_port, minus4A_s_20_port, minus4A_s_19_port, 
      minus4A_s_18_port, minus4A_s_17_port, minus4A_s_16_port, 
      minus4A_s_15_port, minus4A_s_14_port, minus4A_s_13_port, 
      minus4A_s_12_port, minus4A_s_11_port, minus4A_s_10_port, minus4A_s_9_port
      , minus4A_s_8_port, minus4A_s_7_port, minus4A_s_6_port, minus4A_s_5_port,
      minus4A_s_4_port, minus4A_s_3_port, minus4A_s_2_port, minus4A_s_1_port, 
      minus4A_s_0_port, mux_to_adder_63_port, mux_to_adder_62_port, 
      mux_to_adder_61_port, mux_to_adder_60_port, mux_to_adder_59_port, 
      mux_to_adder_58_port, mux_to_adder_57_port, mux_to_adder_56_port, 
      mux_to_adder_55_port, mux_to_adder_54_port, mux_to_adder_53_port, 
      mux_to_adder_52_port, mux_to_adder_51_port, mux_to_adder_50_port, 
      mux_to_adder_49_port, mux_to_adder_48_port, mux_to_adder_47_port, 
      mux_to_adder_46_port, mux_to_adder_45_port, mux_to_adder_44_port, 
      mux_to_adder_43_port, mux_to_adder_42_port, mux_to_adder_41_port, 
      mux_to_adder_40_port, mux_to_adder_39_port, mux_to_adder_38_port, 
      mux_to_adder_37_port, mux_to_adder_36_port, mux_to_adder_35_port, 
      mux_to_adder_34_port, mux_to_adder_33_port, mux_to_adder_32_port, 
      mux_to_adder_31_port, mux_to_adder_30_port, mux_to_adder_29_port, 
      mux_to_adder_28_port, mux_to_adder_27_port, mux_to_adder_26_port, 
      mux_to_adder_25_port, mux_to_adder_24_port, mux_to_adder_23_port, 
      mux_to_adder_22_port, mux_to_adder_21_port, mux_to_adder_20_port, 
      mux_to_adder_19_port, mux_to_adder_18_port, mux_to_adder_17_port, 
      mux_to_adder_16_port, mux_to_adder_15_port, mux_to_adder_14_port, 
      mux_to_adder_13_port, mux_to_adder_12_port, mux_to_adder_11_port, 
      mux_to_adder_10_port, mux_to_adder_9_port, mux_to_adder_8_port, 
      mux_to_adder_7_port, mux_to_adder_6_port, mux_to_adder_5_port, 
      mux_to_adder_4_port, mux_to_adder_3_port, mux_to_adder_2_port, 
      mux_to_adder_1_port, mux_to_adder_0_port, nextA_0_port, nextA_57_port, 
      n_3190, n_3191, n_3192 : std_logic;

begin
   nextA <= ( nextA_63_port, nextA_62_port, nextA_61_port, nextA_60_port, 
      nextA_59_port, nextA_58_port, nextA_57_port, nextA_56_port, nextA_55_port
      , nextA_54_port, nextA_53_port, nextA_52_port, nextA_51_port, 
      nextA_50_port, nextA_49_port, nextA_48_port, nextA_47_port, nextA_46_port
      , nextA_45_port, nextA_44_port, nextA_43_port, nextA_42_port, 
      nextA_41_port, nextA_40_port, nextA_39_port, nextA_38_port, nextA_37_port
      , nextA_36_port, nextA_35_port, nextA_34_port, nextA_33_port, 
      nextA_32_port, nextA_31_port, nextA_30_port, nextA_29_port, nextA_28_port
      , nextA_27_port, nextA_26_port, nextA_25_port, nextA_24_port, 
      nextA_23_port, nextA_22_port, nextA_21_port, nextA_20_port, nextA_19_port
      , nextA_18_port, nextA_17_port, nextA_16_port, nextA_15_port, 
      nextA_14_port, nextA_13_port, nextA_12_port, nextA_11_port, nextA_10_port
      , nextA_9_port, nextA_8_port, nextA_7_port, nextA_6_port, nextA_5_port, 
      nextA_4_port, nextA_3_port, nextA_2_port, nextA_1_port, nextA_0_port );
   
   X_Logic0_port <= '0';
   nextA_0_port <= '0';
   encoder_1 : encoder_N64_RADIX3_6 port map( X(2) => encoderIn(2), X(1) => 
                           encoderIn(1), X(0) => encoderIn(0), Z(2) => 
                           encoder_to_mux_2_port, Z(1) => encoder_to_mux_1_port
                           , Z(0) => encoder_to_mux_0_port);
   ShiftnCompl_1 : ShiftnCompl_N64_6 port map( plusA(63) => prevA(63), 
                           plusA(62) => prevA(62), plusA(61) => prevA(61), 
                           plusA(60) => prevA(60), plusA(59) => prevA(59), 
                           plusA(58) => prevA(58), plusA(57) => prevA(57), 
                           plusA(56) => prevA(56), plusA(55) => prevA(55), 
                           plusA(54) => prevA(54), plusA(53) => prevA(53), 
                           plusA(52) => prevA(52), plusA(51) => prevA(51), 
                           plusA(50) => prevA(50), plusA(49) => prevA(49), 
                           plusA(48) => prevA(48), plusA(47) => prevA(47), 
                           plusA(46) => prevA(46), plusA(45) => prevA(45), 
                           plusA(44) => prevA(44), plusA(43) => prevA(43), 
                           plusA(42) => prevA(42), plusA(41) => prevA(41), 
                           plusA(40) => prevA(40), plusA(39) => prevA(39), 
                           plusA(38) => prevA(38), plusA(37) => prevA(37), 
                           plusA(36) => prevA(36), plusA(35) => prevA(35), 
                           plusA(34) => prevA(34), plusA(33) => prevA(33), 
                           plusA(32) => prevA(32), plusA(31) => prevA(31), 
                           plusA(30) => prevA(30), plusA(29) => prevA(29), 
                           plusA(28) => prevA(28), plusA(27) => prevA(27), 
                           plusA(26) => prevA(26), plusA(25) => prevA(25), 
                           plusA(24) => prevA(24), plusA(23) => prevA(23), 
                           plusA(22) => prevA(22), plusA(21) => prevA(21), 
                           plusA(20) => prevA(20), plusA(19) => prevA(19), 
                           plusA(18) => prevA(18), plusA(17) => prevA(17), 
                           plusA(16) => prevA(16), plusA(15) => prevA(15), 
                           plusA(14) => prevA(14), plusA(13) => prevA(13), 
                           plusA(12) => prevA(12), plusA(11) => prevA(11), 
                           plusA(10) => prevA(10), plusA(9) => prevA(9), 
                           plusA(8) => prevA(8), plusA(7) => prevA(7), plusA(6)
                           => prevA(6), plusA(5) => prevA(5), plusA(4) => 
                           prevA(4), plusA(3) => prevA(3), plusA(2) => prevA(2)
                           , plusA(1) => prevA(1), plusA(0) => prevA(0), 
                           plus2A_out(63) => plus2A_s_63_port, plus2A_out(62) 
                           => plus2A_s_62_port, plus2A_out(61) => 
                           plus2A_s_61_port, plus2A_out(60) => plus2A_s_60_port
                           , plus2A_out(59) => plus2A_s_59_port, plus2A_out(58)
                           => plus2A_s_58_port, plus2A_out(57) => 
                           plus2A_s_57_port, plus2A_out(56) => plus2A_s_56_port
                           , plus2A_out(55) => plus2A_s_55_port, plus2A_out(54)
                           => plus2A_s_54_port, plus2A_out(53) => 
                           plus2A_s_53_port, plus2A_out(52) => plus2A_s_52_port
                           , plus2A_out(51) => plus2A_s_51_port, plus2A_out(50)
                           => plus2A_s_50_port, plus2A_out(49) => 
                           plus2A_s_49_port, plus2A_out(48) => plus2A_s_48_port
                           , plus2A_out(47) => plus2A_s_47_port, plus2A_out(46)
                           => plus2A_s_46_port, plus2A_out(45) => 
                           plus2A_s_45_port, plus2A_out(44) => plus2A_s_44_port
                           , plus2A_out(43) => plus2A_s_43_port, plus2A_out(42)
                           => plus2A_s_42_port, plus2A_out(41) => 
                           plus2A_s_41_port, plus2A_out(40) => plus2A_s_40_port
                           , plus2A_out(39) => plus2A_s_39_port, plus2A_out(38)
                           => plus2A_s_38_port, plus2A_out(37) => 
                           plus2A_s_37_port, plus2A_out(36) => plus2A_s_36_port
                           , plus2A_out(35) => plus2A_s_35_port, plus2A_out(34)
                           => plus2A_s_34_port, plus2A_out(33) => 
                           plus2A_s_33_port, plus2A_out(32) => plus2A_s_32_port
                           , plus2A_out(31) => plus2A_s_31_port, plus2A_out(30)
                           => plus2A_s_30_port, plus2A_out(29) => 
                           plus2A_s_29_port, plus2A_out(28) => plus2A_s_28_port
                           , plus2A_out(27) => plus2A_s_27_port, plus2A_out(26)
                           => plus2A_s_26_port, plus2A_out(25) => 
                           plus2A_s_25_port, plus2A_out(24) => plus2A_s_24_port
                           , plus2A_out(23) => plus2A_s_23_port, plus2A_out(22)
                           => plus2A_s_22_port, plus2A_out(21) => 
                           plus2A_s_21_port, plus2A_out(20) => plus2A_s_20_port
                           , plus2A_out(19) => plus2A_s_19_port, plus2A_out(18)
                           => plus2A_s_18_port, plus2A_out(17) => 
                           plus2A_s_17_port, plus2A_out(16) => plus2A_s_16_port
                           , plus2A_out(15) => plus2A_s_15_port, plus2A_out(14)
                           => plus2A_s_14_port, plus2A_out(13) => 
                           plus2A_s_13_port, plus2A_out(12) => plus2A_s_12_port
                           , plus2A_out(11) => plus2A_s_11_port, plus2A_out(10)
                           => plus2A_s_10_port, plus2A_out(9) => 
                           plus2A_s_9_port, plus2A_out(8) => plus2A_s_8_port, 
                           plus2A_out(7) => plus2A_s_7_port, plus2A_out(6) => 
                           plus2A_s_6_port, plus2A_out(5) => plus2A_s_5_port, 
                           plus2A_out(4) => plus2A_s_4_port, plus2A_out(3) => 
                           plus2A_s_3_port, plus2A_out(2) => plus2A_s_2_port, 
                           plus2A_out(1) => plus2A_s_1_port, plus2A_out(0) => 
                           n_3190, minus2A_out(63) => minus2A_s_63_port, 
                           minus2A_out(62) => minus2A_s_62_port, 
                           minus2A_out(61) => minus2A_s_61_port, 
                           minus2A_out(60) => minus2A_s_60_port, 
                           minus2A_out(59) => minus2A_s_59_port, 
                           minus2A_out(58) => minus2A_s_58_port, 
                           minus2A_out(57) => minus2A_s_57_port, 
                           minus2A_out(56) => minus2A_s_56_port, 
                           minus2A_out(55) => minus2A_s_55_port, 
                           minus2A_out(54) => minus2A_s_54_port, 
                           minus2A_out(53) => minus2A_s_53_port, 
                           minus2A_out(52) => minus2A_s_52_port, 
                           minus2A_out(51) => minus2A_s_51_port, 
                           minus2A_out(50) => minus2A_s_50_port, 
                           minus2A_out(49) => minus2A_s_49_port, 
                           minus2A_out(48) => minus2A_s_48_port, 
                           minus2A_out(47) => minus2A_s_47_port, 
                           minus2A_out(46) => minus2A_s_46_port, 
                           minus2A_out(45) => minus2A_s_45_port, 
                           minus2A_out(44) => minus2A_s_44_port, 
                           minus2A_out(43) => minus2A_s_43_port, 
                           minus2A_out(42) => minus2A_s_42_port, 
                           minus2A_out(41) => minus2A_s_41_port, 
                           minus2A_out(40) => minus2A_s_40_port, 
                           minus2A_out(39) => minus2A_s_39_port, 
                           minus2A_out(38) => minus2A_s_38_port, 
                           minus2A_out(37) => minus2A_s_37_port, 
                           minus2A_out(36) => minus2A_s_36_port, 
                           minus2A_out(35) => minus2A_s_35_port, 
                           minus2A_out(34) => minus2A_s_34_port, 
                           minus2A_out(33) => minus2A_s_33_port, 
                           minus2A_out(32) => minus2A_s_32_port, 
                           minus2A_out(31) => minus2A_s_31_port, 
                           minus2A_out(30) => minus2A_s_30_port, 
                           minus2A_out(29) => minus2A_s_29_port, 
                           minus2A_out(28) => minus2A_s_28_port, 
                           minus2A_out(27) => minus2A_s_27_port, 
                           minus2A_out(26) => minus2A_s_26_port, 
                           minus2A_out(25) => minus2A_s_25_port, 
                           minus2A_out(24) => minus2A_s_24_port, 
                           minus2A_out(23) => minus2A_s_23_port, 
                           minus2A_out(22) => minus2A_s_22_port, 
                           minus2A_out(21) => minus2A_s_21_port, 
                           minus2A_out(20) => minus2A_s_20_port, 
                           minus2A_out(19) => minus2A_s_19_port, 
                           minus2A_out(18) => minus2A_s_18_port, 
                           minus2A_out(17) => minus2A_s_17_port, 
                           minus2A_out(16) => minus2A_s_16_port, 
                           minus2A_out(15) => minus2A_s_15_port, 
                           minus2A_out(14) => minus2A_s_14_port, 
                           minus2A_out(13) => minus2A_s_13_port, 
                           minus2A_out(12) => minus2A_s_12_port, 
                           minus2A_out(11) => minus2A_s_11_port, 
                           minus2A_out(10) => minus2A_s_10_port, minus2A_out(9)
                           => minus2A_s_9_port, minus2A_out(8) => 
                           minus2A_s_8_port, minus2A_out(7) => minus2A_s_7_port
                           , minus2A_out(6) => minus2A_s_6_port, minus2A_out(5)
                           => minus2A_s_5_port, minus2A_out(4) => 
                           minus2A_s_4_port, minus2A_out(3) => minus2A_s_3_port
                           , minus2A_out(2) => minus2A_s_2_port, minus2A_out(1)
                           => minus2A_s_1_port, minus2A_out(0) => 
                           minus2A_s_0_port, plus4A_out(63) => nextA_63_port, 
                           plus4A_out(62) => nextA_62_port, plus4A_out(61) => 
                           nextA_61_port, plus4A_out(60) => nextA_60_port, 
                           plus4A_out(59) => nextA_59_port, plus4A_out(58) => 
                           nextA_58_port, plus4A_out(57) => n3, plus4A_out(56) 
                           => nextA_56_port, plus4A_out(55) => nextA_55_port, 
                           plus4A_out(54) => nextA_54_port, plus4A_out(53) => 
                           nextA_53_port, plus4A_out(52) => nextA_52_port, 
                           plus4A_out(51) => nextA_51_port, plus4A_out(50) => 
                           nextA_50_port, plus4A_out(49) => nextA_49_port, 
                           plus4A_out(48) => nextA_48_port, plus4A_out(47) => 
                           nextA_47_port, plus4A_out(46) => nextA_46_port, 
                           plus4A_out(45) => nextA_45_port, plus4A_out(44) => 
                           nextA_44_port, plus4A_out(43) => nextA_43_port, 
                           plus4A_out(42) => nextA_42_port, plus4A_out(41) => 
                           nextA_41_port, plus4A_out(40) => nextA_40_port, 
                           plus4A_out(39) => nextA_39_port, plus4A_out(38) => 
                           nextA_38_port, plus4A_out(37) => nextA_37_port, 
                           plus4A_out(36) => nextA_36_port, plus4A_out(35) => 
                           nextA_35_port, plus4A_out(34) => nextA_34_port, 
                           plus4A_out(33) => nextA_33_port, plus4A_out(32) => 
                           nextA_32_port, plus4A_out(31) => nextA_31_port, 
                           plus4A_out(30) => nextA_30_port, plus4A_out(29) => 
                           nextA_29_port, plus4A_out(28) => nextA_28_port, 
                           plus4A_out(27) => nextA_27_port, plus4A_out(26) => 
                           nextA_26_port, plus4A_out(25) => nextA_25_port, 
                           plus4A_out(24) => nextA_24_port, plus4A_out(23) => 
                           nextA_23_port, plus4A_out(22) => nextA_22_port, 
                           plus4A_out(21) => nextA_21_port, plus4A_out(20) => 
                           nextA_20_port, plus4A_out(19) => nextA_19_port, 
                           plus4A_out(18) => nextA_18_port, plus4A_out(17) => 
                           nextA_17_port, plus4A_out(16) => nextA_16_port, 
                           plus4A_out(15) => nextA_15_port, plus4A_out(14) => 
                           nextA_14_port, plus4A_out(13) => nextA_13_port, 
                           plus4A_out(12) => nextA_12_port, plus4A_out(11) => 
                           nextA_11_port, plus4A_out(10) => nextA_10_port, 
                           plus4A_out(9) => nextA_9_port, plus4A_out(8) => 
                           nextA_8_port, plus4A_out(7) => nextA_7_port, 
                           plus4A_out(6) => nextA_6_port, plus4A_out(5) => 
                           nextA_5_port, plus4A_out(4) => nextA_4_port, 
                           plus4A_out(3) => nextA_3_port, plus4A_out(2) => 
                           nextA_2_port, plus4A_out(1) => nextA_1_port, 
                           plus4A_out(0) => n_3191, minus4A_out(63) => 
                           minus4A_s_63_port, minus4A_out(62) => 
                           minus4A_s_62_port, minus4A_out(61) => 
                           minus4A_s_61_port, minus4A_out(60) => 
                           minus4A_s_60_port, minus4A_out(59) => 
                           minus4A_s_59_port, minus4A_out(58) => 
                           minus4A_s_58_port, minus4A_out(57) => 
                           minus4A_s_57_port, minus4A_out(56) => 
                           minus4A_s_56_port, minus4A_out(55) => 
                           minus4A_s_55_port, minus4A_out(54) => 
                           minus4A_s_54_port, minus4A_out(53) => 
                           minus4A_s_53_port, minus4A_out(52) => 
                           minus4A_s_52_port, minus4A_out(51) => 
                           minus4A_s_51_port, minus4A_out(50) => 
                           minus4A_s_50_port, minus4A_out(49) => 
                           minus4A_s_49_port, minus4A_out(48) => 
                           minus4A_s_48_port, minus4A_out(47) => 
                           minus4A_s_47_port, minus4A_out(46) => 
                           minus4A_s_46_port, minus4A_out(45) => 
                           minus4A_s_45_port, minus4A_out(44) => 
                           minus4A_s_44_port, minus4A_out(43) => 
                           minus4A_s_43_port, minus4A_out(42) => 
                           minus4A_s_42_port, minus4A_out(41) => 
                           minus4A_s_41_port, minus4A_out(40) => 
                           minus4A_s_40_port, minus4A_out(39) => 
                           minus4A_s_39_port, minus4A_out(38) => 
                           minus4A_s_38_port, minus4A_out(37) => 
                           minus4A_s_37_port, minus4A_out(36) => 
                           minus4A_s_36_port, minus4A_out(35) => 
                           minus4A_s_35_port, minus4A_out(34) => 
                           minus4A_s_34_port, minus4A_out(33) => 
                           minus4A_s_33_port, minus4A_out(32) => 
                           minus4A_s_32_port, minus4A_out(31) => 
                           minus4A_s_31_port, minus4A_out(30) => 
                           minus4A_s_30_port, minus4A_out(29) => 
                           minus4A_s_29_port, minus4A_out(28) => 
                           minus4A_s_28_port, minus4A_out(27) => 
                           minus4A_s_27_port, minus4A_out(26) => 
                           minus4A_s_26_port, minus4A_out(25) => 
                           minus4A_s_25_port, minus4A_out(24) => 
                           minus4A_s_24_port, minus4A_out(23) => 
                           minus4A_s_23_port, minus4A_out(22) => 
                           minus4A_s_22_port, minus4A_out(21) => 
                           minus4A_s_21_port, minus4A_out(20) => 
                           minus4A_s_20_port, minus4A_out(19) => 
                           minus4A_s_19_port, minus4A_out(18) => 
                           minus4A_s_18_port, minus4A_out(17) => 
                           minus4A_s_17_port, minus4A_out(16) => 
                           minus4A_s_16_port, minus4A_out(15) => 
                           minus4A_s_15_port, minus4A_out(14) => 
                           minus4A_s_14_port, minus4A_out(13) => 
                           minus4A_s_13_port, minus4A_out(12) => 
                           minus4A_s_12_port, minus4A_out(11) => 
                           minus4A_s_11_port, minus4A_out(10) => 
                           minus4A_s_10_port, minus4A_out(9) => 
                           minus4A_s_9_port, minus4A_out(8) => minus4A_s_8_port
                           , minus4A_out(7) => minus4A_s_7_port, minus4A_out(6)
                           => minus4A_s_6_port, minus4A_out(5) => 
                           minus4A_s_5_port, minus4A_out(4) => minus4A_s_4_port
                           , minus4A_out(3) => minus4A_s_3_port, minus4A_out(2)
                           => minus4A_s_2_port, minus4A_out(1) => 
                           minus4A_s_1_port, minus4A_out(0) => minus4A_s_0_port
                           );
   mux_1 : MUX_GENERIC_N64_RADIX3_6 port map( plusA(63) => plus2A_s_63_port, 
                           plusA(62) => plus2A_s_62_port, plusA(61) => 
                           plus2A_s_61_port, plusA(60) => plus2A_s_60_port, 
                           plusA(59) => plus2A_s_59_port, plusA(58) => 
                           plus2A_s_58_port, plusA(57) => plus2A_s_57_port, 
                           plusA(56) => plus2A_s_56_port, plusA(55) => 
                           plus2A_s_55_port, plusA(54) => plus2A_s_54_port, 
                           plusA(53) => plus2A_s_53_port, plusA(52) => 
                           plus2A_s_52_port, plusA(51) => plus2A_s_51_port, 
                           plusA(50) => plus2A_s_50_port, plusA(49) => 
                           plus2A_s_49_port, plusA(48) => plus2A_s_48_port, 
                           plusA(47) => plus2A_s_47_port, plusA(46) => 
                           plus2A_s_46_port, plusA(45) => plus2A_s_45_port, 
                           plusA(44) => plus2A_s_44_port, plusA(43) => 
                           plus2A_s_43_port, plusA(42) => plus2A_s_42_port, 
                           plusA(41) => plus2A_s_41_port, plusA(40) => 
                           plus2A_s_40_port, plusA(39) => plus2A_s_39_port, 
                           plusA(38) => plus2A_s_38_port, plusA(37) => 
                           plus2A_s_37_port, plusA(36) => plus2A_s_36_port, 
                           plusA(35) => plus2A_s_35_port, plusA(34) => 
                           plus2A_s_34_port, plusA(33) => plus2A_s_33_port, 
                           plusA(32) => plus2A_s_32_port, plusA(31) => 
                           plus2A_s_31_port, plusA(30) => plus2A_s_30_port, 
                           plusA(29) => plus2A_s_29_port, plusA(28) => 
                           plus2A_s_28_port, plusA(27) => plus2A_s_27_port, 
                           plusA(26) => plus2A_s_26_port, plusA(25) => 
                           plus2A_s_25_port, plusA(24) => plus2A_s_24_port, 
                           plusA(23) => plus2A_s_23_port, plusA(22) => 
                           plus2A_s_22_port, plusA(21) => plus2A_s_21_port, 
                           plusA(20) => plus2A_s_20_port, plusA(19) => 
                           plus2A_s_19_port, plusA(18) => plus2A_s_18_port, 
                           plusA(17) => plus2A_s_17_port, plusA(16) => 
                           plus2A_s_16_port, plusA(15) => plus2A_s_15_port, 
                           plusA(14) => plus2A_s_14_port, plusA(13) => 
                           plus2A_s_13_port, plusA(12) => plus2A_s_12_port, 
                           plusA(11) => plus2A_s_11_port, plusA(10) => 
                           plus2A_s_10_port, plusA(9) => plus2A_s_9_port, 
                           plusA(8) => plus2A_s_8_port, plusA(7) => 
                           plus2A_s_7_port, plusA(6) => plus2A_s_6_port, 
                           plusA(5) => plus2A_s_5_port, plusA(4) => 
                           plus2A_s_4_port, plusA(3) => plus2A_s_3_port, 
                           plusA(2) => plus2A_s_2_port, plusA(1) => 
                           plus2A_s_1_port, plusA(0) => nextA_0_port, 
                           minusA(63) => minus2A_s_63_port, minusA(62) => 
                           minus2A_s_62_port, minusA(61) => minus2A_s_61_port, 
                           minusA(60) => minus2A_s_60_port, minusA(59) => 
                           minus2A_s_59_port, minusA(58) => minus2A_s_58_port, 
                           minusA(57) => minus2A_s_57_port, minusA(56) => 
                           minus2A_s_56_port, minusA(55) => minus2A_s_55_port, 
                           minusA(54) => minus2A_s_54_port, minusA(53) => 
                           minus2A_s_53_port, minusA(52) => minus2A_s_52_port, 
                           minusA(51) => minus2A_s_51_port, minusA(50) => 
                           minus2A_s_50_port, minusA(49) => minus2A_s_49_port, 
                           minusA(48) => minus2A_s_48_port, minusA(47) => 
                           minus2A_s_47_port, minusA(46) => minus2A_s_46_port, 
                           minusA(45) => minus2A_s_45_port, minusA(44) => 
                           minus2A_s_44_port, minusA(43) => minus2A_s_43_port, 
                           minusA(42) => minus2A_s_42_port, minusA(41) => 
                           minus2A_s_41_port, minusA(40) => minus2A_s_40_port, 
                           minusA(39) => minus2A_s_39_port, minusA(38) => 
                           minus2A_s_38_port, minusA(37) => minus2A_s_37_port, 
                           minusA(36) => minus2A_s_36_port, minusA(35) => 
                           minus2A_s_35_port, minusA(34) => minus2A_s_34_port, 
                           minusA(33) => minus2A_s_33_port, minusA(32) => 
                           minus2A_s_32_port, minusA(31) => minus2A_s_31_port, 
                           minusA(30) => minus2A_s_30_port, minusA(29) => 
                           minus2A_s_29_port, minusA(28) => minus2A_s_28_port, 
                           minusA(27) => minus2A_s_27_port, minusA(26) => 
                           minus2A_s_26_port, minusA(25) => minus2A_s_25_port, 
                           minusA(24) => minus2A_s_24_port, minusA(23) => 
                           minus2A_s_23_port, minusA(22) => minus2A_s_22_port, 
                           minusA(21) => minus2A_s_21_port, minusA(20) => 
                           minus2A_s_20_port, minusA(19) => minus2A_s_19_port, 
                           minusA(18) => minus2A_s_18_port, minusA(17) => 
                           minus2A_s_17_port, minusA(16) => minus2A_s_16_port, 
                           minusA(15) => minus2A_s_15_port, minusA(14) => 
                           minus2A_s_14_port, minusA(13) => minus2A_s_13_port, 
                           minusA(12) => minus2A_s_12_port, minusA(11) => 
                           minus2A_s_11_port, minusA(10) => minus2A_s_10_port, 
                           minusA(9) => minus2A_s_9_port, minusA(8) => 
                           minus2A_s_8_port, minusA(7) => minus2A_s_7_port, 
                           minusA(6) => minus2A_s_6_port, minusA(5) => 
                           minus2A_s_5_port, minusA(4) => minus2A_s_4_port, 
                           minusA(3) => minus2A_s_3_port, minusA(2) => 
                           minus2A_s_2_port, minusA(1) => minus2A_s_1_port, 
                           minusA(0) => minus2A_s_0_port, plus2A(63) => 
                           nextA_63_port, plus2A(62) => nextA_62_port, 
                           plus2A(61) => nextA_61_port, plus2A(60) => 
                           nextA_60_port, plus2A(59) => nextA_59_port, 
                           plus2A(58) => nextA_58_port, plus2A(57) => 
                           nextA_57_port, plus2A(56) => nextA_56_port, 
                           plus2A(55) => nextA_55_port, plus2A(54) => 
                           nextA_54_port, plus2A(53) => nextA_53_port, 
                           plus2A(52) => nextA_52_port, plus2A(51) => 
                           nextA_51_port, plus2A(50) => nextA_50_port, 
                           plus2A(49) => nextA_49_port, plus2A(48) => 
                           nextA_48_port, plus2A(47) => nextA_47_port, 
                           plus2A(46) => nextA_46_port, plus2A(45) => 
                           nextA_45_port, plus2A(44) => nextA_44_port, 
                           plus2A(43) => nextA_43_port, plus2A(42) => 
                           nextA_42_port, plus2A(41) => nextA_41_port, 
                           plus2A(40) => nextA_40_port, plus2A(39) => 
                           nextA_39_port, plus2A(38) => nextA_38_port, 
                           plus2A(37) => nextA_37_port, plus2A(36) => 
                           nextA_36_port, plus2A(35) => nextA_35_port, 
                           plus2A(34) => nextA_34_port, plus2A(33) => 
                           nextA_33_port, plus2A(32) => nextA_32_port, 
                           plus2A(31) => nextA_31_port, plus2A(30) => 
                           nextA_30_port, plus2A(29) => nextA_29_port, 
                           plus2A(28) => nextA_28_port, plus2A(27) => 
                           nextA_27_port, plus2A(26) => nextA_26_port, 
                           plus2A(25) => nextA_25_port, plus2A(24) => 
                           nextA_24_port, plus2A(23) => nextA_23_port, 
                           plus2A(22) => nextA_22_port, plus2A(21) => 
                           nextA_21_port, plus2A(20) => nextA_20_port, 
                           plus2A(19) => nextA_19_port, plus2A(18) => 
                           nextA_18_port, plus2A(17) => nextA_17_port, 
                           plus2A(16) => nextA_16_port, plus2A(15) => 
                           nextA_15_port, plus2A(14) => nextA_14_port, 
                           plus2A(13) => nextA_13_port, plus2A(12) => 
                           nextA_12_port, plus2A(11) => nextA_11_port, 
                           plus2A(10) => nextA_10_port, plus2A(9) => 
                           nextA_9_port, plus2A(8) => nextA_8_port, plus2A(7) 
                           => nextA_7_port, plus2A(6) => nextA_6_port, 
                           plus2A(5) => nextA_5_port, plus2A(4) => nextA_4_port
                           , plus2A(3) => nextA_3_port, plus2A(2) => 
                           nextA_2_port, plus2A(1) => nextA_1_port, plus2A(0) 
                           => nextA_0_port, minus2A(63) => minus4A_s_63_port, 
                           minus2A(62) => minus4A_s_62_port, minus2A(61) => 
                           minus4A_s_61_port, minus2A(60) => minus4A_s_60_port,
                           minus2A(59) => minus4A_s_59_port, minus2A(58) => 
                           minus4A_s_58_port, minus2A(57) => minus4A_s_57_port,
                           minus2A(56) => minus4A_s_56_port, minus2A(55) => 
                           minus4A_s_55_port, minus2A(54) => minus4A_s_54_port,
                           minus2A(53) => minus4A_s_53_port, minus2A(52) => 
                           minus4A_s_52_port, minus2A(51) => minus4A_s_51_port,
                           minus2A(50) => minus4A_s_50_port, minus2A(49) => 
                           minus4A_s_49_port, minus2A(48) => minus4A_s_48_port,
                           minus2A(47) => minus4A_s_47_port, minus2A(46) => 
                           minus4A_s_46_port, minus2A(45) => minus4A_s_45_port,
                           minus2A(44) => minus4A_s_44_port, minus2A(43) => 
                           minus4A_s_43_port, minus2A(42) => minus4A_s_42_port,
                           minus2A(41) => minus4A_s_41_port, minus2A(40) => 
                           minus4A_s_40_port, minus2A(39) => minus4A_s_39_port,
                           minus2A(38) => minus4A_s_38_port, minus2A(37) => 
                           minus4A_s_37_port, minus2A(36) => minus4A_s_36_port,
                           minus2A(35) => minus4A_s_35_port, minus2A(34) => 
                           minus4A_s_34_port, minus2A(33) => minus4A_s_33_port,
                           minus2A(32) => minus4A_s_32_port, minus2A(31) => 
                           minus4A_s_31_port, minus2A(30) => minus4A_s_30_port,
                           minus2A(29) => minus4A_s_29_port, minus2A(28) => 
                           minus4A_s_28_port, minus2A(27) => minus4A_s_27_port,
                           minus2A(26) => minus4A_s_26_port, minus2A(25) => 
                           minus4A_s_25_port, minus2A(24) => minus4A_s_24_port,
                           minus2A(23) => minus4A_s_23_port, minus2A(22) => 
                           minus4A_s_22_port, minus2A(21) => minus4A_s_21_port,
                           minus2A(20) => minus4A_s_20_port, minus2A(19) => 
                           minus4A_s_19_port, minus2A(18) => minus4A_s_18_port,
                           minus2A(17) => minus4A_s_17_port, minus2A(16) => 
                           minus4A_s_16_port, minus2A(15) => minus4A_s_15_port,
                           minus2A(14) => minus4A_s_14_port, minus2A(13) => 
                           minus4A_s_13_port, minus2A(12) => minus4A_s_12_port,
                           minus2A(11) => minus4A_s_11_port, minus2A(10) => 
                           minus4A_s_10_port, minus2A(9) => minus4A_s_9_port, 
                           minus2A(8) => minus4A_s_8_port, minus2A(7) => 
                           minus4A_s_7_port, minus2A(6) => minus4A_s_6_port, 
                           minus2A(5) => minus4A_s_5_port, minus2A(4) => 
                           minus4A_s_4_port, minus2A(3) => minus4A_s_3_port, 
                           minus2A(2) => minus4A_s_2_port, minus2A(1) => 
                           minus4A_s_1_port, minus2A(0) => minus4A_s_0_port, 
                           SEL(2) => encoder_to_mux_2_port, SEL(1) => 
                           encoder_to_mux_1_port, SEL(0) => 
                           encoder_to_mux_0_port, Y(63) => mux_to_adder_63_port
                           , Y(62) => mux_to_adder_62_port, Y(61) => 
                           mux_to_adder_61_port, Y(60) => mux_to_adder_60_port,
                           Y(59) => mux_to_adder_59_port, Y(58) => 
                           mux_to_adder_58_port, Y(57) => mux_to_adder_57_port,
                           Y(56) => mux_to_adder_56_port, Y(55) => 
                           mux_to_adder_55_port, Y(54) => mux_to_adder_54_port,
                           Y(53) => mux_to_adder_53_port, Y(52) => 
                           mux_to_adder_52_port, Y(51) => mux_to_adder_51_port,
                           Y(50) => mux_to_adder_50_port, Y(49) => 
                           mux_to_adder_49_port, Y(48) => mux_to_adder_48_port,
                           Y(47) => mux_to_adder_47_port, Y(46) => 
                           mux_to_adder_46_port, Y(45) => mux_to_adder_45_port,
                           Y(44) => mux_to_adder_44_port, Y(43) => 
                           mux_to_adder_43_port, Y(42) => mux_to_adder_42_port,
                           Y(41) => mux_to_adder_41_port, Y(40) => 
                           mux_to_adder_40_port, Y(39) => mux_to_adder_39_port,
                           Y(38) => mux_to_adder_38_port, Y(37) => 
                           mux_to_adder_37_port, Y(36) => mux_to_adder_36_port,
                           Y(35) => mux_to_adder_35_port, Y(34) => 
                           mux_to_adder_34_port, Y(33) => mux_to_adder_33_port,
                           Y(32) => mux_to_adder_32_port, Y(31) => 
                           mux_to_adder_31_port, Y(30) => mux_to_adder_30_port,
                           Y(29) => mux_to_adder_29_port, Y(28) => 
                           mux_to_adder_28_port, Y(27) => mux_to_adder_27_port,
                           Y(26) => mux_to_adder_26_port, Y(25) => 
                           mux_to_adder_25_port, Y(24) => mux_to_adder_24_port,
                           Y(23) => mux_to_adder_23_port, Y(22) => 
                           mux_to_adder_22_port, Y(21) => mux_to_adder_21_port,
                           Y(20) => mux_to_adder_20_port, Y(19) => 
                           mux_to_adder_19_port, Y(18) => mux_to_adder_18_port,
                           Y(17) => mux_to_adder_17_port, Y(16) => 
                           mux_to_adder_16_port, Y(15) => mux_to_adder_15_port,
                           Y(14) => mux_to_adder_14_port, Y(13) => 
                           mux_to_adder_13_port, Y(12) => mux_to_adder_12_port,
                           Y(11) => mux_to_adder_11_port, Y(10) => 
                           mux_to_adder_10_port, Y(9) => mux_to_adder_9_port, 
                           Y(8) => mux_to_adder_8_port, Y(7) => 
                           mux_to_adder_7_port, Y(6) => mux_to_adder_6_port, 
                           Y(5) => mux_to_adder_5_port, Y(4) => 
                           mux_to_adder_4_port, Y(3) => mux_to_adder_3_port, 
                           Y(2) => mux_to_adder_2_port, Y(1) => 
                           mux_to_adder_1_port, Y(0) => mux_to_adder_0_port);
   rca_1 : RCA_N64_6 port map( A(63) => mux_to_adder_63_port, A(62) => 
                           mux_to_adder_62_port, A(61) => mux_to_adder_61_port,
                           A(60) => mux_to_adder_60_port, A(59) => 
                           mux_to_adder_59_port, A(58) => mux_to_adder_58_port,
                           A(57) => mux_to_adder_57_port, A(56) => 
                           mux_to_adder_56_port, A(55) => mux_to_adder_55_port,
                           A(54) => mux_to_adder_54_port, A(53) => 
                           mux_to_adder_53_port, A(52) => mux_to_adder_52_port,
                           A(51) => mux_to_adder_51_port, A(50) => 
                           mux_to_adder_50_port, A(49) => mux_to_adder_49_port,
                           A(48) => mux_to_adder_48_port, A(47) => 
                           mux_to_adder_47_port, A(46) => mux_to_adder_46_port,
                           A(45) => mux_to_adder_45_port, A(44) => 
                           mux_to_adder_44_port, A(43) => mux_to_adder_43_port,
                           A(42) => mux_to_adder_42_port, A(41) => 
                           mux_to_adder_41_port, A(40) => mux_to_adder_40_port,
                           A(39) => mux_to_adder_39_port, A(38) => 
                           mux_to_adder_38_port, A(37) => mux_to_adder_37_port,
                           A(36) => mux_to_adder_36_port, A(35) => 
                           mux_to_adder_35_port, A(34) => mux_to_adder_34_port,
                           A(33) => mux_to_adder_33_port, A(32) => 
                           mux_to_adder_32_port, A(31) => mux_to_adder_31_port,
                           A(30) => mux_to_adder_30_port, A(29) => 
                           mux_to_adder_29_port, A(28) => mux_to_adder_28_port,
                           A(27) => mux_to_adder_27_port, A(26) => 
                           mux_to_adder_26_port, A(25) => mux_to_adder_25_port,
                           A(24) => mux_to_adder_24_port, A(23) => 
                           mux_to_adder_23_port, A(22) => mux_to_adder_22_port,
                           A(21) => mux_to_adder_21_port, A(20) => 
                           mux_to_adder_20_port, A(19) => mux_to_adder_19_port,
                           A(18) => mux_to_adder_18_port, A(17) => 
                           mux_to_adder_17_port, A(16) => mux_to_adder_16_port,
                           A(15) => mux_to_adder_15_port, A(14) => 
                           mux_to_adder_14_port, A(13) => mux_to_adder_13_port,
                           A(12) => mux_to_adder_12_port, A(11) => 
                           mux_to_adder_11_port, A(10) => mux_to_adder_10_port,
                           A(9) => mux_to_adder_9_port, A(8) => 
                           mux_to_adder_8_port, A(7) => mux_to_adder_7_port, 
                           A(6) => mux_to_adder_6_port, A(5) => 
                           mux_to_adder_5_port, A(4) => mux_to_adder_4_port, 
                           A(3) => mux_to_adder_3_port, A(2) => 
                           mux_to_adder_2_port, A(1) => mux_to_adder_1_port, 
                           A(0) => mux_to_adder_0_port, B(63) => prevSum(63), 
                           B(62) => prevSum(62), B(61) => prevSum(61), B(60) =>
                           prevSum(60), B(59) => prevSum(59), B(58) => 
                           prevSum(58), B(57) => prevSum(57), B(56) => 
                           prevSum(56), B(55) => prevSum(55), B(54) => 
                           prevSum(54), B(53) => prevSum(53), B(52) => 
                           prevSum(52), B(51) => prevSum(51), B(50) => 
                           prevSum(50), B(49) => prevSum(49), B(48) => 
                           prevSum(48), B(47) => prevSum(47), B(46) => 
                           prevSum(46), B(45) => prevSum(45), B(44) => 
                           prevSum(44), B(43) => prevSum(43), B(42) => 
                           prevSum(42), B(41) => prevSum(41), B(40) => 
                           prevSum(40), B(39) => prevSum(39), B(38) => 
                           prevSum(38), B(37) => prevSum(37), B(36) => 
                           prevSum(36), B(35) => prevSum(35), B(34) => 
                           prevSum(34), B(33) => prevSum(33), B(32) => 
                           prevSum(32), B(31) => prevSum(31), B(30) => 
                           prevSum(30), B(29) => prevSum(29), B(28) => 
                           prevSum(28), B(27) => prevSum(27), B(26) => 
                           prevSum(26), B(25) => prevSum(25), B(24) => 
                           prevSum(24), B(23) => prevSum(23), B(22) => 
                           prevSum(22), B(21) => prevSum(21), B(20) => 
                           prevSum(20), B(19) => prevSum(19), B(18) => 
                           prevSum(18), B(17) => prevSum(17), B(16) => 
                           prevSum(16), B(15) => prevSum(15), B(14) => 
                           prevSum(14), B(13) => prevSum(13), B(12) => 
                           prevSum(12), B(11) => prevSum(11), B(10) => 
                           prevSum(10), B(9) => prevSum(9), B(8) => prevSum(8),
                           B(7) => prevSum(7), B(6) => prevSum(6), B(5) => 
                           prevSum(5), B(4) => prevSum(4), B(3) => prevSum(3), 
                           B(2) => prevSum(2), B(1) => prevSum(1), B(0) => 
                           prevSum(0), Ci => X_Logic0_port, S(63) => 
                           nextSum(63), S(62) => nextSum(62), S(61) => 
                           nextSum(61), S(60) => nextSum(60), S(59) => 
                           nextSum(59), S(58) => nextSum(58), S(57) => 
                           nextSum(57), S(56) => nextSum(56), S(55) => 
                           nextSum(55), S(54) => nextSum(54), S(53) => 
                           nextSum(53), S(52) => nextSum(52), S(51) => 
                           nextSum(51), S(50) => nextSum(50), S(49) => 
                           nextSum(49), S(48) => nextSum(48), S(47) => 
                           nextSum(47), S(46) => nextSum(46), S(45) => 
                           nextSum(45), S(44) => nextSum(44), S(43) => 
                           nextSum(43), S(42) => nextSum(42), S(41) => 
                           nextSum(41), S(40) => nextSum(40), S(39) => 
                           nextSum(39), S(38) => nextSum(38), S(37) => 
                           nextSum(37), S(36) => nextSum(36), S(35) => 
                           nextSum(35), S(34) => nextSum(34), S(33) => 
                           nextSum(33), S(32) => nextSum(32), S(31) => 
                           nextSum(31), S(30) => nextSum(30), S(29) => 
                           nextSum(29), S(28) => nextSum(28), S(27) => 
                           nextSum(27), S(26) => nextSum(26), S(25) => 
                           nextSum(25), S(24) => nextSum(24), S(23) => 
                           nextSum(23), S(22) => nextSum(22), S(21) => 
                           nextSum(21), S(20) => nextSum(20), S(19) => 
                           nextSum(19), S(18) => nextSum(18), S(17) => 
                           nextSum(17), S(16) => nextSum(16), S(15) => 
                           nextSum(15), S(14) => nextSum(14), S(13) => 
                           nextSum(13), S(12) => nextSum(12), S(11) => 
                           nextSum(11), S(10) => nextSum(10), S(9) => 
                           nextSum(9), S(8) => nextSum(8), S(7) => nextSum(7), 
                           S(6) => nextSum(6), S(5) => nextSum(5), S(4) => 
                           nextSum(4), S(3) => nextSum(3), S(2) => nextSum(2), 
                           S(1) => nextSum(1), S(0) => nextSum(0), Co => n_3192
                           );
   U3 : BUF_X1 port map( A => n3, Z => nextA_57_port);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity booth_mul_row_N64_RADIX3_7 is

   port( prevA, prevSum : in std_logic_vector (63 downto 0);  encoderIn : in 
         std_logic_vector (2 downto 0);  nextA, nextSum : out std_logic_vector 
         (63 downto 0));

end booth_mul_row_N64_RADIX3_7;

architecture SYN_struct of booth_mul_row_N64_RADIX3_7 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component RCA_N64_7
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component MUX_GENERIC_N64_RADIX3_7
      port( plusA, minusA, plus2A, minus2A : in std_logic_vector (63 downto 0);
            SEL : in std_logic_vector (2 downto 0);  Y : out std_logic_vector 
            (63 downto 0));
   end component;
   
   component ShiftnCompl_N64_7
      port( plusA : in std_logic_vector (63 downto 0);  plus2A_out, minus2A_out
            , plus4A_out, minus4A_out : out std_logic_vector (63 downto 0));
   end component;
   
   component encoder_N64_RADIX3_7
      port( X : in std_logic_vector (2 downto 0);  Z : out std_logic_vector (2 
            downto 0));
   end component;
   
   signal X_Logic0_port, nextA_63_port, nextA_62_port, nextA_61_port, 
      nextA_60_port, nextA_59_port, nextA_58_port, n3, nextA_56_port, 
      nextA_55_port, nextA_54_port, nextA_53_port, nextA_52_port, nextA_51_port
      , nextA_50_port, nextA_49_port, nextA_48_port, nextA_47_port, 
      nextA_46_port, nextA_45_port, nextA_44_port, nextA_43_port, nextA_42_port
      , nextA_41_port, nextA_40_port, nextA_39_port, nextA_38_port, 
      nextA_37_port, nextA_36_port, nextA_35_port, nextA_34_port, nextA_33_port
      , nextA_32_port, nextA_31_port, nextA_30_port, nextA_29_port, 
      nextA_28_port, nextA_27_port, nextA_26_port, nextA_25_port, nextA_24_port
      , nextA_23_port, nextA_22_port, nextA_21_port, nextA_20_port, 
      nextA_19_port, nextA_18_port, nextA_17_port, nextA_16_port, nextA_15_port
      , nextA_14_port, nextA_13_port, nextA_12_port, nextA_11_port, 
      nextA_10_port, nextA_9_port, nextA_8_port, nextA_7_port, nextA_6_port, 
      nextA_5_port, nextA_4_port, nextA_3_port, nextA_2_port, nextA_1_port, 
      encoder_to_mux_2_port, encoder_to_mux_1_port, encoder_to_mux_0_port, 
      plus2A_s_63_port, plus2A_s_62_port, plus2A_s_61_port, plus2A_s_60_port, 
      plus2A_s_59_port, plus2A_s_58_port, plus2A_s_57_port, plus2A_s_56_port, 
      plus2A_s_55_port, plus2A_s_54_port, plus2A_s_53_port, plus2A_s_52_port, 
      plus2A_s_51_port, plus2A_s_50_port, plus2A_s_49_port, plus2A_s_48_port, 
      plus2A_s_47_port, plus2A_s_46_port, plus2A_s_45_port, plus2A_s_44_port, 
      plus2A_s_43_port, plus2A_s_42_port, plus2A_s_41_port, plus2A_s_40_port, 
      plus2A_s_39_port, plus2A_s_38_port, plus2A_s_37_port, plus2A_s_36_port, 
      plus2A_s_35_port, plus2A_s_34_port, plus2A_s_33_port, plus2A_s_32_port, 
      plus2A_s_31_port, plus2A_s_30_port, plus2A_s_29_port, plus2A_s_28_port, 
      plus2A_s_27_port, plus2A_s_26_port, plus2A_s_25_port, plus2A_s_24_port, 
      plus2A_s_23_port, plus2A_s_22_port, plus2A_s_21_port, plus2A_s_20_port, 
      plus2A_s_19_port, plus2A_s_18_port, plus2A_s_17_port, plus2A_s_16_port, 
      plus2A_s_15_port, plus2A_s_14_port, plus2A_s_13_port, plus2A_s_12_port, 
      plus2A_s_11_port, plus2A_s_10_port, plus2A_s_9_port, plus2A_s_8_port, 
      plus2A_s_7_port, plus2A_s_6_port, plus2A_s_5_port, plus2A_s_4_port, 
      plus2A_s_3_port, plus2A_s_2_port, plus2A_s_1_port, minus2A_s_63_port, 
      minus2A_s_62_port, minus2A_s_61_port, minus2A_s_60_port, 
      minus2A_s_59_port, minus2A_s_58_port, minus2A_s_57_port, 
      minus2A_s_56_port, minus2A_s_55_port, minus2A_s_54_port, 
      minus2A_s_53_port, minus2A_s_52_port, minus2A_s_51_port, 
      minus2A_s_50_port, minus2A_s_49_port, minus2A_s_48_port, 
      minus2A_s_47_port, minus2A_s_46_port, minus2A_s_45_port, 
      minus2A_s_44_port, minus2A_s_43_port, minus2A_s_42_port, 
      minus2A_s_41_port, minus2A_s_40_port, minus2A_s_39_port, 
      minus2A_s_38_port, minus2A_s_37_port, minus2A_s_36_port, 
      minus2A_s_35_port, minus2A_s_34_port, minus2A_s_33_port, 
      minus2A_s_32_port, minus2A_s_31_port, minus2A_s_30_port, 
      minus2A_s_29_port, minus2A_s_28_port, minus2A_s_27_port, 
      minus2A_s_26_port, minus2A_s_25_port, minus2A_s_24_port, 
      minus2A_s_23_port, minus2A_s_22_port, minus2A_s_21_port, 
      minus2A_s_20_port, minus2A_s_19_port, minus2A_s_18_port, 
      minus2A_s_17_port, minus2A_s_16_port, minus2A_s_15_port, 
      minus2A_s_14_port, minus2A_s_13_port, minus2A_s_12_port, 
      minus2A_s_11_port, minus2A_s_10_port, minus2A_s_9_port, minus2A_s_8_port,
      minus2A_s_7_port, minus2A_s_6_port, minus2A_s_5_port, minus2A_s_4_port, 
      minus2A_s_3_port, minus2A_s_2_port, minus2A_s_1_port, minus2A_s_0_port, 
      minus4A_s_63_port, minus4A_s_62_port, minus4A_s_61_port, 
      minus4A_s_60_port, minus4A_s_59_port, minus4A_s_58_port, 
      minus4A_s_57_port, minus4A_s_56_port, minus4A_s_55_port, 
      minus4A_s_54_port, minus4A_s_53_port, minus4A_s_52_port, 
      minus4A_s_51_port, minus4A_s_50_port, minus4A_s_49_port, 
      minus4A_s_48_port, minus4A_s_47_port, minus4A_s_46_port, 
      minus4A_s_45_port, minus4A_s_44_port, minus4A_s_43_port, 
      minus4A_s_42_port, minus4A_s_41_port, minus4A_s_40_port, 
      minus4A_s_39_port, minus4A_s_38_port, minus4A_s_37_port, 
      minus4A_s_36_port, minus4A_s_35_port, minus4A_s_34_port, 
      minus4A_s_33_port, minus4A_s_32_port, minus4A_s_31_port, 
      minus4A_s_30_port, minus4A_s_29_port, minus4A_s_28_port, 
      minus4A_s_27_port, minus4A_s_26_port, minus4A_s_25_port, 
      minus4A_s_24_port, minus4A_s_23_port, minus4A_s_22_port, 
      minus4A_s_21_port, minus4A_s_20_port, minus4A_s_19_port, 
      minus4A_s_18_port, minus4A_s_17_port, minus4A_s_16_port, 
      minus4A_s_15_port, minus4A_s_14_port, minus4A_s_13_port, 
      minus4A_s_12_port, minus4A_s_11_port, minus4A_s_10_port, minus4A_s_9_port
      , minus4A_s_8_port, minus4A_s_7_port, minus4A_s_6_port, minus4A_s_5_port,
      minus4A_s_4_port, minus4A_s_3_port, minus4A_s_2_port, minus4A_s_1_port, 
      minus4A_s_0_port, mux_to_adder_63_port, mux_to_adder_62_port, 
      mux_to_adder_61_port, mux_to_adder_60_port, mux_to_adder_59_port, 
      mux_to_adder_58_port, mux_to_adder_57_port, mux_to_adder_56_port, 
      mux_to_adder_55_port, mux_to_adder_54_port, mux_to_adder_53_port, 
      mux_to_adder_52_port, mux_to_adder_51_port, mux_to_adder_50_port, 
      mux_to_adder_49_port, mux_to_adder_48_port, mux_to_adder_47_port, 
      mux_to_adder_46_port, mux_to_adder_45_port, mux_to_adder_44_port, 
      mux_to_adder_43_port, mux_to_adder_42_port, mux_to_adder_41_port, 
      mux_to_adder_40_port, mux_to_adder_39_port, mux_to_adder_38_port, 
      mux_to_adder_37_port, mux_to_adder_36_port, mux_to_adder_35_port, 
      mux_to_adder_34_port, mux_to_adder_33_port, mux_to_adder_32_port, 
      mux_to_adder_31_port, mux_to_adder_30_port, mux_to_adder_29_port, 
      mux_to_adder_28_port, mux_to_adder_27_port, mux_to_adder_26_port, 
      mux_to_adder_25_port, mux_to_adder_24_port, mux_to_adder_23_port, 
      mux_to_adder_22_port, mux_to_adder_21_port, mux_to_adder_20_port, 
      mux_to_adder_19_port, mux_to_adder_18_port, mux_to_adder_17_port, 
      mux_to_adder_16_port, mux_to_adder_15_port, mux_to_adder_14_port, 
      mux_to_adder_13_port, mux_to_adder_12_port, mux_to_adder_11_port, 
      mux_to_adder_10_port, mux_to_adder_9_port, mux_to_adder_8_port, 
      mux_to_adder_7_port, mux_to_adder_6_port, mux_to_adder_5_port, 
      mux_to_adder_4_port, mux_to_adder_3_port, mux_to_adder_2_port, 
      mux_to_adder_1_port, mux_to_adder_0_port, nextA_0_port, nextA_57_port, 
      n_3193, n_3194, n_3195 : std_logic;

begin
   nextA <= ( nextA_63_port, nextA_62_port, nextA_61_port, nextA_60_port, 
      nextA_59_port, nextA_58_port, nextA_57_port, nextA_56_port, nextA_55_port
      , nextA_54_port, nextA_53_port, nextA_52_port, nextA_51_port, 
      nextA_50_port, nextA_49_port, nextA_48_port, nextA_47_port, nextA_46_port
      , nextA_45_port, nextA_44_port, nextA_43_port, nextA_42_port, 
      nextA_41_port, nextA_40_port, nextA_39_port, nextA_38_port, nextA_37_port
      , nextA_36_port, nextA_35_port, nextA_34_port, nextA_33_port, 
      nextA_32_port, nextA_31_port, nextA_30_port, nextA_29_port, nextA_28_port
      , nextA_27_port, nextA_26_port, nextA_25_port, nextA_24_port, 
      nextA_23_port, nextA_22_port, nextA_21_port, nextA_20_port, nextA_19_port
      , nextA_18_port, nextA_17_port, nextA_16_port, nextA_15_port, 
      nextA_14_port, nextA_13_port, nextA_12_port, nextA_11_port, nextA_10_port
      , nextA_9_port, nextA_8_port, nextA_7_port, nextA_6_port, nextA_5_port, 
      nextA_4_port, nextA_3_port, nextA_2_port, nextA_1_port, nextA_0_port );
   
   X_Logic0_port <= '0';
   nextA_0_port <= '0';
   encoder_1 : encoder_N64_RADIX3_7 port map( X(2) => encoderIn(2), X(1) => 
                           encoderIn(1), X(0) => encoderIn(0), Z(2) => 
                           encoder_to_mux_2_port, Z(1) => encoder_to_mux_1_port
                           , Z(0) => encoder_to_mux_0_port);
   ShiftnCompl_1 : ShiftnCompl_N64_7 port map( plusA(63) => prevA(63), 
                           plusA(62) => prevA(62), plusA(61) => prevA(61), 
                           plusA(60) => prevA(60), plusA(59) => prevA(59), 
                           plusA(58) => prevA(58), plusA(57) => prevA(57), 
                           plusA(56) => prevA(56), plusA(55) => prevA(55), 
                           plusA(54) => prevA(54), plusA(53) => prevA(53), 
                           plusA(52) => prevA(52), plusA(51) => prevA(51), 
                           plusA(50) => prevA(50), plusA(49) => prevA(49), 
                           plusA(48) => prevA(48), plusA(47) => prevA(47), 
                           plusA(46) => prevA(46), plusA(45) => prevA(45), 
                           plusA(44) => prevA(44), plusA(43) => prevA(43), 
                           plusA(42) => prevA(42), plusA(41) => prevA(41), 
                           plusA(40) => prevA(40), plusA(39) => prevA(39), 
                           plusA(38) => prevA(38), plusA(37) => prevA(37), 
                           plusA(36) => prevA(36), plusA(35) => prevA(35), 
                           plusA(34) => prevA(34), plusA(33) => prevA(33), 
                           plusA(32) => prevA(32), plusA(31) => prevA(31), 
                           plusA(30) => prevA(30), plusA(29) => prevA(29), 
                           plusA(28) => prevA(28), plusA(27) => prevA(27), 
                           plusA(26) => prevA(26), plusA(25) => prevA(25), 
                           plusA(24) => prevA(24), plusA(23) => prevA(23), 
                           plusA(22) => prevA(22), plusA(21) => prevA(21), 
                           plusA(20) => prevA(20), plusA(19) => prevA(19), 
                           plusA(18) => prevA(18), plusA(17) => prevA(17), 
                           plusA(16) => prevA(16), plusA(15) => prevA(15), 
                           plusA(14) => prevA(14), plusA(13) => prevA(13), 
                           plusA(12) => prevA(12), plusA(11) => prevA(11), 
                           plusA(10) => prevA(10), plusA(9) => prevA(9), 
                           plusA(8) => prevA(8), plusA(7) => prevA(7), plusA(6)
                           => prevA(6), plusA(5) => prevA(5), plusA(4) => 
                           prevA(4), plusA(3) => prevA(3), plusA(2) => prevA(2)
                           , plusA(1) => prevA(1), plusA(0) => prevA(0), 
                           plus2A_out(63) => plus2A_s_63_port, plus2A_out(62) 
                           => plus2A_s_62_port, plus2A_out(61) => 
                           plus2A_s_61_port, plus2A_out(60) => plus2A_s_60_port
                           , plus2A_out(59) => plus2A_s_59_port, plus2A_out(58)
                           => plus2A_s_58_port, plus2A_out(57) => 
                           plus2A_s_57_port, plus2A_out(56) => plus2A_s_56_port
                           , plus2A_out(55) => plus2A_s_55_port, plus2A_out(54)
                           => plus2A_s_54_port, plus2A_out(53) => 
                           plus2A_s_53_port, plus2A_out(52) => plus2A_s_52_port
                           , plus2A_out(51) => plus2A_s_51_port, plus2A_out(50)
                           => plus2A_s_50_port, plus2A_out(49) => 
                           plus2A_s_49_port, plus2A_out(48) => plus2A_s_48_port
                           , plus2A_out(47) => plus2A_s_47_port, plus2A_out(46)
                           => plus2A_s_46_port, plus2A_out(45) => 
                           plus2A_s_45_port, plus2A_out(44) => plus2A_s_44_port
                           , plus2A_out(43) => plus2A_s_43_port, plus2A_out(42)
                           => plus2A_s_42_port, plus2A_out(41) => 
                           plus2A_s_41_port, plus2A_out(40) => plus2A_s_40_port
                           , plus2A_out(39) => plus2A_s_39_port, plus2A_out(38)
                           => plus2A_s_38_port, plus2A_out(37) => 
                           plus2A_s_37_port, plus2A_out(36) => plus2A_s_36_port
                           , plus2A_out(35) => plus2A_s_35_port, plus2A_out(34)
                           => plus2A_s_34_port, plus2A_out(33) => 
                           plus2A_s_33_port, plus2A_out(32) => plus2A_s_32_port
                           , plus2A_out(31) => plus2A_s_31_port, plus2A_out(30)
                           => plus2A_s_30_port, plus2A_out(29) => 
                           plus2A_s_29_port, plus2A_out(28) => plus2A_s_28_port
                           , plus2A_out(27) => plus2A_s_27_port, plus2A_out(26)
                           => plus2A_s_26_port, plus2A_out(25) => 
                           plus2A_s_25_port, plus2A_out(24) => plus2A_s_24_port
                           , plus2A_out(23) => plus2A_s_23_port, plus2A_out(22)
                           => plus2A_s_22_port, plus2A_out(21) => 
                           plus2A_s_21_port, plus2A_out(20) => plus2A_s_20_port
                           , plus2A_out(19) => plus2A_s_19_port, plus2A_out(18)
                           => plus2A_s_18_port, plus2A_out(17) => 
                           plus2A_s_17_port, plus2A_out(16) => plus2A_s_16_port
                           , plus2A_out(15) => plus2A_s_15_port, plus2A_out(14)
                           => plus2A_s_14_port, plus2A_out(13) => 
                           plus2A_s_13_port, plus2A_out(12) => plus2A_s_12_port
                           , plus2A_out(11) => plus2A_s_11_port, plus2A_out(10)
                           => plus2A_s_10_port, plus2A_out(9) => 
                           plus2A_s_9_port, plus2A_out(8) => plus2A_s_8_port, 
                           plus2A_out(7) => plus2A_s_7_port, plus2A_out(6) => 
                           plus2A_s_6_port, plus2A_out(5) => plus2A_s_5_port, 
                           plus2A_out(4) => plus2A_s_4_port, plus2A_out(3) => 
                           plus2A_s_3_port, plus2A_out(2) => plus2A_s_2_port, 
                           plus2A_out(1) => plus2A_s_1_port, plus2A_out(0) => 
                           n_3193, minus2A_out(63) => minus2A_s_63_port, 
                           minus2A_out(62) => minus2A_s_62_port, 
                           minus2A_out(61) => minus2A_s_61_port, 
                           minus2A_out(60) => minus2A_s_60_port, 
                           minus2A_out(59) => minus2A_s_59_port, 
                           minus2A_out(58) => minus2A_s_58_port, 
                           minus2A_out(57) => minus2A_s_57_port, 
                           minus2A_out(56) => minus2A_s_56_port, 
                           minus2A_out(55) => minus2A_s_55_port, 
                           minus2A_out(54) => minus2A_s_54_port, 
                           minus2A_out(53) => minus2A_s_53_port, 
                           minus2A_out(52) => minus2A_s_52_port, 
                           minus2A_out(51) => minus2A_s_51_port, 
                           minus2A_out(50) => minus2A_s_50_port, 
                           minus2A_out(49) => minus2A_s_49_port, 
                           minus2A_out(48) => minus2A_s_48_port, 
                           minus2A_out(47) => minus2A_s_47_port, 
                           minus2A_out(46) => minus2A_s_46_port, 
                           minus2A_out(45) => minus2A_s_45_port, 
                           minus2A_out(44) => minus2A_s_44_port, 
                           minus2A_out(43) => minus2A_s_43_port, 
                           minus2A_out(42) => minus2A_s_42_port, 
                           minus2A_out(41) => minus2A_s_41_port, 
                           minus2A_out(40) => minus2A_s_40_port, 
                           minus2A_out(39) => minus2A_s_39_port, 
                           minus2A_out(38) => minus2A_s_38_port, 
                           minus2A_out(37) => minus2A_s_37_port, 
                           minus2A_out(36) => minus2A_s_36_port, 
                           minus2A_out(35) => minus2A_s_35_port, 
                           minus2A_out(34) => minus2A_s_34_port, 
                           minus2A_out(33) => minus2A_s_33_port, 
                           minus2A_out(32) => minus2A_s_32_port, 
                           minus2A_out(31) => minus2A_s_31_port, 
                           minus2A_out(30) => minus2A_s_30_port, 
                           minus2A_out(29) => minus2A_s_29_port, 
                           minus2A_out(28) => minus2A_s_28_port, 
                           minus2A_out(27) => minus2A_s_27_port, 
                           minus2A_out(26) => minus2A_s_26_port, 
                           minus2A_out(25) => minus2A_s_25_port, 
                           minus2A_out(24) => minus2A_s_24_port, 
                           minus2A_out(23) => minus2A_s_23_port, 
                           minus2A_out(22) => minus2A_s_22_port, 
                           minus2A_out(21) => minus2A_s_21_port, 
                           minus2A_out(20) => minus2A_s_20_port, 
                           minus2A_out(19) => minus2A_s_19_port, 
                           minus2A_out(18) => minus2A_s_18_port, 
                           minus2A_out(17) => minus2A_s_17_port, 
                           minus2A_out(16) => minus2A_s_16_port, 
                           minus2A_out(15) => minus2A_s_15_port, 
                           minus2A_out(14) => minus2A_s_14_port, 
                           minus2A_out(13) => minus2A_s_13_port, 
                           minus2A_out(12) => minus2A_s_12_port, 
                           minus2A_out(11) => minus2A_s_11_port, 
                           minus2A_out(10) => minus2A_s_10_port, minus2A_out(9)
                           => minus2A_s_9_port, minus2A_out(8) => 
                           minus2A_s_8_port, minus2A_out(7) => minus2A_s_7_port
                           , minus2A_out(6) => minus2A_s_6_port, minus2A_out(5)
                           => minus2A_s_5_port, minus2A_out(4) => 
                           minus2A_s_4_port, minus2A_out(3) => minus2A_s_3_port
                           , minus2A_out(2) => minus2A_s_2_port, minus2A_out(1)
                           => minus2A_s_1_port, minus2A_out(0) => 
                           minus2A_s_0_port, plus4A_out(63) => nextA_63_port, 
                           plus4A_out(62) => nextA_62_port, plus4A_out(61) => 
                           nextA_61_port, plus4A_out(60) => nextA_60_port, 
                           plus4A_out(59) => nextA_59_port, plus4A_out(58) => 
                           nextA_58_port, plus4A_out(57) => n3, plus4A_out(56) 
                           => nextA_56_port, plus4A_out(55) => nextA_55_port, 
                           plus4A_out(54) => nextA_54_port, plus4A_out(53) => 
                           nextA_53_port, plus4A_out(52) => nextA_52_port, 
                           plus4A_out(51) => nextA_51_port, plus4A_out(50) => 
                           nextA_50_port, plus4A_out(49) => nextA_49_port, 
                           plus4A_out(48) => nextA_48_port, plus4A_out(47) => 
                           nextA_47_port, plus4A_out(46) => nextA_46_port, 
                           plus4A_out(45) => nextA_45_port, plus4A_out(44) => 
                           nextA_44_port, plus4A_out(43) => nextA_43_port, 
                           plus4A_out(42) => nextA_42_port, plus4A_out(41) => 
                           nextA_41_port, plus4A_out(40) => nextA_40_port, 
                           plus4A_out(39) => nextA_39_port, plus4A_out(38) => 
                           nextA_38_port, plus4A_out(37) => nextA_37_port, 
                           plus4A_out(36) => nextA_36_port, plus4A_out(35) => 
                           nextA_35_port, plus4A_out(34) => nextA_34_port, 
                           plus4A_out(33) => nextA_33_port, plus4A_out(32) => 
                           nextA_32_port, plus4A_out(31) => nextA_31_port, 
                           plus4A_out(30) => nextA_30_port, plus4A_out(29) => 
                           nextA_29_port, plus4A_out(28) => nextA_28_port, 
                           plus4A_out(27) => nextA_27_port, plus4A_out(26) => 
                           nextA_26_port, plus4A_out(25) => nextA_25_port, 
                           plus4A_out(24) => nextA_24_port, plus4A_out(23) => 
                           nextA_23_port, plus4A_out(22) => nextA_22_port, 
                           plus4A_out(21) => nextA_21_port, plus4A_out(20) => 
                           nextA_20_port, plus4A_out(19) => nextA_19_port, 
                           plus4A_out(18) => nextA_18_port, plus4A_out(17) => 
                           nextA_17_port, plus4A_out(16) => nextA_16_port, 
                           plus4A_out(15) => nextA_15_port, plus4A_out(14) => 
                           nextA_14_port, plus4A_out(13) => nextA_13_port, 
                           plus4A_out(12) => nextA_12_port, plus4A_out(11) => 
                           nextA_11_port, plus4A_out(10) => nextA_10_port, 
                           plus4A_out(9) => nextA_9_port, plus4A_out(8) => 
                           nextA_8_port, plus4A_out(7) => nextA_7_port, 
                           plus4A_out(6) => nextA_6_port, plus4A_out(5) => 
                           nextA_5_port, plus4A_out(4) => nextA_4_port, 
                           plus4A_out(3) => nextA_3_port, plus4A_out(2) => 
                           nextA_2_port, plus4A_out(1) => nextA_1_port, 
                           plus4A_out(0) => n_3194, minus4A_out(63) => 
                           minus4A_s_63_port, minus4A_out(62) => 
                           minus4A_s_62_port, minus4A_out(61) => 
                           minus4A_s_61_port, minus4A_out(60) => 
                           minus4A_s_60_port, minus4A_out(59) => 
                           minus4A_s_59_port, minus4A_out(58) => 
                           minus4A_s_58_port, minus4A_out(57) => 
                           minus4A_s_57_port, minus4A_out(56) => 
                           minus4A_s_56_port, minus4A_out(55) => 
                           minus4A_s_55_port, minus4A_out(54) => 
                           minus4A_s_54_port, minus4A_out(53) => 
                           minus4A_s_53_port, minus4A_out(52) => 
                           minus4A_s_52_port, minus4A_out(51) => 
                           minus4A_s_51_port, minus4A_out(50) => 
                           minus4A_s_50_port, minus4A_out(49) => 
                           minus4A_s_49_port, minus4A_out(48) => 
                           minus4A_s_48_port, minus4A_out(47) => 
                           minus4A_s_47_port, minus4A_out(46) => 
                           minus4A_s_46_port, minus4A_out(45) => 
                           minus4A_s_45_port, minus4A_out(44) => 
                           minus4A_s_44_port, minus4A_out(43) => 
                           minus4A_s_43_port, minus4A_out(42) => 
                           minus4A_s_42_port, minus4A_out(41) => 
                           minus4A_s_41_port, minus4A_out(40) => 
                           minus4A_s_40_port, minus4A_out(39) => 
                           minus4A_s_39_port, minus4A_out(38) => 
                           minus4A_s_38_port, minus4A_out(37) => 
                           minus4A_s_37_port, minus4A_out(36) => 
                           minus4A_s_36_port, minus4A_out(35) => 
                           minus4A_s_35_port, minus4A_out(34) => 
                           minus4A_s_34_port, minus4A_out(33) => 
                           minus4A_s_33_port, minus4A_out(32) => 
                           minus4A_s_32_port, minus4A_out(31) => 
                           minus4A_s_31_port, minus4A_out(30) => 
                           minus4A_s_30_port, minus4A_out(29) => 
                           minus4A_s_29_port, minus4A_out(28) => 
                           minus4A_s_28_port, minus4A_out(27) => 
                           minus4A_s_27_port, minus4A_out(26) => 
                           minus4A_s_26_port, minus4A_out(25) => 
                           minus4A_s_25_port, minus4A_out(24) => 
                           minus4A_s_24_port, minus4A_out(23) => 
                           minus4A_s_23_port, minus4A_out(22) => 
                           minus4A_s_22_port, minus4A_out(21) => 
                           minus4A_s_21_port, minus4A_out(20) => 
                           minus4A_s_20_port, minus4A_out(19) => 
                           minus4A_s_19_port, minus4A_out(18) => 
                           minus4A_s_18_port, minus4A_out(17) => 
                           minus4A_s_17_port, minus4A_out(16) => 
                           minus4A_s_16_port, minus4A_out(15) => 
                           minus4A_s_15_port, minus4A_out(14) => 
                           minus4A_s_14_port, minus4A_out(13) => 
                           minus4A_s_13_port, minus4A_out(12) => 
                           minus4A_s_12_port, minus4A_out(11) => 
                           minus4A_s_11_port, minus4A_out(10) => 
                           minus4A_s_10_port, minus4A_out(9) => 
                           minus4A_s_9_port, minus4A_out(8) => minus4A_s_8_port
                           , minus4A_out(7) => minus4A_s_7_port, minus4A_out(6)
                           => minus4A_s_6_port, minus4A_out(5) => 
                           minus4A_s_5_port, minus4A_out(4) => minus4A_s_4_port
                           , minus4A_out(3) => minus4A_s_3_port, minus4A_out(2)
                           => minus4A_s_2_port, minus4A_out(1) => 
                           minus4A_s_1_port, minus4A_out(0) => minus4A_s_0_port
                           );
   mux_1 : MUX_GENERIC_N64_RADIX3_7 port map( plusA(63) => plus2A_s_63_port, 
                           plusA(62) => plus2A_s_62_port, plusA(61) => 
                           plus2A_s_61_port, plusA(60) => plus2A_s_60_port, 
                           plusA(59) => plus2A_s_59_port, plusA(58) => 
                           plus2A_s_58_port, plusA(57) => plus2A_s_57_port, 
                           plusA(56) => plus2A_s_56_port, plusA(55) => 
                           plus2A_s_55_port, plusA(54) => plus2A_s_54_port, 
                           plusA(53) => plus2A_s_53_port, plusA(52) => 
                           plus2A_s_52_port, plusA(51) => plus2A_s_51_port, 
                           plusA(50) => plus2A_s_50_port, plusA(49) => 
                           plus2A_s_49_port, plusA(48) => plus2A_s_48_port, 
                           plusA(47) => plus2A_s_47_port, plusA(46) => 
                           plus2A_s_46_port, plusA(45) => plus2A_s_45_port, 
                           plusA(44) => plus2A_s_44_port, plusA(43) => 
                           plus2A_s_43_port, plusA(42) => plus2A_s_42_port, 
                           plusA(41) => plus2A_s_41_port, plusA(40) => 
                           plus2A_s_40_port, plusA(39) => plus2A_s_39_port, 
                           plusA(38) => plus2A_s_38_port, plusA(37) => 
                           plus2A_s_37_port, plusA(36) => plus2A_s_36_port, 
                           plusA(35) => plus2A_s_35_port, plusA(34) => 
                           plus2A_s_34_port, plusA(33) => plus2A_s_33_port, 
                           plusA(32) => plus2A_s_32_port, plusA(31) => 
                           plus2A_s_31_port, plusA(30) => plus2A_s_30_port, 
                           plusA(29) => plus2A_s_29_port, plusA(28) => 
                           plus2A_s_28_port, plusA(27) => plus2A_s_27_port, 
                           plusA(26) => plus2A_s_26_port, plusA(25) => 
                           plus2A_s_25_port, plusA(24) => plus2A_s_24_port, 
                           plusA(23) => plus2A_s_23_port, plusA(22) => 
                           plus2A_s_22_port, plusA(21) => plus2A_s_21_port, 
                           plusA(20) => plus2A_s_20_port, plusA(19) => 
                           plus2A_s_19_port, plusA(18) => plus2A_s_18_port, 
                           plusA(17) => plus2A_s_17_port, plusA(16) => 
                           plus2A_s_16_port, plusA(15) => plus2A_s_15_port, 
                           plusA(14) => plus2A_s_14_port, plusA(13) => 
                           plus2A_s_13_port, plusA(12) => plus2A_s_12_port, 
                           plusA(11) => plus2A_s_11_port, plusA(10) => 
                           plus2A_s_10_port, plusA(9) => plus2A_s_9_port, 
                           plusA(8) => plus2A_s_8_port, plusA(7) => 
                           plus2A_s_7_port, plusA(6) => plus2A_s_6_port, 
                           plusA(5) => plus2A_s_5_port, plusA(4) => 
                           plus2A_s_4_port, plusA(3) => plus2A_s_3_port, 
                           plusA(2) => plus2A_s_2_port, plusA(1) => 
                           plus2A_s_1_port, plusA(0) => nextA_0_port, 
                           minusA(63) => minus2A_s_63_port, minusA(62) => 
                           minus2A_s_62_port, minusA(61) => minus2A_s_61_port, 
                           minusA(60) => minus2A_s_60_port, minusA(59) => 
                           minus2A_s_59_port, minusA(58) => minus2A_s_58_port, 
                           minusA(57) => minus2A_s_57_port, minusA(56) => 
                           minus2A_s_56_port, minusA(55) => minus2A_s_55_port, 
                           minusA(54) => minus2A_s_54_port, minusA(53) => 
                           minus2A_s_53_port, minusA(52) => minus2A_s_52_port, 
                           minusA(51) => minus2A_s_51_port, minusA(50) => 
                           minus2A_s_50_port, minusA(49) => minus2A_s_49_port, 
                           minusA(48) => minus2A_s_48_port, minusA(47) => 
                           minus2A_s_47_port, minusA(46) => minus2A_s_46_port, 
                           minusA(45) => minus2A_s_45_port, minusA(44) => 
                           minus2A_s_44_port, minusA(43) => minus2A_s_43_port, 
                           minusA(42) => minus2A_s_42_port, minusA(41) => 
                           minus2A_s_41_port, minusA(40) => minus2A_s_40_port, 
                           minusA(39) => minus2A_s_39_port, minusA(38) => 
                           minus2A_s_38_port, minusA(37) => minus2A_s_37_port, 
                           minusA(36) => minus2A_s_36_port, minusA(35) => 
                           minus2A_s_35_port, minusA(34) => minus2A_s_34_port, 
                           minusA(33) => minus2A_s_33_port, minusA(32) => 
                           minus2A_s_32_port, minusA(31) => minus2A_s_31_port, 
                           minusA(30) => minus2A_s_30_port, minusA(29) => 
                           minus2A_s_29_port, minusA(28) => minus2A_s_28_port, 
                           minusA(27) => minus2A_s_27_port, minusA(26) => 
                           minus2A_s_26_port, minusA(25) => minus2A_s_25_port, 
                           minusA(24) => minus2A_s_24_port, minusA(23) => 
                           minus2A_s_23_port, minusA(22) => minus2A_s_22_port, 
                           minusA(21) => minus2A_s_21_port, minusA(20) => 
                           minus2A_s_20_port, minusA(19) => minus2A_s_19_port, 
                           minusA(18) => minus2A_s_18_port, minusA(17) => 
                           minus2A_s_17_port, minusA(16) => minus2A_s_16_port, 
                           minusA(15) => minus2A_s_15_port, minusA(14) => 
                           minus2A_s_14_port, minusA(13) => minus2A_s_13_port, 
                           minusA(12) => minus2A_s_12_port, minusA(11) => 
                           minus2A_s_11_port, minusA(10) => minus2A_s_10_port, 
                           minusA(9) => minus2A_s_9_port, minusA(8) => 
                           minus2A_s_8_port, minusA(7) => minus2A_s_7_port, 
                           minusA(6) => minus2A_s_6_port, minusA(5) => 
                           minus2A_s_5_port, minusA(4) => minus2A_s_4_port, 
                           minusA(3) => minus2A_s_3_port, minusA(2) => 
                           minus2A_s_2_port, minusA(1) => minus2A_s_1_port, 
                           minusA(0) => minus2A_s_0_port, plus2A(63) => 
                           nextA_63_port, plus2A(62) => nextA_62_port, 
                           plus2A(61) => nextA_61_port, plus2A(60) => 
                           nextA_60_port, plus2A(59) => nextA_59_port, 
                           plus2A(58) => nextA_58_port, plus2A(57) => 
                           nextA_57_port, plus2A(56) => nextA_56_port, 
                           plus2A(55) => nextA_55_port, plus2A(54) => 
                           nextA_54_port, plus2A(53) => nextA_53_port, 
                           plus2A(52) => nextA_52_port, plus2A(51) => 
                           nextA_51_port, plus2A(50) => nextA_50_port, 
                           plus2A(49) => nextA_49_port, plus2A(48) => 
                           nextA_48_port, plus2A(47) => nextA_47_port, 
                           plus2A(46) => nextA_46_port, plus2A(45) => 
                           nextA_45_port, plus2A(44) => nextA_44_port, 
                           plus2A(43) => nextA_43_port, plus2A(42) => 
                           nextA_42_port, plus2A(41) => nextA_41_port, 
                           plus2A(40) => nextA_40_port, plus2A(39) => 
                           nextA_39_port, plus2A(38) => nextA_38_port, 
                           plus2A(37) => nextA_37_port, plus2A(36) => 
                           nextA_36_port, plus2A(35) => nextA_35_port, 
                           plus2A(34) => nextA_34_port, plus2A(33) => 
                           nextA_33_port, plus2A(32) => nextA_32_port, 
                           plus2A(31) => nextA_31_port, plus2A(30) => 
                           nextA_30_port, plus2A(29) => nextA_29_port, 
                           plus2A(28) => nextA_28_port, plus2A(27) => 
                           nextA_27_port, plus2A(26) => nextA_26_port, 
                           plus2A(25) => nextA_25_port, plus2A(24) => 
                           nextA_24_port, plus2A(23) => nextA_23_port, 
                           plus2A(22) => nextA_22_port, plus2A(21) => 
                           nextA_21_port, plus2A(20) => nextA_20_port, 
                           plus2A(19) => nextA_19_port, plus2A(18) => 
                           nextA_18_port, plus2A(17) => nextA_17_port, 
                           plus2A(16) => nextA_16_port, plus2A(15) => 
                           nextA_15_port, plus2A(14) => nextA_14_port, 
                           plus2A(13) => nextA_13_port, plus2A(12) => 
                           nextA_12_port, plus2A(11) => nextA_11_port, 
                           plus2A(10) => nextA_10_port, plus2A(9) => 
                           nextA_9_port, plus2A(8) => nextA_8_port, plus2A(7) 
                           => nextA_7_port, plus2A(6) => nextA_6_port, 
                           plus2A(5) => nextA_5_port, plus2A(4) => nextA_4_port
                           , plus2A(3) => nextA_3_port, plus2A(2) => 
                           nextA_2_port, plus2A(1) => nextA_1_port, plus2A(0) 
                           => nextA_0_port, minus2A(63) => minus4A_s_63_port, 
                           minus2A(62) => minus4A_s_62_port, minus2A(61) => 
                           minus4A_s_61_port, minus2A(60) => minus4A_s_60_port,
                           minus2A(59) => minus4A_s_59_port, minus2A(58) => 
                           minus4A_s_58_port, minus2A(57) => minus4A_s_57_port,
                           minus2A(56) => minus4A_s_56_port, minus2A(55) => 
                           minus4A_s_55_port, minus2A(54) => minus4A_s_54_port,
                           minus2A(53) => minus4A_s_53_port, minus2A(52) => 
                           minus4A_s_52_port, minus2A(51) => minus4A_s_51_port,
                           minus2A(50) => minus4A_s_50_port, minus2A(49) => 
                           minus4A_s_49_port, minus2A(48) => minus4A_s_48_port,
                           minus2A(47) => minus4A_s_47_port, minus2A(46) => 
                           minus4A_s_46_port, minus2A(45) => minus4A_s_45_port,
                           minus2A(44) => minus4A_s_44_port, minus2A(43) => 
                           minus4A_s_43_port, minus2A(42) => minus4A_s_42_port,
                           minus2A(41) => minus4A_s_41_port, minus2A(40) => 
                           minus4A_s_40_port, minus2A(39) => minus4A_s_39_port,
                           minus2A(38) => minus4A_s_38_port, minus2A(37) => 
                           minus4A_s_37_port, minus2A(36) => minus4A_s_36_port,
                           minus2A(35) => minus4A_s_35_port, minus2A(34) => 
                           minus4A_s_34_port, minus2A(33) => minus4A_s_33_port,
                           minus2A(32) => minus4A_s_32_port, minus2A(31) => 
                           minus4A_s_31_port, minus2A(30) => minus4A_s_30_port,
                           minus2A(29) => minus4A_s_29_port, minus2A(28) => 
                           minus4A_s_28_port, minus2A(27) => minus4A_s_27_port,
                           minus2A(26) => minus4A_s_26_port, minus2A(25) => 
                           minus4A_s_25_port, minus2A(24) => minus4A_s_24_port,
                           minus2A(23) => minus4A_s_23_port, minus2A(22) => 
                           minus4A_s_22_port, minus2A(21) => minus4A_s_21_port,
                           minus2A(20) => minus4A_s_20_port, minus2A(19) => 
                           minus4A_s_19_port, minus2A(18) => minus4A_s_18_port,
                           minus2A(17) => minus4A_s_17_port, minus2A(16) => 
                           minus4A_s_16_port, minus2A(15) => minus4A_s_15_port,
                           minus2A(14) => minus4A_s_14_port, minus2A(13) => 
                           minus4A_s_13_port, minus2A(12) => minus4A_s_12_port,
                           minus2A(11) => minus4A_s_11_port, minus2A(10) => 
                           minus4A_s_10_port, minus2A(9) => minus4A_s_9_port, 
                           minus2A(8) => minus4A_s_8_port, minus2A(7) => 
                           minus4A_s_7_port, minus2A(6) => minus4A_s_6_port, 
                           minus2A(5) => minus4A_s_5_port, minus2A(4) => 
                           minus4A_s_4_port, minus2A(3) => minus4A_s_3_port, 
                           minus2A(2) => minus4A_s_2_port, minus2A(1) => 
                           minus4A_s_1_port, minus2A(0) => minus4A_s_0_port, 
                           SEL(2) => encoder_to_mux_2_port, SEL(1) => 
                           encoder_to_mux_1_port, SEL(0) => 
                           encoder_to_mux_0_port, Y(63) => mux_to_adder_63_port
                           , Y(62) => mux_to_adder_62_port, Y(61) => 
                           mux_to_adder_61_port, Y(60) => mux_to_adder_60_port,
                           Y(59) => mux_to_adder_59_port, Y(58) => 
                           mux_to_adder_58_port, Y(57) => mux_to_adder_57_port,
                           Y(56) => mux_to_adder_56_port, Y(55) => 
                           mux_to_adder_55_port, Y(54) => mux_to_adder_54_port,
                           Y(53) => mux_to_adder_53_port, Y(52) => 
                           mux_to_adder_52_port, Y(51) => mux_to_adder_51_port,
                           Y(50) => mux_to_adder_50_port, Y(49) => 
                           mux_to_adder_49_port, Y(48) => mux_to_adder_48_port,
                           Y(47) => mux_to_adder_47_port, Y(46) => 
                           mux_to_adder_46_port, Y(45) => mux_to_adder_45_port,
                           Y(44) => mux_to_adder_44_port, Y(43) => 
                           mux_to_adder_43_port, Y(42) => mux_to_adder_42_port,
                           Y(41) => mux_to_adder_41_port, Y(40) => 
                           mux_to_adder_40_port, Y(39) => mux_to_adder_39_port,
                           Y(38) => mux_to_adder_38_port, Y(37) => 
                           mux_to_adder_37_port, Y(36) => mux_to_adder_36_port,
                           Y(35) => mux_to_adder_35_port, Y(34) => 
                           mux_to_adder_34_port, Y(33) => mux_to_adder_33_port,
                           Y(32) => mux_to_adder_32_port, Y(31) => 
                           mux_to_adder_31_port, Y(30) => mux_to_adder_30_port,
                           Y(29) => mux_to_adder_29_port, Y(28) => 
                           mux_to_adder_28_port, Y(27) => mux_to_adder_27_port,
                           Y(26) => mux_to_adder_26_port, Y(25) => 
                           mux_to_adder_25_port, Y(24) => mux_to_adder_24_port,
                           Y(23) => mux_to_adder_23_port, Y(22) => 
                           mux_to_adder_22_port, Y(21) => mux_to_adder_21_port,
                           Y(20) => mux_to_adder_20_port, Y(19) => 
                           mux_to_adder_19_port, Y(18) => mux_to_adder_18_port,
                           Y(17) => mux_to_adder_17_port, Y(16) => 
                           mux_to_adder_16_port, Y(15) => mux_to_adder_15_port,
                           Y(14) => mux_to_adder_14_port, Y(13) => 
                           mux_to_adder_13_port, Y(12) => mux_to_adder_12_port,
                           Y(11) => mux_to_adder_11_port, Y(10) => 
                           mux_to_adder_10_port, Y(9) => mux_to_adder_9_port, 
                           Y(8) => mux_to_adder_8_port, Y(7) => 
                           mux_to_adder_7_port, Y(6) => mux_to_adder_6_port, 
                           Y(5) => mux_to_adder_5_port, Y(4) => 
                           mux_to_adder_4_port, Y(3) => mux_to_adder_3_port, 
                           Y(2) => mux_to_adder_2_port, Y(1) => 
                           mux_to_adder_1_port, Y(0) => mux_to_adder_0_port);
   rca_1 : RCA_N64_7 port map( A(63) => mux_to_adder_63_port, A(62) => 
                           mux_to_adder_62_port, A(61) => mux_to_adder_61_port,
                           A(60) => mux_to_adder_60_port, A(59) => 
                           mux_to_adder_59_port, A(58) => mux_to_adder_58_port,
                           A(57) => mux_to_adder_57_port, A(56) => 
                           mux_to_adder_56_port, A(55) => mux_to_adder_55_port,
                           A(54) => mux_to_adder_54_port, A(53) => 
                           mux_to_adder_53_port, A(52) => mux_to_adder_52_port,
                           A(51) => mux_to_adder_51_port, A(50) => 
                           mux_to_adder_50_port, A(49) => mux_to_adder_49_port,
                           A(48) => mux_to_adder_48_port, A(47) => 
                           mux_to_adder_47_port, A(46) => mux_to_adder_46_port,
                           A(45) => mux_to_adder_45_port, A(44) => 
                           mux_to_adder_44_port, A(43) => mux_to_adder_43_port,
                           A(42) => mux_to_adder_42_port, A(41) => 
                           mux_to_adder_41_port, A(40) => mux_to_adder_40_port,
                           A(39) => mux_to_adder_39_port, A(38) => 
                           mux_to_adder_38_port, A(37) => mux_to_adder_37_port,
                           A(36) => mux_to_adder_36_port, A(35) => 
                           mux_to_adder_35_port, A(34) => mux_to_adder_34_port,
                           A(33) => mux_to_adder_33_port, A(32) => 
                           mux_to_adder_32_port, A(31) => mux_to_adder_31_port,
                           A(30) => mux_to_adder_30_port, A(29) => 
                           mux_to_adder_29_port, A(28) => mux_to_adder_28_port,
                           A(27) => mux_to_adder_27_port, A(26) => 
                           mux_to_adder_26_port, A(25) => mux_to_adder_25_port,
                           A(24) => mux_to_adder_24_port, A(23) => 
                           mux_to_adder_23_port, A(22) => mux_to_adder_22_port,
                           A(21) => mux_to_adder_21_port, A(20) => 
                           mux_to_adder_20_port, A(19) => mux_to_adder_19_port,
                           A(18) => mux_to_adder_18_port, A(17) => 
                           mux_to_adder_17_port, A(16) => mux_to_adder_16_port,
                           A(15) => mux_to_adder_15_port, A(14) => 
                           mux_to_adder_14_port, A(13) => mux_to_adder_13_port,
                           A(12) => mux_to_adder_12_port, A(11) => 
                           mux_to_adder_11_port, A(10) => mux_to_adder_10_port,
                           A(9) => mux_to_adder_9_port, A(8) => 
                           mux_to_adder_8_port, A(7) => mux_to_adder_7_port, 
                           A(6) => mux_to_adder_6_port, A(5) => 
                           mux_to_adder_5_port, A(4) => mux_to_adder_4_port, 
                           A(3) => mux_to_adder_3_port, A(2) => 
                           mux_to_adder_2_port, A(1) => mux_to_adder_1_port, 
                           A(0) => mux_to_adder_0_port, B(63) => prevSum(63), 
                           B(62) => prevSum(62), B(61) => prevSum(61), B(60) =>
                           prevSum(60), B(59) => prevSum(59), B(58) => 
                           prevSum(58), B(57) => prevSum(57), B(56) => 
                           prevSum(56), B(55) => prevSum(55), B(54) => 
                           prevSum(54), B(53) => prevSum(53), B(52) => 
                           prevSum(52), B(51) => prevSum(51), B(50) => 
                           prevSum(50), B(49) => prevSum(49), B(48) => 
                           prevSum(48), B(47) => prevSum(47), B(46) => 
                           prevSum(46), B(45) => prevSum(45), B(44) => 
                           prevSum(44), B(43) => prevSum(43), B(42) => 
                           prevSum(42), B(41) => prevSum(41), B(40) => 
                           prevSum(40), B(39) => prevSum(39), B(38) => 
                           prevSum(38), B(37) => prevSum(37), B(36) => 
                           prevSum(36), B(35) => prevSum(35), B(34) => 
                           prevSum(34), B(33) => prevSum(33), B(32) => 
                           prevSum(32), B(31) => prevSum(31), B(30) => 
                           prevSum(30), B(29) => prevSum(29), B(28) => 
                           prevSum(28), B(27) => prevSum(27), B(26) => 
                           prevSum(26), B(25) => prevSum(25), B(24) => 
                           prevSum(24), B(23) => prevSum(23), B(22) => 
                           prevSum(22), B(21) => prevSum(21), B(20) => 
                           prevSum(20), B(19) => prevSum(19), B(18) => 
                           prevSum(18), B(17) => prevSum(17), B(16) => 
                           prevSum(16), B(15) => prevSum(15), B(14) => 
                           prevSum(14), B(13) => prevSum(13), B(12) => 
                           prevSum(12), B(11) => prevSum(11), B(10) => 
                           prevSum(10), B(9) => prevSum(9), B(8) => prevSum(8),
                           B(7) => prevSum(7), B(6) => prevSum(6), B(5) => 
                           prevSum(5), B(4) => prevSum(4), B(3) => prevSum(3), 
                           B(2) => prevSum(2), B(1) => prevSum(1), B(0) => 
                           prevSum(0), Ci => X_Logic0_port, S(63) => 
                           nextSum(63), S(62) => nextSum(62), S(61) => 
                           nextSum(61), S(60) => nextSum(60), S(59) => 
                           nextSum(59), S(58) => nextSum(58), S(57) => 
                           nextSum(57), S(56) => nextSum(56), S(55) => 
                           nextSum(55), S(54) => nextSum(54), S(53) => 
                           nextSum(53), S(52) => nextSum(52), S(51) => 
                           nextSum(51), S(50) => nextSum(50), S(49) => 
                           nextSum(49), S(48) => nextSum(48), S(47) => 
                           nextSum(47), S(46) => nextSum(46), S(45) => 
                           nextSum(45), S(44) => nextSum(44), S(43) => 
                           nextSum(43), S(42) => nextSum(42), S(41) => 
                           nextSum(41), S(40) => nextSum(40), S(39) => 
                           nextSum(39), S(38) => nextSum(38), S(37) => 
                           nextSum(37), S(36) => nextSum(36), S(35) => 
                           nextSum(35), S(34) => nextSum(34), S(33) => 
                           nextSum(33), S(32) => nextSum(32), S(31) => 
                           nextSum(31), S(30) => nextSum(30), S(29) => 
                           nextSum(29), S(28) => nextSum(28), S(27) => 
                           nextSum(27), S(26) => nextSum(26), S(25) => 
                           nextSum(25), S(24) => nextSum(24), S(23) => 
                           nextSum(23), S(22) => nextSum(22), S(21) => 
                           nextSum(21), S(20) => nextSum(20), S(19) => 
                           nextSum(19), S(18) => nextSum(18), S(17) => 
                           nextSum(17), S(16) => nextSum(16), S(15) => 
                           nextSum(15), S(14) => nextSum(14), S(13) => 
                           nextSum(13), S(12) => nextSum(12), S(11) => 
                           nextSum(11), S(10) => nextSum(10), S(9) => 
                           nextSum(9), S(8) => nextSum(8), S(7) => nextSum(7), 
                           S(6) => nextSum(6), S(5) => nextSum(5), S(4) => 
                           nextSum(4), S(3) => nextSum(3), S(2) => nextSum(2), 
                           S(1) => nextSum(1), S(0) => nextSum(0), Co => n_3195
                           );
   U3 : BUF_X1 port map( A => n3, Z => nextA_57_port);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity booth_mul_row_N64_RADIX3_8 is

   port( prevA, prevSum : in std_logic_vector (63 downto 0);  encoderIn : in 
         std_logic_vector (2 downto 0);  nextA, nextSum : out std_logic_vector 
         (63 downto 0));

end booth_mul_row_N64_RADIX3_8;

architecture SYN_struct of booth_mul_row_N64_RADIX3_8 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component RCA_N64_8
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component MUX_GENERIC_N64_RADIX3_8
      port( plusA, minusA, plus2A, minus2A : in std_logic_vector (63 downto 0);
            SEL : in std_logic_vector (2 downto 0);  Y : out std_logic_vector 
            (63 downto 0));
   end component;
   
   component ShiftnCompl_N64_8
      port( plusA : in std_logic_vector (63 downto 0);  plus2A_out, minus2A_out
            , plus4A_out, minus4A_out : out std_logic_vector (63 downto 0));
   end component;
   
   component encoder_N64_RADIX3_8
      port( X : in std_logic_vector (2 downto 0);  Z : out std_logic_vector (2 
            downto 0));
   end component;
   
   signal X_Logic0_port, nextA_63_port, nextA_62_port, nextA_61_port, 
      nextA_60_port, nextA_59_port, nextA_58_port, n3, nextA_56_port, 
      nextA_55_port, nextA_54_port, nextA_53_port, nextA_52_port, nextA_51_port
      , nextA_50_port, nextA_49_port, nextA_48_port, nextA_47_port, 
      nextA_46_port, nextA_45_port, nextA_44_port, nextA_43_port, nextA_42_port
      , nextA_41_port, nextA_40_port, nextA_39_port, nextA_38_port, 
      nextA_37_port, nextA_36_port, nextA_35_port, nextA_34_port, nextA_33_port
      , nextA_32_port, nextA_31_port, nextA_30_port, nextA_29_port, 
      nextA_28_port, nextA_27_port, nextA_26_port, nextA_25_port, nextA_24_port
      , nextA_23_port, nextA_22_port, nextA_21_port, nextA_20_port, 
      nextA_19_port, nextA_18_port, nextA_17_port, nextA_16_port, nextA_15_port
      , nextA_14_port, nextA_13_port, nextA_12_port, nextA_11_port, 
      nextA_10_port, nextA_9_port, nextA_8_port, nextA_7_port, nextA_6_port, 
      nextA_5_port, nextA_4_port, nextA_3_port, nextA_2_port, nextA_1_port, 
      encoder_to_mux_2_port, encoder_to_mux_1_port, encoder_to_mux_0_port, 
      plus2A_s_63_port, plus2A_s_62_port, plus2A_s_61_port, plus2A_s_60_port, 
      plus2A_s_59_port, plus2A_s_58_port, plus2A_s_57_port, plus2A_s_56_port, 
      plus2A_s_55_port, plus2A_s_54_port, plus2A_s_53_port, plus2A_s_52_port, 
      plus2A_s_51_port, plus2A_s_50_port, plus2A_s_49_port, plus2A_s_48_port, 
      plus2A_s_47_port, plus2A_s_46_port, plus2A_s_45_port, plus2A_s_44_port, 
      plus2A_s_43_port, plus2A_s_42_port, plus2A_s_41_port, plus2A_s_40_port, 
      plus2A_s_39_port, plus2A_s_38_port, plus2A_s_37_port, plus2A_s_36_port, 
      plus2A_s_35_port, plus2A_s_34_port, plus2A_s_33_port, plus2A_s_32_port, 
      plus2A_s_31_port, plus2A_s_30_port, plus2A_s_29_port, plus2A_s_28_port, 
      plus2A_s_27_port, plus2A_s_26_port, plus2A_s_25_port, plus2A_s_24_port, 
      plus2A_s_23_port, plus2A_s_22_port, plus2A_s_21_port, plus2A_s_20_port, 
      plus2A_s_19_port, plus2A_s_18_port, plus2A_s_17_port, plus2A_s_16_port, 
      plus2A_s_15_port, plus2A_s_14_port, plus2A_s_13_port, plus2A_s_12_port, 
      plus2A_s_11_port, plus2A_s_10_port, plus2A_s_9_port, plus2A_s_8_port, 
      plus2A_s_7_port, plus2A_s_6_port, plus2A_s_5_port, plus2A_s_4_port, 
      plus2A_s_3_port, plus2A_s_2_port, plus2A_s_1_port, minus2A_s_63_port, 
      minus2A_s_62_port, minus2A_s_61_port, minus2A_s_60_port, 
      minus2A_s_59_port, minus2A_s_58_port, minus2A_s_57_port, 
      minus2A_s_56_port, minus2A_s_55_port, minus2A_s_54_port, 
      minus2A_s_53_port, minus2A_s_52_port, minus2A_s_51_port, 
      minus2A_s_50_port, minus2A_s_49_port, minus2A_s_48_port, 
      minus2A_s_47_port, minus2A_s_46_port, minus2A_s_45_port, 
      minus2A_s_44_port, minus2A_s_43_port, minus2A_s_42_port, 
      minus2A_s_41_port, minus2A_s_40_port, minus2A_s_39_port, 
      minus2A_s_38_port, minus2A_s_37_port, minus2A_s_36_port, 
      minus2A_s_35_port, minus2A_s_34_port, minus2A_s_33_port, 
      minus2A_s_32_port, minus2A_s_31_port, minus2A_s_30_port, 
      minus2A_s_29_port, minus2A_s_28_port, minus2A_s_27_port, 
      minus2A_s_26_port, minus2A_s_25_port, minus2A_s_24_port, 
      minus2A_s_23_port, minus2A_s_22_port, minus2A_s_21_port, 
      minus2A_s_20_port, minus2A_s_19_port, minus2A_s_18_port, 
      minus2A_s_17_port, minus2A_s_16_port, minus2A_s_15_port, 
      minus2A_s_14_port, minus2A_s_13_port, minus2A_s_12_port, 
      minus2A_s_11_port, minus2A_s_10_port, minus2A_s_9_port, minus2A_s_8_port,
      minus2A_s_7_port, minus2A_s_6_port, minus2A_s_5_port, minus2A_s_4_port, 
      minus2A_s_3_port, minus2A_s_2_port, minus2A_s_1_port, minus2A_s_0_port, 
      minus4A_s_63_port, minus4A_s_62_port, minus4A_s_61_port, 
      minus4A_s_60_port, minus4A_s_59_port, minus4A_s_58_port, 
      minus4A_s_57_port, minus4A_s_56_port, minus4A_s_55_port, 
      minus4A_s_54_port, minus4A_s_53_port, minus4A_s_52_port, 
      minus4A_s_51_port, minus4A_s_50_port, minus4A_s_49_port, 
      minus4A_s_48_port, minus4A_s_47_port, minus4A_s_46_port, 
      minus4A_s_45_port, minus4A_s_44_port, minus4A_s_43_port, 
      minus4A_s_42_port, minus4A_s_41_port, minus4A_s_40_port, 
      minus4A_s_39_port, minus4A_s_38_port, minus4A_s_37_port, 
      minus4A_s_36_port, minus4A_s_35_port, minus4A_s_34_port, 
      minus4A_s_33_port, minus4A_s_32_port, minus4A_s_31_port, 
      minus4A_s_30_port, minus4A_s_29_port, minus4A_s_28_port, 
      minus4A_s_27_port, minus4A_s_26_port, minus4A_s_25_port, 
      minus4A_s_24_port, minus4A_s_23_port, minus4A_s_22_port, 
      minus4A_s_21_port, minus4A_s_20_port, minus4A_s_19_port, 
      minus4A_s_18_port, minus4A_s_17_port, minus4A_s_16_port, 
      minus4A_s_15_port, minus4A_s_14_port, minus4A_s_13_port, 
      minus4A_s_12_port, minus4A_s_11_port, minus4A_s_10_port, minus4A_s_9_port
      , minus4A_s_8_port, minus4A_s_7_port, minus4A_s_6_port, minus4A_s_5_port,
      minus4A_s_4_port, minus4A_s_3_port, minus4A_s_2_port, minus4A_s_1_port, 
      minus4A_s_0_port, mux_to_adder_63_port, mux_to_adder_62_port, 
      mux_to_adder_61_port, mux_to_adder_60_port, mux_to_adder_59_port, 
      mux_to_adder_58_port, mux_to_adder_57_port, mux_to_adder_56_port, 
      mux_to_adder_55_port, mux_to_adder_54_port, mux_to_adder_53_port, 
      mux_to_adder_52_port, mux_to_adder_51_port, mux_to_adder_50_port, 
      mux_to_adder_49_port, mux_to_adder_48_port, mux_to_adder_47_port, 
      mux_to_adder_46_port, mux_to_adder_45_port, mux_to_adder_44_port, 
      mux_to_adder_43_port, mux_to_adder_42_port, mux_to_adder_41_port, 
      mux_to_adder_40_port, mux_to_adder_39_port, mux_to_adder_38_port, 
      mux_to_adder_37_port, mux_to_adder_36_port, mux_to_adder_35_port, 
      mux_to_adder_34_port, mux_to_adder_33_port, mux_to_adder_32_port, 
      mux_to_adder_31_port, mux_to_adder_30_port, mux_to_adder_29_port, 
      mux_to_adder_28_port, mux_to_adder_27_port, mux_to_adder_26_port, 
      mux_to_adder_25_port, mux_to_adder_24_port, mux_to_adder_23_port, 
      mux_to_adder_22_port, mux_to_adder_21_port, mux_to_adder_20_port, 
      mux_to_adder_19_port, mux_to_adder_18_port, mux_to_adder_17_port, 
      mux_to_adder_16_port, mux_to_adder_15_port, mux_to_adder_14_port, 
      mux_to_adder_13_port, mux_to_adder_12_port, mux_to_adder_11_port, 
      mux_to_adder_10_port, mux_to_adder_9_port, mux_to_adder_8_port, 
      mux_to_adder_7_port, mux_to_adder_6_port, mux_to_adder_5_port, 
      mux_to_adder_4_port, mux_to_adder_3_port, mux_to_adder_2_port, 
      mux_to_adder_1_port, mux_to_adder_0_port, nextA_0_port, nextA_57_port, 
      n_3196, n_3197, n_3198 : std_logic;

begin
   nextA <= ( nextA_63_port, nextA_62_port, nextA_61_port, nextA_60_port, 
      nextA_59_port, nextA_58_port, nextA_57_port, nextA_56_port, nextA_55_port
      , nextA_54_port, nextA_53_port, nextA_52_port, nextA_51_port, 
      nextA_50_port, nextA_49_port, nextA_48_port, nextA_47_port, nextA_46_port
      , nextA_45_port, nextA_44_port, nextA_43_port, nextA_42_port, 
      nextA_41_port, nextA_40_port, nextA_39_port, nextA_38_port, nextA_37_port
      , nextA_36_port, nextA_35_port, nextA_34_port, nextA_33_port, 
      nextA_32_port, nextA_31_port, nextA_30_port, nextA_29_port, nextA_28_port
      , nextA_27_port, nextA_26_port, nextA_25_port, nextA_24_port, 
      nextA_23_port, nextA_22_port, nextA_21_port, nextA_20_port, nextA_19_port
      , nextA_18_port, nextA_17_port, nextA_16_port, nextA_15_port, 
      nextA_14_port, nextA_13_port, nextA_12_port, nextA_11_port, nextA_10_port
      , nextA_9_port, nextA_8_port, nextA_7_port, nextA_6_port, nextA_5_port, 
      nextA_4_port, nextA_3_port, nextA_2_port, nextA_1_port, nextA_0_port );
   
   X_Logic0_port <= '0';
   nextA_0_port <= '0';
   encoder_1 : encoder_N64_RADIX3_8 port map( X(2) => encoderIn(2), X(1) => 
                           encoderIn(1), X(0) => encoderIn(0), Z(2) => 
                           encoder_to_mux_2_port, Z(1) => encoder_to_mux_1_port
                           , Z(0) => encoder_to_mux_0_port);
   ShiftnCompl_1 : ShiftnCompl_N64_8 port map( plusA(63) => prevA(63), 
                           plusA(62) => prevA(62), plusA(61) => prevA(61), 
                           plusA(60) => prevA(60), plusA(59) => prevA(59), 
                           plusA(58) => prevA(58), plusA(57) => prevA(57), 
                           plusA(56) => prevA(56), plusA(55) => prevA(55), 
                           plusA(54) => prevA(54), plusA(53) => prevA(53), 
                           plusA(52) => prevA(52), plusA(51) => prevA(51), 
                           plusA(50) => prevA(50), plusA(49) => prevA(49), 
                           plusA(48) => prevA(48), plusA(47) => prevA(47), 
                           plusA(46) => prevA(46), plusA(45) => prevA(45), 
                           plusA(44) => prevA(44), plusA(43) => prevA(43), 
                           plusA(42) => prevA(42), plusA(41) => prevA(41), 
                           plusA(40) => prevA(40), plusA(39) => prevA(39), 
                           plusA(38) => prevA(38), plusA(37) => prevA(37), 
                           plusA(36) => prevA(36), plusA(35) => prevA(35), 
                           plusA(34) => prevA(34), plusA(33) => prevA(33), 
                           plusA(32) => prevA(32), plusA(31) => prevA(31), 
                           plusA(30) => prevA(30), plusA(29) => prevA(29), 
                           plusA(28) => prevA(28), plusA(27) => prevA(27), 
                           plusA(26) => prevA(26), plusA(25) => prevA(25), 
                           plusA(24) => prevA(24), plusA(23) => prevA(23), 
                           plusA(22) => prevA(22), plusA(21) => prevA(21), 
                           plusA(20) => prevA(20), plusA(19) => prevA(19), 
                           plusA(18) => prevA(18), plusA(17) => prevA(17), 
                           plusA(16) => prevA(16), plusA(15) => prevA(15), 
                           plusA(14) => prevA(14), plusA(13) => prevA(13), 
                           plusA(12) => prevA(12), plusA(11) => prevA(11), 
                           plusA(10) => prevA(10), plusA(9) => prevA(9), 
                           plusA(8) => prevA(8), plusA(7) => prevA(7), plusA(6)
                           => prevA(6), plusA(5) => prevA(5), plusA(4) => 
                           prevA(4), plusA(3) => prevA(3), plusA(2) => prevA(2)
                           , plusA(1) => prevA(1), plusA(0) => prevA(0), 
                           plus2A_out(63) => plus2A_s_63_port, plus2A_out(62) 
                           => plus2A_s_62_port, plus2A_out(61) => 
                           plus2A_s_61_port, plus2A_out(60) => plus2A_s_60_port
                           , plus2A_out(59) => plus2A_s_59_port, plus2A_out(58)
                           => plus2A_s_58_port, plus2A_out(57) => 
                           plus2A_s_57_port, plus2A_out(56) => plus2A_s_56_port
                           , plus2A_out(55) => plus2A_s_55_port, plus2A_out(54)
                           => plus2A_s_54_port, plus2A_out(53) => 
                           plus2A_s_53_port, plus2A_out(52) => plus2A_s_52_port
                           , plus2A_out(51) => plus2A_s_51_port, plus2A_out(50)
                           => plus2A_s_50_port, plus2A_out(49) => 
                           plus2A_s_49_port, plus2A_out(48) => plus2A_s_48_port
                           , plus2A_out(47) => plus2A_s_47_port, plus2A_out(46)
                           => plus2A_s_46_port, plus2A_out(45) => 
                           plus2A_s_45_port, plus2A_out(44) => plus2A_s_44_port
                           , plus2A_out(43) => plus2A_s_43_port, plus2A_out(42)
                           => plus2A_s_42_port, plus2A_out(41) => 
                           plus2A_s_41_port, plus2A_out(40) => plus2A_s_40_port
                           , plus2A_out(39) => plus2A_s_39_port, plus2A_out(38)
                           => plus2A_s_38_port, plus2A_out(37) => 
                           plus2A_s_37_port, plus2A_out(36) => plus2A_s_36_port
                           , plus2A_out(35) => plus2A_s_35_port, plus2A_out(34)
                           => plus2A_s_34_port, plus2A_out(33) => 
                           plus2A_s_33_port, plus2A_out(32) => plus2A_s_32_port
                           , plus2A_out(31) => plus2A_s_31_port, plus2A_out(30)
                           => plus2A_s_30_port, plus2A_out(29) => 
                           plus2A_s_29_port, plus2A_out(28) => plus2A_s_28_port
                           , plus2A_out(27) => plus2A_s_27_port, plus2A_out(26)
                           => plus2A_s_26_port, plus2A_out(25) => 
                           plus2A_s_25_port, plus2A_out(24) => plus2A_s_24_port
                           , plus2A_out(23) => plus2A_s_23_port, plus2A_out(22)
                           => plus2A_s_22_port, plus2A_out(21) => 
                           plus2A_s_21_port, plus2A_out(20) => plus2A_s_20_port
                           , plus2A_out(19) => plus2A_s_19_port, plus2A_out(18)
                           => plus2A_s_18_port, plus2A_out(17) => 
                           plus2A_s_17_port, plus2A_out(16) => plus2A_s_16_port
                           , plus2A_out(15) => plus2A_s_15_port, plus2A_out(14)
                           => plus2A_s_14_port, plus2A_out(13) => 
                           plus2A_s_13_port, plus2A_out(12) => plus2A_s_12_port
                           , plus2A_out(11) => plus2A_s_11_port, plus2A_out(10)
                           => plus2A_s_10_port, plus2A_out(9) => 
                           plus2A_s_9_port, plus2A_out(8) => plus2A_s_8_port, 
                           plus2A_out(7) => plus2A_s_7_port, plus2A_out(6) => 
                           plus2A_s_6_port, plus2A_out(5) => plus2A_s_5_port, 
                           plus2A_out(4) => plus2A_s_4_port, plus2A_out(3) => 
                           plus2A_s_3_port, plus2A_out(2) => plus2A_s_2_port, 
                           plus2A_out(1) => plus2A_s_1_port, plus2A_out(0) => 
                           n_3196, minus2A_out(63) => minus2A_s_63_port, 
                           minus2A_out(62) => minus2A_s_62_port, 
                           minus2A_out(61) => minus2A_s_61_port, 
                           minus2A_out(60) => minus2A_s_60_port, 
                           minus2A_out(59) => minus2A_s_59_port, 
                           minus2A_out(58) => minus2A_s_58_port, 
                           minus2A_out(57) => minus2A_s_57_port, 
                           minus2A_out(56) => minus2A_s_56_port, 
                           minus2A_out(55) => minus2A_s_55_port, 
                           minus2A_out(54) => minus2A_s_54_port, 
                           minus2A_out(53) => minus2A_s_53_port, 
                           minus2A_out(52) => minus2A_s_52_port, 
                           minus2A_out(51) => minus2A_s_51_port, 
                           minus2A_out(50) => minus2A_s_50_port, 
                           minus2A_out(49) => minus2A_s_49_port, 
                           minus2A_out(48) => minus2A_s_48_port, 
                           minus2A_out(47) => minus2A_s_47_port, 
                           minus2A_out(46) => minus2A_s_46_port, 
                           minus2A_out(45) => minus2A_s_45_port, 
                           minus2A_out(44) => minus2A_s_44_port, 
                           minus2A_out(43) => minus2A_s_43_port, 
                           minus2A_out(42) => minus2A_s_42_port, 
                           minus2A_out(41) => minus2A_s_41_port, 
                           minus2A_out(40) => minus2A_s_40_port, 
                           minus2A_out(39) => minus2A_s_39_port, 
                           minus2A_out(38) => minus2A_s_38_port, 
                           minus2A_out(37) => minus2A_s_37_port, 
                           minus2A_out(36) => minus2A_s_36_port, 
                           minus2A_out(35) => minus2A_s_35_port, 
                           minus2A_out(34) => minus2A_s_34_port, 
                           minus2A_out(33) => minus2A_s_33_port, 
                           minus2A_out(32) => minus2A_s_32_port, 
                           minus2A_out(31) => minus2A_s_31_port, 
                           minus2A_out(30) => minus2A_s_30_port, 
                           minus2A_out(29) => minus2A_s_29_port, 
                           minus2A_out(28) => minus2A_s_28_port, 
                           minus2A_out(27) => minus2A_s_27_port, 
                           minus2A_out(26) => minus2A_s_26_port, 
                           minus2A_out(25) => minus2A_s_25_port, 
                           minus2A_out(24) => minus2A_s_24_port, 
                           minus2A_out(23) => minus2A_s_23_port, 
                           minus2A_out(22) => minus2A_s_22_port, 
                           minus2A_out(21) => minus2A_s_21_port, 
                           minus2A_out(20) => minus2A_s_20_port, 
                           minus2A_out(19) => minus2A_s_19_port, 
                           minus2A_out(18) => minus2A_s_18_port, 
                           minus2A_out(17) => minus2A_s_17_port, 
                           minus2A_out(16) => minus2A_s_16_port, 
                           minus2A_out(15) => minus2A_s_15_port, 
                           minus2A_out(14) => minus2A_s_14_port, 
                           minus2A_out(13) => minus2A_s_13_port, 
                           minus2A_out(12) => minus2A_s_12_port, 
                           minus2A_out(11) => minus2A_s_11_port, 
                           minus2A_out(10) => minus2A_s_10_port, minus2A_out(9)
                           => minus2A_s_9_port, minus2A_out(8) => 
                           minus2A_s_8_port, minus2A_out(7) => minus2A_s_7_port
                           , minus2A_out(6) => minus2A_s_6_port, minus2A_out(5)
                           => minus2A_s_5_port, minus2A_out(4) => 
                           minus2A_s_4_port, minus2A_out(3) => minus2A_s_3_port
                           , minus2A_out(2) => minus2A_s_2_port, minus2A_out(1)
                           => minus2A_s_1_port, minus2A_out(0) => 
                           minus2A_s_0_port, plus4A_out(63) => nextA_63_port, 
                           plus4A_out(62) => nextA_62_port, plus4A_out(61) => 
                           nextA_61_port, plus4A_out(60) => nextA_60_port, 
                           plus4A_out(59) => nextA_59_port, plus4A_out(58) => 
                           nextA_58_port, plus4A_out(57) => n3, plus4A_out(56) 
                           => nextA_56_port, plus4A_out(55) => nextA_55_port, 
                           plus4A_out(54) => nextA_54_port, plus4A_out(53) => 
                           nextA_53_port, plus4A_out(52) => nextA_52_port, 
                           plus4A_out(51) => nextA_51_port, plus4A_out(50) => 
                           nextA_50_port, plus4A_out(49) => nextA_49_port, 
                           plus4A_out(48) => nextA_48_port, plus4A_out(47) => 
                           nextA_47_port, plus4A_out(46) => nextA_46_port, 
                           plus4A_out(45) => nextA_45_port, plus4A_out(44) => 
                           nextA_44_port, plus4A_out(43) => nextA_43_port, 
                           plus4A_out(42) => nextA_42_port, plus4A_out(41) => 
                           nextA_41_port, plus4A_out(40) => nextA_40_port, 
                           plus4A_out(39) => nextA_39_port, plus4A_out(38) => 
                           nextA_38_port, plus4A_out(37) => nextA_37_port, 
                           plus4A_out(36) => nextA_36_port, plus4A_out(35) => 
                           nextA_35_port, plus4A_out(34) => nextA_34_port, 
                           plus4A_out(33) => nextA_33_port, plus4A_out(32) => 
                           nextA_32_port, plus4A_out(31) => nextA_31_port, 
                           plus4A_out(30) => nextA_30_port, plus4A_out(29) => 
                           nextA_29_port, plus4A_out(28) => nextA_28_port, 
                           plus4A_out(27) => nextA_27_port, plus4A_out(26) => 
                           nextA_26_port, plus4A_out(25) => nextA_25_port, 
                           plus4A_out(24) => nextA_24_port, plus4A_out(23) => 
                           nextA_23_port, plus4A_out(22) => nextA_22_port, 
                           plus4A_out(21) => nextA_21_port, plus4A_out(20) => 
                           nextA_20_port, plus4A_out(19) => nextA_19_port, 
                           plus4A_out(18) => nextA_18_port, plus4A_out(17) => 
                           nextA_17_port, plus4A_out(16) => nextA_16_port, 
                           plus4A_out(15) => nextA_15_port, plus4A_out(14) => 
                           nextA_14_port, plus4A_out(13) => nextA_13_port, 
                           plus4A_out(12) => nextA_12_port, plus4A_out(11) => 
                           nextA_11_port, plus4A_out(10) => nextA_10_port, 
                           plus4A_out(9) => nextA_9_port, plus4A_out(8) => 
                           nextA_8_port, plus4A_out(7) => nextA_7_port, 
                           plus4A_out(6) => nextA_6_port, plus4A_out(5) => 
                           nextA_5_port, plus4A_out(4) => nextA_4_port, 
                           plus4A_out(3) => nextA_3_port, plus4A_out(2) => 
                           nextA_2_port, plus4A_out(1) => nextA_1_port, 
                           plus4A_out(0) => n_3197, minus4A_out(63) => 
                           minus4A_s_63_port, minus4A_out(62) => 
                           minus4A_s_62_port, minus4A_out(61) => 
                           minus4A_s_61_port, minus4A_out(60) => 
                           minus4A_s_60_port, minus4A_out(59) => 
                           minus4A_s_59_port, minus4A_out(58) => 
                           minus4A_s_58_port, minus4A_out(57) => 
                           minus4A_s_57_port, minus4A_out(56) => 
                           minus4A_s_56_port, minus4A_out(55) => 
                           minus4A_s_55_port, minus4A_out(54) => 
                           minus4A_s_54_port, minus4A_out(53) => 
                           minus4A_s_53_port, minus4A_out(52) => 
                           minus4A_s_52_port, minus4A_out(51) => 
                           minus4A_s_51_port, minus4A_out(50) => 
                           minus4A_s_50_port, minus4A_out(49) => 
                           minus4A_s_49_port, minus4A_out(48) => 
                           minus4A_s_48_port, minus4A_out(47) => 
                           minus4A_s_47_port, minus4A_out(46) => 
                           minus4A_s_46_port, minus4A_out(45) => 
                           minus4A_s_45_port, minus4A_out(44) => 
                           minus4A_s_44_port, minus4A_out(43) => 
                           minus4A_s_43_port, minus4A_out(42) => 
                           minus4A_s_42_port, minus4A_out(41) => 
                           minus4A_s_41_port, minus4A_out(40) => 
                           minus4A_s_40_port, minus4A_out(39) => 
                           minus4A_s_39_port, minus4A_out(38) => 
                           minus4A_s_38_port, minus4A_out(37) => 
                           minus4A_s_37_port, minus4A_out(36) => 
                           minus4A_s_36_port, minus4A_out(35) => 
                           minus4A_s_35_port, minus4A_out(34) => 
                           minus4A_s_34_port, minus4A_out(33) => 
                           minus4A_s_33_port, minus4A_out(32) => 
                           minus4A_s_32_port, minus4A_out(31) => 
                           minus4A_s_31_port, minus4A_out(30) => 
                           minus4A_s_30_port, minus4A_out(29) => 
                           minus4A_s_29_port, minus4A_out(28) => 
                           minus4A_s_28_port, minus4A_out(27) => 
                           minus4A_s_27_port, minus4A_out(26) => 
                           minus4A_s_26_port, minus4A_out(25) => 
                           minus4A_s_25_port, minus4A_out(24) => 
                           minus4A_s_24_port, minus4A_out(23) => 
                           minus4A_s_23_port, minus4A_out(22) => 
                           minus4A_s_22_port, minus4A_out(21) => 
                           minus4A_s_21_port, minus4A_out(20) => 
                           minus4A_s_20_port, minus4A_out(19) => 
                           minus4A_s_19_port, minus4A_out(18) => 
                           minus4A_s_18_port, minus4A_out(17) => 
                           minus4A_s_17_port, minus4A_out(16) => 
                           minus4A_s_16_port, minus4A_out(15) => 
                           minus4A_s_15_port, minus4A_out(14) => 
                           minus4A_s_14_port, minus4A_out(13) => 
                           minus4A_s_13_port, minus4A_out(12) => 
                           minus4A_s_12_port, minus4A_out(11) => 
                           minus4A_s_11_port, minus4A_out(10) => 
                           minus4A_s_10_port, minus4A_out(9) => 
                           minus4A_s_9_port, minus4A_out(8) => minus4A_s_8_port
                           , minus4A_out(7) => minus4A_s_7_port, minus4A_out(6)
                           => minus4A_s_6_port, minus4A_out(5) => 
                           minus4A_s_5_port, minus4A_out(4) => minus4A_s_4_port
                           , minus4A_out(3) => minus4A_s_3_port, minus4A_out(2)
                           => minus4A_s_2_port, minus4A_out(1) => 
                           minus4A_s_1_port, minus4A_out(0) => minus4A_s_0_port
                           );
   mux_1 : MUX_GENERIC_N64_RADIX3_8 port map( plusA(63) => plus2A_s_63_port, 
                           plusA(62) => plus2A_s_62_port, plusA(61) => 
                           plus2A_s_61_port, plusA(60) => plus2A_s_60_port, 
                           plusA(59) => plus2A_s_59_port, plusA(58) => 
                           plus2A_s_58_port, plusA(57) => plus2A_s_57_port, 
                           plusA(56) => plus2A_s_56_port, plusA(55) => 
                           plus2A_s_55_port, plusA(54) => plus2A_s_54_port, 
                           plusA(53) => plus2A_s_53_port, plusA(52) => 
                           plus2A_s_52_port, plusA(51) => plus2A_s_51_port, 
                           plusA(50) => plus2A_s_50_port, plusA(49) => 
                           plus2A_s_49_port, plusA(48) => plus2A_s_48_port, 
                           plusA(47) => plus2A_s_47_port, plusA(46) => 
                           plus2A_s_46_port, plusA(45) => plus2A_s_45_port, 
                           plusA(44) => plus2A_s_44_port, plusA(43) => 
                           plus2A_s_43_port, plusA(42) => plus2A_s_42_port, 
                           plusA(41) => plus2A_s_41_port, plusA(40) => 
                           plus2A_s_40_port, plusA(39) => plus2A_s_39_port, 
                           plusA(38) => plus2A_s_38_port, plusA(37) => 
                           plus2A_s_37_port, plusA(36) => plus2A_s_36_port, 
                           plusA(35) => plus2A_s_35_port, plusA(34) => 
                           plus2A_s_34_port, plusA(33) => plus2A_s_33_port, 
                           plusA(32) => plus2A_s_32_port, plusA(31) => 
                           plus2A_s_31_port, plusA(30) => plus2A_s_30_port, 
                           plusA(29) => plus2A_s_29_port, plusA(28) => 
                           plus2A_s_28_port, plusA(27) => plus2A_s_27_port, 
                           plusA(26) => plus2A_s_26_port, plusA(25) => 
                           plus2A_s_25_port, plusA(24) => plus2A_s_24_port, 
                           plusA(23) => plus2A_s_23_port, plusA(22) => 
                           plus2A_s_22_port, plusA(21) => plus2A_s_21_port, 
                           plusA(20) => plus2A_s_20_port, plusA(19) => 
                           plus2A_s_19_port, plusA(18) => plus2A_s_18_port, 
                           plusA(17) => plus2A_s_17_port, plusA(16) => 
                           plus2A_s_16_port, plusA(15) => plus2A_s_15_port, 
                           plusA(14) => plus2A_s_14_port, plusA(13) => 
                           plus2A_s_13_port, plusA(12) => plus2A_s_12_port, 
                           plusA(11) => plus2A_s_11_port, plusA(10) => 
                           plus2A_s_10_port, plusA(9) => plus2A_s_9_port, 
                           plusA(8) => plus2A_s_8_port, plusA(7) => 
                           plus2A_s_7_port, plusA(6) => plus2A_s_6_port, 
                           plusA(5) => plus2A_s_5_port, plusA(4) => 
                           plus2A_s_4_port, plusA(3) => plus2A_s_3_port, 
                           plusA(2) => plus2A_s_2_port, plusA(1) => 
                           plus2A_s_1_port, plusA(0) => nextA_0_port, 
                           minusA(63) => minus2A_s_63_port, minusA(62) => 
                           minus2A_s_62_port, minusA(61) => minus2A_s_61_port, 
                           minusA(60) => minus2A_s_60_port, minusA(59) => 
                           minus2A_s_59_port, minusA(58) => minus2A_s_58_port, 
                           minusA(57) => minus2A_s_57_port, minusA(56) => 
                           minus2A_s_56_port, minusA(55) => minus2A_s_55_port, 
                           minusA(54) => minus2A_s_54_port, minusA(53) => 
                           minus2A_s_53_port, minusA(52) => minus2A_s_52_port, 
                           minusA(51) => minus2A_s_51_port, minusA(50) => 
                           minus2A_s_50_port, minusA(49) => minus2A_s_49_port, 
                           minusA(48) => minus2A_s_48_port, minusA(47) => 
                           minus2A_s_47_port, minusA(46) => minus2A_s_46_port, 
                           minusA(45) => minus2A_s_45_port, minusA(44) => 
                           minus2A_s_44_port, minusA(43) => minus2A_s_43_port, 
                           minusA(42) => minus2A_s_42_port, minusA(41) => 
                           minus2A_s_41_port, minusA(40) => minus2A_s_40_port, 
                           minusA(39) => minus2A_s_39_port, minusA(38) => 
                           minus2A_s_38_port, minusA(37) => minus2A_s_37_port, 
                           minusA(36) => minus2A_s_36_port, minusA(35) => 
                           minus2A_s_35_port, minusA(34) => minus2A_s_34_port, 
                           minusA(33) => minus2A_s_33_port, minusA(32) => 
                           minus2A_s_32_port, minusA(31) => minus2A_s_31_port, 
                           minusA(30) => minus2A_s_30_port, minusA(29) => 
                           minus2A_s_29_port, minusA(28) => minus2A_s_28_port, 
                           minusA(27) => minus2A_s_27_port, minusA(26) => 
                           minus2A_s_26_port, minusA(25) => minus2A_s_25_port, 
                           minusA(24) => minus2A_s_24_port, minusA(23) => 
                           minus2A_s_23_port, minusA(22) => minus2A_s_22_port, 
                           minusA(21) => minus2A_s_21_port, minusA(20) => 
                           minus2A_s_20_port, minusA(19) => minus2A_s_19_port, 
                           minusA(18) => minus2A_s_18_port, minusA(17) => 
                           minus2A_s_17_port, minusA(16) => minus2A_s_16_port, 
                           minusA(15) => minus2A_s_15_port, minusA(14) => 
                           minus2A_s_14_port, minusA(13) => minus2A_s_13_port, 
                           minusA(12) => minus2A_s_12_port, minusA(11) => 
                           minus2A_s_11_port, minusA(10) => minus2A_s_10_port, 
                           minusA(9) => minus2A_s_9_port, minusA(8) => 
                           minus2A_s_8_port, minusA(7) => minus2A_s_7_port, 
                           minusA(6) => minus2A_s_6_port, minusA(5) => 
                           minus2A_s_5_port, minusA(4) => minus2A_s_4_port, 
                           minusA(3) => minus2A_s_3_port, minusA(2) => 
                           minus2A_s_2_port, minusA(1) => minus2A_s_1_port, 
                           minusA(0) => minus2A_s_0_port, plus2A(63) => 
                           nextA_63_port, plus2A(62) => nextA_62_port, 
                           plus2A(61) => nextA_61_port, plus2A(60) => 
                           nextA_60_port, plus2A(59) => nextA_59_port, 
                           plus2A(58) => nextA_58_port, plus2A(57) => 
                           nextA_57_port, plus2A(56) => nextA_56_port, 
                           plus2A(55) => nextA_55_port, plus2A(54) => 
                           nextA_54_port, plus2A(53) => nextA_53_port, 
                           plus2A(52) => nextA_52_port, plus2A(51) => 
                           nextA_51_port, plus2A(50) => nextA_50_port, 
                           plus2A(49) => nextA_49_port, plus2A(48) => 
                           nextA_48_port, plus2A(47) => nextA_47_port, 
                           plus2A(46) => nextA_46_port, plus2A(45) => 
                           nextA_45_port, plus2A(44) => nextA_44_port, 
                           plus2A(43) => nextA_43_port, plus2A(42) => 
                           nextA_42_port, plus2A(41) => nextA_41_port, 
                           plus2A(40) => nextA_40_port, plus2A(39) => 
                           nextA_39_port, plus2A(38) => nextA_38_port, 
                           plus2A(37) => nextA_37_port, plus2A(36) => 
                           nextA_36_port, plus2A(35) => nextA_35_port, 
                           plus2A(34) => nextA_34_port, plus2A(33) => 
                           nextA_33_port, plus2A(32) => nextA_32_port, 
                           plus2A(31) => nextA_31_port, plus2A(30) => 
                           nextA_30_port, plus2A(29) => nextA_29_port, 
                           plus2A(28) => nextA_28_port, plus2A(27) => 
                           nextA_27_port, plus2A(26) => nextA_26_port, 
                           plus2A(25) => nextA_25_port, plus2A(24) => 
                           nextA_24_port, plus2A(23) => nextA_23_port, 
                           plus2A(22) => nextA_22_port, plus2A(21) => 
                           nextA_21_port, plus2A(20) => nextA_20_port, 
                           plus2A(19) => nextA_19_port, plus2A(18) => 
                           nextA_18_port, plus2A(17) => nextA_17_port, 
                           plus2A(16) => nextA_16_port, plus2A(15) => 
                           nextA_15_port, plus2A(14) => nextA_14_port, 
                           plus2A(13) => nextA_13_port, plus2A(12) => 
                           nextA_12_port, plus2A(11) => nextA_11_port, 
                           plus2A(10) => nextA_10_port, plus2A(9) => 
                           nextA_9_port, plus2A(8) => nextA_8_port, plus2A(7) 
                           => nextA_7_port, plus2A(6) => nextA_6_port, 
                           plus2A(5) => nextA_5_port, plus2A(4) => nextA_4_port
                           , plus2A(3) => nextA_3_port, plus2A(2) => 
                           nextA_2_port, plus2A(1) => nextA_1_port, plus2A(0) 
                           => nextA_0_port, minus2A(63) => minus4A_s_63_port, 
                           minus2A(62) => minus4A_s_62_port, minus2A(61) => 
                           minus4A_s_61_port, minus2A(60) => minus4A_s_60_port,
                           minus2A(59) => minus4A_s_59_port, minus2A(58) => 
                           minus4A_s_58_port, minus2A(57) => minus4A_s_57_port,
                           minus2A(56) => minus4A_s_56_port, minus2A(55) => 
                           minus4A_s_55_port, minus2A(54) => minus4A_s_54_port,
                           minus2A(53) => minus4A_s_53_port, minus2A(52) => 
                           minus4A_s_52_port, minus2A(51) => minus4A_s_51_port,
                           minus2A(50) => minus4A_s_50_port, minus2A(49) => 
                           minus4A_s_49_port, minus2A(48) => minus4A_s_48_port,
                           minus2A(47) => minus4A_s_47_port, minus2A(46) => 
                           minus4A_s_46_port, minus2A(45) => minus4A_s_45_port,
                           minus2A(44) => minus4A_s_44_port, minus2A(43) => 
                           minus4A_s_43_port, minus2A(42) => minus4A_s_42_port,
                           minus2A(41) => minus4A_s_41_port, minus2A(40) => 
                           minus4A_s_40_port, minus2A(39) => minus4A_s_39_port,
                           minus2A(38) => minus4A_s_38_port, minus2A(37) => 
                           minus4A_s_37_port, minus2A(36) => minus4A_s_36_port,
                           minus2A(35) => minus4A_s_35_port, minus2A(34) => 
                           minus4A_s_34_port, minus2A(33) => minus4A_s_33_port,
                           minus2A(32) => minus4A_s_32_port, minus2A(31) => 
                           minus4A_s_31_port, minus2A(30) => minus4A_s_30_port,
                           minus2A(29) => minus4A_s_29_port, minus2A(28) => 
                           minus4A_s_28_port, minus2A(27) => minus4A_s_27_port,
                           minus2A(26) => minus4A_s_26_port, minus2A(25) => 
                           minus4A_s_25_port, minus2A(24) => minus4A_s_24_port,
                           minus2A(23) => minus4A_s_23_port, minus2A(22) => 
                           minus4A_s_22_port, minus2A(21) => minus4A_s_21_port,
                           minus2A(20) => minus4A_s_20_port, minus2A(19) => 
                           minus4A_s_19_port, minus2A(18) => minus4A_s_18_port,
                           minus2A(17) => minus4A_s_17_port, minus2A(16) => 
                           minus4A_s_16_port, minus2A(15) => minus4A_s_15_port,
                           minus2A(14) => minus4A_s_14_port, minus2A(13) => 
                           minus4A_s_13_port, minus2A(12) => minus4A_s_12_port,
                           minus2A(11) => minus4A_s_11_port, minus2A(10) => 
                           minus4A_s_10_port, minus2A(9) => minus4A_s_9_port, 
                           minus2A(8) => minus4A_s_8_port, minus2A(7) => 
                           minus4A_s_7_port, minus2A(6) => minus4A_s_6_port, 
                           minus2A(5) => minus4A_s_5_port, minus2A(4) => 
                           minus4A_s_4_port, minus2A(3) => minus4A_s_3_port, 
                           minus2A(2) => minus4A_s_2_port, minus2A(1) => 
                           minus4A_s_1_port, minus2A(0) => minus4A_s_0_port, 
                           SEL(2) => encoder_to_mux_2_port, SEL(1) => 
                           encoder_to_mux_1_port, SEL(0) => 
                           encoder_to_mux_0_port, Y(63) => mux_to_adder_63_port
                           , Y(62) => mux_to_adder_62_port, Y(61) => 
                           mux_to_adder_61_port, Y(60) => mux_to_adder_60_port,
                           Y(59) => mux_to_adder_59_port, Y(58) => 
                           mux_to_adder_58_port, Y(57) => mux_to_adder_57_port,
                           Y(56) => mux_to_adder_56_port, Y(55) => 
                           mux_to_adder_55_port, Y(54) => mux_to_adder_54_port,
                           Y(53) => mux_to_adder_53_port, Y(52) => 
                           mux_to_adder_52_port, Y(51) => mux_to_adder_51_port,
                           Y(50) => mux_to_adder_50_port, Y(49) => 
                           mux_to_adder_49_port, Y(48) => mux_to_adder_48_port,
                           Y(47) => mux_to_adder_47_port, Y(46) => 
                           mux_to_adder_46_port, Y(45) => mux_to_adder_45_port,
                           Y(44) => mux_to_adder_44_port, Y(43) => 
                           mux_to_adder_43_port, Y(42) => mux_to_adder_42_port,
                           Y(41) => mux_to_adder_41_port, Y(40) => 
                           mux_to_adder_40_port, Y(39) => mux_to_adder_39_port,
                           Y(38) => mux_to_adder_38_port, Y(37) => 
                           mux_to_adder_37_port, Y(36) => mux_to_adder_36_port,
                           Y(35) => mux_to_adder_35_port, Y(34) => 
                           mux_to_adder_34_port, Y(33) => mux_to_adder_33_port,
                           Y(32) => mux_to_adder_32_port, Y(31) => 
                           mux_to_adder_31_port, Y(30) => mux_to_adder_30_port,
                           Y(29) => mux_to_adder_29_port, Y(28) => 
                           mux_to_adder_28_port, Y(27) => mux_to_adder_27_port,
                           Y(26) => mux_to_adder_26_port, Y(25) => 
                           mux_to_adder_25_port, Y(24) => mux_to_adder_24_port,
                           Y(23) => mux_to_adder_23_port, Y(22) => 
                           mux_to_adder_22_port, Y(21) => mux_to_adder_21_port,
                           Y(20) => mux_to_adder_20_port, Y(19) => 
                           mux_to_adder_19_port, Y(18) => mux_to_adder_18_port,
                           Y(17) => mux_to_adder_17_port, Y(16) => 
                           mux_to_adder_16_port, Y(15) => mux_to_adder_15_port,
                           Y(14) => mux_to_adder_14_port, Y(13) => 
                           mux_to_adder_13_port, Y(12) => mux_to_adder_12_port,
                           Y(11) => mux_to_adder_11_port, Y(10) => 
                           mux_to_adder_10_port, Y(9) => mux_to_adder_9_port, 
                           Y(8) => mux_to_adder_8_port, Y(7) => 
                           mux_to_adder_7_port, Y(6) => mux_to_adder_6_port, 
                           Y(5) => mux_to_adder_5_port, Y(4) => 
                           mux_to_adder_4_port, Y(3) => mux_to_adder_3_port, 
                           Y(2) => mux_to_adder_2_port, Y(1) => 
                           mux_to_adder_1_port, Y(0) => mux_to_adder_0_port);
   rca_1 : RCA_N64_8 port map( A(63) => mux_to_adder_63_port, A(62) => 
                           mux_to_adder_62_port, A(61) => mux_to_adder_61_port,
                           A(60) => mux_to_adder_60_port, A(59) => 
                           mux_to_adder_59_port, A(58) => mux_to_adder_58_port,
                           A(57) => mux_to_adder_57_port, A(56) => 
                           mux_to_adder_56_port, A(55) => mux_to_adder_55_port,
                           A(54) => mux_to_adder_54_port, A(53) => 
                           mux_to_adder_53_port, A(52) => mux_to_adder_52_port,
                           A(51) => mux_to_adder_51_port, A(50) => 
                           mux_to_adder_50_port, A(49) => mux_to_adder_49_port,
                           A(48) => mux_to_adder_48_port, A(47) => 
                           mux_to_adder_47_port, A(46) => mux_to_adder_46_port,
                           A(45) => mux_to_adder_45_port, A(44) => 
                           mux_to_adder_44_port, A(43) => mux_to_adder_43_port,
                           A(42) => mux_to_adder_42_port, A(41) => 
                           mux_to_adder_41_port, A(40) => mux_to_adder_40_port,
                           A(39) => mux_to_adder_39_port, A(38) => 
                           mux_to_adder_38_port, A(37) => mux_to_adder_37_port,
                           A(36) => mux_to_adder_36_port, A(35) => 
                           mux_to_adder_35_port, A(34) => mux_to_adder_34_port,
                           A(33) => mux_to_adder_33_port, A(32) => 
                           mux_to_adder_32_port, A(31) => mux_to_adder_31_port,
                           A(30) => mux_to_adder_30_port, A(29) => 
                           mux_to_adder_29_port, A(28) => mux_to_adder_28_port,
                           A(27) => mux_to_adder_27_port, A(26) => 
                           mux_to_adder_26_port, A(25) => mux_to_adder_25_port,
                           A(24) => mux_to_adder_24_port, A(23) => 
                           mux_to_adder_23_port, A(22) => mux_to_adder_22_port,
                           A(21) => mux_to_adder_21_port, A(20) => 
                           mux_to_adder_20_port, A(19) => mux_to_adder_19_port,
                           A(18) => mux_to_adder_18_port, A(17) => 
                           mux_to_adder_17_port, A(16) => mux_to_adder_16_port,
                           A(15) => mux_to_adder_15_port, A(14) => 
                           mux_to_adder_14_port, A(13) => mux_to_adder_13_port,
                           A(12) => mux_to_adder_12_port, A(11) => 
                           mux_to_adder_11_port, A(10) => mux_to_adder_10_port,
                           A(9) => mux_to_adder_9_port, A(8) => 
                           mux_to_adder_8_port, A(7) => mux_to_adder_7_port, 
                           A(6) => mux_to_adder_6_port, A(5) => 
                           mux_to_adder_5_port, A(4) => mux_to_adder_4_port, 
                           A(3) => mux_to_adder_3_port, A(2) => 
                           mux_to_adder_2_port, A(1) => mux_to_adder_1_port, 
                           A(0) => mux_to_adder_0_port, B(63) => prevSum(63), 
                           B(62) => prevSum(62), B(61) => prevSum(61), B(60) =>
                           prevSum(60), B(59) => prevSum(59), B(58) => 
                           prevSum(58), B(57) => prevSum(57), B(56) => 
                           prevSum(56), B(55) => prevSum(55), B(54) => 
                           prevSum(54), B(53) => prevSum(53), B(52) => 
                           prevSum(52), B(51) => prevSum(51), B(50) => 
                           prevSum(50), B(49) => prevSum(49), B(48) => 
                           prevSum(48), B(47) => prevSum(47), B(46) => 
                           prevSum(46), B(45) => prevSum(45), B(44) => 
                           prevSum(44), B(43) => prevSum(43), B(42) => 
                           prevSum(42), B(41) => prevSum(41), B(40) => 
                           prevSum(40), B(39) => prevSum(39), B(38) => 
                           prevSum(38), B(37) => prevSum(37), B(36) => 
                           prevSum(36), B(35) => prevSum(35), B(34) => 
                           prevSum(34), B(33) => prevSum(33), B(32) => 
                           prevSum(32), B(31) => prevSum(31), B(30) => 
                           prevSum(30), B(29) => prevSum(29), B(28) => 
                           prevSum(28), B(27) => prevSum(27), B(26) => 
                           prevSum(26), B(25) => prevSum(25), B(24) => 
                           prevSum(24), B(23) => prevSum(23), B(22) => 
                           prevSum(22), B(21) => prevSum(21), B(20) => 
                           prevSum(20), B(19) => prevSum(19), B(18) => 
                           prevSum(18), B(17) => prevSum(17), B(16) => 
                           prevSum(16), B(15) => prevSum(15), B(14) => 
                           prevSum(14), B(13) => prevSum(13), B(12) => 
                           prevSum(12), B(11) => prevSum(11), B(10) => 
                           prevSum(10), B(9) => prevSum(9), B(8) => prevSum(8),
                           B(7) => prevSum(7), B(6) => prevSum(6), B(5) => 
                           prevSum(5), B(4) => prevSum(4), B(3) => prevSum(3), 
                           B(2) => prevSum(2), B(1) => prevSum(1), B(0) => 
                           prevSum(0), Ci => X_Logic0_port, S(63) => 
                           nextSum(63), S(62) => nextSum(62), S(61) => 
                           nextSum(61), S(60) => nextSum(60), S(59) => 
                           nextSum(59), S(58) => nextSum(58), S(57) => 
                           nextSum(57), S(56) => nextSum(56), S(55) => 
                           nextSum(55), S(54) => nextSum(54), S(53) => 
                           nextSum(53), S(52) => nextSum(52), S(51) => 
                           nextSum(51), S(50) => nextSum(50), S(49) => 
                           nextSum(49), S(48) => nextSum(48), S(47) => 
                           nextSum(47), S(46) => nextSum(46), S(45) => 
                           nextSum(45), S(44) => nextSum(44), S(43) => 
                           nextSum(43), S(42) => nextSum(42), S(41) => 
                           nextSum(41), S(40) => nextSum(40), S(39) => 
                           nextSum(39), S(38) => nextSum(38), S(37) => 
                           nextSum(37), S(36) => nextSum(36), S(35) => 
                           nextSum(35), S(34) => nextSum(34), S(33) => 
                           nextSum(33), S(32) => nextSum(32), S(31) => 
                           nextSum(31), S(30) => nextSum(30), S(29) => 
                           nextSum(29), S(28) => nextSum(28), S(27) => 
                           nextSum(27), S(26) => nextSum(26), S(25) => 
                           nextSum(25), S(24) => nextSum(24), S(23) => 
                           nextSum(23), S(22) => nextSum(22), S(21) => 
                           nextSum(21), S(20) => nextSum(20), S(19) => 
                           nextSum(19), S(18) => nextSum(18), S(17) => 
                           nextSum(17), S(16) => nextSum(16), S(15) => 
                           nextSum(15), S(14) => nextSum(14), S(13) => 
                           nextSum(13), S(12) => nextSum(12), S(11) => 
                           nextSum(11), S(10) => nextSum(10), S(9) => 
                           nextSum(9), S(8) => nextSum(8), S(7) => nextSum(7), 
                           S(6) => nextSum(6), S(5) => nextSum(5), S(4) => 
                           nextSum(4), S(3) => nextSum(3), S(2) => nextSum(2), 
                           S(1) => nextSum(1), S(0) => nextSum(0), Co => n_3198
                           );
   U3 : BUF_X1 port map( A => n3, Z => nextA_57_port);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity booth_mul_row_N64_RADIX3_9 is

   port( prevA, prevSum : in std_logic_vector (63 downto 0);  encoderIn : in 
         std_logic_vector (2 downto 0);  nextA, nextSum : out std_logic_vector 
         (63 downto 0));

end booth_mul_row_N64_RADIX3_9;

architecture SYN_struct of booth_mul_row_N64_RADIX3_9 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component RCA_N64_9
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component MUX_GENERIC_N64_RADIX3_9
      port( plusA, minusA, plus2A, minus2A : in std_logic_vector (63 downto 0);
            SEL : in std_logic_vector (2 downto 0);  Y : out std_logic_vector 
            (63 downto 0));
   end component;
   
   component ShiftnCompl_N64_9
      port( plusA : in std_logic_vector (63 downto 0);  plus2A_out, minus2A_out
            , plus4A_out, minus4A_out : out std_logic_vector (63 downto 0));
   end component;
   
   component encoder_N64_RADIX3_9
      port( X : in std_logic_vector (2 downto 0);  Z : out std_logic_vector (2 
            downto 0));
   end component;
   
   signal X_Logic0_port, nextA_63_port, nextA_62_port, nextA_61_port, 
      nextA_60_port, nextA_59_port, nextA_58_port, n3, nextA_56_port, 
      nextA_55_port, nextA_54_port, nextA_53_port, nextA_52_port, nextA_51_port
      , nextA_50_port, nextA_49_port, nextA_48_port, nextA_47_port, 
      nextA_46_port, nextA_45_port, nextA_44_port, nextA_43_port, nextA_42_port
      , nextA_41_port, nextA_40_port, nextA_39_port, nextA_38_port, 
      nextA_37_port, nextA_36_port, nextA_35_port, nextA_34_port, nextA_33_port
      , nextA_32_port, nextA_31_port, nextA_30_port, nextA_29_port, 
      nextA_28_port, nextA_27_port, nextA_26_port, nextA_25_port, nextA_24_port
      , nextA_23_port, nextA_22_port, nextA_21_port, nextA_20_port, 
      nextA_19_port, nextA_18_port, nextA_17_port, nextA_16_port, nextA_15_port
      , nextA_14_port, nextA_13_port, nextA_12_port, nextA_11_port, 
      nextA_10_port, nextA_9_port, nextA_8_port, nextA_7_port, nextA_6_port, 
      nextA_5_port, nextA_4_port, nextA_3_port, nextA_2_port, nextA_1_port, 
      encoder_to_mux_2_port, encoder_to_mux_1_port, encoder_to_mux_0_port, 
      plus2A_s_63_port, plus2A_s_62_port, plus2A_s_61_port, plus2A_s_60_port, 
      plus2A_s_59_port, plus2A_s_58_port, plus2A_s_57_port, plus2A_s_56_port, 
      plus2A_s_55_port, plus2A_s_54_port, plus2A_s_53_port, plus2A_s_52_port, 
      plus2A_s_51_port, plus2A_s_50_port, plus2A_s_49_port, plus2A_s_48_port, 
      plus2A_s_47_port, plus2A_s_46_port, plus2A_s_45_port, plus2A_s_44_port, 
      plus2A_s_43_port, plus2A_s_42_port, plus2A_s_41_port, plus2A_s_40_port, 
      plus2A_s_39_port, plus2A_s_38_port, plus2A_s_37_port, plus2A_s_36_port, 
      plus2A_s_35_port, plus2A_s_34_port, plus2A_s_33_port, plus2A_s_32_port, 
      plus2A_s_31_port, plus2A_s_30_port, plus2A_s_29_port, plus2A_s_28_port, 
      plus2A_s_27_port, plus2A_s_26_port, plus2A_s_25_port, plus2A_s_24_port, 
      plus2A_s_23_port, plus2A_s_22_port, plus2A_s_21_port, plus2A_s_20_port, 
      plus2A_s_19_port, plus2A_s_18_port, plus2A_s_17_port, plus2A_s_16_port, 
      plus2A_s_15_port, plus2A_s_14_port, plus2A_s_13_port, plus2A_s_12_port, 
      plus2A_s_11_port, plus2A_s_10_port, plus2A_s_9_port, plus2A_s_8_port, 
      plus2A_s_7_port, plus2A_s_6_port, plus2A_s_5_port, plus2A_s_4_port, 
      plus2A_s_3_port, plus2A_s_2_port, plus2A_s_1_port, minus2A_s_63_port, 
      minus2A_s_62_port, minus2A_s_61_port, minus2A_s_60_port, 
      minus2A_s_59_port, minus2A_s_58_port, minus2A_s_57_port, 
      minus2A_s_56_port, minus2A_s_55_port, minus2A_s_54_port, 
      minus2A_s_53_port, minus2A_s_52_port, minus2A_s_51_port, 
      minus2A_s_50_port, minus2A_s_49_port, minus2A_s_48_port, 
      minus2A_s_47_port, minus2A_s_46_port, minus2A_s_45_port, 
      minus2A_s_44_port, minus2A_s_43_port, minus2A_s_42_port, 
      minus2A_s_41_port, minus2A_s_40_port, minus2A_s_39_port, 
      minus2A_s_38_port, minus2A_s_37_port, minus2A_s_36_port, 
      minus2A_s_35_port, minus2A_s_34_port, minus2A_s_33_port, 
      minus2A_s_32_port, minus2A_s_31_port, minus2A_s_30_port, 
      minus2A_s_29_port, minus2A_s_28_port, minus2A_s_27_port, 
      minus2A_s_26_port, minus2A_s_25_port, minus2A_s_24_port, 
      minus2A_s_23_port, minus2A_s_22_port, minus2A_s_21_port, 
      minus2A_s_20_port, minus2A_s_19_port, minus2A_s_18_port, 
      minus2A_s_17_port, minus2A_s_16_port, minus2A_s_15_port, 
      minus2A_s_14_port, minus2A_s_13_port, minus2A_s_12_port, 
      minus2A_s_11_port, minus2A_s_10_port, minus2A_s_9_port, minus2A_s_8_port,
      minus2A_s_7_port, minus2A_s_6_port, minus2A_s_5_port, minus2A_s_4_port, 
      minus2A_s_3_port, minus2A_s_2_port, minus2A_s_1_port, minus2A_s_0_port, 
      minus4A_s_63_port, minus4A_s_62_port, minus4A_s_61_port, 
      minus4A_s_60_port, minus4A_s_59_port, minus4A_s_58_port, 
      minus4A_s_57_port, minus4A_s_56_port, minus4A_s_55_port, 
      minus4A_s_54_port, minus4A_s_53_port, minus4A_s_52_port, 
      minus4A_s_51_port, minus4A_s_50_port, minus4A_s_49_port, 
      minus4A_s_48_port, minus4A_s_47_port, minus4A_s_46_port, 
      minus4A_s_45_port, minus4A_s_44_port, minus4A_s_43_port, 
      minus4A_s_42_port, minus4A_s_41_port, minus4A_s_40_port, 
      minus4A_s_39_port, minus4A_s_38_port, minus4A_s_37_port, 
      minus4A_s_36_port, minus4A_s_35_port, minus4A_s_34_port, 
      minus4A_s_33_port, minus4A_s_32_port, minus4A_s_31_port, 
      minus4A_s_30_port, minus4A_s_29_port, minus4A_s_28_port, 
      minus4A_s_27_port, minus4A_s_26_port, minus4A_s_25_port, 
      minus4A_s_24_port, minus4A_s_23_port, minus4A_s_22_port, 
      minus4A_s_21_port, minus4A_s_20_port, minus4A_s_19_port, 
      minus4A_s_18_port, minus4A_s_17_port, minus4A_s_16_port, 
      minus4A_s_15_port, minus4A_s_14_port, minus4A_s_13_port, 
      minus4A_s_12_port, minus4A_s_11_port, minus4A_s_10_port, minus4A_s_9_port
      , minus4A_s_8_port, minus4A_s_7_port, minus4A_s_6_port, minus4A_s_5_port,
      minus4A_s_4_port, minus4A_s_3_port, minus4A_s_2_port, minus4A_s_1_port, 
      minus4A_s_0_port, mux_to_adder_63_port, mux_to_adder_62_port, 
      mux_to_adder_61_port, mux_to_adder_60_port, mux_to_adder_59_port, 
      mux_to_adder_58_port, mux_to_adder_57_port, mux_to_adder_56_port, 
      mux_to_adder_55_port, mux_to_adder_54_port, mux_to_adder_53_port, 
      mux_to_adder_52_port, mux_to_adder_51_port, mux_to_adder_50_port, 
      mux_to_adder_49_port, mux_to_adder_48_port, mux_to_adder_47_port, 
      mux_to_adder_46_port, mux_to_adder_45_port, mux_to_adder_44_port, 
      mux_to_adder_43_port, mux_to_adder_42_port, mux_to_adder_41_port, 
      mux_to_adder_40_port, mux_to_adder_39_port, mux_to_adder_38_port, 
      mux_to_adder_37_port, mux_to_adder_36_port, mux_to_adder_35_port, 
      mux_to_adder_34_port, mux_to_adder_33_port, mux_to_adder_32_port, 
      mux_to_adder_31_port, mux_to_adder_30_port, mux_to_adder_29_port, 
      mux_to_adder_28_port, mux_to_adder_27_port, mux_to_adder_26_port, 
      mux_to_adder_25_port, mux_to_adder_24_port, mux_to_adder_23_port, 
      mux_to_adder_22_port, mux_to_adder_21_port, mux_to_adder_20_port, 
      mux_to_adder_19_port, mux_to_adder_18_port, mux_to_adder_17_port, 
      mux_to_adder_16_port, mux_to_adder_15_port, mux_to_adder_14_port, 
      mux_to_adder_13_port, mux_to_adder_12_port, mux_to_adder_11_port, 
      mux_to_adder_10_port, mux_to_adder_9_port, mux_to_adder_8_port, 
      mux_to_adder_7_port, mux_to_adder_6_port, mux_to_adder_5_port, 
      mux_to_adder_4_port, mux_to_adder_3_port, mux_to_adder_2_port, 
      mux_to_adder_1_port, mux_to_adder_0_port, nextA_0_port, nextA_57_port, 
      n_3199, n_3200, n_3201 : std_logic;

begin
   nextA <= ( nextA_63_port, nextA_62_port, nextA_61_port, nextA_60_port, 
      nextA_59_port, nextA_58_port, nextA_57_port, nextA_56_port, nextA_55_port
      , nextA_54_port, nextA_53_port, nextA_52_port, nextA_51_port, 
      nextA_50_port, nextA_49_port, nextA_48_port, nextA_47_port, nextA_46_port
      , nextA_45_port, nextA_44_port, nextA_43_port, nextA_42_port, 
      nextA_41_port, nextA_40_port, nextA_39_port, nextA_38_port, nextA_37_port
      , nextA_36_port, nextA_35_port, nextA_34_port, nextA_33_port, 
      nextA_32_port, nextA_31_port, nextA_30_port, nextA_29_port, nextA_28_port
      , nextA_27_port, nextA_26_port, nextA_25_port, nextA_24_port, 
      nextA_23_port, nextA_22_port, nextA_21_port, nextA_20_port, nextA_19_port
      , nextA_18_port, nextA_17_port, nextA_16_port, nextA_15_port, 
      nextA_14_port, nextA_13_port, nextA_12_port, nextA_11_port, nextA_10_port
      , nextA_9_port, nextA_8_port, nextA_7_port, nextA_6_port, nextA_5_port, 
      nextA_4_port, nextA_3_port, nextA_2_port, nextA_1_port, nextA_0_port );
   
   X_Logic0_port <= '0';
   nextA_0_port <= '0';
   encoder_1 : encoder_N64_RADIX3_9 port map( X(2) => encoderIn(2), X(1) => 
                           encoderIn(1), X(0) => encoderIn(0), Z(2) => 
                           encoder_to_mux_2_port, Z(1) => encoder_to_mux_1_port
                           , Z(0) => encoder_to_mux_0_port);
   ShiftnCompl_1 : ShiftnCompl_N64_9 port map( plusA(63) => prevA(63), 
                           plusA(62) => prevA(62), plusA(61) => prevA(61), 
                           plusA(60) => prevA(60), plusA(59) => prevA(59), 
                           plusA(58) => prevA(58), plusA(57) => prevA(57), 
                           plusA(56) => prevA(56), plusA(55) => prevA(55), 
                           plusA(54) => prevA(54), plusA(53) => prevA(53), 
                           plusA(52) => prevA(52), plusA(51) => prevA(51), 
                           plusA(50) => prevA(50), plusA(49) => prevA(49), 
                           plusA(48) => prevA(48), plusA(47) => prevA(47), 
                           plusA(46) => prevA(46), plusA(45) => prevA(45), 
                           plusA(44) => prevA(44), plusA(43) => prevA(43), 
                           plusA(42) => prevA(42), plusA(41) => prevA(41), 
                           plusA(40) => prevA(40), plusA(39) => prevA(39), 
                           plusA(38) => prevA(38), plusA(37) => prevA(37), 
                           plusA(36) => prevA(36), plusA(35) => prevA(35), 
                           plusA(34) => prevA(34), plusA(33) => prevA(33), 
                           plusA(32) => prevA(32), plusA(31) => prevA(31), 
                           plusA(30) => prevA(30), plusA(29) => prevA(29), 
                           plusA(28) => prevA(28), plusA(27) => prevA(27), 
                           plusA(26) => prevA(26), plusA(25) => prevA(25), 
                           plusA(24) => prevA(24), plusA(23) => prevA(23), 
                           plusA(22) => prevA(22), plusA(21) => prevA(21), 
                           plusA(20) => prevA(20), plusA(19) => prevA(19), 
                           plusA(18) => prevA(18), plusA(17) => prevA(17), 
                           plusA(16) => prevA(16), plusA(15) => prevA(15), 
                           plusA(14) => prevA(14), plusA(13) => prevA(13), 
                           plusA(12) => prevA(12), plusA(11) => prevA(11), 
                           plusA(10) => prevA(10), plusA(9) => prevA(9), 
                           plusA(8) => prevA(8), plusA(7) => prevA(7), plusA(6)
                           => prevA(6), plusA(5) => prevA(5), plusA(4) => 
                           prevA(4), plusA(3) => prevA(3), plusA(2) => prevA(2)
                           , plusA(1) => prevA(1), plusA(0) => prevA(0), 
                           plus2A_out(63) => plus2A_s_63_port, plus2A_out(62) 
                           => plus2A_s_62_port, plus2A_out(61) => 
                           plus2A_s_61_port, plus2A_out(60) => plus2A_s_60_port
                           , plus2A_out(59) => plus2A_s_59_port, plus2A_out(58)
                           => plus2A_s_58_port, plus2A_out(57) => 
                           plus2A_s_57_port, plus2A_out(56) => plus2A_s_56_port
                           , plus2A_out(55) => plus2A_s_55_port, plus2A_out(54)
                           => plus2A_s_54_port, plus2A_out(53) => 
                           plus2A_s_53_port, plus2A_out(52) => plus2A_s_52_port
                           , plus2A_out(51) => plus2A_s_51_port, plus2A_out(50)
                           => plus2A_s_50_port, plus2A_out(49) => 
                           plus2A_s_49_port, plus2A_out(48) => plus2A_s_48_port
                           , plus2A_out(47) => plus2A_s_47_port, plus2A_out(46)
                           => plus2A_s_46_port, plus2A_out(45) => 
                           plus2A_s_45_port, plus2A_out(44) => plus2A_s_44_port
                           , plus2A_out(43) => plus2A_s_43_port, plus2A_out(42)
                           => plus2A_s_42_port, plus2A_out(41) => 
                           plus2A_s_41_port, plus2A_out(40) => plus2A_s_40_port
                           , plus2A_out(39) => plus2A_s_39_port, plus2A_out(38)
                           => plus2A_s_38_port, plus2A_out(37) => 
                           plus2A_s_37_port, plus2A_out(36) => plus2A_s_36_port
                           , plus2A_out(35) => plus2A_s_35_port, plus2A_out(34)
                           => plus2A_s_34_port, plus2A_out(33) => 
                           plus2A_s_33_port, plus2A_out(32) => plus2A_s_32_port
                           , plus2A_out(31) => plus2A_s_31_port, plus2A_out(30)
                           => plus2A_s_30_port, plus2A_out(29) => 
                           plus2A_s_29_port, plus2A_out(28) => plus2A_s_28_port
                           , plus2A_out(27) => plus2A_s_27_port, plus2A_out(26)
                           => plus2A_s_26_port, plus2A_out(25) => 
                           plus2A_s_25_port, plus2A_out(24) => plus2A_s_24_port
                           , plus2A_out(23) => plus2A_s_23_port, plus2A_out(22)
                           => plus2A_s_22_port, plus2A_out(21) => 
                           plus2A_s_21_port, plus2A_out(20) => plus2A_s_20_port
                           , plus2A_out(19) => plus2A_s_19_port, plus2A_out(18)
                           => plus2A_s_18_port, plus2A_out(17) => 
                           plus2A_s_17_port, plus2A_out(16) => plus2A_s_16_port
                           , plus2A_out(15) => plus2A_s_15_port, plus2A_out(14)
                           => plus2A_s_14_port, plus2A_out(13) => 
                           plus2A_s_13_port, plus2A_out(12) => plus2A_s_12_port
                           , plus2A_out(11) => plus2A_s_11_port, plus2A_out(10)
                           => plus2A_s_10_port, plus2A_out(9) => 
                           plus2A_s_9_port, plus2A_out(8) => plus2A_s_8_port, 
                           plus2A_out(7) => plus2A_s_7_port, plus2A_out(6) => 
                           plus2A_s_6_port, plus2A_out(5) => plus2A_s_5_port, 
                           plus2A_out(4) => plus2A_s_4_port, plus2A_out(3) => 
                           plus2A_s_3_port, plus2A_out(2) => plus2A_s_2_port, 
                           plus2A_out(1) => plus2A_s_1_port, plus2A_out(0) => 
                           n_3199, minus2A_out(63) => minus2A_s_63_port, 
                           minus2A_out(62) => minus2A_s_62_port, 
                           minus2A_out(61) => minus2A_s_61_port, 
                           minus2A_out(60) => minus2A_s_60_port, 
                           minus2A_out(59) => minus2A_s_59_port, 
                           minus2A_out(58) => minus2A_s_58_port, 
                           minus2A_out(57) => minus2A_s_57_port, 
                           minus2A_out(56) => minus2A_s_56_port, 
                           minus2A_out(55) => minus2A_s_55_port, 
                           minus2A_out(54) => minus2A_s_54_port, 
                           minus2A_out(53) => minus2A_s_53_port, 
                           minus2A_out(52) => minus2A_s_52_port, 
                           minus2A_out(51) => minus2A_s_51_port, 
                           minus2A_out(50) => minus2A_s_50_port, 
                           minus2A_out(49) => minus2A_s_49_port, 
                           minus2A_out(48) => minus2A_s_48_port, 
                           minus2A_out(47) => minus2A_s_47_port, 
                           minus2A_out(46) => minus2A_s_46_port, 
                           minus2A_out(45) => minus2A_s_45_port, 
                           minus2A_out(44) => minus2A_s_44_port, 
                           minus2A_out(43) => minus2A_s_43_port, 
                           minus2A_out(42) => minus2A_s_42_port, 
                           minus2A_out(41) => minus2A_s_41_port, 
                           minus2A_out(40) => minus2A_s_40_port, 
                           minus2A_out(39) => minus2A_s_39_port, 
                           minus2A_out(38) => minus2A_s_38_port, 
                           minus2A_out(37) => minus2A_s_37_port, 
                           minus2A_out(36) => minus2A_s_36_port, 
                           minus2A_out(35) => minus2A_s_35_port, 
                           minus2A_out(34) => minus2A_s_34_port, 
                           minus2A_out(33) => minus2A_s_33_port, 
                           minus2A_out(32) => minus2A_s_32_port, 
                           minus2A_out(31) => minus2A_s_31_port, 
                           minus2A_out(30) => minus2A_s_30_port, 
                           minus2A_out(29) => minus2A_s_29_port, 
                           minus2A_out(28) => minus2A_s_28_port, 
                           minus2A_out(27) => minus2A_s_27_port, 
                           minus2A_out(26) => minus2A_s_26_port, 
                           minus2A_out(25) => minus2A_s_25_port, 
                           minus2A_out(24) => minus2A_s_24_port, 
                           minus2A_out(23) => minus2A_s_23_port, 
                           minus2A_out(22) => minus2A_s_22_port, 
                           minus2A_out(21) => minus2A_s_21_port, 
                           minus2A_out(20) => minus2A_s_20_port, 
                           minus2A_out(19) => minus2A_s_19_port, 
                           minus2A_out(18) => minus2A_s_18_port, 
                           minus2A_out(17) => minus2A_s_17_port, 
                           minus2A_out(16) => minus2A_s_16_port, 
                           minus2A_out(15) => minus2A_s_15_port, 
                           minus2A_out(14) => minus2A_s_14_port, 
                           minus2A_out(13) => minus2A_s_13_port, 
                           minus2A_out(12) => minus2A_s_12_port, 
                           minus2A_out(11) => minus2A_s_11_port, 
                           minus2A_out(10) => minus2A_s_10_port, minus2A_out(9)
                           => minus2A_s_9_port, minus2A_out(8) => 
                           minus2A_s_8_port, minus2A_out(7) => minus2A_s_7_port
                           , minus2A_out(6) => minus2A_s_6_port, minus2A_out(5)
                           => minus2A_s_5_port, minus2A_out(4) => 
                           minus2A_s_4_port, minus2A_out(3) => minus2A_s_3_port
                           , minus2A_out(2) => minus2A_s_2_port, minus2A_out(1)
                           => minus2A_s_1_port, minus2A_out(0) => 
                           minus2A_s_0_port, plus4A_out(63) => nextA_63_port, 
                           plus4A_out(62) => nextA_62_port, plus4A_out(61) => 
                           nextA_61_port, plus4A_out(60) => nextA_60_port, 
                           plus4A_out(59) => nextA_59_port, plus4A_out(58) => 
                           nextA_58_port, plus4A_out(57) => n3, plus4A_out(56) 
                           => nextA_56_port, plus4A_out(55) => nextA_55_port, 
                           plus4A_out(54) => nextA_54_port, plus4A_out(53) => 
                           nextA_53_port, plus4A_out(52) => nextA_52_port, 
                           plus4A_out(51) => nextA_51_port, plus4A_out(50) => 
                           nextA_50_port, plus4A_out(49) => nextA_49_port, 
                           plus4A_out(48) => nextA_48_port, plus4A_out(47) => 
                           nextA_47_port, plus4A_out(46) => nextA_46_port, 
                           plus4A_out(45) => nextA_45_port, plus4A_out(44) => 
                           nextA_44_port, plus4A_out(43) => nextA_43_port, 
                           plus4A_out(42) => nextA_42_port, plus4A_out(41) => 
                           nextA_41_port, plus4A_out(40) => nextA_40_port, 
                           plus4A_out(39) => nextA_39_port, plus4A_out(38) => 
                           nextA_38_port, plus4A_out(37) => nextA_37_port, 
                           plus4A_out(36) => nextA_36_port, plus4A_out(35) => 
                           nextA_35_port, plus4A_out(34) => nextA_34_port, 
                           plus4A_out(33) => nextA_33_port, plus4A_out(32) => 
                           nextA_32_port, plus4A_out(31) => nextA_31_port, 
                           plus4A_out(30) => nextA_30_port, plus4A_out(29) => 
                           nextA_29_port, plus4A_out(28) => nextA_28_port, 
                           plus4A_out(27) => nextA_27_port, plus4A_out(26) => 
                           nextA_26_port, plus4A_out(25) => nextA_25_port, 
                           plus4A_out(24) => nextA_24_port, plus4A_out(23) => 
                           nextA_23_port, plus4A_out(22) => nextA_22_port, 
                           plus4A_out(21) => nextA_21_port, plus4A_out(20) => 
                           nextA_20_port, plus4A_out(19) => nextA_19_port, 
                           plus4A_out(18) => nextA_18_port, plus4A_out(17) => 
                           nextA_17_port, plus4A_out(16) => nextA_16_port, 
                           plus4A_out(15) => nextA_15_port, plus4A_out(14) => 
                           nextA_14_port, plus4A_out(13) => nextA_13_port, 
                           plus4A_out(12) => nextA_12_port, plus4A_out(11) => 
                           nextA_11_port, plus4A_out(10) => nextA_10_port, 
                           plus4A_out(9) => nextA_9_port, plus4A_out(8) => 
                           nextA_8_port, plus4A_out(7) => nextA_7_port, 
                           plus4A_out(6) => nextA_6_port, plus4A_out(5) => 
                           nextA_5_port, plus4A_out(4) => nextA_4_port, 
                           plus4A_out(3) => nextA_3_port, plus4A_out(2) => 
                           nextA_2_port, plus4A_out(1) => nextA_1_port, 
                           plus4A_out(0) => n_3200, minus4A_out(63) => 
                           minus4A_s_63_port, minus4A_out(62) => 
                           minus4A_s_62_port, minus4A_out(61) => 
                           minus4A_s_61_port, minus4A_out(60) => 
                           minus4A_s_60_port, minus4A_out(59) => 
                           minus4A_s_59_port, minus4A_out(58) => 
                           minus4A_s_58_port, minus4A_out(57) => 
                           minus4A_s_57_port, minus4A_out(56) => 
                           minus4A_s_56_port, minus4A_out(55) => 
                           minus4A_s_55_port, minus4A_out(54) => 
                           minus4A_s_54_port, minus4A_out(53) => 
                           minus4A_s_53_port, minus4A_out(52) => 
                           minus4A_s_52_port, minus4A_out(51) => 
                           minus4A_s_51_port, minus4A_out(50) => 
                           minus4A_s_50_port, minus4A_out(49) => 
                           minus4A_s_49_port, minus4A_out(48) => 
                           minus4A_s_48_port, minus4A_out(47) => 
                           minus4A_s_47_port, minus4A_out(46) => 
                           minus4A_s_46_port, minus4A_out(45) => 
                           minus4A_s_45_port, minus4A_out(44) => 
                           minus4A_s_44_port, minus4A_out(43) => 
                           minus4A_s_43_port, minus4A_out(42) => 
                           minus4A_s_42_port, minus4A_out(41) => 
                           minus4A_s_41_port, minus4A_out(40) => 
                           minus4A_s_40_port, minus4A_out(39) => 
                           minus4A_s_39_port, minus4A_out(38) => 
                           minus4A_s_38_port, minus4A_out(37) => 
                           minus4A_s_37_port, minus4A_out(36) => 
                           minus4A_s_36_port, minus4A_out(35) => 
                           minus4A_s_35_port, minus4A_out(34) => 
                           minus4A_s_34_port, minus4A_out(33) => 
                           minus4A_s_33_port, minus4A_out(32) => 
                           minus4A_s_32_port, minus4A_out(31) => 
                           minus4A_s_31_port, minus4A_out(30) => 
                           minus4A_s_30_port, minus4A_out(29) => 
                           minus4A_s_29_port, minus4A_out(28) => 
                           minus4A_s_28_port, minus4A_out(27) => 
                           minus4A_s_27_port, minus4A_out(26) => 
                           minus4A_s_26_port, minus4A_out(25) => 
                           minus4A_s_25_port, minus4A_out(24) => 
                           minus4A_s_24_port, minus4A_out(23) => 
                           minus4A_s_23_port, minus4A_out(22) => 
                           minus4A_s_22_port, minus4A_out(21) => 
                           minus4A_s_21_port, minus4A_out(20) => 
                           minus4A_s_20_port, minus4A_out(19) => 
                           minus4A_s_19_port, minus4A_out(18) => 
                           minus4A_s_18_port, minus4A_out(17) => 
                           minus4A_s_17_port, minus4A_out(16) => 
                           minus4A_s_16_port, minus4A_out(15) => 
                           minus4A_s_15_port, minus4A_out(14) => 
                           minus4A_s_14_port, minus4A_out(13) => 
                           minus4A_s_13_port, minus4A_out(12) => 
                           minus4A_s_12_port, minus4A_out(11) => 
                           minus4A_s_11_port, minus4A_out(10) => 
                           minus4A_s_10_port, minus4A_out(9) => 
                           minus4A_s_9_port, minus4A_out(8) => minus4A_s_8_port
                           , minus4A_out(7) => minus4A_s_7_port, minus4A_out(6)
                           => minus4A_s_6_port, minus4A_out(5) => 
                           minus4A_s_5_port, minus4A_out(4) => minus4A_s_4_port
                           , minus4A_out(3) => minus4A_s_3_port, minus4A_out(2)
                           => minus4A_s_2_port, minus4A_out(1) => 
                           minus4A_s_1_port, minus4A_out(0) => minus4A_s_0_port
                           );
   mux_1 : MUX_GENERIC_N64_RADIX3_9 port map( plusA(63) => plus2A_s_63_port, 
                           plusA(62) => plus2A_s_62_port, plusA(61) => 
                           plus2A_s_61_port, plusA(60) => plus2A_s_60_port, 
                           plusA(59) => plus2A_s_59_port, plusA(58) => 
                           plus2A_s_58_port, plusA(57) => plus2A_s_57_port, 
                           plusA(56) => plus2A_s_56_port, plusA(55) => 
                           plus2A_s_55_port, plusA(54) => plus2A_s_54_port, 
                           plusA(53) => plus2A_s_53_port, plusA(52) => 
                           plus2A_s_52_port, plusA(51) => plus2A_s_51_port, 
                           plusA(50) => plus2A_s_50_port, plusA(49) => 
                           plus2A_s_49_port, plusA(48) => plus2A_s_48_port, 
                           plusA(47) => plus2A_s_47_port, plusA(46) => 
                           plus2A_s_46_port, plusA(45) => plus2A_s_45_port, 
                           plusA(44) => plus2A_s_44_port, plusA(43) => 
                           plus2A_s_43_port, plusA(42) => plus2A_s_42_port, 
                           plusA(41) => plus2A_s_41_port, plusA(40) => 
                           plus2A_s_40_port, plusA(39) => plus2A_s_39_port, 
                           plusA(38) => plus2A_s_38_port, plusA(37) => 
                           plus2A_s_37_port, plusA(36) => plus2A_s_36_port, 
                           plusA(35) => plus2A_s_35_port, plusA(34) => 
                           plus2A_s_34_port, plusA(33) => plus2A_s_33_port, 
                           plusA(32) => plus2A_s_32_port, plusA(31) => 
                           plus2A_s_31_port, plusA(30) => plus2A_s_30_port, 
                           plusA(29) => plus2A_s_29_port, plusA(28) => 
                           plus2A_s_28_port, plusA(27) => plus2A_s_27_port, 
                           plusA(26) => plus2A_s_26_port, plusA(25) => 
                           plus2A_s_25_port, plusA(24) => plus2A_s_24_port, 
                           plusA(23) => plus2A_s_23_port, plusA(22) => 
                           plus2A_s_22_port, plusA(21) => plus2A_s_21_port, 
                           plusA(20) => plus2A_s_20_port, plusA(19) => 
                           plus2A_s_19_port, plusA(18) => plus2A_s_18_port, 
                           plusA(17) => plus2A_s_17_port, plusA(16) => 
                           plus2A_s_16_port, plusA(15) => plus2A_s_15_port, 
                           plusA(14) => plus2A_s_14_port, plusA(13) => 
                           plus2A_s_13_port, plusA(12) => plus2A_s_12_port, 
                           plusA(11) => plus2A_s_11_port, plusA(10) => 
                           plus2A_s_10_port, plusA(9) => plus2A_s_9_port, 
                           plusA(8) => plus2A_s_8_port, plusA(7) => 
                           plus2A_s_7_port, plusA(6) => plus2A_s_6_port, 
                           plusA(5) => plus2A_s_5_port, plusA(4) => 
                           plus2A_s_4_port, plusA(3) => plus2A_s_3_port, 
                           plusA(2) => plus2A_s_2_port, plusA(1) => 
                           plus2A_s_1_port, plusA(0) => nextA_0_port, 
                           minusA(63) => minus2A_s_63_port, minusA(62) => 
                           minus2A_s_62_port, minusA(61) => minus2A_s_61_port, 
                           minusA(60) => minus2A_s_60_port, minusA(59) => 
                           minus2A_s_59_port, minusA(58) => minus2A_s_58_port, 
                           minusA(57) => minus2A_s_57_port, minusA(56) => 
                           minus2A_s_56_port, minusA(55) => minus2A_s_55_port, 
                           minusA(54) => minus2A_s_54_port, minusA(53) => 
                           minus2A_s_53_port, minusA(52) => minus2A_s_52_port, 
                           minusA(51) => minus2A_s_51_port, minusA(50) => 
                           minus2A_s_50_port, minusA(49) => minus2A_s_49_port, 
                           minusA(48) => minus2A_s_48_port, minusA(47) => 
                           minus2A_s_47_port, minusA(46) => minus2A_s_46_port, 
                           minusA(45) => minus2A_s_45_port, minusA(44) => 
                           minus2A_s_44_port, minusA(43) => minus2A_s_43_port, 
                           minusA(42) => minus2A_s_42_port, minusA(41) => 
                           minus2A_s_41_port, minusA(40) => minus2A_s_40_port, 
                           minusA(39) => minus2A_s_39_port, minusA(38) => 
                           minus2A_s_38_port, minusA(37) => minus2A_s_37_port, 
                           minusA(36) => minus2A_s_36_port, minusA(35) => 
                           minus2A_s_35_port, minusA(34) => minus2A_s_34_port, 
                           minusA(33) => minus2A_s_33_port, minusA(32) => 
                           minus2A_s_32_port, minusA(31) => minus2A_s_31_port, 
                           minusA(30) => minus2A_s_30_port, minusA(29) => 
                           minus2A_s_29_port, minusA(28) => minus2A_s_28_port, 
                           minusA(27) => minus2A_s_27_port, minusA(26) => 
                           minus2A_s_26_port, minusA(25) => minus2A_s_25_port, 
                           minusA(24) => minus2A_s_24_port, minusA(23) => 
                           minus2A_s_23_port, minusA(22) => minus2A_s_22_port, 
                           minusA(21) => minus2A_s_21_port, minusA(20) => 
                           minus2A_s_20_port, minusA(19) => minus2A_s_19_port, 
                           minusA(18) => minus2A_s_18_port, minusA(17) => 
                           minus2A_s_17_port, minusA(16) => minus2A_s_16_port, 
                           minusA(15) => minus2A_s_15_port, minusA(14) => 
                           minus2A_s_14_port, minusA(13) => minus2A_s_13_port, 
                           minusA(12) => minus2A_s_12_port, minusA(11) => 
                           minus2A_s_11_port, minusA(10) => minus2A_s_10_port, 
                           minusA(9) => minus2A_s_9_port, minusA(8) => 
                           minus2A_s_8_port, minusA(7) => minus2A_s_7_port, 
                           minusA(6) => minus2A_s_6_port, minusA(5) => 
                           minus2A_s_5_port, minusA(4) => minus2A_s_4_port, 
                           minusA(3) => minus2A_s_3_port, minusA(2) => 
                           minus2A_s_2_port, minusA(1) => minus2A_s_1_port, 
                           minusA(0) => minus2A_s_0_port, plus2A(63) => 
                           nextA_63_port, plus2A(62) => nextA_62_port, 
                           plus2A(61) => nextA_61_port, plus2A(60) => 
                           nextA_60_port, plus2A(59) => nextA_59_port, 
                           plus2A(58) => nextA_58_port, plus2A(57) => 
                           nextA_57_port, plus2A(56) => nextA_56_port, 
                           plus2A(55) => nextA_55_port, plus2A(54) => 
                           nextA_54_port, plus2A(53) => nextA_53_port, 
                           plus2A(52) => nextA_52_port, plus2A(51) => 
                           nextA_51_port, plus2A(50) => nextA_50_port, 
                           plus2A(49) => nextA_49_port, plus2A(48) => 
                           nextA_48_port, plus2A(47) => nextA_47_port, 
                           plus2A(46) => nextA_46_port, plus2A(45) => 
                           nextA_45_port, plus2A(44) => nextA_44_port, 
                           plus2A(43) => nextA_43_port, plus2A(42) => 
                           nextA_42_port, plus2A(41) => nextA_41_port, 
                           plus2A(40) => nextA_40_port, plus2A(39) => 
                           nextA_39_port, plus2A(38) => nextA_38_port, 
                           plus2A(37) => nextA_37_port, plus2A(36) => 
                           nextA_36_port, plus2A(35) => nextA_35_port, 
                           plus2A(34) => nextA_34_port, plus2A(33) => 
                           nextA_33_port, plus2A(32) => nextA_32_port, 
                           plus2A(31) => nextA_31_port, plus2A(30) => 
                           nextA_30_port, plus2A(29) => nextA_29_port, 
                           plus2A(28) => nextA_28_port, plus2A(27) => 
                           nextA_27_port, plus2A(26) => nextA_26_port, 
                           plus2A(25) => nextA_25_port, plus2A(24) => 
                           nextA_24_port, plus2A(23) => nextA_23_port, 
                           plus2A(22) => nextA_22_port, plus2A(21) => 
                           nextA_21_port, plus2A(20) => nextA_20_port, 
                           plus2A(19) => nextA_19_port, plus2A(18) => 
                           nextA_18_port, plus2A(17) => nextA_17_port, 
                           plus2A(16) => nextA_16_port, plus2A(15) => 
                           nextA_15_port, plus2A(14) => nextA_14_port, 
                           plus2A(13) => nextA_13_port, plus2A(12) => 
                           nextA_12_port, plus2A(11) => nextA_11_port, 
                           plus2A(10) => nextA_10_port, plus2A(9) => 
                           nextA_9_port, plus2A(8) => nextA_8_port, plus2A(7) 
                           => nextA_7_port, plus2A(6) => nextA_6_port, 
                           plus2A(5) => nextA_5_port, plus2A(4) => nextA_4_port
                           , plus2A(3) => nextA_3_port, plus2A(2) => 
                           nextA_2_port, plus2A(1) => nextA_1_port, plus2A(0) 
                           => nextA_0_port, minus2A(63) => minus4A_s_63_port, 
                           minus2A(62) => minus4A_s_62_port, minus2A(61) => 
                           minus4A_s_61_port, minus2A(60) => minus4A_s_60_port,
                           minus2A(59) => minus4A_s_59_port, minus2A(58) => 
                           minus4A_s_58_port, minus2A(57) => minus4A_s_57_port,
                           minus2A(56) => minus4A_s_56_port, minus2A(55) => 
                           minus4A_s_55_port, minus2A(54) => minus4A_s_54_port,
                           minus2A(53) => minus4A_s_53_port, minus2A(52) => 
                           minus4A_s_52_port, minus2A(51) => minus4A_s_51_port,
                           minus2A(50) => minus4A_s_50_port, minus2A(49) => 
                           minus4A_s_49_port, minus2A(48) => minus4A_s_48_port,
                           minus2A(47) => minus4A_s_47_port, minus2A(46) => 
                           minus4A_s_46_port, minus2A(45) => minus4A_s_45_port,
                           minus2A(44) => minus4A_s_44_port, minus2A(43) => 
                           minus4A_s_43_port, minus2A(42) => minus4A_s_42_port,
                           minus2A(41) => minus4A_s_41_port, minus2A(40) => 
                           minus4A_s_40_port, minus2A(39) => minus4A_s_39_port,
                           minus2A(38) => minus4A_s_38_port, minus2A(37) => 
                           minus4A_s_37_port, minus2A(36) => minus4A_s_36_port,
                           minus2A(35) => minus4A_s_35_port, minus2A(34) => 
                           minus4A_s_34_port, minus2A(33) => minus4A_s_33_port,
                           minus2A(32) => minus4A_s_32_port, minus2A(31) => 
                           minus4A_s_31_port, minus2A(30) => minus4A_s_30_port,
                           minus2A(29) => minus4A_s_29_port, minus2A(28) => 
                           minus4A_s_28_port, minus2A(27) => minus4A_s_27_port,
                           minus2A(26) => minus4A_s_26_port, minus2A(25) => 
                           minus4A_s_25_port, minus2A(24) => minus4A_s_24_port,
                           minus2A(23) => minus4A_s_23_port, minus2A(22) => 
                           minus4A_s_22_port, minus2A(21) => minus4A_s_21_port,
                           minus2A(20) => minus4A_s_20_port, minus2A(19) => 
                           minus4A_s_19_port, minus2A(18) => minus4A_s_18_port,
                           minus2A(17) => minus4A_s_17_port, minus2A(16) => 
                           minus4A_s_16_port, minus2A(15) => minus4A_s_15_port,
                           minus2A(14) => minus4A_s_14_port, minus2A(13) => 
                           minus4A_s_13_port, minus2A(12) => minus4A_s_12_port,
                           minus2A(11) => minus4A_s_11_port, minus2A(10) => 
                           minus4A_s_10_port, minus2A(9) => minus4A_s_9_port, 
                           minus2A(8) => minus4A_s_8_port, minus2A(7) => 
                           minus4A_s_7_port, minus2A(6) => minus4A_s_6_port, 
                           minus2A(5) => minus4A_s_5_port, minus2A(4) => 
                           minus4A_s_4_port, minus2A(3) => minus4A_s_3_port, 
                           minus2A(2) => minus4A_s_2_port, minus2A(1) => 
                           minus4A_s_1_port, minus2A(0) => minus4A_s_0_port, 
                           SEL(2) => encoder_to_mux_2_port, SEL(1) => 
                           encoder_to_mux_1_port, SEL(0) => 
                           encoder_to_mux_0_port, Y(63) => mux_to_adder_63_port
                           , Y(62) => mux_to_adder_62_port, Y(61) => 
                           mux_to_adder_61_port, Y(60) => mux_to_adder_60_port,
                           Y(59) => mux_to_adder_59_port, Y(58) => 
                           mux_to_adder_58_port, Y(57) => mux_to_adder_57_port,
                           Y(56) => mux_to_adder_56_port, Y(55) => 
                           mux_to_adder_55_port, Y(54) => mux_to_adder_54_port,
                           Y(53) => mux_to_adder_53_port, Y(52) => 
                           mux_to_adder_52_port, Y(51) => mux_to_adder_51_port,
                           Y(50) => mux_to_adder_50_port, Y(49) => 
                           mux_to_adder_49_port, Y(48) => mux_to_adder_48_port,
                           Y(47) => mux_to_adder_47_port, Y(46) => 
                           mux_to_adder_46_port, Y(45) => mux_to_adder_45_port,
                           Y(44) => mux_to_adder_44_port, Y(43) => 
                           mux_to_adder_43_port, Y(42) => mux_to_adder_42_port,
                           Y(41) => mux_to_adder_41_port, Y(40) => 
                           mux_to_adder_40_port, Y(39) => mux_to_adder_39_port,
                           Y(38) => mux_to_adder_38_port, Y(37) => 
                           mux_to_adder_37_port, Y(36) => mux_to_adder_36_port,
                           Y(35) => mux_to_adder_35_port, Y(34) => 
                           mux_to_adder_34_port, Y(33) => mux_to_adder_33_port,
                           Y(32) => mux_to_adder_32_port, Y(31) => 
                           mux_to_adder_31_port, Y(30) => mux_to_adder_30_port,
                           Y(29) => mux_to_adder_29_port, Y(28) => 
                           mux_to_adder_28_port, Y(27) => mux_to_adder_27_port,
                           Y(26) => mux_to_adder_26_port, Y(25) => 
                           mux_to_adder_25_port, Y(24) => mux_to_adder_24_port,
                           Y(23) => mux_to_adder_23_port, Y(22) => 
                           mux_to_adder_22_port, Y(21) => mux_to_adder_21_port,
                           Y(20) => mux_to_adder_20_port, Y(19) => 
                           mux_to_adder_19_port, Y(18) => mux_to_adder_18_port,
                           Y(17) => mux_to_adder_17_port, Y(16) => 
                           mux_to_adder_16_port, Y(15) => mux_to_adder_15_port,
                           Y(14) => mux_to_adder_14_port, Y(13) => 
                           mux_to_adder_13_port, Y(12) => mux_to_adder_12_port,
                           Y(11) => mux_to_adder_11_port, Y(10) => 
                           mux_to_adder_10_port, Y(9) => mux_to_adder_9_port, 
                           Y(8) => mux_to_adder_8_port, Y(7) => 
                           mux_to_adder_7_port, Y(6) => mux_to_adder_6_port, 
                           Y(5) => mux_to_adder_5_port, Y(4) => 
                           mux_to_adder_4_port, Y(3) => mux_to_adder_3_port, 
                           Y(2) => mux_to_adder_2_port, Y(1) => 
                           mux_to_adder_1_port, Y(0) => mux_to_adder_0_port);
   rca_1 : RCA_N64_9 port map( A(63) => mux_to_adder_63_port, A(62) => 
                           mux_to_adder_62_port, A(61) => mux_to_adder_61_port,
                           A(60) => mux_to_adder_60_port, A(59) => 
                           mux_to_adder_59_port, A(58) => mux_to_adder_58_port,
                           A(57) => mux_to_adder_57_port, A(56) => 
                           mux_to_adder_56_port, A(55) => mux_to_adder_55_port,
                           A(54) => mux_to_adder_54_port, A(53) => 
                           mux_to_adder_53_port, A(52) => mux_to_adder_52_port,
                           A(51) => mux_to_adder_51_port, A(50) => 
                           mux_to_adder_50_port, A(49) => mux_to_adder_49_port,
                           A(48) => mux_to_adder_48_port, A(47) => 
                           mux_to_adder_47_port, A(46) => mux_to_adder_46_port,
                           A(45) => mux_to_adder_45_port, A(44) => 
                           mux_to_adder_44_port, A(43) => mux_to_adder_43_port,
                           A(42) => mux_to_adder_42_port, A(41) => 
                           mux_to_adder_41_port, A(40) => mux_to_adder_40_port,
                           A(39) => mux_to_adder_39_port, A(38) => 
                           mux_to_adder_38_port, A(37) => mux_to_adder_37_port,
                           A(36) => mux_to_adder_36_port, A(35) => 
                           mux_to_adder_35_port, A(34) => mux_to_adder_34_port,
                           A(33) => mux_to_adder_33_port, A(32) => 
                           mux_to_adder_32_port, A(31) => mux_to_adder_31_port,
                           A(30) => mux_to_adder_30_port, A(29) => 
                           mux_to_adder_29_port, A(28) => mux_to_adder_28_port,
                           A(27) => mux_to_adder_27_port, A(26) => 
                           mux_to_adder_26_port, A(25) => mux_to_adder_25_port,
                           A(24) => mux_to_adder_24_port, A(23) => 
                           mux_to_adder_23_port, A(22) => mux_to_adder_22_port,
                           A(21) => mux_to_adder_21_port, A(20) => 
                           mux_to_adder_20_port, A(19) => mux_to_adder_19_port,
                           A(18) => mux_to_adder_18_port, A(17) => 
                           mux_to_adder_17_port, A(16) => mux_to_adder_16_port,
                           A(15) => mux_to_adder_15_port, A(14) => 
                           mux_to_adder_14_port, A(13) => mux_to_adder_13_port,
                           A(12) => mux_to_adder_12_port, A(11) => 
                           mux_to_adder_11_port, A(10) => mux_to_adder_10_port,
                           A(9) => mux_to_adder_9_port, A(8) => 
                           mux_to_adder_8_port, A(7) => mux_to_adder_7_port, 
                           A(6) => mux_to_adder_6_port, A(5) => 
                           mux_to_adder_5_port, A(4) => mux_to_adder_4_port, 
                           A(3) => mux_to_adder_3_port, A(2) => 
                           mux_to_adder_2_port, A(1) => mux_to_adder_1_port, 
                           A(0) => mux_to_adder_0_port, B(63) => prevSum(63), 
                           B(62) => prevSum(62), B(61) => prevSum(61), B(60) =>
                           prevSum(60), B(59) => prevSum(59), B(58) => 
                           prevSum(58), B(57) => prevSum(57), B(56) => 
                           prevSum(56), B(55) => prevSum(55), B(54) => 
                           prevSum(54), B(53) => prevSum(53), B(52) => 
                           prevSum(52), B(51) => prevSum(51), B(50) => 
                           prevSum(50), B(49) => prevSum(49), B(48) => 
                           prevSum(48), B(47) => prevSum(47), B(46) => 
                           prevSum(46), B(45) => prevSum(45), B(44) => 
                           prevSum(44), B(43) => prevSum(43), B(42) => 
                           prevSum(42), B(41) => prevSum(41), B(40) => 
                           prevSum(40), B(39) => prevSum(39), B(38) => 
                           prevSum(38), B(37) => prevSum(37), B(36) => 
                           prevSum(36), B(35) => prevSum(35), B(34) => 
                           prevSum(34), B(33) => prevSum(33), B(32) => 
                           prevSum(32), B(31) => prevSum(31), B(30) => 
                           prevSum(30), B(29) => prevSum(29), B(28) => 
                           prevSum(28), B(27) => prevSum(27), B(26) => 
                           prevSum(26), B(25) => prevSum(25), B(24) => 
                           prevSum(24), B(23) => prevSum(23), B(22) => 
                           prevSum(22), B(21) => prevSum(21), B(20) => 
                           prevSum(20), B(19) => prevSum(19), B(18) => 
                           prevSum(18), B(17) => prevSum(17), B(16) => 
                           prevSum(16), B(15) => prevSum(15), B(14) => 
                           prevSum(14), B(13) => prevSum(13), B(12) => 
                           prevSum(12), B(11) => prevSum(11), B(10) => 
                           prevSum(10), B(9) => prevSum(9), B(8) => prevSum(8),
                           B(7) => prevSum(7), B(6) => prevSum(6), B(5) => 
                           prevSum(5), B(4) => prevSum(4), B(3) => prevSum(3), 
                           B(2) => prevSum(2), B(1) => prevSum(1), B(0) => 
                           prevSum(0), Ci => X_Logic0_port, S(63) => 
                           nextSum(63), S(62) => nextSum(62), S(61) => 
                           nextSum(61), S(60) => nextSum(60), S(59) => 
                           nextSum(59), S(58) => nextSum(58), S(57) => 
                           nextSum(57), S(56) => nextSum(56), S(55) => 
                           nextSum(55), S(54) => nextSum(54), S(53) => 
                           nextSum(53), S(52) => nextSum(52), S(51) => 
                           nextSum(51), S(50) => nextSum(50), S(49) => 
                           nextSum(49), S(48) => nextSum(48), S(47) => 
                           nextSum(47), S(46) => nextSum(46), S(45) => 
                           nextSum(45), S(44) => nextSum(44), S(43) => 
                           nextSum(43), S(42) => nextSum(42), S(41) => 
                           nextSum(41), S(40) => nextSum(40), S(39) => 
                           nextSum(39), S(38) => nextSum(38), S(37) => 
                           nextSum(37), S(36) => nextSum(36), S(35) => 
                           nextSum(35), S(34) => nextSum(34), S(33) => 
                           nextSum(33), S(32) => nextSum(32), S(31) => 
                           nextSum(31), S(30) => nextSum(30), S(29) => 
                           nextSum(29), S(28) => nextSum(28), S(27) => 
                           nextSum(27), S(26) => nextSum(26), S(25) => 
                           nextSum(25), S(24) => nextSum(24), S(23) => 
                           nextSum(23), S(22) => nextSum(22), S(21) => 
                           nextSum(21), S(20) => nextSum(20), S(19) => 
                           nextSum(19), S(18) => nextSum(18), S(17) => 
                           nextSum(17), S(16) => nextSum(16), S(15) => 
                           nextSum(15), S(14) => nextSum(14), S(13) => 
                           nextSum(13), S(12) => nextSum(12), S(11) => 
                           nextSum(11), S(10) => nextSum(10), S(9) => 
                           nextSum(9), S(8) => nextSum(8), S(7) => nextSum(7), 
                           S(6) => nextSum(6), S(5) => nextSum(5), S(4) => 
                           nextSum(4), S(3) => nextSum(3), S(2) => nextSum(2), 
                           S(1) => nextSum(1), S(0) => nextSum(0), Co => n_3201
                           );
   U3 : BUF_X1 port map( A => n3, Z => nextA_57_port);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity booth_mul_row_N64_RADIX3_10 is

   port( prevA, prevSum : in std_logic_vector (63 downto 0);  encoderIn : in 
         std_logic_vector (2 downto 0);  nextA, nextSum : out std_logic_vector 
         (63 downto 0));

end booth_mul_row_N64_RADIX3_10;

architecture SYN_struct of booth_mul_row_N64_RADIX3_10 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component RCA_N64_10
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component MUX_GENERIC_N64_RADIX3_10
      port( plusA, minusA, plus2A, minus2A : in std_logic_vector (63 downto 0);
            SEL : in std_logic_vector (2 downto 0);  Y : out std_logic_vector 
            (63 downto 0));
   end component;
   
   component ShiftnCompl_N64_10
      port( plusA : in std_logic_vector (63 downto 0);  plus2A_out, minus2A_out
            , plus4A_out, minus4A_out : out std_logic_vector (63 downto 0));
   end component;
   
   component encoder_N64_RADIX3_10
      port( X : in std_logic_vector (2 downto 0);  Z : out std_logic_vector (2 
            downto 0));
   end component;
   
   signal X_Logic0_port, nextA_63_port, nextA_62_port, nextA_61_port, 
      nextA_60_port, nextA_59_port, nextA_58_port, n3, nextA_56_port, 
      nextA_55_port, nextA_54_port, nextA_53_port, nextA_52_port, nextA_51_port
      , nextA_50_port, nextA_49_port, nextA_48_port, nextA_47_port, 
      nextA_46_port, nextA_45_port, nextA_44_port, nextA_43_port, nextA_42_port
      , nextA_41_port, nextA_40_port, nextA_39_port, nextA_38_port, 
      nextA_37_port, nextA_36_port, nextA_35_port, nextA_34_port, nextA_33_port
      , nextA_32_port, nextA_31_port, nextA_30_port, nextA_29_port, 
      nextA_28_port, nextA_27_port, nextA_26_port, nextA_25_port, nextA_24_port
      , nextA_23_port, nextA_22_port, nextA_21_port, nextA_20_port, 
      nextA_19_port, nextA_18_port, nextA_17_port, nextA_16_port, nextA_15_port
      , nextA_14_port, nextA_13_port, nextA_12_port, nextA_11_port, 
      nextA_10_port, nextA_9_port, nextA_8_port, nextA_7_port, nextA_6_port, 
      nextA_5_port, nextA_4_port, nextA_3_port, nextA_2_port, nextA_1_port, 
      encoder_to_mux_2_port, encoder_to_mux_1_port, encoder_to_mux_0_port, 
      plus2A_s_63_port, plus2A_s_62_port, plus2A_s_61_port, plus2A_s_60_port, 
      plus2A_s_59_port, plus2A_s_58_port, plus2A_s_57_port, plus2A_s_56_port, 
      plus2A_s_55_port, plus2A_s_54_port, plus2A_s_53_port, plus2A_s_52_port, 
      plus2A_s_51_port, plus2A_s_50_port, plus2A_s_49_port, plus2A_s_48_port, 
      plus2A_s_47_port, plus2A_s_46_port, plus2A_s_45_port, plus2A_s_44_port, 
      plus2A_s_43_port, plus2A_s_42_port, plus2A_s_41_port, plus2A_s_40_port, 
      plus2A_s_39_port, plus2A_s_38_port, plus2A_s_37_port, plus2A_s_36_port, 
      plus2A_s_35_port, plus2A_s_34_port, plus2A_s_33_port, plus2A_s_32_port, 
      plus2A_s_31_port, plus2A_s_30_port, plus2A_s_29_port, plus2A_s_28_port, 
      plus2A_s_27_port, plus2A_s_26_port, plus2A_s_25_port, plus2A_s_24_port, 
      plus2A_s_23_port, plus2A_s_22_port, plus2A_s_21_port, plus2A_s_20_port, 
      plus2A_s_19_port, plus2A_s_18_port, plus2A_s_17_port, plus2A_s_16_port, 
      plus2A_s_15_port, plus2A_s_14_port, plus2A_s_13_port, plus2A_s_12_port, 
      plus2A_s_11_port, plus2A_s_10_port, plus2A_s_9_port, plus2A_s_8_port, 
      plus2A_s_7_port, plus2A_s_6_port, plus2A_s_5_port, plus2A_s_4_port, 
      plus2A_s_3_port, plus2A_s_2_port, plus2A_s_1_port, minus2A_s_63_port, 
      minus2A_s_62_port, minus2A_s_61_port, minus2A_s_60_port, 
      minus2A_s_59_port, minus2A_s_58_port, minus2A_s_57_port, 
      minus2A_s_56_port, minus2A_s_55_port, minus2A_s_54_port, 
      minus2A_s_53_port, minus2A_s_52_port, minus2A_s_51_port, 
      minus2A_s_50_port, minus2A_s_49_port, minus2A_s_48_port, 
      minus2A_s_47_port, minus2A_s_46_port, minus2A_s_45_port, 
      minus2A_s_44_port, minus2A_s_43_port, minus2A_s_42_port, 
      minus2A_s_41_port, minus2A_s_40_port, minus2A_s_39_port, 
      minus2A_s_38_port, minus2A_s_37_port, minus2A_s_36_port, 
      minus2A_s_35_port, minus2A_s_34_port, minus2A_s_33_port, 
      minus2A_s_32_port, minus2A_s_31_port, minus2A_s_30_port, 
      minus2A_s_29_port, minus2A_s_28_port, minus2A_s_27_port, 
      minus2A_s_26_port, minus2A_s_25_port, minus2A_s_24_port, 
      minus2A_s_23_port, minus2A_s_22_port, minus2A_s_21_port, 
      minus2A_s_20_port, minus2A_s_19_port, minus2A_s_18_port, 
      minus2A_s_17_port, minus2A_s_16_port, minus2A_s_15_port, 
      minus2A_s_14_port, minus2A_s_13_port, minus2A_s_12_port, 
      minus2A_s_11_port, minus2A_s_10_port, minus2A_s_9_port, minus2A_s_8_port,
      minus2A_s_7_port, minus2A_s_6_port, minus2A_s_5_port, minus2A_s_4_port, 
      minus2A_s_3_port, minus2A_s_2_port, minus2A_s_1_port, minus2A_s_0_port, 
      minus4A_s_63_port, minus4A_s_62_port, minus4A_s_61_port, 
      minus4A_s_60_port, minus4A_s_59_port, minus4A_s_58_port, 
      minus4A_s_57_port, minus4A_s_56_port, minus4A_s_55_port, 
      minus4A_s_54_port, minus4A_s_53_port, minus4A_s_52_port, 
      minus4A_s_51_port, minus4A_s_50_port, minus4A_s_49_port, 
      minus4A_s_48_port, minus4A_s_47_port, minus4A_s_46_port, 
      minus4A_s_45_port, minus4A_s_44_port, minus4A_s_43_port, 
      minus4A_s_42_port, minus4A_s_41_port, minus4A_s_40_port, 
      minus4A_s_39_port, minus4A_s_38_port, minus4A_s_37_port, 
      minus4A_s_36_port, minus4A_s_35_port, minus4A_s_34_port, 
      minus4A_s_33_port, minus4A_s_32_port, minus4A_s_31_port, 
      minus4A_s_30_port, minus4A_s_29_port, minus4A_s_28_port, 
      minus4A_s_27_port, minus4A_s_26_port, minus4A_s_25_port, 
      minus4A_s_24_port, minus4A_s_23_port, minus4A_s_22_port, 
      minus4A_s_21_port, minus4A_s_20_port, minus4A_s_19_port, 
      minus4A_s_18_port, minus4A_s_17_port, minus4A_s_16_port, 
      minus4A_s_15_port, minus4A_s_14_port, minus4A_s_13_port, 
      minus4A_s_12_port, minus4A_s_11_port, minus4A_s_10_port, minus4A_s_9_port
      , minus4A_s_8_port, minus4A_s_7_port, minus4A_s_6_port, minus4A_s_5_port,
      minus4A_s_4_port, minus4A_s_3_port, minus4A_s_2_port, minus4A_s_1_port, 
      minus4A_s_0_port, mux_to_adder_63_port, mux_to_adder_62_port, 
      mux_to_adder_61_port, mux_to_adder_60_port, mux_to_adder_59_port, 
      mux_to_adder_58_port, mux_to_adder_57_port, mux_to_adder_56_port, 
      mux_to_adder_55_port, mux_to_adder_54_port, mux_to_adder_53_port, 
      mux_to_adder_52_port, mux_to_adder_51_port, mux_to_adder_50_port, 
      mux_to_adder_49_port, mux_to_adder_48_port, mux_to_adder_47_port, 
      mux_to_adder_46_port, mux_to_adder_45_port, mux_to_adder_44_port, 
      mux_to_adder_43_port, mux_to_adder_42_port, mux_to_adder_41_port, 
      mux_to_adder_40_port, mux_to_adder_39_port, mux_to_adder_38_port, 
      mux_to_adder_37_port, mux_to_adder_36_port, mux_to_adder_35_port, 
      mux_to_adder_34_port, mux_to_adder_33_port, mux_to_adder_32_port, 
      mux_to_adder_31_port, mux_to_adder_30_port, mux_to_adder_29_port, 
      mux_to_adder_28_port, mux_to_adder_27_port, mux_to_adder_26_port, 
      mux_to_adder_25_port, mux_to_adder_24_port, mux_to_adder_23_port, 
      mux_to_adder_22_port, mux_to_adder_21_port, mux_to_adder_20_port, 
      mux_to_adder_19_port, mux_to_adder_18_port, mux_to_adder_17_port, 
      mux_to_adder_16_port, mux_to_adder_15_port, mux_to_adder_14_port, 
      mux_to_adder_13_port, mux_to_adder_12_port, mux_to_adder_11_port, 
      mux_to_adder_10_port, mux_to_adder_9_port, mux_to_adder_8_port, 
      mux_to_adder_7_port, mux_to_adder_6_port, mux_to_adder_5_port, 
      mux_to_adder_4_port, mux_to_adder_3_port, mux_to_adder_2_port, 
      mux_to_adder_1_port, mux_to_adder_0_port, nextA_0_port, nextA_57_port, 
      n_3202, n_3203, n_3204 : std_logic;

begin
   nextA <= ( nextA_63_port, nextA_62_port, nextA_61_port, nextA_60_port, 
      nextA_59_port, nextA_58_port, nextA_57_port, nextA_56_port, nextA_55_port
      , nextA_54_port, nextA_53_port, nextA_52_port, nextA_51_port, 
      nextA_50_port, nextA_49_port, nextA_48_port, nextA_47_port, nextA_46_port
      , nextA_45_port, nextA_44_port, nextA_43_port, nextA_42_port, 
      nextA_41_port, nextA_40_port, nextA_39_port, nextA_38_port, nextA_37_port
      , nextA_36_port, nextA_35_port, nextA_34_port, nextA_33_port, 
      nextA_32_port, nextA_31_port, nextA_30_port, nextA_29_port, nextA_28_port
      , nextA_27_port, nextA_26_port, nextA_25_port, nextA_24_port, 
      nextA_23_port, nextA_22_port, nextA_21_port, nextA_20_port, nextA_19_port
      , nextA_18_port, nextA_17_port, nextA_16_port, nextA_15_port, 
      nextA_14_port, nextA_13_port, nextA_12_port, nextA_11_port, nextA_10_port
      , nextA_9_port, nextA_8_port, nextA_7_port, nextA_6_port, nextA_5_port, 
      nextA_4_port, nextA_3_port, nextA_2_port, nextA_1_port, nextA_0_port );
   
   X_Logic0_port <= '0';
   nextA_0_port <= '0';
   encoder_1 : encoder_N64_RADIX3_10 port map( X(2) => encoderIn(2), X(1) => 
                           encoderIn(1), X(0) => encoderIn(0), Z(2) => 
                           encoder_to_mux_2_port, Z(1) => encoder_to_mux_1_port
                           , Z(0) => encoder_to_mux_0_port);
   ShiftnCompl_1 : ShiftnCompl_N64_10 port map( plusA(63) => prevA(63), 
                           plusA(62) => prevA(62), plusA(61) => prevA(61), 
                           plusA(60) => prevA(60), plusA(59) => prevA(59), 
                           plusA(58) => prevA(58), plusA(57) => prevA(57), 
                           plusA(56) => prevA(56), plusA(55) => prevA(55), 
                           plusA(54) => prevA(54), plusA(53) => prevA(53), 
                           plusA(52) => prevA(52), plusA(51) => prevA(51), 
                           plusA(50) => prevA(50), plusA(49) => prevA(49), 
                           plusA(48) => prevA(48), plusA(47) => prevA(47), 
                           plusA(46) => prevA(46), plusA(45) => prevA(45), 
                           plusA(44) => prevA(44), plusA(43) => prevA(43), 
                           plusA(42) => prevA(42), plusA(41) => prevA(41), 
                           plusA(40) => prevA(40), plusA(39) => prevA(39), 
                           plusA(38) => prevA(38), plusA(37) => prevA(37), 
                           plusA(36) => prevA(36), plusA(35) => prevA(35), 
                           plusA(34) => prevA(34), plusA(33) => prevA(33), 
                           plusA(32) => prevA(32), plusA(31) => prevA(31), 
                           plusA(30) => prevA(30), plusA(29) => prevA(29), 
                           plusA(28) => prevA(28), plusA(27) => prevA(27), 
                           plusA(26) => prevA(26), plusA(25) => prevA(25), 
                           plusA(24) => prevA(24), plusA(23) => prevA(23), 
                           plusA(22) => prevA(22), plusA(21) => prevA(21), 
                           plusA(20) => prevA(20), plusA(19) => prevA(19), 
                           plusA(18) => prevA(18), plusA(17) => prevA(17), 
                           plusA(16) => prevA(16), plusA(15) => prevA(15), 
                           plusA(14) => prevA(14), plusA(13) => prevA(13), 
                           plusA(12) => prevA(12), plusA(11) => prevA(11), 
                           plusA(10) => prevA(10), plusA(9) => prevA(9), 
                           plusA(8) => prevA(8), plusA(7) => prevA(7), plusA(6)
                           => prevA(6), plusA(5) => prevA(5), plusA(4) => 
                           prevA(4), plusA(3) => prevA(3), plusA(2) => prevA(2)
                           , plusA(1) => prevA(1), plusA(0) => prevA(0), 
                           plus2A_out(63) => plus2A_s_63_port, plus2A_out(62) 
                           => plus2A_s_62_port, plus2A_out(61) => 
                           plus2A_s_61_port, plus2A_out(60) => plus2A_s_60_port
                           , plus2A_out(59) => plus2A_s_59_port, plus2A_out(58)
                           => plus2A_s_58_port, plus2A_out(57) => 
                           plus2A_s_57_port, plus2A_out(56) => plus2A_s_56_port
                           , plus2A_out(55) => plus2A_s_55_port, plus2A_out(54)
                           => plus2A_s_54_port, plus2A_out(53) => 
                           plus2A_s_53_port, plus2A_out(52) => plus2A_s_52_port
                           , plus2A_out(51) => plus2A_s_51_port, plus2A_out(50)
                           => plus2A_s_50_port, plus2A_out(49) => 
                           plus2A_s_49_port, plus2A_out(48) => plus2A_s_48_port
                           , plus2A_out(47) => plus2A_s_47_port, plus2A_out(46)
                           => plus2A_s_46_port, plus2A_out(45) => 
                           plus2A_s_45_port, plus2A_out(44) => plus2A_s_44_port
                           , plus2A_out(43) => plus2A_s_43_port, plus2A_out(42)
                           => plus2A_s_42_port, plus2A_out(41) => 
                           plus2A_s_41_port, plus2A_out(40) => plus2A_s_40_port
                           , plus2A_out(39) => plus2A_s_39_port, plus2A_out(38)
                           => plus2A_s_38_port, plus2A_out(37) => 
                           plus2A_s_37_port, plus2A_out(36) => plus2A_s_36_port
                           , plus2A_out(35) => plus2A_s_35_port, plus2A_out(34)
                           => plus2A_s_34_port, plus2A_out(33) => 
                           plus2A_s_33_port, plus2A_out(32) => plus2A_s_32_port
                           , plus2A_out(31) => plus2A_s_31_port, plus2A_out(30)
                           => plus2A_s_30_port, plus2A_out(29) => 
                           plus2A_s_29_port, plus2A_out(28) => plus2A_s_28_port
                           , plus2A_out(27) => plus2A_s_27_port, plus2A_out(26)
                           => plus2A_s_26_port, plus2A_out(25) => 
                           plus2A_s_25_port, plus2A_out(24) => plus2A_s_24_port
                           , plus2A_out(23) => plus2A_s_23_port, plus2A_out(22)
                           => plus2A_s_22_port, plus2A_out(21) => 
                           plus2A_s_21_port, plus2A_out(20) => plus2A_s_20_port
                           , plus2A_out(19) => plus2A_s_19_port, plus2A_out(18)
                           => plus2A_s_18_port, plus2A_out(17) => 
                           plus2A_s_17_port, plus2A_out(16) => plus2A_s_16_port
                           , plus2A_out(15) => plus2A_s_15_port, plus2A_out(14)
                           => plus2A_s_14_port, plus2A_out(13) => 
                           plus2A_s_13_port, plus2A_out(12) => plus2A_s_12_port
                           , plus2A_out(11) => plus2A_s_11_port, plus2A_out(10)
                           => plus2A_s_10_port, plus2A_out(9) => 
                           plus2A_s_9_port, plus2A_out(8) => plus2A_s_8_port, 
                           plus2A_out(7) => plus2A_s_7_port, plus2A_out(6) => 
                           plus2A_s_6_port, plus2A_out(5) => plus2A_s_5_port, 
                           plus2A_out(4) => plus2A_s_4_port, plus2A_out(3) => 
                           plus2A_s_3_port, plus2A_out(2) => plus2A_s_2_port, 
                           plus2A_out(1) => plus2A_s_1_port, plus2A_out(0) => 
                           n_3202, minus2A_out(63) => minus2A_s_63_port, 
                           minus2A_out(62) => minus2A_s_62_port, 
                           minus2A_out(61) => minus2A_s_61_port, 
                           minus2A_out(60) => minus2A_s_60_port, 
                           minus2A_out(59) => minus2A_s_59_port, 
                           minus2A_out(58) => minus2A_s_58_port, 
                           minus2A_out(57) => minus2A_s_57_port, 
                           minus2A_out(56) => minus2A_s_56_port, 
                           minus2A_out(55) => minus2A_s_55_port, 
                           minus2A_out(54) => minus2A_s_54_port, 
                           minus2A_out(53) => minus2A_s_53_port, 
                           minus2A_out(52) => minus2A_s_52_port, 
                           minus2A_out(51) => minus2A_s_51_port, 
                           minus2A_out(50) => minus2A_s_50_port, 
                           minus2A_out(49) => minus2A_s_49_port, 
                           minus2A_out(48) => minus2A_s_48_port, 
                           minus2A_out(47) => minus2A_s_47_port, 
                           minus2A_out(46) => minus2A_s_46_port, 
                           minus2A_out(45) => minus2A_s_45_port, 
                           minus2A_out(44) => minus2A_s_44_port, 
                           minus2A_out(43) => minus2A_s_43_port, 
                           minus2A_out(42) => minus2A_s_42_port, 
                           minus2A_out(41) => minus2A_s_41_port, 
                           minus2A_out(40) => minus2A_s_40_port, 
                           minus2A_out(39) => minus2A_s_39_port, 
                           minus2A_out(38) => minus2A_s_38_port, 
                           minus2A_out(37) => minus2A_s_37_port, 
                           minus2A_out(36) => minus2A_s_36_port, 
                           minus2A_out(35) => minus2A_s_35_port, 
                           minus2A_out(34) => minus2A_s_34_port, 
                           minus2A_out(33) => minus2A_s_33_port, 
                           minus2A_out(32) => minus2A_s_32_port, 
                           minus2A_out(31) => minus2A_s_31_port, 
                           minus2A_out(30) => minus2A_s_30_port, 
                           minus2A_out(29) => minus2A_s_29_port, 
                           minus2A_out(28) => minus2A_s_28_port, 
                           minus2A_out(27) => minus2A_s_27_port, 
                           minus2A_out(26) => minus2A_s_26_port, 
                           minus2A_out(25) => minus2A_s_25_port, 
                           minus2A_out(24) => minus2A_s_24_port, 
                           minus2A_out(23) => minus2A_s_23_port, 
                           minus2A_out(22) => minus2A_s_22_port, 
                           minus2A_out(21) => minus2A_s_21_port, 
                           minus2A_out(20) => minus2A_s_20_port, 
                           minus2A_out(19) => minus2A_s_19_port, 
                           minus2A_out(18) => minus2A_s_18_port, 
                           minus2A_out(17) => minus2A_s_17_port, 
                           minus2A_out(16) => minus2A_s_16_port, 
                           minus2A_out(15) => minus2A_s_15_port, 
                           minus2A_out(14) => minus2A_s_14_port, 
                           minus2A_out(13) => minus2A_s_13_port, 
                           minus2A_out(12) => minus2A_s_12_port, 
                           minus2A_out(11) => minus2A_s_11_port, 
                           minus2A_out(10) => minus2A_s_10_port, minus2A_out(9)
                           => minus2A_s_9_port, minus2A_out(8) => 
                           minus2A_s_8_port, minus2A_out(7) => minus2A_s_7_port
                           , minus2A_out(6) => minus2A_s_6_port, minus2A_out(5)
                           => minus2A_s_5_port, minus2A_out(4) => 
                           minus2A_s_4_port, minus2A_out(3) => minus2A_s_3_port
                           , minus2A_out(2) => minus2A_s_2_port, minus2A_out(1)
                           => minus2A_s_1_port, minus2A_out(0) => 
                           minus2A_s_0_port, plus4A_out(63) => nextA_63_port, 
                           plus4A_out(62) => nextA_62_port, plus4A_out(61) => 
                           nextA_61_port, plus4A_out(60) => nextA_60_port, 
                           plus4A_out(59) => nextA_59_port, plus4A_out(58) => 
                           nextA_58_port, plus4A_out(57) => n3, plus4A_out(56) 
                           => nextA_56_port, plus4A_out(55) => nextA_55_port, 
                           plus4A_out(54) => nextA_54_port, plus4A_out(53) => 
                           nextA_53_port, plus4A_out(52) => nextA_52_port, 
                           plus4A_out(51) => nextA_51_port, plus4A_out(50) => 
                           nextA_50_port, plus4A_out(49) => nextA_49_port, 
                           plus4A_out(48) => nextA_48_port, plus4A_out(47) => 
                           nextA_47_port, plus4A_out(46) => nextA_46_port, 
                           plus4A_out(45) => nextA_45_port, plus4A_out(44) => 
                           nextA_44_port, plus4A_out(43) => nextA_43_port, 
                           plus4A_out(42) => nextA_42_port, plus4A_out(41) => 
                           nextA_41_port, plus4A_out(40) => nextA_40_port, 
                           plus4A_out(39) => nextA_39_port, plus4A_out(38) => 
                           nextA_38_port, plus4A_out(37) => nextA_37_port, 
                           plus4A_out(36) => nextA_36_port, plus4A_out(35) => 
                           nextA_35_port, plus4A_out(34) => nextA_34_port, 
                           plus4A_out(33) => nextA_33_port, plus4A_out(32) => 
                           nextA_32_port, plus4A_out(31) => nextA_31_port, 
                           plus4A_out(30) => nextA_30_port, plus4A_out(29) => 
                           nextA_29_port, plus4A_out(28) => nextA_28_port, 
                           plus4A_out(27) => nextA_27_port, plus4A_out(26) => 
                           nextA_26_port, plus4A_out(25) => nextA_25_port, 
                           plus4A_out(24) => nextA_24_port, plus4A_out(23) => 
                           nextA_23_port, plus4A_out(22) => nextA_22_port, 
                           plus4A_out(21) => nextA_21_port, plus4A_out(20) => 
                           nextA_20_port, plus4A_out(19) => nextA_19_port, 
                           plus4A_out(18) => nextA_18_port, plus4A_out(17) => 
                           nextA_17_port, plus4A_out(16) => nextA_16_port, 
                           plus4A_out(15) => nextA_15_port, plus4A_out(14) => 
                           nextA_14_port, plus4A_out(13) => nextA_13_port, 
                           plus4A_out(12) => nextA_12_port, plus4A_out(11) => 
                           nextA_11_port, plus4A_out(10) => nextA_10_port, 
                           plus4A_out(9) => nextA_9_port, plus4A_out(8) => 
                           nextA_8_port, plus4A_out(7) => nextA_7_port, 
                           plus4A_out(6) => nextA_6_port, plus4A_out(5) => 
                           nextA_5_port, plus4A_out(4) => nextA_4_port, 
                           plus4A_out(3) => nextA_3_port, plus4A_out(2) => 
                           nextA_2_port, plus4A_out(1) => nextA_1_port, 
                           plus4A_out(0) => n_3203, minus4A_out(63) => 
                           minus4A_s_63_port, minus4A_out(62) => 
                           minus4A_s_62_port, minus4A_out(61) => 
                           minus4A_s_61_port, minus4A_out(60) => 
                           minus4A_s_60_port, minus4A_out(59) => 
                           minus4A_s_59_port, minus4A_out(58) => 
                           minus4A_s_58_port, minus4A_out(57) => 
                           minus4A_s_57_port, minus4A_out(56) => 
                           minus4A_s_56_port, minus4A_out(55) => 
                           minus4A_s_55_port, minus4A_out(54) => 
                           minus4A_s_54_port, minus4A_out(53) => 
                           minus4A_s_53_port, minus4A_out(52) => 
                           minus4A_s_52_port, minus4A_out(51) => 
                           minus4A_s_51_port, minus4A_out(50) => 
                           minus4A_s_50_port, minus4A_out(49) => 
                           minus4A_s_49_port, minus4A_out(48) => 
                           minus4A_s_48_port, minus4A_out(47) => 
                           minus4A_s_47_port, minus4A_out(46) => 
                           minus4A_s_46_port, minus4A_out(45) => 
                           minus4A_s_45_port, minus4A_out(44) => 
                           minus4A_s_44_port, minus4A_out(43) => 
                           minus4A_s_43_port, minus4A_out(42) => 
                           minus4A_s_42_port, minus4A_out(41) => 
                           minus4A_s_41_port, minus4A_out(40) => 
                           minus4A_s_40_port, minus4A_out(39) => 
                           minus4A_s_39_port, minus4A_out(38) => 
                           minus4A_s_38_port, minus4A_out(37) => 
                           minus4A_s_37_port, minus4A_out(36) => 
                           minus4A_s_36_port, minus4A_out(35) => 
                           minus4A_s_35_port, minus4A_out(34) => 
                           minus4A_s_34_port, minus4A_out(33) => 
                           minus4A_s_33_port, minus4A_out(32) => 
                           minus4A_s_32_port, minus4A_out(31) => 
                           minus4A_s_31_port, minus4A_out(30) => 
                           minus4A_s_30_port, minus4A_out(29) => 
                           minus4A_s_29_port, minus4A_out(28) => 
                           minus4A_s_28_port, minus4A_out(27) => 
                           minus4A_s_27_port, minus4A_out(26) => 
                           minus4A_s_26_port, minus4A_out(25) => 
                           minus4A_s_25_port, minus4A_out(24) => 
                           minus4A_s_24_port, minus4A_out(23) => 
                           minus4A_s_23_port, minus4A_out(22) => 
                           minus4A_s_22_port, minus4A_out(21) => 
                           minus4A_s_21_port, minus4A_out(20) => 
                           minus4A_s_20_port, minus4A_out(19) => 
                           minus4A_s_19_port, minus4A_out(18) => 
                           minus4A_s_18_port, minus4A_out(17) => 
                           minus4A_s_17_port, minus4A_out(16) => 
                           minus4A_s_16_port, minus4A_out(15) => 
                           minus4A_s_15_port, minus4A_out(14) => 
                           minus4A_s_14_port, minus4A_out(13) => 
                           minus4A_s_13_port, minus4A_out(12) => 
                           minus4A_s_12_port, minus4A_out(11) => 
                           minus4A_s_11_port, minus4A_out(10) => 
                           minus4A_s_10_port, minus4A_out(9) => 
                           minus4A_s_9_port, minus4A_out(8) => minus4A_s_8_port
                           , minus4A_out(7) => minus4A_s_7_port, minus4A_out(6)
                           => minus4A_s_6_port, minus4A_out(5) => 
                           minus4A_s_5_port, minus4A_out(4) => minus4A_s_4_port
                           , minus4A_out(3) => minus4A_s_3_port, minus4A_out(2)
                           => minus4A_s_2_port, minus4A_out(1) => 
                           minus4A_s_1_port, minus4A_out(0) => minus4A_s_0_port
                           );
   mux_1 : MUX_GENERIC_N64_RADIX3_10 port map( plusA(63) => plus2A_s_63_port, 
                           plusA(62) => plus2A_s_62_port, plusA(61) => 
                           plus2A_s_61_port, plusA(60) => plus2A_s_60_port, 
                           plusA(59) => plus2A_s_59_port, plusA(58) => 
                           plus2A_s_58_port, plusA(57) => plus2A_s_57_port, 
                           plusA(56) => plus2A_s_56_port, plusA(55) => 
                           plus2A_s_55_port, plusA(54) => plus2A_s_54_port, 
                           plusA(53) => plus2A_s_53_port, plusA(52) => 
                           plus2A_s_52_port, plusA(51) => plus2A_s_51_port, 
                           plusA(50) => plus2A_s_50_port, plusA(49) => 
                           plus2A_s_49_port, plusA(48) => plus2A_s_48_port, 
                           plusA(47) => plus2A_s_47_port, plusA(46) => 
                           plus2A_s_46_port, plusA(45) => plus2A_s_45_port, 
                           plusA(44) => plus2A_s_44_port, plusA(43) => 
                           plus2A_s_43_port, plusA(42) => plus2A_s_42_port, 
                           plusA(41) => plus2A_s_41_port, plusA(40) => 
                           plus2A_s_40_port, plusA(39) => plus2A_s_39_port, 
                           plusA(38) => plus2A_s_38_port, plusA(37) => 
                           plus2A_s_37_port, plusA(36) => plus2A_s_36_port, 
                           plusA(35) => plus2A_s_35_port, plusA(34) => 
                           plus2A_s_34_port, plusA(33) => plus2A_s_33_port, 
                           plusA(32) => plus2A_s_32_port, plusA(31) => 
                           plus2A_s_31_port, plusA(30) => plus2A_s_30_port, 
                           plusA(29) => plus2A_s_29_port, plusA(28) => 
                           plus2A_s_28_port, plusA(27) => plus2A_s_27_port, 
                           plusA(26) => plus2A_s_26_port, plusA(25) => 
                           plus2A_s_25_port, plusA(24) => plus2A_s_24_port, 
                           plusA(23) => plus2A_s_23_port, plusA(22) => 
                           plus2A_s_22_port, plusA(21) => plus2A_s_21_port, 
                           plusA(20) => plus2A_s_20_port, plusA(19) => 
                           plus2A_s_19_port, plusA(18) => plus2A_s_18_port, 
                           plusA(17) => plus2A_s_17_port, plusA(16) => 
                           plus2A_s_16_port, plusA(15) => plus2A_s_15_port, 
                           plusA(14) => plus2A_s_14_port, plusA(13) => 
                           plus2A_s_13_port, plusA(12) => plus2A_s_12_port, 
                           plusA(11) => plus2A_s_11_port, plusA(10) => 
                           plus2A_s_10_port, plusA(9) => plus2A_s_9_port, 
                           plusA(8) => plus2A_s_8_port, plusA(7) => 
                           plus2A_s_7_port, plusA(6) => plus2A_s_6_port, 
                           plusA(5) => plus2A_s_5_port, plusA(4) => 
                           plus2A_s_4_port, plusA(3) => plus2A_s_3_port, 
                           plusA(2) => plus2A_s_2_port, plusA(1) => 
                           plus2A_s_1_port, plusA(0) => nextA_0_port, 
                           minusA(63) => minus2A_s_63_port, minusA(62) => 
                           minus2A_s_62_port, minusA(61) => minus2A_s_61_port, 
                           minusA(60) => minus2A_s_60_port, minusA(59) => 
                           minus2A_s_59_port, minusA(58) => minus2A_s_58_port, 
                           minusA(57) => minus2A_s_57_port, minusA(56) => 
                           minus2A_s_56_port, minusA(55) => minus2A_s_55_port, 
                           minusA(54) => minus2A_s_54_port, minusA(53) => 
                           minus2A_s_53_port, minusA(52) => minus2A_s_52_port, 
                           minusA(51) => minus2A_s_51_port, minusA(50) => 
                           minus2A_s_50_port, minusA(49) => minus2A_s_49_port, 
                           minusA(48) => minus2A_s_48_port, minusA(47) => 
                           minus2A_s_47_port, minusA(46) => minus2A_s_46_port, 
                           minusA(45) => minus2A_s_45_port, minusA(44) => 
                           minus2A_s_44_port, minusA(43) => minus2A_s_43_port, 
                           minusA(42) => minus2A_s_42_port, minusA(41) => 
                           minus2A_s_41_port, minusA(40) => minus2A_s_40_port, 
                           minusA(39) => minus2A_s_39_port, minusA(38) => 
                           minus2A_s_38_port, minusA(37) => minus2A_s_37_port, 
                           minusA(36) => minus2A_s_36_port, minusA(35) => 
                           minus2A_s_35_port, minusA(34) => minus2A_s_34_port, 
                           minusA(33) => minus2A_s_33_port, minusA(32) => 
                           minus2A_s_32_port, minusA(31) => minus2A_s_31_port, 
                           minusA(30) => minus2A_s_30_port, minusA(29) => 
                           minus2A_s_29_port, minusA(28) => minus2A_s_28_port, 
                           minusA(27) => minus2A_s_27_port, minusA(26) => 
                           minus2A_s_26_port, minusA(25) => minus2A_s_25_port, 
                           minusA(24) => minus2A_s_24_port, minusA(23) => 
                           minus2A_s_23_port, minusA(22) => minus2A_s_22_port, 
                           minusA(21) => minus2A_s_21_port, minusA(20) => 
                           minus2A_s_20_port, minusA(19) => minus2A_s_19_port, 
                           minusA(18) => minus2A_s_18_port, minusA(17) => 
                           minus2A_s_17_port, minusA(16) => minus2A_s_16_port, 
                           minusA(15) => minus2A_s_15_port, minusA(14) => 
                           minus2A_s_14_port, minusA(13) => minus2A_s_13_port, 
                           minusA(12) => minus2A_s_12_port, minusA(11) => 
                           minus2A_s_11_port, minusA(10) => minus2A_s_10_port, 
                           minusA(9) => minus2A_s_9_port, minusA(8) => 
                           minus2A_s_8_port, minusA(7) => minus2A_s_7_port, 
                           minusA(6) => minus2A_s_6_port, minusA(5) => 
                           minus2A_s_5_port, minusA(4) => minus2A_s_4_port, 
                           minusA(3) => minus2A_s_3_port, minusA(2) => 
                           minus2A_s_2_port, minusA(1) => minus2A_s_1_port, 
                           minusA(0) => minus2A_s_0_port, plus2A(63) => 
                           nextA_63_port, plus2A(62) => nextA_62_port, 
                           plus2A(61) => nextA_61_port, plus2A(60) => 
                           nextA_60_port, plus2A(59) => nextA_59_port, 
                           plus2A(58) => nextA_58_port, plus2A(57) => 
                           nextA_57_port, plus2A(56) => nextA_56_port, 
                           plus2A(55) => nextA_55_port, plus2A(54) => 
                           nextA_54_port, plus2A(53) => nextA_53_port, 
                           plus2A(52) => nextA_52_port, plus2A(51) => 
                           nextA_51_port, plus2A(50) => nextA_50_port, 
                           plus2A(49) => nextA_49_port, plus2A(48) => 
                           nextA_48_port, plus2A(47) => nextA_47_port, 
                           plus2A(46) => nextA_46_port, plus2A(45) => 
                           nextA_45_port, plus2A(44) => nextA_44_port, 
                           plus2A(43) => nextA_43_port, plus2A(42) => 
                           nextA_42_port, plus2A(41) => nextA_41_port, 
                           plus2A(40) => nextA_40_port, plus2A(39) => 
                           nextA_39_port, plus2A(38) => nextA_38_port, 
                           plus2A(37) => nextA_37_port, plus2A(36) => 
                           nextA_36_port, plus2A(35) => nextA_35_port, 
                           plus2A(34) => nextA_34_port, plus2A(33) => 
                           nextA_33_port, plus2A(32) => nextA_32_port, 
                           plus2A(31) => nextA_31_port, plus2A(30) => 
                           nextA_30_port, plus2A(29) => nextA_29_port, 
                           plus2A(28) => nextA_28_port, plus2A(27) => 
                           nextA_27_port, plus2A(26) => nextA_26_port, 
                           plus2A(25) => nextA_25_port, plus2A(24) => 
                           nextA_24_port, plus2A(23) => nextA_23_port, 
                           plus2A(22) => nextA_22_port, plus2A(21) => 
                           nextA_21_port, plus2A(20) => nextA_20_port, 
                           plus2A(19) => nextA_19_port, plus2A(18) => 
                           nextA_18_port, plus2A(17) => nextA_17_port, 
                           plus2A(16) => nextA_16_port, plus2A(15) => 
                           nextA_15_port, plus2A(14) => nextA_14_port, 
                           plus2A(13) => nextA_13_port, plus2A(12) => 
                           nextA_12_port, plus2A(11) => nextA_11_port, 
                           plus2A(10) => nextA_10_port, plus2A(9) => 
                           nextA_9_port, plus2A(8) => nextA_8_port, plus2A(7) 
                           => nextA_7_port, plus2A(6) => nextA_6_port, 
                           plus2A(5) => nextA_5_port, plus2A(4) => nextA_4_port
                           , plus2A(3) => nextA_3_port, plus2A(2) => 
                           nextA_2_port, plus2A(1) => nextA_1_port, plus2A(0) 
                           => nextA_0_port, minus2A(63) => minus4A_s_63_port, 
                           minus2A(62) => minus4A_s_62_port, minus2A(61) => 
                           minus4A_s_61_port, minus2A(60) => minus4A_s_60_port,
                           minus2A(59) => minus4A_s_59_port, minus2A(58) => 
                           minus4A_s_58_port, minus2A(57) => minus4A_s_57_port,
                           minus2A(56) => minus4A_s_56_port, minus2A(55) => 
                           minus4A_s_55_port, minus2A(54) => minus4A_s_54_port,
                           minus2A(53) => minus4A_s_53_port, minus2A(52) => 
                           minus4A_s_52_port, minus2A(51) => minus4A_s_51_port,
                           minus2A(50) => minus4A_s_50_port, minus2A(49) => 
                           minus4A_s_49_port, minus2A(48) => minus4A_s_48_port,
                           minus2A(47) => minus4A_s_47_port, minus2A(46) => 
                           minus4A_s_46_port, minus2A(45) => minus4A_s_45_port,
                           minus2A(44) => minus4A_s_44_port, minus2A(43) => 
                           minus4A_s_43_port, minus2A(42) => minus4A_s_42_port,
                           minus2A(41) => minus4A_s_41_port, minus2A(40) => 
                           minus4A_s_40_port, minus2A(39) => minus4A_s_39_port,
                           minus2A(38) => minus4A_s_38_port, minus2A(37) => 
                           minus4A_s_37_port, minus2A(36) => minus4A_s_36_port,
                           minus2A(35) => minus4A_s_35_port, minus2A(34) => 
                           minus4A_s_34_port, minus2A(33) => minus4A_s_33_port,
                           minus2A(32) => minus4A_s_32_port, minus2A(31) => 
                           minus4A_s_31_port, minus2A(30) => minus4A_s_30_port,
                           minus2A(29) => minus4A_s_29_port, minus2A(28) => 
                           minus4A_s_28_port, minus2A(27) => minus4A_s_27_port,
                           minus2A(26) => minus4A_s_26_port, minus2A(25) => 
                           minus4A_s_25_port, minus2A(24) => minus4A_s_24_port,
                           minus2A(23) => minus4A_s_23_port, minus2A(22) => 
                           minus4A_s_22_port, minus2A(21) => minus4A_s_21_port,
                           minus2A(20) => minus4A_s_20_port, minus2A(19) => 
                           minus4A_s_19_port, minus2A(18) => minus4A_s_18_port,
                           minus2A(17) => minus4A_s_17_port, minus2A(16) => 
                           minus4A_s_16_port, minus2A(15) => minus4A_s_15_port,
                           minus2A(14) => minus4A_s_14_port, minus2A(13) => 
                           minus4A_s_13_port, minus2A(12) => minus4A_s_12_port,
                           minus2A(11) => minus4A_s_11_port, minus2A(10) => 
                           minus4A_s_10_port, minus2A(9) => minus4A_s_9_port, 
                           minus2A(8) => minus4A_s_8_port, minus2A(7) => 
                           minus4A_s_7_port, minus2A(6) => minus4A_s_6_port, 
                           minus2A(5) => minus4A_s_5_port, minus2A(4) => 
                           minus4A_s_4_port, minus2A(3) => minus4A_s_3_port, 
                           minus2A(2) => minus4A_s_2_port, minus2A(1) => 
                           minus4A_s_1_port, minus2A(0) => minus4A_s_0_port, 
                           SEL(2) => encoder_to_mux_2_port, SEL(1) => 
                           encoder_to_mux_1_port, SEL(0) => 
                           encoder_to_mux_0_port, Y(63) => mux_to_adder_63_port
                           , Y(62) => mux_to_adder_62_port, Y(61) => 
                           mux_to_adder_61_port, Y(60) => mux_to_adder_60_port,
                           Y(59) => mux_to_adder_59_port, Y(58) => 
                           mux_to_adder_58_port, Y(57) => mux_to_adder_57_port,
                           Y(56) => mux_to_adder_56_port, Y(55) => 
                           mux_to_adder_55_port, Y(54) => mux_to_adder_54_port,
                           Y(53) => mux_to_adder_53_port, Y(52) => 
                           mux_to_adder_52_port, Y(51) => mux_to_adder_51_port,
                           Y(50) => mux_to_adder_50_port, Y(49) => 
                           mux_to_adder_49_port, Y(48) => mux_to_adder_48_port,
                           Y(47) => mux_to_adder_47_port, Y(46) => 
                           mux_to_adder_46_port, Y(45) => mux_to_adder_45_port,
                           Y(44) => mux_to_adder_44_port, Y(43) => 
                           mux_to_adder_43_port, Y(42) => mux_to_adder_42_port,
                           Y(41) => mux_to_adder_41_port, Y(40) => 
                           mux_to_adder_40_port, Y(39) => mux_to_adder_39_port,
                           Y(38) => mux_to_adder_38_port, Y(37) => 
                           mux_to_adder_37_port, Y(36) => mux_to_adder_36_port,
                           Y(35) => mux_to_adder_35_port, Y(34) => 
                           mux_to_adder_34_port, Y(33) => mux_to_adder_33_port,
                           Y(32) => mux_to_adder_32_port, Y(31) => 
                           mux_to_adder_31_port, Y(30) => mux_to_adder_30_port,
                           Y(29) => mux_to_adder_29_port, Y(28) => 
                           mux_to_adder_28_port, Y(27) => mux_to_adder_27_port,
                           Y(26) => mux_to_adder_26_port, Y(25) => 
                           mux_to_adder_25_port, Y(24) => mux_to_adder_24_port,
                           Y(23) => mux_to_adder_23_port, Y(22) => 
                           mux_to_adder_22_port, Y(21) => mux_to_adder_21_port,
                           Y(20) => mux_to_adder_20_port, Y(19) => 
                           mux_to_adder_19_port, Y(18) => mux_to_adder_18_port,
                           Y(17) => mux_to_adder_17_port, Y(16) => 
                           mux_to_adder_16_port, Y(15) => mux_to_adder_15_port,
                           Y(14) => mux_to_adder_14_port, Y(13) => 
                           mux_to_adder_13_port, Y(12) => mux_to_adder_12_port,
                           Y(11) => mux_to_adder_11_port, Y(10) => 
                           mux_to_adder_10_port, Y(9) => mux_to_adder_9_port, 
                           Y(8) => mux_to_adder_8_port, Y(7) => 
                           mux_to_adder_7_port, Y(6) => mux_to_adder_6_port, 
                           Y(5) => mux_to_adder_5_port, Y(4) => 
                           mux_to_adder_4_port, Y(3) => mux_to_adder_3_port, 
                           Y(2) => mux_to_adder_2_port, Y(1) => 
                           mux_to_adder_1_port, Y(0) => mux_to_adder_0_port);
   rca_1 : RCA_N64_10 port map( A(63) => mux_to_adder_63_port, A(62) => 
                           mux_to_adder_62_port, A(61) => mux_to_adder_61_port,
                           A(60) => mux_to_adder_60_port, A(59) => 
                           mux_to_adder_59_port, A(58) => mux_to_adder_58_port,
                           A(57) => mux_to_adder_57_port, A(56) => 
                           mux_to_adder_56_port, A(55) => mux_to_adder_55_port,
                           A(54) => mux_to_adder_54_port, A(53) => 
                           mux_to_adder_53_port, A(52) => mux_to_adder_52_port,
                           A(51) => mux_to_adder_51_port, A(50) => 
                           mux_to_adder_50_port, A(49) => mux_to_adder_49_port,
                           A(48) => mux_to_adder_48_port, A(47) => 
                           mux_to_adder_47_port, A(46) => mux_to_adder_46_port,
                           A(45) => mux_to_adder_45_port, A(44) => 
                           mux_to_adder_44_port, A(43) => mux_to_adder_43_port,
                           A(42) => mux_to_adder_42_port, A(41) => 
                           mux_to_adder_41_port, A(40) => mux_to_adder_40_port,
                           A(39) => mux_to_adder_39_port, A(38) => 
                           mux_to_adder_38_port, A(37) => mux_to_adder_37_port,
                           A(36) => mux_to_adder_36_port, A(35) => 
                           mux_to_adder_35_port, A(34) => mux_to_adder_34_port,
                           A(33) => mux_to_adder_33_port, A(32) => 
                           mux_to_adder_32_port, A(31) => mux_to_adder_31_port,
                           A(30) => mux_to_adder_30_port, A(29) => 
                           mux_to_adder_29_port, A(28) => mux_to_adder_28_port,
                           A(27) => mux_to_adder_27_port, A(26) => 
                           mux_to_adder_26_port, A(25) => mux_to_adder_25_port,
                           A(24) => mux_to_adder_24_port, A(23) => 
                           mux_to_adder_23_port, A(22) => mux_to_adder_22_port,
                           A(21) => mux_to_adder_21_port, A(20) => 
                           mux_to_adder_20_port, A(19) => mux_to_adder_19_port,
                           A(18) => mux_to_adder_18_port, A(17) => 
                           mux_to_adder_17_port, A(16) => mux_to_adder_16_port,
                           A(15) => mux_to_adder_15_port, A(14) => 
                           mux_to_adder_14_port, A(13) => mux_to_adder_13_port,
                           A(12) => mux_to_adder_12_port, A(11) => 
                           mux_to_adder_11_port, A(10) => mux_to_adder_10_port,
                           A(9) => mux_to_adder_9_port, A(8) => 
                           mux_to_adder_8_port, A(7) => mux_to_adder_7_port, 
                           A(6) => mux_to_adder_6_port, A(5) => 
                           mux_to_adder_5_port, A(4) => mux_to_adder_4_port, 
                           A(3) => mux_to_adder_3_port, A(2) => 
                           mux_to_adder_2_port, A(1) => mux_to_adder_1_port, 
                           A(0) => mux_to_adder_0_port, B(63) => prevSum(63), 
                           B(62) => prevSum(62), B(61) => prevSum(61), B(60) =>
                           prevSum(60), B(59) => prevSum(59), B(58) => 
                           prevSum(58), B(57) => prevSum(57), B(56) => 
                           prevSum(56), B(55) => prevSum(55), B(54) => 
                           prevSum(54), B(53) => prevSum(53), B(52) => 
                           prevSum(52), B(51) => prevSum(51), B(50) => 
                           prevSum(50), B(49) => prevSum(49), B(48) => 
                           prevSum(48), B(47) => prevSum(47), B(46) => 
                           prevSum(46), B(45) => prevSum(45), B(44) => 
                           prevSum(44), B(43) => prevSum(43), B(42) => 
                           prevSum(42), B(41) => prevSum(41), B(40) => 
                           prevSum(40), B(39) => prevSum(39), B(38) => 
                           prevSum(38), B(37) => prevSum(37), B(36) => 
                           prevSum(36), B(35) => prevSum(35), B(34) => 
                           prevSum(34), B(33) => prevSum(33), B(32) => 
                           prevSum(32), B(31) => prevSum(31), B(30) => 
                           prevSum(30), B(29) => prevSum(29), B(28) => 
                           prevSum(28), B(27) => prevSum(27), B(26) => 
                           prevSum(26), B(25) => prevSum(25), B(24) => 
                           prevSum(24), B(23) => prevSum(23), B(22) => 
                           prevSum(22), B(21) => prevSum(21), B(20) => 
                           prevSum(20), B(19) => prevSum(19), B(18) => 
                           prevSum(18), B(17) => prevSum(17), B(16) => 
                           prevSum(16), B(15) => prevSum(15), B(14) => 
                           prevSum(14), B(13) => prevSum(13), B(12) => 
                           prevSum(12), B(11) => prevSum(11), B(10) => 
                           prevSum(10), B(9) => prevSum(9), B(8) => prevSum(8),
                           B(7) => prevSum(7), B(6) => prevSum(6), B(5) => 
                           prevSum(5), B(4) => prevSum(4), B(3) => prevSum(3), 
                           B(2) => prevSum(2), B(1) => prevSum(1), B(0) => 
                           prevSum(0), Ci => X_Logic0_port, S(63) => 
                           nextSum(63), S(62) => nextSum(62), S(61) => 
                           nextSum(61), S(60) => nextSum(60), S(59) => 
                           nextSum(59), S(58) => nextSum(58), S(57) => 
                           nextSum(57), S(56) => nextSum(56), S(55) => 
                           nextSum(55), S(54) => nextSum(54), S(53) => 
                           nextSum(53), S(52) => nextSum(52), S(51) => 
                           nextSum(51), S(50) => nextSum(50), S(49) => 
                           nextSum(49), S(48) => nextSum(48), S(47) => 
                           nextSum(47), S(46) => nextSum(46), S(45) => 
                           nextSum(45), S(44) => nextSum(44), S(43) => 
                           nextSum(43), S(42) => nextSum(42), S(41) => 
                           nextSum(41), S(40) => nextSum(40), S(39) => 
                           nextSum(39), S(38) => nextSum(38), S(37) => 
                           nextSum(37), S(36) => nextSum(36), S(35) => 
                           nextSum(35), S(34) => nextSum(34), S(33) => 
                           nextSum(33), S(32) => nextSum(32), S(31) => 
                           nextSum(31), S(30) => nextSum(30), S(29) => 
                           nextSum(29), S(28) => nextSum(28), S(27) => 
                           nextSum(27), S(26) => nextSum(26), S(25) => 
                           nextSum(25), S(24) => nextSum(24), S(23) => 
                           nextSum(23), S(22) => nextSum(22), S(21) => 
                           nextSum(21), S(20) => nextSum(20), S(19) => 
                           nextSum(19), S(18) => nextSum(18), S(17) => 
                           nextSum(17), S(16) => nextSum(16), S(15) => 
                           nextSum(15), S(14) => nextSum(14), S(13) => 
                           nextSum(13), S(12) => nextSum(12), S(11) => 
                           nextSum(11), S(10) => nextSum(10), S(9) => 
                           nextSum(9), S(8) => nextSum(8), S(7) => nextSum(7), 
                           S(6) => nextSum(6), S(5) => nextSum(5), S(4) => 
                           nextSum(4), S(3) => nextSum(3), S(2) => nextSum(2), 
                           S(1) => nextSum(1), S(0) => nextSum(0), Co => n_3204
                           );
   U3 : BUF_X1 port map( A => n3, Z => nextA_57_port);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity booth_mul_row_N64_RADIX3_11 is

   port( prevA, prevSum : in std_logic_vector (63 downto 0);  encoderIn : in 
         std_logic_vector (2 downto 0);  nextA, nextSum : out std_logic_vector 
         (63 downto 0));

end booth_mul_row_N64_RADIX3_11;

architecture SYN_struct of booth_mul_row_N64_RADIX3_11 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component RCA_N64_11
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component MUX_GENERIC_N64_RADIX3_11
      port( plusA, minusA, plus2A, minus2A : in std_logic_vector (63 downto 0);
            SEL : in std_logic_vector (2 downto 0);  Y : out std_logic_vector 
            (63 downto 0));
   end component;
   
   component ShiftnCompl_N64_11
      port( plusA : in std_logic_vector (63 downto 0);  plus2A_out, minus2A_out
            , plus4A_out, minus4A_out : out std_logic_vector (63 downto 0));
   end component;
   
   component encoder_N64_RADIX3_11
      port( X : in std_logic_vector (2 downto 0);  Z : out std_logic_vector (2 
            downto 0));
   end component;
   
   signal X_Logic0_port, nextA_63_port, nextA_62_port, nextA_61_port, 
      nextA_60_port, nextA_59_port, nextA_58_port, n3, nextA_56_port, 
      nextA_55_port, nextA_54_port, nextA_53_port, nextA_52_port, nextA_51_port
      , nextA_50_port, nextA_49_port, nextA_48_port, nextA_47_port, 
      nextA_46_port, nextA_45_port, nextA_44_port, nextA_43_port, nextA_42_port
      , nextA_41_port, nextA_40_port, nextA_39_port, nextA_38_port, 
      nextA_37_port, nextA_36_port, nextA_35_port, nextA_34_port, nextA_33_port
      , nextA_32_port, nextA_31_port, nextA_30_port, nextA_29_port, 
      nextA_28_port, nextA_27_port, nextA_26_port, nextA_25_port, nextA_24_port
      , nextA_23_port, nextA_22_port, nextA_21_port, nextA_20_port, 
      nextA_19_port, nextA_18_port, nextA_17_port, nextA_16_port, nextA_15_port
      , nextA_14_port, nextA_13_port, nextA_12_port, nextA_11_port, 
      nextA_10_port, nextA_9_port, nextA_8_port, nextA_7_port, nextA_6_port, 
      nextA_5_port, nextA_4_port, nextA_3_port, nextA_2_port, nextA_1_port, 
      encoder_to_mux_2_port, encoder_to_mux_1_port, encoder_to_mux_0_port, 
      plus2A_s_63_port, plus2A_s_62_port, plus2A_s_61_port, plus2A_s_60_port, 
      plus2A_s_59_port, plus2A_s_58_port, plus2A_s_57_port, plus2A_s_56_port, 
      plus2A_s_55_port, plus2A_s_54_port, plus2A_s_53_port, plus2A_s_52_port, 
      plus2A_s_51_port, plus2A_s_50_port, plus2A_s_49_port, plus2A_s_48_port, 
      plus2A_s_47_port, plus2A_s_46_port, plus2A_s_45_port, plus2A_s_44_port, 
      plus2A_s_43_port, plus2A_s_42_port, plus2A_s_41_port, plus2A_s_40_port, 
      plus2A_s_39_port, plus2A_s_38_port, plus2A_s_37_port, plus2A_s_36_port, 
      plus2A_s_35_port, plus2A_s_34_port, plus2A_s_33_port, plus2A_s_32_port, 
      plus2A_s_31_port, plus2A_s_30_port, plus2A_s_29_port, plus2A_s_28_port, 
      plus2A_s_27_port, plus2A_s_26_port, plus2A_s_25_port, plus2A_s_24_port, 
      plus2A_s_23_port, plus2A_s_22_port, plus2A_s_21_port, plus2A_s_20_port, 
      plus2A_s_19_port, plus2A_s_18_port, plus2A_s_17_port, plus2A_s_16_port, 
      plus2A_s_15_port, plus2A_s_14_port, plus2A_s_13_port, plus2A_s_12_port, 
      plus2A_s_11_port, plus2A_s_10_port, plus2A_s_9_port, plus2A_s_8_port, 
      plus2A_s_7_port, plus2A_s_6_port, plus2A_s_5_port, plus2A_s_4_port, 
      plus2A_s_3_port, plus2A_s_2_port, plus2A_s_1_port, minus2A_s_63_port, 
      minus2A_s_62_port, minus2A_s_61_port, minus2A_s_60_port, 
      minus2A_s_59_port, minus2A_s_58_port, minus2A_s_57_port, 
      minus2A_s_56_port, minus2A_s_55_port, minus2A_s_54_port, 
      minus2A_s_53_port, minus2A_s_52_port, minus2A_s_51_port, 
      minus2A_s_50_port, minus2A_s_49_port, minus2A_s_48_port, 
      minus2A_s_47_port, minus2A_s_46_port, minus2A_s_45_port, 
      minus2A_s_44_port, minus2A_s_43_port, minus2A_s_42_port, 
      minus2A_s_41_port, minus2A_s_40_port, minus2A_s_39_port, 
      minus2A_s_38_port, minus2A_s_37_port, minus2A_s_36_port, 
      minus2A_s_35_port, minus2A_s_34_port, minus2A_s_33_port, 
      minus2A_s_32_port, minus2A_s_31_port, minus2A_s_30_port, 
      minus2A_s_29_port, minus2A_s_28_port, minus2A_s_27_port, 
      minus2A_s_26_port, minus2A_s_25_port, minus2A_s_24_port, 
      minus2A_s_23_port, minus2A_s_22_port, minus2A_s_21_port, 
      minus2A_s_20_port, minus2A_s_19_port, minus2A_s_18_port, 
      minus2A_s_17_port, minus2A_s_16_port, minus2A_s_15_port, 
      minus2A_s_14_port, minus2A_s_13_port, minus2A_s_12_port, 
      minus2A_s_11_port, minus2A_s_10_port, minus2A_s_9_port, minus2A_s_8_port,
      minus2A_s_7_port, minus2A_s_6_port, minus2A_s_5_port, minus2A_s_4_port, 
      minus2A_s_3_port, minus2A_s_2_port, minus2A_s_1_port, minus2A_s_0_port, 
      minus4A_s_63_port, minus4A_s_62_port, minus4A_s_61_port, 
      minus4A_s_60_port, minus4A_s_59_port, minus4A_s_58_port, 
      minus4A_s_57_port, minus4A_s_56_port, minus4A_s_55_port, 
      minus4A_s_54_port, minus4A_s_53_port, minus4A_s_52_port, 
      minus4A_s_51_port, minus4A_s_50_port, minus4A_s_49_port, 
      minus4A_s_48_port, minus4A_s_47_port, minus4A_s_46_port, 
      minus4A_s_45_port, minus4A_s_44_port, minus4A_s_43_port, 
      minus4A_s_42_port, minus4A_s_41_port, minus4A_s_40_port, 
      minus4A_s_39_port, minus4A_s_38_port, minus4A_s_37_port, 
      minus4A_s_36_port, minus4A_s_35_port, minus4A_s_34_port, 
      minus4A_s_33_port, minus4A_s_32_port, minus4A_s_31_port, 
      minus4A_s_30_port, minus4A_s_29_port, minus4A_s_28_port, 
      minus4A_s_27_port, minus4A_s_26_port, minus4A_s_25_port, 
      minus4A_s_24_port, minus4A_s_23_port, minus4A_s_22_port, 
      minus4A_s_21_port, minus4A_s_20_port, minus4A_s_19_port, 
      minus4A_s_18_port, minus4A_s_17_port, minus4A_s_16_port, 
      minus4A_s_15_port, minus4A_s_14_port, minus4A_s_13_port, 
      minus4A_s_12_port, minus4A_s_11_port, minus4A_s_10_port, minus4A_s_9_port
      , minus4A_s_8_port, minus4A_s_7_port, minus4A_s_6_port, minus4A_s_5_port,
      minus4A_s_4_port, minus4A_s_3_port, minus4A_s_2_port, minus4A_s_1_port, 
      minus4A_s_0_port, mux_to_adder_63_port, mux_to_adder_62_port, 
      mux_to_adder_61_port, mux_to_adder_60_port, mux_to_adder_59_port, 
      mux_to_adder_58_port, mux_to_adder_57_port, mux_to_adder_56_port, 
      mux_to_adder_55_port, mux_to_adder_54_port, mux_to_adder_53_port, 
      mux_to_adder_52_port, mux_to_adder_51_port, mux_to_adder_50_port, 
      mux_to_adder_49_port, mux_to_adder_48_port, mux_to_adder_47_port, 
      mux_to_adder_46_port, mux_to_adder_45_port, mux_to_adder_44_port, 
      mux_to_adder_43_port, mux_to_adder_42_port, mux_to_adder_41_port, 
      mux_to_adder_40_port, mux_to_adder_39_port, mux_to_adder_38_port, 
      mux_to_adder_37_port, mux_to_adder_36_port, mux_to_adder_35_port, 
      mux_to_adder_34_port, mux_to_adder_33_port, mux_to_adder_32_port, 
      mux_to_adder_31_port, mux_to_adder_30_port, mux_to_adder_29_port, 
      mux_to_adder_28_port, mux_to_adder_27_port, mux_to_adder_26_port, 
      mux_to_adder_25_port, mux_to_adder_24_port, mux_to_adder_23_port, 
      mux_to_adder_22_port, mux_to_adder_21_port, mux_to_adder_20_port, 
      mux_to_adder_19_port, mux_to_adder_18_port, mux_to_adder_17_port, 
      mux_to_adder_16_port, mux_to_adder_15_port, mux_to_adder_14_port, 
      mux_to_adder_13_port, mux_to_adder_12_port, mux_to_adder_11_port, 
      mux_to_adder_10_port, mux_to_adder_9_port, mux_to_adder_8_port, 
      mux_to_adder_7_port, mux_to_adder_6_port, mux_to_adder_5_port, 
      mux_to_adder_4_port, mux_to_adder_3_port, mux_to_adder_2_port, 
      mux_to_adder_1_port, mux_to_adder_0_port, nextA_0_port, nextA_57_port, 
      n_3205, n_3206, n_3207 : std_logic;

begin
   nextA <= ( nextA_63_port, nextA_62_port, nextA_61_port, nextA_60_port, 
      nextA_59_port, nextA_58_port, nextA_57_port, nextA_56_port, nextA_55_port
      , nextA_54_port, nextA_53_port, nextA_52_port, nextA_51_port, 
      nextA_50_port, nextA_49_port, nextA_48_port, nextA_47_port, nextA_46_port
      , nextA_45_port, nextA_44_port, nextA_43_port, nextA_42_port, 
      nextA_41_port, nextA_40_port, nextA_39_port, nextA_38_port, nextA_37_port
      , nextA_36_port, nextA_35_port, nextA_34_port, nextA_33_port, 
      nextA_32_port, nextA_31_port, nextA_30_port, nextA_29_port, nextA_28_port
      , nextA_27_port, nextA_26_port, nextA_25_port, nextA_24_port, 
      nextA_23_port, nextA_22_port, nextA_21_port, nextA_20_port, nextA_19_port
      , nextA_18_port, nextA_17_port, nextA_16_port, nextA_15_port, 
      nextA_14_port, nextA_13_port, nextA_12_port, nextA_11_port, nextA_10_port
      , nextA_9_port, nextA_8_port, nextA_7_port, nextA_6_port, nextA_5_port, 
      nextA_4_port, nextA_3_port, nextA_2_port, nextA_1_port, nextA_0_port );
   
   X_Logic0_port <= '0';
   nextA_0_port <= '0';
   encoder_1 : encoder_N64_RADIX3_11 port map( X(2) => encoderIn(2), X(1) => 
                           encoderIn(1), X(0) => encoderIn(0), Z(2) => 
                           encoder_to_mux_2_port, Z(1) => encoder_to_mux_1_port
                           , Z(0) => encoder_to_mux_0_port);
   ShiftnCompl_1 : ShiftnCompl_N64_11 port map( plusA(63) => prevA(63), 
                           plusA(62) => prevA(62), plusA(61) => prevA(61), 
                           plusA(60) => prevA(60), plusA(59) => prevA(59), 
                           plusA(58) => prevA(58), plusA(57) => prevA(57), 
                           plusA(56) => prevA(56), plusA(55) => prevA(55), 
                           plusA(54) => prevA(54), plusA(53) => prevA(53), 
                           plusA(52) => prevA(52), plusA(51) => prevA(51), 
                           plusA(50) => prevA(50), plusA(49) => prevA(49), 
                           plusA(48) => prevA(48), plusA(47) => prevA(47), 
                           plusA(46) => prevA(46), plusA(45) => prevA(45), 
                           plusA(44) => prevA(44), plusA(43) => prevA(43), 
                           plusA(42) => prevA(42), plusA(41) => prevA(41), 
                           plusA(40) => prevA(40), plusA(39) => prevA(39), 
                           plusA(38) => prevA(38), plusA(37) => prevA(37), 
                           plusA(36) => prevA(36), plusA(35) => prevA(35), 
                           plusA(34) => prevA(34), plusA(33) => prevA(33), 
                           plusA(32) => prevA(32), plusA(31) => prevA(31), 
                           plusA(30) => prevA(30), plusA(29) => prevA(29), 
                           plusA(28) => prevA(28), plusA(27) => prevA(27), 
                           plusA(26) => prevA(26), plusA(25) => prevA(25), 
                           plusA(24) => prevA(24), plusA(23) => prevA(23), 
                           plusA(22) => prevA(22), plusA(21) => prevA(21), 
                           plusA(20) => prevA(20), plusA(19) => prevA(19), 
                           plusA(18) => prevA(18), plusA(17) => prevA(17), 
                           plusA(16) => prevA(16), plusA(15) => prevA(15), 
                           plusA(14) => prevA(14), plusA(13) => prevA(13), 
                           plusA(12) => prevA(12), plusA(11) => prevA(11), 
                           plusA(10) => prevA(10), plusA(9) => prevA(9), 
                           plusA(8) => prevA(8), plusA(7) => prevA(7), plusA(6)
                           => prevA(6), plusA(5) => prevA(5), plusA(4) => 
                           prevA(4), plusA(3) => prevA(3), plusA(2) => prevA(2)
                           , plusA(1) => prevA(1), plusA(0) => prevA(0), 
                           plus2A_out(63) => plus2A_s_63_port, plus2A_out(62) 
                           => plus2A_s_62_port, plus2A_out(61) => 
                           plus2A_s_61_port, plus2A_out(60) => plus2A_s_60_port
                           , plus2A_out(59) => plus2A_s_59_port, plus2A_out(58)
                           => plus2A_s_58_port, plus2A_out(57) => 
                           plus2A_s_57_port, plus2A_out(56) => plus2A_s_56_port
                           , plus2A_out(55) => plus2A_s_55_port, plus2A_out(54)
                           => plus2A_s_54_port, plus2A_out(53) => 
                           plus2A_s_53_port, plus2A_out(52) => plus2A_s_52_port
                           , plus2A_out(51) => plus2A_s_51_port, plus2A_out(50)
                           => plus2A_s_50_port, plus2A_out(49) => 
                           plus2A_s_49_port, plus2A_out(48) => plus2A_s_48_port
                           , plus2A_out(47) => plus2A_s_47_port, plus2A_out(46)
                           => plus2A_s_46_port, plus2A_out(45) => 
                           plus2A_s_45_port, plus2A_out(44) => plus2A_s_44_port
                           , plus2A_out(43) => plus2A_s_43_port, plus2A_out(42)
                           => plus2A_s_42_port, plus2A_out(41) => 
                           plus2A_s_41_port, plus2A_out(40) => plus2A_s_40_port
                           , plus2A_out(39) => plus2A_s_39_port, plus2A_out(38)
                           => plus2A_s_38_port, plus2A_out(37) => 
                           plus2A_s_37_port, plus2A_out(36) => plus2A_s_36_port
                           , plus2A_out(35) => plus2A_s_35_port, plus2A_out(34)
                           => plus2A_s_34_port, plus2A_out(33) => 
                           plus2A_s_33_port, plus2A_out(32) => plus2A_s_32_port
                           , plus2A_out(31) => plus2A_s_31_port, plus2A_out(30)
                           => plus2A_s_30_port, plus2A_out(29) => 
                           plus2A_s_29_port, plus2A_out(28) => plus2A_s_28_port
                           , plus2A_out(27) => plus2A_s_27_port, plus2A_out(26)
                           => plus2A_s_26_port, plus2A_out(25) => 
                           plus2A_s_25_port, plus2A_out(24) => plus2A_s_24_port
                           , plus2A_out(23) => plus2A_s_23_port, plus2A_out(22)
                           => plus2A_s_22_port, plus2A_out(21) => 
                           plus2A_s_21_port, plus2A_out(20) => plus2A_s_20_port
                           , plus2A_out(19) => plus2A_s_19_port, plus2A_out(18)
                           => plus2A_s_18_port, plus2A_out(17) => 
                           plus2A_s_17_port, plus2A_out(16) => plus2A_s_16_port
                           , plus2A_out(15) => plus2A_s_15_port, plus2A_out(14)
                           => plus2A_s_14_port, plus2A_out(13) => 
                           plus2A_s_13_port, plus2A_out(12) => plus2A_s_12_port
                           , plus2A_out(11) => plus2A_s_11_port, plus2A_out(10)
                           => plus2A_s_10_port, plus2A_out(9) => 
                           plus2A_s_9_port, plus2A_out(8) => plus2A_s_8_port, 
                           plus2A_out(7) => plus2A_s_7_port, plus2A_out(6) => 
                           plus2A_s_6_port, plus2A_out(5) => plus2A_s_5_port, 
                           plus2A_out(4) => plus2A_s_4_port, plus2A_out(3) => 
                           plus2A_s_3_port, plus2A_out(2) => plus2A_s_2_port, 
                           plus2A_out(1) => plus2A_s_1_port, plus2A_out(0) => 
                           n_3205, minus2A_out(63) => minus2A_s_63_port, 
                           minus2A_out(62) => minus2A_s_62_port, 
                           minus2A_out(61) => minus2A_s_61_port, 
                           minus2A_out(60) => minus2A_s_60_port, 
                           minus2A_out(59) => minus2A_s_59_port, 
                           minus2A_out(58) => minus2A_s_58_port, 
                           minus2A_out(57) => minus2A_s_57_port, 
                           minus2A_out(56) => minus2A_s_56_port, 
                           minus2A_out(55) => minus2A_s_55_port, 
                           minus2A_out(54) => minus2A_s_54_port, 
                           minus2A_out(53) => minus2A_s_53_port, 
                           minus2A_out(52) => minus2A_s_52_port, 
                           minus2A_out(51) => minus2A_s_51_port, 
                           minus2A_out(50) => minus2A_s_50_port, 
                           minus2A_out(49) => minus2A_s_49_port, 
                           minus2A_out(48) => minus2A_s_48_port, 
                           minus2A_out(47) => minus2A_s_47_port, 
                           minus2A_out(46) => minus2A_s_46_port, 
                           minus2A_out(45) => minus2A_s_45_port, 
                           minus2A_out(44) => minus2A_s_44_port, 
                           minus2A_out(43) => minus2A_s_43_port, 
                           minus2A_out(42) => minus2A_s_42_port, 
                           minus2A_out(41) => minus2A_s_41_port, 
                           minus2A_out(40) => minus2A_s_40_port, 
                           minus2A_out(39) => minus2A_s_39_port, 
                           minus2A_out(38) => minus2A_s_38_port, 
                           minus2A_out(37) => minus2A_s_37_port, 
                           minus2A_out(36) => minus2A_s_36_port, 
                           minus2A_out(35) => minus2A_s_35_port, 
                           minus2A_out(34) => minus2A_s_34_port, 
                           minus2A_out(33) => minus2A_s_33_port, 
                           minus2A_out(32) => minus2A_s_32_port, 
                           minus2A_out(31) => minus2A_s_31_port, 
                           minus2A_out(30) => minus2A_s_30_port, 
                           minus2A_out(29) => minus2A_s_29_port, 
                           minus2A_out(28) => minus2A_s_28_port, 
                           minus2A_out(27) => minus2A_s_27_port, 
                           minus2A_out(26) => minus2A_s_26_port, 
                           minus2A_out(25) => minus2A_s_25_port, 
                           minus2A_out(24) => minus2A_s_24_port, 
                           minus2A_out(23) => minus2A_s_23_port, 
                           minus2A_out(22) => minus2A_s_22_port, 
                           minus2A_out(21) => minus2A_s_21_port, 
                           minus2A_out(20) => minus2A_s_20_port, 
                           minus2A_out(19) => minus2A_s_19_port, 
                           minus2A_out(18) => minus2A_s_18_port, 
                           minus2A_out(17) => minus2A_s_17_port, 
                           minus2A_out(16) => minus2A_s_16_port, 
                           minus2A_out(15) => minus2A_s_15_port, 
                           minus2A_out(14) => minus2A_s_14_port, 
                           minus2A_out(13) => minus2A_s_13_port, 
                           minus2A_out(12) => minus2A_s_12_port, 
                           minus2A_out(11) => minus2A_s_11_port, 
                           minus2A_out(10) => minus2A_s_10_port, minus2A_out(9)
                           => minus2A_s_9_port, minus2A_out(8) => 
                           minus2A_s_8_port, minus2A_out(7) => minus2A_s_7_port
                           , minus2A_out(6) => minus2A_s_6_port, minus2A_out(5)
                           => minus2A_s_5_port, minus2A_out(4) => 
                           minus2A_s_4_port, minus2A_out(3) => minus2A_s_3_port
                           , minus2A_out(2) => minus2A_s_2_port, minus2A_out(1)
                           => minus2A_s_1_port, minus2A_out(0) => 
                           minus2A_s_0_port, plus4A_out(63) => nextA_63_port, 
                           plus4A_out(62) => nextA_62_port, plus4A_out(61) => 
                           nextA_61_port, plus4A_out(60) => nextA_60_port, 
                           plus4A_out(59) => nextA_59_port, plus4A_out(58) => 
                           nextA_58_port, plus4A_out(57) => n3, plus4A_out(56) 
                           => nextA_56_port, plus4A_out(55) => nextA_55_port, 
                           plus4A_out(54) => nextA_54_port, plus4A_out(53) => 
                           nextA_53_port, plus4A_out(52) => nextA_52_port, 
                           plus4A_out(51) => nextA_51_port, plus4A_out(50) => 
                           nextA_50_port, plus4A_out(49) => nextA_49_port, 
                           plus4A_out(48) => nextA_48_port, plus4A_out(47) => 
                           nextA_47_port, plus4A_out(46) => nextA_46_port, 
                           plus4A_out(45) => nextA_45_port, plus4A_out(44) => 
                           nextA_44_port, plus4A_out(43) => nextA_43_port, 
                           plus4A_out(42) => nextA_42_port, plus4A_out(41) => 
                           nextA_41_port, plus4A_out(40) => nextA_40_port, 
                           plus4A_out(39) => nextA_39_port, plus4A_out(38) => 
                           nextA_38_port, plus4A_out(37) => nextA_37_port, 
                           plus4A_out(36) => nextA_36_port, plus4A_out(35) => 
                           nextA_35_port, plus4A_out(34) => nextA_34_port, 
                           plus4A_out(33) => nextA_33_port, plus4A_out(32) => 
                           nextA_32_port, plus4A_out(31) => nextA_31_port, 
                           plus4A_out(30) => nextA_30_port, plus4A_out(29) => 
                           nextA_29_port, plus4A_out(28) => nextA_28_port, 
                           plus4A_out(27) => nextA_27_port, plus4A_out(26) => 
                           nextA_26_port, plus4A_out(25) => nextA_25_port, 
                           plus4A_out(24) => nextA_24_port, plus4A_out(23) => 
                           nextA_23_port, plus4A_out(22) => nextA_22_port, 
                           plus4A_out(21) => nextA_21_port, plus4A_out(20) => 
                           nextA_20_port, plus4A_out(19) => nextA_19_port, 
                           plus4A_out(18) => nextA_18_port, plus4A_out(17) => 
                           nextA_17_port, plus4A_out(16) => nextA_16_port, 
                           plus4A_out(15) => nextA_15_port, plus4A_out(14) => 
                           nextA_14_port, plus4A_out(13) => nextA_13_port, 
                           plus4A_out(12) => nextA_12_port, plus4A_out(11) => 
                           nextA_11_port, plus4A_out(10) => nextA_10_port, 
                           plus4A_out(9) => nextA_9_port, plus4A_out(8) => 
                           nextA_8_port, plus4A_out(7) => nextA_7_port, 
                           plus4A_out(6) => nextA_6_port, plus4A_out(5) => 
                           nextA_5_port, plus4A_out(4) => nextA_4_port, 
                           plus4A_out(3) => nextA_3_port, plus4A_out(2) => 
                           nextA_2_port, plus4A_out(1) => nextA_1_port, 
                           plus4A_out(0) => n_3206, minus4A_out(63) => 
                           minus4A_s_63_port, minus4A_out(62) => 
                           minus4A_s_62_port, minus4A_out(61) => 
                           minus4A_s_61_port, minus4A_out(60) => 
                           minus4A_s_60_port, minus4A_out(59) => 
                           minus4A_s_59_port, minus4A_out(58) => 
                           minus4A_s_58_port, minus4A_out(57) => 
                           minus4A_s_57_port, minus4A_out(56) => 
                           minus4A_s_56_port, minus4A_out(55) => 
                           minus4A_s_55_port, minus4A_out(54) => 
                           minus4A_s_54_port, minus4A_out(53) => 
                           minus4A_s_53_port, minus4A_out(52) => 
                           minus4A_s_52_port, minus4A_out(51) => 
                           minus4A_s_51_port, minus4A_out(50) => 
                           minus4A_s_50_port, minus4A_out(49) => 
                           minus4A_s_49_port, minus4A_out(48) => 
                           minus4A_s_48_port, minus4A_out(47) => 
                           minus4A_s_47_port, minus4A_out(46) => 
                           minus4A_s_46_port, minus4A_out(45) => 
                           minus4A_s_45_port, minus4A_out(44) => 
                           minus4A_s_44_port, minus4A_out(43) => 
                           minus4A_s_43_port, minus4A_out(42) => 
                           minus4A_s_42_port, minus4A_out(41) => 
                           minus4A_s_41_port, minus4A_out(40) => 
                           minus4A_s_40_port, minus4A_out(39) => 
                           minus4A_s_39_port, minus4A_out(38) => 
                           minus4A_s_38_port, minus4A_out(37) => 
                           minus4A_s_37_port, minus4A_out(36) => 
                           minus4A_s_36_port, minus4A_out(35) => 
                           minus4A_s_35_port, minus4A_out(34) => 
                           minus4A_s_34_port, minus4A_out(33) => 
                           minus4A_s_33_port, minus4A_out(32) => 
                           minus4A_s_32_port, minus4A_out(31) => 
                           minus4A_s_31_port, minus4A_out(30) => 
                           minus4A_s_30_port, minus4A_out(29) => 
                           minus4A_s_29_port, minus4A_out(28) => 
                           minus4A_s_28_port, minus4A_out(27) => 
                           minus4A_s_27_port, minus4A_out(26) => 
                           minus4A_s_26_port, minus4A_out(25) => 
                           minus4A_s_25_port, minus4A_out(24) => 
                           minus4A_s_24_port, minus4A_out(23) => 
                           minus4A_s_23_port, minus4A_out(22) => 
                           minus4A_s_22_port, minus4A_out(21) => 
                           minus4A_s_21_port, minus4A_out(20) => 
                           minus4A_s_20_port, minus4A_out(19) => 
                           minus4A_s_19_port, minus4A_out(18) => 
                           minus4A_s_18_port, minus4A_out(17) => 
                           minus4A_s_17_port, minus4A_out(16) => 
                           minus4A_s_16_port, minus4A_out(15) => 
                           minus4A_s_15_port, minus4A_out(14) => 
                           minus4A_s_14_port, minus4A_out(13) => 
                           minus4A_s_13_port, minus4A_out(12) => 
                           minus4A_s_12_port, minus4A_out(11) => 
                           minus4A_s_11_port, minus4A_out(10) => 
                           minus4A_s_10_port, minus4A_out(9) => 
                           minus4A_s_9_port, minus4A_out(8) => minus4A_s_8_port
                           , minus4A_out(7) => minus4A_s_7_port, minus4A_out(6)
                           => minus4A_s_6_port, minus4A_out(5) => 
                           minus4A_s_5_port, minus4A_out(4) => minus4A_s_4_port
                           , minus4A_out(3) => minus4A_s_3_port, minus4A_out(2)
                           => minus4A_s_2_port, minus4A_out(1) => 
                           minus4A_s_1_port, minus4A_out(0) => minus4A_s_0_port
                           );
   mux_1 : MUX_GENERIC_N64_RADIX3_11 port map( plusA(63) => plus2A_s_63_port, 
                           plusA(62) => plus2A_s_62_port, plusA(61) => 
                           plus2A_s_61_port, plusA(60) => plus2A_s_60_port, 
                           plusA(59) => plus2A_s_59_port, plusA(58) => 
                           plus2A_s_58_port, plusA(57) => plus2A_s_57_port, 
                           plusA(56) => plus2A_s_56_port, plusA(55) => 
                           plus2A_s_55_port, plusA(54) => plus2A_s_54_port, 
                           plusA(53) => plus2A_s_53_port, plusA(52) => 
                           plus2A_s_52_port, plusA(51) => plus2A_s_51_port, 
                           plusA(50) => plus2A_s_50_port, plusA(49) => 
                           plus2A_s_49_port, plusA(48) => plus2A_s_48_port, 
                           plusA(47) => plus2A_s_47_port, plusA(46) => 
                           plus2A_s_46_port, plusA(45) => plus2A_s_45_port, 
                           plusA(44) => plus2A_s_44_port, plusA(43) => 
                           plus2A_s_43_port, plusA(42) => plus2A_s_42_port, 
                           plusA(41) => plus2A_s_41_port, plusA(40) => 
                           plus2A_s_40_port, plusA(39) => plus2A_s_39_port, 
                           plusA(38) => plus2A_s_38_port, plusA(37) => 
                           plus2A_s_37_port, plusA(36) => plus2A_s_36_port, 
                           plusA(35) => plus2A_s_35_port, plusA(34) => 
                           plus2A_s_34_port, plusA(33) => plus2A_s_33_port, 
                           plusA(32) => plus2A_s_32_port, plusA(31) => 
                           plus2A_s_31_port, plusA(30) => plus2A_s_30_port, 
                           plusA(29) => plus2A_s_29_port, plusA(28) => 
                           plus2A_s_28_port, plusA(27) => plus2A_s_27_port, 
                           plusA(26) => plus2A_s_26_port, plusA(25) => 
                           plus2A_s_25_port, plusA(24) => plus2A_s_24_port, 
                           plusA(23) => plus2A_s_23_port, plusA(22) => 
                           plus2A_s_22_port, plusA(21) => plus2A_s_21_port, 
                           plusA(20) => plus2A_s_20_port, plusA(19) => 
                           plus2A_s_19_port, plusA(18) => plus2A_s_18_port, 
                           plusA(17) => plus2A_s_17_port, plusA(16) => 
                           plus2A_s_16_port, plusA(15) => plus2A_s_15_port, 
                           plusA(14) => plus2A_s_14_port, plusA(13) => 
                           plus2A_s_13_port, plusA(12) => plus2A_s_12_port, 
                           plusA(11) => plus2A_s_11_port, plusA(10) => 
                           plus2A_s_10_port, plusA(9) => plus2A_s_9_port, 
                           plusA(8) => plus2A_s_8_port, plusA(7) => 
                           plus2A_s_7_port, plusA(6) => plus2A_s_6_port, 
                           plusA(5) => plus2A_s_5_port, plusA(4) => 
                           plus2A_s_4_port, plusA(3) => plus2A_s_3_port, 
                           plusA(2) => plus2A_s_2_port, plusA(1) => 
                           plus2A_s_1_port, plusA(0) => nextA_0_port, 
                           minusA(63) => minus2A_s_63_port, minusA(62) => 
                           minus2A_s_62_port, minusA(61) => minus2A_s_61_port, 
                           minusA(60) => minus2A_s_60_port, minusA(59) => 
                           minus2A_s_59_port, minusA(58) => minus2A_s_58_port, 
                           minusA(57) => minus2A_s_57_port, minusA(56) => 
                           minus2A_s_56_port, minusA(55) => minus2A_s_55_port, 
                           minusA(54) => minus2A_s_54_port, minusA(53) => 
                           minus2A_s_53_port, minusA(52) => minus2A_s_52_port, 
                           minusA(51) => minus2A_s_51_port, minusA(50) => 
                           minus2A_s_50_port, minusA(49) => minus2A_s_49_port, 
                           minusA(48) => minus2A_s_48_port, minusA(47) => 
                           minus2A_s_47_port, minusA(46) => minus2A_s_46_port, 
                           minusA(45) => minus2A_s_45_port, minusA(44) => 
                           minus2A_s_44_port, minusA(43) => minus2A_s_43_port, 
                           minusA(42) => minus2A_s_42_port, minusA(41) => 
                           minus2A_s_41_port, minusA(40) => minus2A_s_40_port, 
                           minusA(39) => minus2A_s_39_port, minusA(38) => 
                           minus2A_s_38_port, minusA(37) => minus2A_s_37_port, 
                           minusA(36) => minus2A_s_36_port, minusA(35) => 
                           minus2A_s_35_port, minusA(34) => minus2A_s_34_port, 
                           minusA(33) => minus2A_s_33_port, minusA(32) => 
                           minus2A_s_32_port, minusA(31) => minus2A_s_31_port, 
                           minusA(30) => minus2A_s_30_port, minusA(29) => 
                           minus2A_s_29_port, minusA(28) => minus2A_s_28_port, 
                           minusA(27) => minus2A_s_27_port, minusA(26) => 
                           minus2A_s_26_port, minusA(25) => minus2A_s_25_port, 
                           minusA(24) => minus2A_s_24_port, minusA(23) => 
                           minus2A_s_23_port, minusA(22) => minus2A_s_22_port, 
                           minusA(21) => minus2A_s_21_port, minusA(20) => 
                           minus2A_s_20_port, minusA(19) => minus2A_s_19_port, 
                           minusA(18) => minus2A_s_18_port, minusA(17) => 
                           minus2A_s_17_port, minusA(16) => minus2A_s_16_port, 
                           minusA(15) => minus2A_s_15_port, minusA(14) => 
                           minus2A_s_14_port, minusA(13) => minus2A_s_13_port, 
                           minusA(12) => minus2A_s_12_port, minusA(11) => 
                           minus2A_s_11_port, minusA(10) => minus2A_s_10_port, 
                           minusA(9) => minus2A_s_9_port, minusA(8) => 
                           minus2A_s_8_port, minusA(7) => minus2A_s_7_port, 
                           minusA(6) => minus2A_s_6_port, minusA(5) => 
                           minus2A_s_5_port, minusA(4) => minus2A_s_4_port, 
                           minusA(3) => minus2A_s_3_port, minusA(2) => 
                           minus2A_s_2_port, minusA(1) => minus2A_s_1_port, 
                           minusA(0) => minus2A_s_0_port, plus2A(63) => 
                           nextA_63_port, plus2A(62) => nextA_62_port, 
                           plus2A(61) => nextA_61_port, plus2A(60) => 
                           nextA_60_port, plus2A(59) => nextA_59_port, 
                           plus2A(58) => nextA_58_port, plus2A(57) => 
                           nextA_57_port, plus2A(56) => nextA_56_port, 
                           plus2A(55) => nextA_55_port, plus2A(54) => 
                           nextA_54_port, plus2A(53) => nextA_53_port, 
                           plus2A(52) => nextA_52_port, plus2A(51) => 
                           nextA_51_port, plus2A(50) => nextA_50_port, 
                           plus2A(49) => nextA_49_port, plus2A(48) => 
                           nextA_48_port, plus2A(47) => nextA_47_port, 
                           plus2A(46) => nextA_46_port, plus2A(45) => 
                           nextA_45_port, plus2A(44) => nextA_44_port, 
                           plus2A(43) => nextA_43_port, plus2A(42) => 
                           nextA_42_port, plus2A(41) => nextA_41_port, 
                           plus2A(40) => nextA_40_port, plus2A(39) => 
                           nextA_39_port, plus2A(38) => nextA_38_port, 
                           plus2A(37) => nextA_37_port, plus2A(36) => 
                           nextA_36_port, plus2A(35) => nextA_35_port, 
                           plus2A(34) => nextA_34_port, plus2A(33) => 
                           nextA_33_port, plus2A(32) => nextA_32_port, 
                           plus2A(31) => nextA_31_port, plus2A(30) => 
                           nextA_30_port, plus2A(29) => nextA_29_port, 
                           plus2A(28) => nextA_28_port, plus2A(27) => 
                           nextA_27_port, plus2A(26) => nextA_26_port, 
                           plus2A(25) => nextA_25_port, plus2A(24) => 
                           nextA_24_port, plus2A(23) => nextA_23_port, 
                           plus2A(22) => nextA_22_port, plus2A(21) => 
                           nextA_21_port, plus2A(20) => nextA_20_port, 
                           plus2A(19) => nextA_19_port, plus2A(18) => 
                           nextA_18_port, plus2A(17) => nextA_17_port, 
                           plus2A(16) => nextA_16_port, plus2A(15) => 
                           nextA_15_port, plus2A(14) => nextA_14_port, 
                           plus2A(13) => nextA_13_port, plus2A(12) => 
                           nextA_12_port, plus2A(11) => nextA_11_port, 
                           plus2A(10) => nextA_10_port, plus2A(9) => 
                           nextA_9_port, plus2A(8) => nextA_8_port, plus2A(7) 
                           => nextA_7_port, plus2A(6) => nextA_6_port, 
                           plus2A(5) => nextA_5_port, plus2A(4) => nextA_4_port
                           , plus2A(3) => nextA_3_port, plus2A(2) => 
                           nextA_2_port, plus2A(1) => nextA_1_port, plus2A(0) 
                           => nextA_0_port, minus2A(63) => minus4A_s_63_port, 
                           minus2A(62) => minus4A_s_62_port, minus2A(61) => 
                           minus4A_s_61_port, minus2A(60) => minus4A_s_60_port,
                           minus2A(59) => minus4A_s_59_port, minus2A(58) => 
                           minus4A_s_58_port, minus2A(57) => minus4A_s_57_port,
                           minus2A(56) => minus4A_s_56_port, minus2A(55) => 
                           minus4A_s_55_port, minus2A(54) => minus4A_s_54_port,
                           minus2A(53) => minus4A_s_53_port, minus2A(52) => 
                           minus4A_s_52_port, minus2A(51) => minus4A_s_51_port,
                           minus2A(50) => minus4A_s_50_port, minus2A(49) => 
                           minus4A_s_49_port, minus2A(48) => minus4A_s_48_port,
                           minus2A(47) => minus4A_s_47_port, minus2A(46) => 
                           minus4A_s_46_port, minus2A(45) => minus4A_s_45_port,
                           minus2A(44) => minus4A_s_44_port, minus2A(43) => 
                           minus4A_s_43_port, minus2A(42) => minus4A_s_42_port,
                           minus2A(41) => minus4A_s_41_port, minus2A(40) => 
                           minus4A_s_40_port, minus2A(39) => minus4A_s_39_port,
                           minus2A(38) => minus4A_s_38_port, minus2A(37) => 
                           minus4A_s_37_port, minus2A(36) => minus4A_s_36_port,
                           minus2A(35) => minus4A_s_35_port, minus2A(34) => 
                           minus4A_s_34_port, minus2A(33) => minus4A_s_33_port,
                           minus2A(32) => minus4A_s_32_port, minus2A(31) => 
                           minus4A_s_31_port, minus2A(30) => minus4A_s_30_port,
                           minus2A(29) => minus4A_s_29_port, minus2A(28) => 
                           minus4A_s_28_port, minus2A(27) => minus4A_s_27_port,
                           minus2A(26) => minus4A_s_26_port, minus2A(25) => 
                           minus4A_s_25_port, minus2A(24) => minus4A_s_24_port,
                           minus2A(23) => minus4A_s_23_port, minus2A(22) => 
                           minus4A_s_22_port, minus2A(21) => minus4A_s_21_port,
                           minus2A(20) => minus4A_s_20_port, minus2A(19) => 
                           minus4A_s_19_port, minus2A(18) => minus4A_s_18_port,
                           minus2A(17) => minus4A_s_17_port, minus2A(16) => 
                           minus4A_s_16_port, minus2A(15) => minus4A_s_15_port,
                           minus2A(14) => minus4A_s_14_port, minus2A(13) => 
                           minus4A_s_13_port, minus2A(12) => minus4A_s_12_port,
                           minus2A(11) => minus4A_s_11_port, minus2A(10) => 
                           minus4A_s_10_port, minus2A(9) => minus4A_s_9_port, 
                           minus2A(8) => minus4A_s_8_port, minus2A(7) => 
                           minus4A_s_7_port, minus2A(6) => minus4A_s_6_port, 
                           minus2A(5) => minus4A_s_5_port, minus2A(4) => 
                           minus4A_s_4_port, minus2A(3) => minus4A_s_3_port, 
                           minus2A(2) => minus4A_s_2_port, minus2A(1) => 
                           minus4A_s_1_port, minus2A(0) => minus4A_s_0_port, 
                           SEL(2) => encoder_to_mux_2_port, SEL(1) => 
                           encoder_to_mux_1_port, SEL(0) => 
                           encoder_to_mux_0_port, Y(63) => mux_to_adder_63_port
                           , Y(62) => mux_to_adder_62_port, Y(61) => 
                           mux_to_adder_61_port, Y(60) => mux_to_adder_60_port,
                           Y(59) => mux_to_adder_59_port, Y(58) => 
                           mux_to_adder_58_port, Y(57) => mux_to_adder_57_port,
                           Y(56) => mux_to_adder_56_port, Y(55) => 
                           mux_to_adder_55_port, Y(54) => mux_to_adder_54_port,
                           Y(53) => mux_to_adder_53_port, Y(52) => 
                           mux_to_adder_52_port, Y(51) => mux_to_adder_51_port,
                           Y(50) => mux_to_adder_50_port, Y(49) => 
                           mux_to_adder_49_port, Y(48) => mux_to_adder_48_port,
                           Y(47) => mux_to_adder_47_port, Y(46) => 
                           mux_to_adder_46_port, Y(45) => mux_to_adder_45_port,
                           Y(44) => mux_to_adder_44_port, Y(43) => 
                           mux_to_adder_43_port, Y(42) => mux_to_adder_42_port,
                           Y(41) => mux_to_adder_41_port, Y(40) => 
                           mux_to_adder_40_port, Y(39) => mux_to_adder_39_port,
                           Y(38) => mux_to_adder_38_port, Y(37) => 
                           mux_to_adder_37_port, Y(36) => mux_to_adder_36_port,
                           Y(35) => mux_to_adder_35_port, Y(34) => 
                           mux_to_adder_34_port, Y(33) => mux_to_adder_33_port,
                           Y(32) => mux_to_adder_32_port, Y(31) => 
                           mux_to_adder_31_port, Y(30) => mux_to_adder_30_port,
                           Y(29) => mux_to_adder_29_port, Y(28) => 
                           mux_to_adder_28_port, Y(27) => mux_to_adder_27_port,
                           Y(26) => mux_to_adder_26_port, Y(25) => 
                           mux_to_adder_25_port, Y(24) => mux_to_adder_24_port,
                           Y(23) => mux_to_adder_23_port, Y(22) => 
                           mux_to_adder_22_port, Y(21) => mux_to_adder_21_port,
                           Y(20) => mux_to_adder_20_port, Y(19) => 
                           mux_to_adder_19_port, Y(18) => mux_to_adder_18_port,
                           Y(17) => mux_to_adder_17_port, Y(16) => 
                           mux_to_adder_16_port, Y(15) => mux_to_adder_15_port,
                           Y(14) => mux_to_adder_14_port, Y(13) => 
                           mux_to_adder_13_port, Y(12) => mux_to_adder_12_port,
                           Y(11) => mux_to_adder_11_port, Y(10) => 
                           mux_to_adder_10_port, Y(9) => mux_to_adder_9_port, 
                           Y(8) => mux_to_adder_8_port, Y(7) => 
                           mux_to_adder_7_port, Y(6) => mux_to_adder_6_port, 
                           Y(5) => mux_to_adder_5_port, Y(4) => 
                           mux_to_adder_4_port, Y(3) => mux_to_adder_3_port, 
                           Y(2) => mux_to_adder_2_port, Y(1) => 
                           mux_to_adder_1_port, Y(0) => mux_to_adder_0_port);
   rca_1 : RCA_N64_11 port map( A(63) => mux_to_adder_63_port, A(62) => 
                           mux_to_adder_62_port, A(61) => mux_to_adder_61_port,
                           A(60) => mux_to_adder_60_port, A(59) => 
                           mux_to_adder_59_port, A(58) => mux_to_adder_58_port,
                           A(57) => mux_to_adder_57_port, A(56) => 
                           mux_to_adder_56_port, A(55) => mux_to_adder_55_port,
                           A(54) => mux_to_adder_54_port, A(53) => 
                           mux_to_adder_53_port, A(52) => mux_to_adder_52_port,
                           A(51) => mux_to_adder_51_port, A(50) => 
                           mux_to_adder_50_port, A(49) => mux_to_adder_49_port,
                           A(48) => mux_to_adder_48_port, A(47) => 
                           mux_to_adder_47_port, A(46) => mux_to_adder_46_port,
                           A(45) => mux_to_adder_45_port, A(44) => 
                           mux_to_adder_44_port, A(43) => mux_to_adder_43_port,
                           A(42) => mux_to_adder_42_port, A(41) => 
                           mux_to_adder_41_port, A(40) => mux_to_adder_40_port,
                           A(39) => mux_to_adder_39_port, A(38) => 
                           mux_to_adder_38_port, A(37) => mux_to_adder_37_port,
                           A(36) => mux_to_adder_36_port, A(35) => 
                           mux_to_adder_35_port, A(34) => mux_to_adder_34_port,
                           A(33) => mux_to_adder_33_port, A(32) => 
                           mux_to_adder_32_port, A(31) => mux_to_adder_31_port,
                           A(30) => mux_to_adder_30_port, A(29) => 
                           mux_to_adder_29_port, A(28) => mux_to_adder_28_port,
                           A(27) => mux_to_adder_27_port, A(26) => 
                           mux_to_adder_26_port, A(25) => mux_to_adder_25_port,
                           A(24) => mux_to_adder_24_port, A(23) => 
                           mux_to_adder_23_port, A(22) => mux_to_adder_22_port,
                           A(21) => mux_to_adder_21_port, A(20) => 
                           mux_to_adder_20_port, A(19) => mux_to_adder_19_port,
                           A(18) => mux_to_adder_18_port, A(17) => 
                           mux_to_adder_17_port, A(16) => mux_to_adder_16_port,
                           A(15) => mux_to_adder_15_port, A(14) => 
                           mux_to_adder_14_port, A(13) => mux_to_adder_13_port,
                           A(12) => mux_to_adder_12_port, A(11) => 
                           mux_to_adder_11_port, A(10) => mux_to_adder_10_port,
                           A(9) => mux_to_adder_9_port, A(8) => 
                           mux_to_adder_8_port, A(7) => mux_to_adder_7_port, 
                           A(6) => mux_to_adder_6_port, A(5) => 
                           mux_to_adder_5_port, A(4) => mux_to_adder_4_port, 
                           A(3) => mux_to_adder_3_port, A(2) => 
                           mux_to_adder_2_port, A(1) => mux_to_adder_1_port, 
                           A(0) => mux_to_adder_0_port, B(63) => prevSum(63), 
                           B(62) => prevSum(62), B(61) => prevSum(61), B(60) =>
                           prevSum(60), B(59) => prevSum(59), B(58) => 
                           prevSum(58), B(57) => prevSum(57), B(56) => 
                           prevSum(56), B(55) => prevSum(55), B(54) => 
                           prevSum(54), B(53) => prevSum(53), B(52) => 
                           prevSum(52), B(51) => prevSum(51), B(50) => 
                           prevSum(50), B(49) => prevSum(49), B(48) => 
                           prevSum(48), B(47) => prevSum(47), B(46) => 
                           prevSum(46), B(45) => prevSum(45), B(44) => 
                           prevSum(44), B(43) => prevSum(43), B(42) => 
                           prevSum(42), B(41) => prevSum(41), B(40) => 
                           prevSum(40), B(39) => prevSum(39), B(38) => 
                           prevSum(38), B(37) => prevSum(37), B(36) => 
                           prevSum(36), B(35) => prevSum(35), B(34) => 
                           prevSum(34), B(33) => prevSum(33), B(32) => 
                           prevSum(32), B(31) => prevSum(31), B(30) => 
                           prevSum(30), B(29) => prevSum(29), B(28) => 
                           prevSum(28), B(27) => prevSum(27), B(26) => 
                           prevSum(26), B(25) => prevSum(25), B(24) => 
                           prevSum(24), B(23) => prevSum(23), B(22) => 
                           prevSum(22), B(21) => prevSum(21), B(20) => 
                           prevSum(20), B(19) => prevSum(19), B(18) => 
                           prevSum(18), B(17) => prevSum(17), B(16) => 
                           prevSum(16), B(15) => prevSum(15), B(14) => 
                           prevSum(14), B(13) => prevSum(13), B(12) => 
                           prevSum(12), B(11) => prevSum(11), B(10) => 
                           prevSum(10), B(9) => prevSum(9), B(8) => prevSum(8),
                           B(7) => prevSum(7), B(6) => prevSum(6), B(5) => 
                           prevSum(5), B(4) => prevSum(4), B(3) => prevSum(3), 
                           B(2) => prevSum(2), B(1) => prevSum(1), B(0) => 
                           prevSum(0), Ci => X_Logic0_port, S(63) => 
                           nextSum(63), S(62) => nextSum(62), S(61) => 
                           nextSum(61), S(60) => nextSum(60), S(59) => 
                           nextSum(59), S(58) => nextSum(58), S(57) => 
                           nextSum(57), S(56) => nextSum(56), S(55) => 
                           nextSum(55), S(54) => nextSum(54), S(53) => 
                           nextSum(53), S(52) => nextSum(52), S(51) => 
                           nextSum(51), S(50) => nextSum(50), S(49) => 
                           nextSum(49), S(48) => nextSum(48), S(47) => 
                           nextSum(47), S(46) => nextSum(46), S(45) => 
                           nextSum(45), S(44) => nextSum(44), S(43) => 
                           nextSum(43), S(42) => nextSum(42), S(41) => 
                           nextSum(41), S(40) => nextSum(40), S(39) => 
                           nextSum(39), S(38) => nextSum(38), S(37) => 
                           nextSum(37), S(36) => nextSum(36), S(35) => 
                           nextSum(35), S(34) => nextSum(34), S(33) => 
                           nextSum(33), S(32) => nextSum(32), S(31) => 
                           nextSum(31), S(30) => nextSum(30), S(29) => 
                           nextSum(29), S(28) => nextSum(28), S(27) => 
                           nextSum(27), S(26) => nextSum(26), S(25) => 
                           nextSum(25), S(24) => nextSum(24), S(23) => 
                           nextSum(23), S(22) => nextSum(22), S(21) => 
                           nextSum(21), S(20) => nextSum(20), S(19) => 
                           nextSum(19), S(18) => nextSum(18), S(17) => 
                           nextSum(17), S(16) => nextSum(16), S(15) => 
                           nextSum(15), S(14) => nextSum(14), S(13) => 
                           nextSum(13), S(12) => nextSum(12), S(11) => 
                           nextSum(11), S(10) => nextSum(10), S(9) => 
                           nextSum(9), S(8) => nextSum(8), S(7) => nextSum(7), 
                           S(6) => nextSum(6), S(5) => nextSum(5), S(4) => 
                           nextSum(4), S(3) => nextSum(3), S(2) => nextSum(2), 
                           S(1) => nextSum(1), S(0) => nextSum(0), Co => n_3207
                           );
   U3 : BUF_X1 port map( A => n3, Z => nextA_57_port);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity booth_mul_row_N64_RADIX3_12 is

   port( prevA, prevSum : in std_logic_vector (63 downto 0);  encoderIn : in 
         std_logic_vector (2 downto 0);  nextA, nextSum : out std_logic_vector 
         (63 downto 0));

end booth_mul_row_N64_RADIX3_12;

architecture SYN_struct of booth_mul_row_N64_RADIX3_12 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component RCA_N64_12
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component MUX_GENERIC_N64_RADIX3_12
      port( plusA, minusA, plus2A, minus2A : in std_logic_vector (63 downto 0);
            SEL : in std_logic_vector (2 downto 0);  Y : out std_logic_vector 
            (63 downto 0));
   end component;
   
   component ShiftnCompl_N64_12
      port( plusA : in std_logic_vector (63 downto 0);  plus2A_out, minus2A_out
            , plus4A_out, minus4A_out : out std_logic_vector (63 downto 0));
   end component;
   
   component encoder_N64_RADIX3_12
      port( X : in std_logic_vector (2 downto 0);  Z : out std_logic_vector (2 
            downto 0));
   end component;
   
   signal X_Logic0_port, nextA_63_port, nextA_62_port, nextA_61_port, 
      nextA_60_port, nextA_59_port, nextA_58_port, n3, nextA_56_port, 
      nextA_55_port, nextA_54_port, nextA_53_port, nextA_52_port, nextA_51_port
      , nextA_50_port, nextA_49_port, nextA_48_port, nextA_47_port, 
      nextA_46_port, nextA_45_port, nextA_44_port, nextA_43_port, nextA_42_port
      , nextA_41_port, nextA_40_port, nextA_39_port, nextA_38_port, 
      nextA_37_port, nextA_36_port, nextA_35_port, nextA_34_port, nextA_33_port
      , nextA_32_port, nextA_31_port, nextA_30_port, nextA_29_port, 
      nextA_28_port, nextA_27_port, nextA_26_port, nextA_25_port, nextA_24_port
      , nextA_23_port, nextA_22_port, nextA_21_port, nextA_20_port, 
      nextA_19_port, nextA_18_port, nextA_17_port, nextA_16_port, nextA_15_port
      , nextA_14_port, nextA_13_port, nextA_12_port, nextA_11_port, 
      nextA_10_port, nextA_9_port, nextA_8_port, nextA_7_port, nextA_6_port, 
      nextA_5_port, nextA_4_port, nextA_3_port, nextA_2_port, nextA_1_port, 
      encoder_to_mux_2_port, encoder_to_mux_1_port, encoder_to_mux_0_port, 
      plus2A_s_63_port, plus2A_s_62_port, plus2A_s_61_port, plus2A_s_60_port, 
      plus2A_s_59_port, plus2A_s_58_port, plus2A_s_57_port, plus2A_s_56_port, 
      plus2A_s_55_port, plus2A_s_54_port, plus2A_s_53_port, plus2A_s_52_port, 
      plus2A_s_51_port, plus2A_s_50_port, plus2A_s_49_port, plus2A_s_48_port, 
      plus2A_s_47_port, plus2A_s_46_port, plus2A_s_45_port, plus2A_s_44_port, 
      plus2A_s_43_port, plus2A_s_42_port, plus2A_s_41_port, plus2A_s_40_port, 
      plus2A_s_39_port, plus2A_s_38_port, plus2A_s_37_port, plus2A_s_36_port, 
      plus2A_s_35_port, plus2A_s_34_port, plus2A_s_33_port, plus2A_s_32_port, 
      plus2A_s_31_port, plus2A_s_30_port, plus2A_s_29_port, plus2A_s_28_port, 
      plus2A_s_27_port, plus2A_s_26_port, plus2A_s_25_port, plus2A_s_24_port, 
      plus2A_s_23_port, plus2A_s_22_port, plus2A_s_21_port, plus2A_s_20_port, 
      plus2A_s_19_port, plus2A_s_18_port, plus2A_s_17_port, plus2A_s_16_port, 
      plus2A_s_15_port, plus2A_s_14_port, plus2A_s_13_port, plus2A_s_12_port, 
      plus2A_s_11_port, plus2A_s_10_port, plus2A_s_9_port, plus2A_s_8_port, 
      plus2A_s_7_port, plus2A_s_6_port, plus2A_s_5_port, plus2A_s_4_port, 
      plus2A_s_3_port, plus2A_s_2_port, plus2A_s_1_port, minus2A_s_63_port, 
      minus2A_s_62_port, minus2A_s_61_port, minus2A_s_60_port, 
      minus2A_s_59_port, minus2A_s_58_port, minus2A_s_57_port, 
      minus2A_s_56_port, minus2A_s_55_port, minus2A_s_54_port, 
      minus2A_s_53_port, minus2A_s_52_port, minus2A_s_51_port, 
      minus2A_s_50_port, minus2A_s_49_port, minus2A_s_48_port, 
      minus2A_s_47_port, minus2A_s_46_port, minus2A_s_45_port, 
      minus2A_s_44_port, minus2A_s_43_port, minus2A_s_42_port, 
      minus2A_s_41_port, minus2A_s_40_port, minus2A_s_39_port, 
      minus2A_s_38_port, minus2A_s_37_port, minus2A_s_36_port, 
      minus2A_s_35_port, minus2A_s_34_port, minus2A_s_33_port, 
      minus2A_s_32_port, minus2A_s_31_port, minus2A_s_30_port, 
      minus2A_s_29_port, minus2A_s_28_port, minus2A_s_27_port, 
      minus2A_s_26_port, minus2A_s_25_port, minus2A_s_24_port, 
      minus2A_s_23_port, minus2A_s_22_port, minus2A_s_21_port, 
      minus2A_s_20_port, minus2A_s_19_port, minus2A_s_18_port, 
      minus2A_s_17_port, minus2A_s_16_port, minus2A_s_15_port, 
      minus2A_s_14_port, minus2A_s_13_port, minus2A_s_12_port, 
      minus2A_s_11_port, minus2A_s_10_port, minus2A_s_9_port, minus2A_s_8_port,
      minus2A_s_7_port, minus2A_s_6_port, minus2A_s_5_port, minus2A_s_4_port, 
      minus2A_s_3_port, minus2A_s_2_port, minus2A_s_1_port, minus2A_s_0_port, 
      minus4A_s_63_port, minus4A_s_62_port, minus4A_s_61_port, 
      minus4A_s_60_port, minus4A_s_59_port, minus4A_s_58_port, 
      minus4A_s_57_port, minus4A_s_56_port, minus4A_s_55_port, 
      minus4A_s_54_port, minus4A_s_53_port, minus4A_s_52_port, 
      minus4A_s_51_port, minus4A_s_50_port, minus4A_s_49_port, 
      minus4A_s_48_port, minus4A_s_47_port, minus4A_s_46_port, 
      minus4A_s_45_port, minus4A_s_44_port, minus4A_s_43_port, 
      minus4A_s_42_port, minus4A_s_41_port, minus4A_s_40_port, 
      minus4A_s_39_port, minus4A_s_38_port, minus4A_s_37_port, 
      minus4A_s_36_port, minus4A_s_35_port, minus4A_s_34_port, 
      minus4A_s_33_port, minus4A_s_32_port, minus4A_s_31_port, 
      minus4A_s_30_port, minus4A_s_29_port, minus4A_s_28_port, 
      minus4A_s_27_port, minus4A_s_26_port, minus4A_s_25_port, 
      minus4A_s_24_port, minus4A_s_23_port, minus4A_s_22_port, 
      minus4A_s_21_port, minus4A_s_20_port, minus4A_s_19_port, 
      minus4A_s_18_port, minus4A_s_17_port, minus4A_s_16_port, 
      minus4A_s_15_port, minus4A_s_14_port, minus4A_s_13_port, 
      minus4A_s_12_port, minus4A_s_11_port, minus4A_s_10_port, minus4A_s_9_port
      , minus4A_s_8_port, minus4A_s_7_port, minus4A_s_6_port, minus4A_s_5_port,
      minus4A_s_4_port, minus4A_s_3_port, minus4A_s_2_port, minus4A_s_1_port, 
      minus4A_s_0_port, mux_to_adder_63_port, mux_to_adder_62_port, 
      mux_to_adder_61_port, mux_to_adder_60_port, mux_to_adder_59_port, 
      mux_to_adder_58_port, mux_to_adder_57_port, mux_to_adder_56_port, 
      mux_to_adder_55_port, mux_to_adder_54_port, mux_to_adder_53_port, 
      mux_to_adder_52_port, mux_to_adder_51_port, mux_to_adder_50_port, 
      mux_to_adder_49_port, mux_to_adder_48_port, mux_to_adder_47_port, 
      mux_to_adder_46_port, mux_to_adder_45_port, mux_to_adder_44_port, 
      mux_to_adder_43_port, mux_to_adder_42_port, mux_to_adder_41_port, 
      mux_to_adder_40_port, mux_to_adder_39_port, mux_to_adder_38_port, 
      mux_to_adder_37_port, mux_to_adder_36_port, mux_to_adder_35_port, 
      mux_to_adder_34_port, mux_to_adder_33_port, mux_to_adder_32_port, 
      mux_to_adder_31_port, mux_to_adder_30_port, mux_to_adder_29_port, 
      mux_to_adder_28_port, mux_to_adder_27_port, mux_to_adder_26_port, 
      mux_to_adder_25_port, mux_to_adder_24_port, mux_to_adder_23_port, 
      mux_to_adder_22_port, mux_to_adder_21_port, mux_to_adder_20_port, 
      mux_to_adder_19_port, mux_to_adder_18_port, mux_to_adder_17_port, 
      mux_to_adder_16_port, mux_to_adder_15_port, mux_to_adder_14_port, 
      mux_to_adder_13_port, mux_to_adder_12_port, mux_to_adder_11_port, 
      mux_to_adder_10_port, mux_to_adder_9_port, mux_to_adder_8_port, 
      mux_to_adder_7_port, mux_to_adder_6_port, mux_to_adder_5_port, 
      mux_to_adder_4_port, mux_to_adder_3_port, mux_to_adder_2_port, 
      mux_to_adder_1_port, mux_to_adder_0_port, nextA_0_port, nextA_57_port, 
      n_3208, n_3209, n_3210 : std_logic;

begin
   nextA <= ( nextA_63_port, nextA_62_port, nextA_61_port, nextA_60_port, 
      nextA_59_port, nextA_58_port, nextA_57_port, nextA_56_port, nextA_55_port
      , nextA_54_port, nextA_53_port, nextA_52_port, nextA_51_port, 
      nextA_50_port, nextA_49_port, nextA_48_port, nextA_47_port, nextA_46_port
      , nextA_45_port, nextA_44_port, nextA_43_port, nextA_42_port, 
      nextA_41_port, nextA_40_port, nextA_39_port, nextA_38_port, nextA_37_port
      , nextA_36_port, nextA_35_port, nextA_34_port, nextA_33_port, 
      nextA_32_port, nextA_31_port, nextA_30_port, nextA_29_port, nextA_28_port
      , nextA_27_port, nextA_26_port, nextA_25_port, nextA_24_port, 
      nextA_23_port, nextA_22_port, nextA_21_port, nextA_20_port, nextA_19_port
      , nextA_18_port, nextA_17_port, nextA_16_port, nextA_15_port, 
      nextA_14_port, nextA_13_port, nextA_12_port, nextA_11_port, nextA_10_port
      , nextA_9_port, nextA_8_port, nextA_7_port, nextA_6_port, nextA_5_port, 
      nextA_4_port, nextA_3_port, nextA_2_port, nextA_1_port, nextA_0_port );
   
   X_Logic0_port <= '0';
   nextA_0_port <= '0';
   encoder_1 : encoder_N64_RADIX3_12 port map( X(2) => encoderIn(2), X(1) => 
                           encoderIn(1), X(0) => encoderIn(0), Z(2) => 
                           encoder_to_mux_2_port, Z(1) => encoder_to_mux_1_port
                           , Z(0) => encoder_to_mux_0_port);
   ShiftnCompl_1 : ShiftnCompl_N64_12 port map( plusA(63) => prevA(63), 
                           plusA(62) => prevA(62), plusA(61) => prevA(61), 
                           plusA(60) => prevA(60), plusA(59) => prevA(59), 
                           plusA(58) => prevA(58), plusA(57) => prevA(57), 
                           plusA(56) => prevA(56), plusA(55) => prevA(55), 
                           plusA(54) => prevA(54), plusA(53) => prevA(53), 
                           plusA(52) => prevA(52), plusA(51) => prevA(51), 
                           plusA(50) => prevA(50), plusA(49) => prevA(49), 
                           plusA(48) => prevA(48), plusA(47) => prevA(47), 
                           plusA(46) => prevA(46), plusA(45) => prevA(45), 
                           plusA(44) => prevA(44), plusA(43) => prevA(43), 
                           plusA(42) => prevA(42), plusA(41) => prevA(41), 
                           plusA(40) => prevA(40), plusA(39) => prevA(39), 
                           plusA(38) => prevA(38), plusA(37) => prevA(37), 
                           plusA(36) => prevA(36), plusA(35) => prevA(35), 
                           plusA(34) => prevA(34), plusA(33) => prevA(33), 
                           plusA(32) => prevA(32), plusA(31) => prevA(31), 
                           plusA(30) => prevA(30), plusA(29) => prevA(29), 
                           plusA(28) => prevA(28), plusA(27) => prevA(27), 
                           plusA(26) => prevA(26), plusA(25) => prevA(25), 
                           plusA(24) => prevA(24), plusA(23) => prevA(23), 
                           plusA(22) => prevA(22), plusA(21) => prevA(21), 
                           plusA(20) => prevA(20), plusA(19) => prevA(19), 
                           plusA(18) => prevA(18), plusA(17) => prevA(17), 
                           plusA(16) => prevA(16), plusA(15) => prevA(15), 
                           plusA(14) => prevA(14), plusA(13) => prevA(13), 
                           plusA(12) => prevA(12), plusA(11) => prevA(11), 
                           plusA(10) => prevA(10), plusA(9) => prevA(9), 
                           plusA(8) => prevA(8), plusA(7) => prevA(7), plusA(6)
                           => prevA(6), plusA(5) => prevA(5), plusA(4) => 
                           prevA(4), plusA(3) => prevA(3), plusA(2) => prevA(2)
                           , plusA(1) => prevA(1), plusA(0) => prevA(0), 
                           plus2A_out(63) => plus2A_s_63_port, plus2A_out(62) 
                           => plus2A_s_62_port, plus2A_out(61) => 
                           plus2A_s_61_port, plus2A_out(60) => plus2A_s_60_port
                           , plus2A_out(59) => plus2A_s_59_port, plus2A_out(58)
                           => plus2A_s_58_port, plus2A_out(57) => 
                           plus2A_s_57_port, plus2A_out(56) => plus2A_s_56_port
                           , plus2A_out(55) => plus2A_s_55_port, plus2A_out(54)
                           => plus2A_s_54_port, plus2A_out(53) => 
                           plus2A_s_53_port, plus2A_out(52) => plus2A_s_52_port
                           , plus2A_out(51) => plus2A_s_51_port, plus2A_out(50)
                           => plus2A_s_50_port, plus2A_out(49) => 
                           plus2A_s_49_port, plus2A_out(48) => plus2A_s_48_port
                           , plus2A_out(47) => plus2A_s_47_port, plus2A_out(46)
                           => plus2A_s_46_port, plus2A_out(45) => 
                           plus2A_s_45_port, plus2A_out(44) => plus2A_s_44_port
                           , plus2A_out(43) => plus2A_s_43_port, plus2A_out(42)
                           => plus2A_s_42_port, plus2A_out(41) => 
                           plus2A_s_41_port, plus2A_out(40) => plus2A_s_40_port
                           , plus2A_out(39) => plus2A_s_39_port, plus2A_out(38)
                           => plus2A_s_38_port, plus2A_out(37) => 
                           plus2A_s_37_port, plus2A_out(36) => plus2A_s_36_port
                           , plus2A_out(35) => plus2A_s_35_port, plus2A_out(34)
                           => plus2A_s_34_port, plus2A_out(33) => 
                           plus2A_s_33_port, plus2A_out(32) => plus2A_s_32_port
                           , plus2A_out(31) => plus2A_s_31_port, plus2A_out(30)
                           => plus2A_s_30_port, plus2A_out(29) => 
                           plus2A_s_29_port, plus2A_out(28) => plus2A_s_28_port
                           , plus2A_out(27) => plus2A_s_27_port, plus2A_out(26)
                           => plus2A_s_26_port, plus2A_out(25) => 
                           plus2A_s_25_port, plus2A_out(24) => plus2A_s_24_port
                           , plus2A_out(23) => plus2A_s_23_port, plus2A_out(22)
                           => plus2A_s_22_port, plus2A_out(21) => 
                           plus2A_s_21_port, plus2A_out(20) => plus2A_s_20_port
                           , plus2A_out(19) => plus2A_s_19_port, plus2A_out(18)
                           => plus2A_s_18_port, plus2A_out(17) => 
                           plus2A_s_17_port, plus2A_out(16) => plus2A_s_16_port
                           , plus2A_out(15) => plus2A_s_15_port, plus2A_out(14)
                           => plus2A_s_14_port, plus2A_out(13) => 
                           plus2A_s_13_port, plus2A_out(12) => plus2A_s_12_port
                           , plus2A_out(11) => plus2A_s_11_port, plus2A_out(10)
                           => plus2A_s_10_port, plus2A_out(9) => 
                           plus2A_s_9_port, plus2A_out(8) => plus2A_s_8_port, 
                           plus2A_out(7) => plus2A_s_7_port, plus2A_out(6) => 
                           plus2A_s_6_port, plus2A_out(5) => plus2A_s_5_port, 
                           plus2A_out(4) => plus2A_s_4_port, plus2A_out(3) => 
                           plus2A_s_3_port, plus2A_out(2) => plus2A_s_2_port, 
                           plus2A_out(1) => plus2A_s_1_port, plus2A_out(0) => 
                           n_3208, minus2A_out(63) => minus2A_s_63_port, 
                           minus2A_out(62) => minus2A_s_62_port, 
                           minus2A_out(61) => minus2A_s_61_port, 
                           minus2A_out(60) => minus2A_s_60_port, 
                           minus2A_out(59) => minus2A_s_59_port, 
                           minus2A_out(58) => minus2A_s_58_port, 
                           minus2A_out(57) => minus2A_s_57_port, 
                           minus2A_out(56) => minus2A_s_56_port, 
                           minus2A_out(55) => minus2A_s_55_port, 
                           minus2A_out(54) => minus2A_s_54_port, 
                           minus2A_out(53) => minus2A_s_53_port, 
                           minus2A_out(52) => minus2A_s_52_port, 
                           minus2A_out(51) => minus2A_s_51_port, 
                           minus2A_out(50) => minus2A_s_50_port, 
                           minus2A_out(49) => minus2A_s_49_port, 
                           minus2A_out(48) => minus2A_s_48_port, 
                           minus2A_out(47) => minus2A_s_47_port, 
                           minus2A_out(46) => minus2A_s_46_port, 
                           minus2A_out(45) => minus2A_s_45_port, 
                           minus2A_out(44) => minus2A_s_44_port, 
                           minus2A_out(43) => minus2A_s_43_port, 
                           minus2A_out(42) => minus2A_s_42_port, 
                           minus2A_out(41) => minus2A_s_41_port, 
                           minus2A_out(40) => minus2A_s_40_port, 
                           minus2A_out(39) => minus2A_s_39_port, 
                           minus2A_out(38) => minus2A_s_38_port, 
                           minus2A_out(37) => minus2A_s_37_port, 
                           minus2A_out(36) => minus2A_s_36_port, 
                           minus2A_out(35) => minus2A_s_35_port, 
                           minus2A_out(34) => minus2A_s_34_port, 
                           minus2A_out(33) => minus2A_s_33_port, 
                           minus2A_out(32) => minus2A_s_32_port, 
                           minus2A_out(31) => minus2A_s_31_port, 
                           minus2A_out(30) => minus2A_s_30_port, 
                           minus2A_out(29) => minus2A_s_29_port, 
                           minus2A_out(28) => minus2A_s_28_port, 
                           minus2A_out(27) => minus2A_s_27_port, 
                           minus2A_out(26) => minus2A_s_26_port, 
                           minus2A_out(25) => minus2A_s_25_port, 
                           minus2A_out(24) => minus2A_s_24_port, 
                           minus2A_out(23) => minus2A_s_23_port, 
                           minus2A_out(22) => minus2A_s_22_port, 
                           minus2A_out(21) => minus2A_s_21_port, 
                           minus2A_out(20) => minus2A_s_20_port, 
                           minus2A_out(19) => minus2A_s_19_port, 
                           minus2A_out(18) => minus2A_s_18_port, 
                           minus2A_out(17) => minus2A_s_17_port, 
                           minus2A_out(16) => minus2A_s_16_port, 
                           minus2A_out(15) => minus2A_s_15_port, 
                           minus2A_out(14) => minus2A_s_14_port, 
                           minus2A_out(13) => minus2A_s_13_port, 
                           minus2A_out(12) => minus2A_s_12_port, 
                           minus2A_out(11) => minus2A_s_11_port, 
                           minus2A_out(10) => minus2A_s_10_port, minus2A_out(9)
                           => minus2A_s_9_port, minus2A_out(8) => 
                           minus2A_s_8_port, minus2A_out(7) => minus2A_s_7_port
                           , minus2A_out(6) => minus2A_s_6_port, minus2A_out(5)
                           => minus2A_s_5_port, minus2A_out(4) => 
                           minus2A_s_4_port, minus2A_out(3) => minus2A_s_3_port
                           , minus2A_out(2) => minus2A_s_2_port, minus2A_out(1)
                           => minus2A_s_1_port, minus2A_out(0) => 
                           minus2A_s_0_port, plus4A_out(63) => nextA_63_port, 
                           plus4A_out(62) => nextA_62_port, plus4A_out(61) => 
                           nextA_61_port, plus4A_out(60) => nextA_60_port, 
                           plus4A_out(59) => nextA_59_port, plus4A_out(58) => 
                           nextA_58_port, plus4A_out(57) => n3, plus4A_out(56) 
                           => nextA_56_port, plus4A_out(55) => nextA_55_port, 
                           plus4A_out(54) => nextA_54_port, plus4A_out(53) => 
                           nextA_53_port, plus4A_out(52) => nextA_52_port, 
                           plus4A_out(51) => nextA_51_port, plus4A_out(50) => 
                           nextA_50_port, plus4A_out(49) => nextA_49_port, 
                           plus4A_out(48) => nextA_48_port, plus4A_out(47) => 
                           nextA_47_port, plus4A_out(46) => nextA_46_port, 
                           plus4A_out(45) => nextA_45_port, plus4A_out(44) => 
                           nextA_44_port, plus4A_out(43) => nextA_43_port, 
                           plus4A_out(42) => nextA_42_port, plus4A_out(41) => 
                           nextA_41_port, plus4A_out(40) => nextA_40_port, 
                           plus4A_out(39) => nextA_39_port, plus4A_out(38) => 
                           nextA_38_port, plus4A_out(37) => nextA_37_port, 
                           plus4A_out(36) => nextA_36_port, plus4A_out(35) => 
                           nextA_35_port, plus4A_out(34) => nextA_34_port, 
                           plus4A_out(33) => nextA_33_port, plus4A_out(32) => 
                           nextA_32_port, plus4A_out(31) => nextA_31_port, 
                           plus4A_out(30) => nextA_30_port, plus4A_out(29) => 
                           nextA_29_port, plus4A_out(28) => nextA_28_port, 
                           plus4A_out(27) => nextA_27_port, plus4A_out(26) => 
                           nextA_26_port, plus4A_out(25) => nextA_25_port, 
                           plus4A_out(24) => nextA_24_port, plus4A_out(23) => 
                           nextA_23_port, plus4A_out(22) => nextA_22_port, 
                           plus4A_out(21) => nextA_21_port, plus4A_out(20) => 
                           nextA_20_port, plus4A_out(19) => nextA_19_port, 
                           plus4A_out(18) => nextA_18_port, plus4A_out(17) => 
                           nextA_17_port, plus4A_out(16) => nextA_16_port, 
                           plus4A_out(15) => nextA_15_port, plus4A_out(14) => 
                           nextA_14_port, plus4A_out(13) => nextA_13_port, 
                           plus4A_out(12) => nextA_12_port, plus4A_out(11) => 
                           nextA_11_port, plus4A_out(10) => nextA_10_port, 
                           plus4A_out(9) => nextA_9_port, plus4A_out(8) => 
                           nextA_8_port, plus4A_out(7) => nextA_7_port, 
                           plus4A_out(6) => nextA_6_port, plus4A_out(5) => 
                           nextA_5_port, plus4A_out(4) => nextA_4_port, 
                           plus4A_out(3) => nextA_3_port, plus4A_out(2) => 
                           nextA_2_port, plus4A_out(1) => nextA_1_port, 
                           plus4A_out(0) => n_3209, minus4A_out(63) => 
                           minus4A_s_63_port, minus4A_out(62) => 
                           minus4A_s_62_port, minus4A_out(61) => 
                           minus4A_s_61_port, minus4A_out(60) => 
                           minus4A_s_60_port, minus4A_out(59) => 
                           minus4A_s_59_port, minus4A_out(58) => 
                           minus4A_s_58_port, minus4A_out(57) => 
                           minus4A_s_57_port, minus4A_out(56) => 
                           minus4A_s_56_port, minus4A_out(55) => 
                           minus4A_s_55_port, minus4A_out(54) => 
                           minus4A_s_54_port, minus4A_out(53) => 
                           minus4A_s_53_port, minus4A_out(52) => 
                           minus4A_s_52_port, minus4A_out(51) => 
                           minus4A_s_51_port, minus4A_out(50) => 
                           minus4A_s_50_port, minus4A_out(49) => 
                           minus4A_s_49_port, minus4A_out(48) => 
                           minus4A_s_48_port, minus4A_out(47) => 
                           minus4A_s_47_port, minus4A_out(46) => 
                           minus4A_s_46_port, minus4A_out(45) => 
                           minus4A_s_45_port, minus4A_out(44) => 
                           minus4A_s_44_port, minus4A_out(43) => 
                           minus4A_s_43_port, minus4A_out(42) => 
                           minus4A_s_42_port, minus4A_out(41) => 
                           minus4A_s_41_port, minus4A_out(40) => 
                           minus4A_s_40_port, minus4A_out(39) => 
                           minus4A_s_39_port, minus4A_out(38) => 
                           minus4A_s_38_port, minus4A_out(37) => 
                           minus4A_s_37_port, minus4A_out(36) => 
                           minus4A_s_36_port, minus4A_out(35) => 
                           minus4A_s_35_port, minus4A_out(34) => 
                           minus4A_s_34_port, minus4A_out(33) => 
                           minus4A_s_33_port, minus4A_out(32) => 
                           minus4A_s_32_port, minus4A_out(31) => 
                           minus4A_s_31_port, minus4A_out(30) => 
                           minus4A_s_30_port, minus4A_out(29) => 
                           minus4A_s_29_port, minus4A_out(28) => 
                           minus4A_s_28_port, minus4A_out(27) => 
                           minus4A_s_27_port, minus4A_out(26) => 
                           minus4A_s_26_port, minus4A_out(25) => 
                           minus4A_s_25_port, minus4A_out(24) => 
                           minus4A_s_24_port, minus4A_out(23) => 
                           minus4A_s_23_port, minus4A_out(22) => 
                           minus4A_s_22_port, minus4A_out(21) => 
                           minus4A_s_21_port, minus4A_out(20) => 
                           minus4A_s_20_port, minus4A_out(19) => 
                           minus4A_s_19_port, minus4A_out(18) => 
                           minus4A_s_18_port, minus4A_out(17) => 
                           minus4A_s_17_port, minus4A_out(16) => 
                           minus4A_s_16_port, minus4A_out(15) => 
                           minus4A_s_15_port, minus4A_out(14) => 
                           minus4A_s_14_port, minus4A_out(13) => 
                           minus4A_s_13_port, minus4A_out(12) => 
                           minus4A_s_12_port, minus4A_out(11) => 
                           minus4A_s_11_port, minus4A_out(10) => 
                           minus4A_s_10_port, minus4A_out(9) => 
                           minus4A_s_9_port, minus4A_out(8) => minus4A_s_8_port
                           , minus4A_out(7) => minus4A_s_7_port, minus4A_out(6)
                           => minus4A_s_6_port, minus4A_out(5) => 
                           minus4A_s_5_port, minus4A_out(4) => minus4A_s_4_port
                           , minus4A_out(3) => minus4A_s_3_port, minus4A_out(2)
                           => minus4A_s_2_port, minus4A_out(1) => 
                           minus4A_s_1_port, minus4A_out(0) => minus4A_s_0_port
                           );
   mux_1 : MUX_GENERIC_N64_RADIX3_12 port map( plusA(63) => plus2A_s_63_port, 
                           plusA(62) => plus2A_s_62_port, plusA(61) => 
                           plus2A_s_61_port, plusA(60) => plus2A_s_60_port, 
                           plusA(59) => plus2A_s_59_port, plusA(58) => 
                           plus2A_s_58_port, plusA(57) => plus2A_s_57_port, 
                           plusA(56) => plus2A_s_56_port, plusA(55) => 
                           plus2A_s_55_port, plusA(54) => plus2A_s_54_port, 
                           plusA(53) => plus2A_s_53_port, plusA(52) => 
                           plus2A_s_52_port, plusA(51) => plus2A_s_51_port, 
                           plusA(50) => plus2A_s_50_port, plusA(49) => 
                           plus2A_s_49_port, plusA(48) => plus2A_s_48_port, 
                           plusA(47) => plus2A_s_47_port, plusA(46) => 
                           plus2A_s_46_port, plusA(45) => plus2A_s_45_port, 
                           plusA(44) => plus2A_s_44_port, plusA(43) => 
                           plus2A_s_43_port, plusA(42) => plus2A_s_42_port, 
                           plusA(41) => plus2A_s_41_port, plusA(40) => 
                           plus2A_s_40_port, plusA(39) => plus2A_s_39_port, 
                           plusA(38) => plus2A_s_38_port, plusA(37) => 
                           plus2A_s_37_port, plusA(36) => plus2A_s_36_port, 
                           plusA(35) => plus2A_s_35_port, plusA(34) => 
                           plus2A_s_34_port, plusA(33) => plus2A_s_33_port, 
                           plusA(32) => plus2A_s_32_port, plusA(31) => 
                           plus2A_s_31_port, plusA(30) => plus2A_s_30_port, 
                           plusA(29) => plus2A_s_29_port, plusA(28) => 
                           plus2A_s_28_port, plusA(27) => plus2A_s_27_port, 
                           plusA(26) => plus2A_s_26_port, plusA(25) => 
                           plus2A_s_25_port, plusA(24) => plus2A_s_24_port, 
                           plusA(23) => plus2A_s_23_port, plusA(22) => 
                           plus2A_s_22_port, plusA(21) => plus2A_s_21_port, 
                           plusA(20) => plus2A_s_20_port, plusA(19) => 
                           plus2A_s_19_port, plusA(18) => plus2A_s_18_port, 
                           plusA(17) => plus2A_s_17_port, plusA(16) => 
                           plus2A_s_16_port, plusA(15) => plus2A_s_15_port, 
                           plusA(14) => plus2A_s_14_port, plusA(13) => 
                           plus2A_s_13_port, plusA(12) => plus2A_s_12_port, 
                           plusA(11) => plus2A_s_11_port, plusA(10) => 
                           plus2A_s_10_port, plusA(9) => plus2A_s_9_port, 
                           plusA(8) => plus2A_s_8_port, plusA(7) => 
                           plus2A_s_7_port, plusA(6) => plus2A_s_6_port, 
                           plusA(5) => plus2A_s_5_port, plusA(4) => 
                           plus2A_s_4_port, plusA(3) => plus2A_s_3_port, 
                           plusA(2) => plus2A_s_2_port, plusA(1) => 
                           plus2A_s_1_port, plusA(0) => nextA_0_port, 
                           minusA(63) => minus2A_s_63_port, minusA(62) => 
                           minus2A_s_62_port, minusA(61) => minus2A_s_61_port, 
                           minusA(60) => minus2A_s_60_port, minusA(59) => 
                           minus2A_s_59_port, minusA(58) => minus2A_s_58_port, 
                           minusA(57) => minus2A_s_57_port, minusA(56) => 
                           minus2A_s_56_port, minusA(55) => minus2A_s_55_port, 
                           minusA(54) => minus2A_s_54_port, minusA(53) => 
                           minus2A_s_53_port, minusA(52) => minus2A_s_52_port, 
                           minusA(51) => minus2A_s_51_port, minusA(50) => 
                           minus2A_s_50_port, minusA(49) => minus2A_s_49_port, 
                           minusA(48) => minus2A_s_48_port, minusA(47) => 
                           minus2A_s_47_port, minusA(46) => minus2A_s_46_port, 
                           minusA(45) => minus2A_s_45_port, minusA(44) => 
                           minus2A_s_44_port, minusA(43) => minus2A_s_43_port, 
                           minusA(42) => minus2A_s_42_port, minusA(41) => 
                           minus2A_s_41_port, minusA(40) => minus2A_s_40_port, 
                           minusA(39) => minus2A_s_39_port, minusA(38) => 
                           minus2A_s_38_port, minusA(37) => minus2A_s_37_port, 
                           minusA(36) => minus2A_s_36_port, minusA(35) => 
                           minus2A_s_35_port, minusA(34) => minus2A_s_34_port, 
                           minusA(33) => minus2A_s_33_port, minusA(32) => 
                           minus2A_s_32_port, minusA(31) => minus2A_s_31_port, 
                           minusA(30) => minus2A_s_30_port, minusA(29) => 
                           minus2A_s_29_port, minusA(28) => minus2A_s_28_port, 
                           minusA(27) => minus2A_s_27_port, minusA(26) => 
                           minus2A_s_26_port, minusA(25) => minus2A_s_25_port, 
                           minusA(24) => minus2A_s_24_port, minusA(23) => 
                           minus2A_s_23_port, minusA(22) => minus2A_s_22_port, 
                           minusA(21) => minus2A_s_21_port, minusA(20) => 
                           minus2A_s_20_port, minusA(19) => minus2A_s_19_port, 
                           minusA(18) => minus2A_s_18_port, minusA(17) => 
                           minus2A_s_17_port, minusA(16) => minus2A_s_16_port, 
                           minusA(15) => minus2A_s_15_port, minusA(14) => 
                           minus2A_s_14_port, minusA(13) => minus2A_s_13_port, 
                           minusA(12) => minus2A_s_12_port, minusA(11) => 
                           minus2A_s_11_port, minusA(10) => minus2A_s_10_port, 
                           minusA(9) => minus2A_s_9_port, minusA(8) => 
                           minus2A_s_8_port, minusA(7) => minus2A_s_7_port, 
                           minusA(6) => minus2A_s_6_port, minusA(5) => 
                           minus2A_s_5_port, minusA(4) => minus2A_s_4_port, 
                           minusA(3) => minus2A_s_3_port, minusA(2) => 
                           minus2A_s_2_port, minusA(1) => minus2A_s_1_port, 
                           minusA(0) => minus2A_s_0_port, plus2A(63) => 
                           nextA_63_port, plus2A(62) => nextA_62_port, 
                           plus2A(61) => nextA_61_port, plus2A(60) => 
                           nextA_60_port, plus2A(59) => nextA_59_port, 
                           plus2A(58) => nextA_58_port, plus2A(57) => 
                           nextA_57_port, plus2A(56) => nextA_56_port, 
                           plus2A(55) => nextA_55_port, plus2A(54) => 
                           nextA_54_port, plus2A(53) => nextA_53_port, 
                           plus2A(52) => nextA_52_port, plus2A(51) => 
                           nextA_51_port, plus2A(50) => nextA_50_port, 
                           plus2A(49) => nextA_49_port, plus2A(48) => 
                           nextA_48_port, plus2A(47) => nextA_47_port, 
                           plus2A(46) => nextA_46_port, plus2A(45) => 
                           nextA_45_port, plus2A(44) => nextA_44_port, 
                           plus2A(43) => nextA_43_port, plus2A(42) => 
                           nextA_42_port, plus2A(41) => nextA_41_port, 
                           plus2A(40) => nextA_40_port, plus2A(39) => 
                           nextA_39_port, plus2A(38) => nextA_38_port, 
                           plus2A(37) => nextA_37_port, plus2A(36) => 
                           nextA_36_port, plus2A(35) => nextA_35_port, 
                           plus2A(34) => nextA_34_port, plus2A(33) => 
                           nextA_33_port, plus2A(32) => nextA_32_port, 
                           plus2A(31) => nextA_31_port, plus2A(30) => 
                           nextA_30_port, plus2A(29) => nextA_29_port, 
                           plus2A(28) => nextA_28_port, plus2A(27) => 
                           nextA_27_port, plus2A(26) => nextA_26_port, 
                           plus2A(25) => nextA_25_port, plus2A(24) => 
                           nextA_24_port, plus2A(23) => nextA_23_port, 
                           plus2A(22) => nextA_22_port, plus2A(21) => 
                           nextA_21_port, plus2A(20) => nextA_20_port, 
                           plus2A(19) => nextA_19_port, plus2A(18) => 
                           nextA_18_port, plus2A(17) => nextA_17_port, 
                           plus2A(16) => nextA_16_port, plus2A(15) => 
                           nextA_15_port, plus2A(14) => nextA_14_port, 
                           plus2A(13) => nextA_13_port, plus2A(12) => 
                           nextA_12_port, plus2A(11) => nextA_11_port, 
                           plus2A(10) => nextA_10_port, plus2A(9) => 
                           nextA_9_port, plus2A(8) => nextA_8_port, plus2A(7) 
                           => nextA_7_port, plus2A(6) => nextA_6_port, 
                           plus2A(5) => nextA_5_port, plus2A(4) => nextA_4_port
                           , plus2A(3) => nextA_3_port, plus2A(2) => 
                           nextA_2_port, plus2A(1) => nextA_1_port, plus2A(0) 
                           => nextA_0_port, minus2A(63) => minus4A_s_63_port, 
                           minus2A(62) => minus4A_s_62_port, minus2A(61) => 
                           minus4A_s_61_port, minus2A(60) => minus4A_s_60_port,
                           minus2A(59) => minus4A_s_59_port, minus2A(58) => 
                           minus4A_s_58_port, minus2A(57) => minus4A_s_57_port,
                           minus2A(56) => minus4A_s_56_port, minus2A(55) => 
                           minus4A_s_55_port, minus2A(54) => minus4A_s_54_port,
                           minus2A(53) => minus4A_s_53_port, minus2A(52) => 
                           minus4A_s_52_port, minus2A(51) => minus4A_s_51_port,
                           minus2A(50) => minus4A_s_50_port, minus2A(49) => 
                           minus4A_s_49_port, minus2A(48) => minus4A_s_48_port,
                           minus2A(47) => minus4A_s_47_port, minus2A(46) => 
                           minus4A_s_46_port, minus2A(45) => minus4A_s_45_port,
                           minus2A(44) => minus4A_s_44_port, minus2A(43) => 
                           minus4A_s_43_port, minus2A(42) => minus4A_s_42_port,
                           minus2A(41) => minus4A_s_41_port, minus2A(40) => 
                           minus4A_s_40_port, minus2A(39) => minus4A_s_39_port,
                           minus2A(38) => minus4A_s_38_port, minus2A(37) => 
                           minus4A_s_37_port, minus2A(36) => minus4A_s_36_port,
                           minus2A(35) => minus4A_s_35_port, minus2A(34) => 
                           minus4A_s_34_port, minus2A(33) => minus4A_s_33_port,
                           minus2A(32) => minus4A_s_32_port, minus2A(31) => 
                           minus4A_s_31_port, minus2A(30) => minus4A_s_30_port,
                           minus2A(29) => minus4A_s_29_port, minus2A(28) => 
                           minus4A_s_28_port, minus2A(27) => minus4A_s_27_port,
                           minus2A(26) => minus4A_s_26_port, minus2A(25) => 
                           minus4A_s_25_port, minus2A(24) => minus4A_s_24_port,
                           minus2A(23) => minus4A_s_23_port, minus2A(22) => 
                           minus4A_s_22_port, minus2A(21) => minus4A_s_21_port,
                           minus2A(20) => minus4A_s_20_port, minus2A(19) => 
                           minus4A_s_19_port, minus2A(18) => minus4A_s_18_port,
                           minus2A(17) => minus4A_s_17_port, minus2A(16) => 
                           minus4A_s_16_port, minus2A(15) => minus4A_s_15_port,
                           minus2A(14) => minus4A_s_14_port, minus2A(13) => 
                           minus4A_s_13_port, minus2A(12) => minus4A_s_12_port,
                           minus2A(11) => minus4A_s_11_port, minus2A(10) => 
                           minus4A_s_10_port, minus2A(9) => minus4A_s_9_port, 
                           minus2A(8) => minus4A_s_8_port, minus2A(7) => 
                           minus4A_s_7_port, minus2A(6) => minus4A_s_6_port, 
                           minus2A(5) => minus4A_s_5_port, minus2A(4) => 
                           minus4A_s_4_port, minus2A(3) => minus4A_s_3_port, 
                           minus2A(2) => minus4A_s_2_port, minus2A(1) => 
                           minus4A_s_1_port, minus2A(0) => minus4A_s_0_port, 
                           SEL(2) => encoder_to_mux_2_port, SEL(1) => 
                           encoder_to_mux_1_port, SEL(0) => 
                           encoder_to_mux_0_port, Y(63) => mux_to_adder_63_port
                           , Y(62) => mux_to_adder_62_port, Y(61) => 
                           mux_to_adder_61_port, Y(60) => mux_to_adder_60_port,
                           Y(59) => mux_to_adder_59_port, Y(58) => 
                           mux_to_adder_58_port, Y(57) => mux_to_adder_57_port,
                           Y(56) => mux_to_adder_56_port, Y(55) => 
                           mux_to_adder_55_port, Y(54) => mux_to_adder_54_port,
                           Y(53) => mux_to_adder_53_port, Y(52) => 
                           mux_to_adder_52_port, Y(51) => mux_to_adder_51_port,
                           Y(50) => mux_to_adder_50_port, Y(49) => 
                           mux_to_adder_49_port, Y(48) => mux_to_adder_48_port,
                           Y(47) => mux_to_adder_47_port, Y(46) => 
                           mux_to_adder_46_port, Y(45) => mux_to_adder_45_port,
                           Y(44) => mux_to_adder_44_port, Y(43) => 
                           mux_to_adder_43_port, Y(42) => mux_to_adder_42_port,
                           Y(41) => mux_to_adder_41_port, Y(40) => 
                           mux_to_adder_40_port, Y(39) => mux_to_adder_39_port,
                           Y(38) => mux_to_adder_38_port, Y(37) => 
                           mux_to_adder_37_port, Y(36) => mux_to_adder_36_port,
                           Y(35) => mux_to_adder_35_port, Y(34) => 
                           mux_to_adder_34_port, Y(33) => mux_to_adder_33_port,
                           Y(32) => mux_to_adder_32_port, Y(31) => 
                           mux_to_adder_31_port, Y(30) => mux_to_adder_30_port,
                           Y(29) => mux_to_adder_29_port, Y(28) => 
                           mux_to_adder_28_port, Y(27) => mux_to_adder_27_port,
                           Y(26) => mux_to_adder_26_port, Y(25) => 
                           mux_to_adder_25_port, Y(24) => mux_to_adder_24_port,
                           Y(23) => mux_to_adder_23_port, Y(22) => 
                           mux_to_adder_22_port, Y(21) => mux_to_adder_21_port,
                           Y(20) => mux_to_adder_20_port, Y(19) => 
                           mux_to_adder_19_port, Y(18) => mux_to_adder_18_port,
                           Y(17) => mux_to_adder_17_port, Y(16) => 
                           mux_to_adder_16_port, Y(15) => mux_to_adder_15_port,
                           Y(14) => mux_to_adder_14_port, Y(13) => 
                           mux_to_adder_13_port, Y(12) => mux_to_adder_12_port,
                           Y(11) => mux_to_adder_11_port, Y(10) => 
                           mux_to_adder_10_port, Y(9) => mux_to_adder_9_port, 
                           Y(8) => mux_to_adder_8_port, Y(7) => 
                           mux_to_adder_7_port, Y(6) => mux_to_adder_6_port, 
                           Y(5) => mux_to_adder_5_port, Y(4) => 
                           mux_to_adder_4_port, Y(3) => mux_to_adder_3_port, 
                           Y(2) => mux_to_adder_2_port, Y(1) => 
                           mux_to_adder_1_port, Y(0) => mux_to_adder_0_port);
   rca_1 : RCA_N64_12 port map( A(63) => mux_to_adder_63_port, A(62) => 
                           mux_to_adder_62_port, A(61) => mux_to_adder_61_port,
                           A(60) => mux_to_adder_60_port, A(59) => 
                           mux_to_adder_59_port, A(58) => mux_to_adder_58_port,
                           A(57) => mux_to_adder_57_port, A(56) => 
                           mux_to_adder_56_port, A(55) => mux_to_adder_55_port,
                           A(54) => mux_to_adder_54_port, A(53) => 
                           mux_to_adder_53_port, A(52) => mux_to_adder_52_port,
                           A(51) => mux_to_adder_51_port, A(50) => 
                           mux_to_adder_50_port, A(49) => mux_to_adder_49_port,
                           A(48) => mux_to_adder_48_port, A(47) => 
                           mux_to_adder_47_port, A(46) => mux_to_adder_46_port,
                           A(45) => mux_to_adder_45_port, A(44) => 
                           mux_to_adder_44_port, A(43) => mux_to_adder_43_port,
                           A(42) => mux_to_adder_42_port, A(41) => 
                           mux_to_adder_41_port, A(40) => mux_to_adder_40_port,
                           A(39) => mux_to_adder_39_port, A(38) => 
                           mux_to_adder_38_port, A(37) => mux_to_adder_37_port,
                           A(36) => mux_to_adder_36_port, A(35) => 
                           mux_to_adder_35_port, A(34) => mux_to_adder_34_port,
                           A(33) => mux_to_adder_33_port, A(32) => 
                           mux_to_adder_32_port, A(31) => mux_to_adder_31_port,
                           A(30) => mux_to_adder_30_port, A(29) => 
                           mux_to_adder_29_port, A(28) => mux_to_adder_28_port,
                           A(27) => mux_to_adder_27_port, A(26) => 
                           mux_to_adder_26_port, A(25) => mux_to_adder_25_port,
                           A(24) => mux_to_adder_24_port, A(23) => 
                           mux_to_adder_23_port, A(22) => mux_to_adder_22_port,
                           A(21) => mux_to_adder_21_port, A(20) => 
                           mux_to_adder_20_port, A(19) => mux_to_adder_19_port,
                           A(18) => mux_to_adder_18_port, A(17) => 
                           mux_to_adder_17_port, A(16) => mux_to_adder_16_port,
                           A(15) => mux_to_adder_15_port, A(14) => 
                           mux_to_adder_14_port, A(13) => mux_to_adder_13_port,
                           A(12) => mux_to_adder_12_port, A(11) => 
                           mux_to_adder_11_port, A(10) => mux_to_adder_10_port,
                           A(9) => mux_to_adder_9_port, A(8) => 
                           mux_to_adder_8_port, A(7) => mux_to_adder_7_port, 
                           A(6) => mux_to_adder_6_port, A(5) => 
                           mux_to_adder_5_port, A(4) => mux_to_adder_4_port, 
                           A(3) => mux_to_adder_3_port, A(2) => 
                           mux_to_adder_2_port, A(1) => mux_to_adder_1_port, 
                           A(0) => mux_to_adder_0_port, B(63) => prevSum(63), 
                           B(62) => prevSum(62), B(61) => prevSum(61), B(60) =>
                           prevSum(60), B(59) => prevSum(59), B(58) => 
                           prevSum(58), B(57) => prevSum(57), B(56) => 
                           prevSum(56), B(55) => prevSum(55), B(54) => 
                           prevSum(54), B(53) => prevSum(53), B(52) => 
                           prevSum(52), B(51) => prevSum(51), B(50) => 
                           prevSum(50), B(49) => prevSum(49), B(48) => 
                           prevSum(48), B(47) => prevSum(47), B(46) => 
                           prevSum(46), B(45) => prevSum(45), B(44) => 
                           prevSum(44), B(43) => prevSum(43), B(42) => 
                           prevSum(42), B(41) => prevSum(41), B(40) => 
                           prevSum(40), B(39) => prevSum(39), B(38) => 
                           prevSum(38), B(37) => prevSum(37), B(36) => 
                           prevSum(36), B(35) => prevSum(35), B(34) => 
                           prevSum(34), B(33) => prevSum(33), B(32) => 
                           prevSum(32), B(31) => prevSum(31), B(30) => 
                           prevSum(30), B(29) => prevSum(29), B(28) => 
                           prevSum(28), B(27) => prevSum(27), B(26) => 
                           prevSum(26), B(25) => prevSum(25), B(24) => 
                           prevSum(24), B(23) => prevSum(23), B(22) => 
                           prevSum(22), B(21) => prevSum(21), B(20) => 
                           prevSum(20), B(19) => prevSum(19), B(18) => 
                           prevSum(18), B(17) => prevSum(17), B(16) => 
                           prevSum(16), B(15) => prevSum(15), B(14) => 
                           prevSum(14), B(13) => prevSum(13), B(12) => 
                           prevSum(12), B(11) => prevSum(11), B(10) => 
                           prevSum(10), B(9) => prevSum(9), B(8) => prevSum(8),
                           B(7) => prevSum(7), B(6) => prevSum(6), B(5) => 
                           prevSum(5), B(4) => prevSum(4), B(3) => prevSum(3), 
                           B(2) => prevSum(2), B(1) => prevSum(1), B(0) => 
                           prevSum(0), Ci => X_Logic0_port, S(63) => 
                           nextSum(63), S(62) => nextSum(62), S(61) => 
                           nextSum(61), S(60) => nextSum(60), S(59) => 
                           nextSum(59), S(58) => nextSum(58), S(57) => 
                           nextSum(57), S(56) => nextSum(56), S(55) => 
                           nextSum(55), S(54) => nextSum(54), S(53) => 
                           nextSum(53), S(52) => nextSum(52), S(51) => 
                           nextSum(51), S(50) => nextSum(50), S(49) => 
                           nextSum(49), S(48) => nextSum(48), S(47) => 
                           nextSum(47), S(46) => nextSum(46), S(45) => 
                           nextSum(45), S(44) => nextSum(44), S(43) => 
                           nextSum(43), S(42) => nextSum(42), S(41) => 
                           nextSum(41), S(40) => nextSum(40), S(39) => 
                           nextSum(39), S(38) => nextSum(38), S(37) => 
                           nextSum(37), S(36) => nextSum(36), S(35) => 
                           nextSum(35), S(34) => nextSum(34), S(33) => 
                           nextSum(33), S(32) => nextSum(32), S(31) => 
                           nextSum(31), S(30) => nextSum(30), S(29) => 
                           nextSum(29), S(28) => nextSum(28), S(27) => 
                           nextSum(27), S(26) => nextSum(26), S(25) => 
                           nextSum(25), S(24) => nextSum(24), S(23) => 
                           nextSum(23), S(22) => nextSum(22), S(21) => 
                           nextSum(21), S(20) => nextSum(20), S(19) => 
                           nextSum(19), S(18) => nextSum(18), S(17) => 
                           nextSum(17), S(16) => nextSum(16), S(15) => 
                           nextSum(15), S(14) => nextSum(14), S(13) => 
                           nextSum(13), S(12) => nextSum(12), S(11) => 
                           nextSum(11), S(10) => nextSum(10), S(9) => 
                           nextSum(9), S(8) => nextSum(8), S(7) => nextSum(7), 
                           S(6) => nextSum(6), S(5) => nextSum(5), S(4) => 
                           nextSum(4), S(3) => nextSum(3), S(2) => nextSum(2), 
                           S(1) => nextSum(1), S(0) => nextSum(0), Co => n_3210
                           );
   U3 : BUF_X1 port map( A => n3, Z => nextA_57_port);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity booth_mul_row_N64_RADIX3_13 is

   port( prevA, prevSum : in std_logic_vector (63 downto 0);  encoderIn : in 
         std_logic_vector (2 downto 0);  nextA, nextSum : out std_logic_vector 
         (63 downto 0));

end booth_mul_row_N64_RADIX3_13;

architecture SYN_struct of booth_mul_row_N64_RADIX3_13 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component RCA_N64_13
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component MUX_GENERIC_N64_RADIX3_13
      port( plusA, minusA, plus2A, minus2A : in std_logic_vector (63 downto 0);
            SEL : in std_logic_vector (2 downto 0);  Y : out std_logic_vector 
            (63 downto 0));
   end component;
   
   component ShiftnCompl_N64_13
      port( plusA : in std_logic_vector (63 downto 0);  plus2A_out, minus2A_out
            , plus4A_out, minus4A_out : out std_logic_vector (63 downto 0));
   end component;
   
   component encoder_N64_RADIX3_13
      port( X : in std_logic_vector (2 downto 0);  Z : out std_logic_vector (2 
            downto 0));
   end component;
   
   signal X_Logic0_port, nextA_63_port, nextA_62_port, nextA_61_port, 
      nextA_60_port, nextA_59_port, nextA_58_port, n3, nextA_56_port, 
      nextA_55_port, nextA_54_port, nextA_53_port, nextA_52_port, nextA_51_port
      , nextA_50_port, nextA_49_port, nextA_48_port, nextA_47_port, 
      nextA_46_port, nextA_45_port, nextA_44_port, nextA_43_port, nextA_42_port
      , nextA_41_port, nextA_40_port, nextA_39_port, nextA_38_port, 
      nextA_37_port, nextA_36_port, nextA_35_port, nextA_34_port, nextA_33_port
      , nextA_32_port, nextA_31_port, nextA_30_port, nextA_29_port, 
      nextA_28_port, nextA_27_port, nextA_26_port, nextA_25_port, nextA_24_port
      , nextA_23_port, nextA_22_port, nextA_21_port, nextA_20_port, 
      nextA_19_port, nextA_18_port, nextA_17_port, nextA_16_port, nextA_15_port
      , nextA_14_port, nextA_13_port, nextA_12_port, nextA_11_port, 
      nextA_10_port, nextA_9_port, nextA_8_port, nextA_7_port, nextA_6_port, 
      nextA_5_port, nextA_4_port, nextA_3_port, nextA_2_port, nextA_1_port, 
      encoder_to_mux_2_port, encoder_to_mux_1_port, encoder_to_mux_0_port, 
      plus2A_s_63_port, plus2A_s_62_port, plus2A_s_61_port, plus2A_s_60_port, 
      plus2A_s_59_port, plus2A_s_58_port, plus2A_s_57_port, plus2A_s_56_port, 
      plus2A_s_55_port, plus2A_s_54_port, plus2A_s_53_port, plus2A_s_52_port, 
      plus2A_s_51_port, plus2A_s_50_port, plus2A_s_49_port, plus2A_s_48_port, 
      plus2A_s_47_port, plus2A_s_46_port, plus2A_s_45_port, plus2A_s_44_port, 
      plus2A_s_43_port, plus2A_s_42_port, plus2A_s_41_port, plus2A_s_40_port, 
      plus2A_s_39_port, plus2A_s_38_port, plus2A_s_37_port, plus2A_s_36_port, 
      plus2A_s_35_port, plus2A_s_34_port, plus2A_s_33_port, plus2A_s_32_port, 
      plus2A_s_31_port, plus2A_s_30_port, plus2A_s_29_port, plus2A_s_28_port, 
      plus2A_s_27_port, plus2A_s_26_port, plus2A_s_25_port, plus2A_s_24_port, 
      plus2A_s_23_port, plus2A_s_22_port, plus2A_s_21_port, plus2A_s_20_port, 
      plus2A_s_19_port, plus2A_s_18_port, plus2A_s_17_port, plus2A_s_16_port, 
      plus2A_s_15_port, plus2A_s_14_port, plus2A_s_13_port, plus2A_s_12_port, 
      plus2A_s_11_port, plus2A_s_10_port, plus2A_s_9_port, plus2A_s_8_port, 
      plus2A_s_7_port, plus2A_s_6_port, plus2A_s_5_port, plus2A_s_4_port, 
      plus2A_s_3_port, plus2A_s_2_port, plus2A_s_1_port, minus2A_s_63_port, 
      minus2A_s_62_port, minus2A_s_61_port, minus2A_s_60_port, 
      minus2A_s_59_port, minus2A_s_58_port, minus2A_s_57_port, 
      minus2A_s_56_port, minus2A_s_55_port, minus2A_s_54_port, 
      minus2A_s_53_port, minus2A_s_52_port, minus2A_s_51_port, 
      minus2A_s_50_port, minus2A_s_49_port, minus2A_s_48_port, 
      minus2A_s_47_port, minus2A_s_46_port, minus2A_s_45_port, 
      minus2A_s_44_port, minus2A_s_43_port, minus2A_s_42_port, 
      minus2A_s_41_port, minus2A_s_40_port, minus2A_s_39_port, 
      minus2A_s_38_port, minus2A_s_37_port, minus2A_s_36_port, 
      minus2A_s_35_port, minus2A_s_34_port, minus2A_s_33_port, 
      minus2A_s_32_port, minus2A_s_31_port, minus2A_s_30_port, 
      minus2A_s_29_port, minus2A_s_28_port, minus2A_s_27_port, 
      minus2A_s_26_port, minus2A_s_25_port, minus2A_s_24_port, 
      minus2A_s_23_port, minus2A_s_22_port, minus2A_s_21_port, 
      minus2A_s_20_port, minus2A_s_19_port, minus2A_s_18_port, 
      minus2A_s_17_port, minus2A_s_16_port, minus2A_s_15_port, 
      minus2A_s_14_port, minus2A_s_13_port, minus2A_s_12_port, 
      minus2A_s_11_port, minus2A_s_10_port, minus2A_s_9_port, minus2A_s_8_port,
      minus2A_s_7_port, minus2A_s_6_port, minus2A_s_5_port, minus2A_s_4_port, 
      minus2A_s_3_port, minus2A_s_2_port, minus2A_s_1_port, minus2A_s_0_port, 
      minus4A_s_63_port, minus4A_s_62_port, minus4A_s_61_port, 
      minus4A_s_60_port, minus4A_s_59_port, minus4A_s_58_port, 
      minus4A_s_57_port, minus4A_s_56_port, minus4A_s_55_port, 
      minus4A_s_54_port, minus4A_s_53_port, minus4A_s_52_port, 
      minus4A_s_51_port, minus4A_s_50_port, minus4A_s_49_port, 
      minus4A_s_48_port, minus4A_s_47_port, minus4A_s_46_port, 
      minus4A_s_45_port, minus4A_s_44_port, minus4A_s_43_port, 
      minus4A_s_42_port, minus4A_s_41_port, minus4A_s_40_port, 
      minus4A_s_39_port, minus4A_s_38_port, minus4A_s_37_port, 
      minus4A_s_36_port, minus4A_s_35_port, minus4A_s_34_port, 
      minus4A_s_33_port, minus4A_s_32_port, minus4A_s_31_port, 
      minus4A_s_30_port, minus4A_s_29_port, minus4A_s_28_port, 
      minus4A_s_27_port, minus4A_s_26_port, minus4A_s_25_port, 
      minus4A_s_24_port, minus4A_s_23_port, minus4A_s_22_port, 
      minus4A_s_21_port, minus4A_s_20_port, minus4A_s_19_port, 
      minus4A_s_18_port, minus4A_s_17_port, minus4A_s_16_port, 
      minus4A_s_15_port, minus4A_s_14_port, minus4A_s_13_port, 
      minus4A_s_12_port, minus4A_s_11_port, minus4A_s_10_port, minus4A_s_9_port
      , minus4A_s_8_port, minus4A_s_7_port, minus4A_s_6_port, minus4A_s_5_port,
      minus4A_s_4_port, minus4A_s_3_port, minus4A_s_2_port, minus4A_s_1_port, 
      minus4A_s_0_port, mux_to_adder_63_port, mux_to_adder_62_port, 
      mux_to_adder_61_port, mux_to_adder_60_port, mux_to_adder_59_port, 
      mux_to_adder_58_port, mux_to_adder_57_port, mux_to_adder_56_port, 
      mux_to_adder_55_port, mux_to_adder_54_port, mux_to_adder_53_port, 
      mux_to_adder_52_port, mux_to_adder_51_port, mux_to_adder_50_port, 
      mux_to_adder_49_port, mux_to_adder_48_port, mux_to_adder_47_port, 
      mux_to_adder_46_port, mux_to_adder_45_port, mux_to_adder_44_port, 
      mux_to_adder_43_port, mux_to_adder_42_port, mux_to_adder_41_port, 
      mux_to_adder_40_port, mux_to_adder_39_port, mux_to_adder_38_port, 
      mux_to_adder_37_port, mux_to_adder_36_port, mux_to_adder_35_port, 
      mux_to_adder_34_port, mux_to_adder_33_port, mux_to_adder_32_port, 
      mux_to_adder_31_port, mux_to_adder_30_port, mux_to_adder_29_port, 
      mux_to_adder_28_port, mux_to_adder_27_port, mux_to_adder_26_port, 
      mux_to_adder_25_port, mux_to_adder_24_port, mux_to_adder_23_port, 
      mux_to_adder_22_port, mux_to_adder_21_port, mux_to_adder_20_port, 
      mux_to_adder_19_port, mux_to_adder_18_port, mux_to_adder_17_port, 
      mux_to_adder_16_port, mux_to_adder_15_port, mux_to_adder_14_port, 
      mux_to_adder_13_port, mux_to_adder_12_port, mux_to_adder_11_port, 
      mux_to_adder_10_port, mux_to_adder_9_port, mux_to_adder_8_port, 
      mux_to_adder_7_port, mux_to_adder_6_port, mux_to_adder_5_port, 
      mux_to_adder_4_port, mux_to_adder_3_port, mux_to_adder_2_port, 
      mux_to_adder_1_port, mux_to_adder_0_port, nextA_0_port, nextA_57_port, 
      n_3211, n_3212, n_3213 : std_logic;

begin
   nextA <= ( nextA_63_port, nextA_62_port, nextA_61_port, nextA_60_port, 
      nextA_59_port, nextA_58_port, nextA_57_port, nextA_56_port, nextA_55_port
      , nextA_54_port, nextA_53_port, nextA_52_port, nextA_51_port, 
      nextA_50_port, nextA_49_port, nextA_48_port, nextA_47_port, nextA_46_port
      , nextA_45_port, nextA_44_port, nextA_43_port, nextA_42_port, 
      nextA_41_port, nextA_40_port, nextA_39_port, nextA_38_port, nextA_37_port
      , nextA_36_port, nextA_35_port, nextA_34_port, nextA_33_port, 
      nextA_32_port, nextA_31_port, nextA_30_port, nextA_29_port, nextA_28_port
      , nextA_27_port, nextA_26_port, nextA_25_port, nextA_24_port, 
      nextA_23_port, nextA_22_port, nextA_21_port, nextA_20_port, nextA_19_port
      , nextA_18_port, nextA_17_port, nextA_16_port, nextA_15_port, 
      nextA_14_port, nextA_13_port, nextA_12_port, nextA_11_port, nextA_10_port
      , nextA_9_port, nextA_8_port, nextA_7_port, nextA_6_port, nextA_5_port, 
      nextA_4_port, nextA_3_port, nextA_2_port, nextA_1_port, nextA_0_port );
   
   X_Logic0_port <= '0';
   nextA_0_port <= '0';
   encoder_1 : encoder_N64_RADIX3_13 port map( X(2) => encoderIn(2), X(1) => 
                           encoderIn(1), X(0) => encoderIn(0), Z(2) => 
                           encoder_to_mux_2_port, Z(1) => encoder_to_mux_1_port
                           , Z(0) => encoder_to_mux_0_port);
   ShiftnCompl_1 : ShiftnCompl_N64_13 port map( plusA(63) => prevA(63), 
                           plusA(62) => prevA(62), plusA(61) => prevA(61), 
                           plusA(60) => prevA(60), plusA(59) => prevA(59), 
                           plusA(58) => prevA(58), plusA(57) => prevA(57), 
                           plusA(56) => prevA(56), plusA(55) => prevA(55), 
                           plusA(54) => prevA(54), plusA(53) => prevA(53), 
                           plusA(52) => prevA(52), plusA(51) => prevA(51), 
                           plusA(50) => prevA(50), plusA(49) => prevA(49), 
                           plusA(48) => prevA(48), plusA(47) => prevA(47), 
                           plusA(46) => prevA(46), plusA(45) => prevA(45), 
                           plusA(44) => prevA(44), plusA(43) => prevA(43), 
                           plusA(42) => prevA(42), plusA(41) => prevA(41), 
                           plusA(40) => prevA(40), plusA(39) => prevA(39), 
                           plusA(38) => prevA(38), plusA(37) => prevA(37), 
                           plusA(36) => prevA(36), plusA(35) => prevA(35), 
                           plusA(34) => prevA(34), plusA(33) => prevA(33), 
                           plusA(32) => prevA(32), plusA(31) => prevA(31), 
                           plusA(30) => prevA(30), plusA(29) => prevA(29), 
                           plusA(28) => prevA(28), plusA(27) => prevA(27), 
                           plusA(26) => prevA(26), plusA(25) => prevA(25), 
                           plusA(24) => prevA(24), plusA(23) => prevA(23), 
                           plusA(22) => prevA(22), plusA(21) => prevA(21), 
                           plusA(20) => prevA(20), plusA(19) => prevA(19), 
                           plusA(18) => prevA(18), plusA(17) => prevA(17), 
                           plusA(16) => prevA(16), plusA(15) => prevA(15), 
                           plusA(14) => prevA(14), plusA(13) => prevA(13), 
                           plusA(12) => prevA(12), plusA(11) => prevA(11), 
                           plusA(10) => prevA(10), plusA(9) => prevA(9), 
                           plusA(8) => prevA(8), plusA(7) => prevA(7), plusA(6)
                           => prevA(6), plusA(5) => prevA(5), plusA(4) => 
                           prevA(4), plusA(3) => prevA(3), plusA(2) => prevA(2)
                           , plusA(1) => prevA(1), plusA(0) => prevA(0), 
                           plus2A_out(63) => plus2A_s_63_port, plus2A_out(62) 
                           => plus2A_s_62_port, plus2A_out(61) => 
                           plus2A_s_61_port, plus2A_out(60) => plus2A_s_60_port
                           , plus2A_out(59) => plus2A_s_59_port, plus2A_out(58)
                           => plus2A_s_58_port, plus2A_out(57) => 
                           plus2A_s_57_port, plus2A_out(56) => plus2A_s_56_port
                           , plus2A_out(55) => plus2A_s_55_port, plus2A_out(54)
                           => plus2A_s_54_port, plus2A_out(53) => 
                           plus2A_s_53_port, plus2A_out(52) => plus2A_s_52_port
                           , plus2A_out(51) => plus2A_s_51_port, plus2A_out(50)
                           => plus2A_s_50_port, plus2A_out(49) => 
                           plus2A_s_49_port, plus2A_out(48) => plus2A_s_48_port
                           , plus2A_out(47) => plus2A_s_47_port, plus2A_out(46)
                           => plus2A_s_46_port, plus2A_out(45) => 
                           plus2A_s_45_port, plus2A_out(44) => plus2A_s_44_port
                           , plus2A_out(43) => plus2A_s_43_port, plus2A_out(42)
                           => plus2A_s_42_port, plus2A_out(41) => 
                           plus2A_s_41_port, plus2A_out(40) => plus2A_s_40_port
                           , plus2A_out(39) => plus2A_s_39_port, plus2A_out(38)
                           => plus2A_s_38_port, plus2A_out(37) => 
                           plus2A_s_37_port, plus2A_out(36) => plus2A_s_36_port
                           , plus2A_out(35) => plus2A_s_35_port, plus2A_out(34)
                           => plus2A_s_34_port, plus2A_out(33) => 
                           plus2A_s_33_port, plus2A_out(32) => plus2A_s_32_port
                           , plus2A_out(31) => plus2A_s_31_port, plus2A_out(30)
                           => plus2A_s_30_port, plus2A_out(29) => 
                           plus2A_s_29_port, plus2A_out(28) => plus2A_s_28_port
                           , plus2A_out(27) => plus2A_s_27_port, plus2A_out(26)
                           => plus2A_s_26_port, plus2A_out(25) => 
                           plus2A_s_25_port, plus2A_out(24) => plus2A_s_24_port
                           , plus2A_out(23) => plus2A_s_23_port, plus2A_out(22)
                           => plus2A_s_22_port, plus2A_out(21) => 
                           plus2A_s_21_port, plus2A_out(20) => plus2A_s_20_port
                           , plus2A_out(19) => plus2A_s_19_port, plus2A_out(18)
                           => plus2A_s_18_port, plus2A_out(17) => 
                           plus2A_s_17_port, plus2A_out(16) => plus2A_s_16_port
                           , plus2A_out(15) => plus2A_s_15_port, plus2A_out(14)
                           => plus2A_s_14_port, plus2A_out(13) => 
                           plus2A_s_13_port, plus2A_out(12) => plus2A_s_12_port
                           , plus2A_out(11) => plus2A_s_11_port, plus2A_out(10)
                           => plus2A_s_10_port, plus2A_out(9) => 
                           plus2A_s_9_port, plus2A_out(8) => plus2A_s_8_port, 
                           plus2A_out(7) => plus2A_s_7_port, plus2A_out(6) => 
                           plus2A_s_6_port, plus2A_out(5) => plus2A_s_5_port, 
                           plus2A_out(4) => plus2A_s_4_port, plus2A_out(3) => 
                           plus2A_s_3_port, plus2A_out(2) => plus2A_s_2_port, 
                           plus2A_out(1) => plus2A_s_1_port, plus2A_out(0) => 
                           n_3211, minus2A_out(63) => minus2A_s_63_port, 
                           minus2A_out(62) => minus2A_s_62_port, 
                           minus2A_out(61) => minus2A_s_61_port, 
                           minus2A_out(60) => minus2A_s_60_port, 
                           minus2A_out(59) => minus2A_s_59_port, 
                           minus2A_out(58) => minus2A_s_58_port, 
                           minus2A_out(57) => minus2A_s_57_port, 
                           minus2A_out(56) => minus2A_s_56_port, 
                           minus2A_out(55) => minus2A_s_55_port, 
                           minus2A_out(54) => minus2A_s_54_port, 
                           minus2A_out(53) => minus2A_s_53_port, 
                           minus2A_out(52) => minus2A_s_52_port, 
                           minus2A_out(51) => minus2A_s_51_port, 
                           minus2A_out(50) => minus2A_s_50_port, 
                           minus2A_out(49) => minus2A_s_49_port, 
                           minus2A_out(48) => minus2A_s_48_port, 
                           minus2A_out(47) => minus2A_s_47_port, 
                           minus2A_out(46) => minus2A_s_46_port, 
                           minus2A_out(45) => minus2A_s_45_port, 
                           minus2A_out(44) => minus2A_s_44_port, 
                           minus2A_out(43) => minus2A_s_43_port, 
                           minus2A_out(42) => minus2A_s_42_port, 
                           minus2A_out(41) => minus2A_s_41_port, 
                           minus2A_out(40) => minus2A_s_40_port, 
                           minus2A_out(39) => minus2A_s_39_port, 
                           minus2A_out(38) => minus2A_s_38_port, 
                           minus2A_out(37) => minus2A_s_37_port, 
                           minus2A_out(36) => minus2A_s_36_port, 
                           minus2A_out(35) => minus2A_s_35_port, 
                           minus2A_out(34) => minus2A_s_34_port, 
                           minus2A_out(33) => minus2A_s_33_port, 
                           minus2A_out(32) => minus2A_s_32_port, 
                           minus2A_out(31) => minus2A_s_31_port, 
                           minus2A_out(30) => minus2A_s_30_port, 
                           minus2A_out(29) => minus2A_s_29_port, 
                           minus2A_out(28) => minus2A_s_28_port, 
                           minus2A_out(27) => minus2A_s_27_port, 
                           minus2A_out(26) => minus2A_s_26_port, 
                           minus2A_out(25) => minus2A_s_25_port, 
                           minus2A_out(24) => minus2A_s_24_port, 
                           minus2A_out(23) => minus2A_s_23_port, 
                           minus2A_out(22) => minus2A_s_22_port, 
                           minus2A_out(21) => minus2A_s_21_port, 
                           minus2A_out(20) => minus2A_s_20_port, 
                           minus2A_out(19) => minus2A_s_19_port, 
                           minus2A_out(18) => minus2A_s_18_port, 
                           minus2A_out(17) => minus2A_s_17_port, 
                           minus2A_out(16) => minus2A_s_16_port, 
                           minus2A_out(15) => minus2A_s_15_port, 
                           minus2A_out(14) => minus2A_s_14_port, 
                           minus2A_out(13) => minus2A_s_13_port, 
                           minus2A_out(12) => minus2A_s_12_port, 
                           minus2A_out(11) => minus2A_s_11_port, 
                           minus2A_out(10) => minus2A_s_10_port, minus2A_out(9)
                           => minus2A_s_9_port, minus2A_out(8) => 
                           minus2A_s_8_port, minus2A_out(7) => minus2A_s_7_port
                           , minus2A_out(6) => minus2A_s_6_port, minus2A_out(5)
                           => minus2A_s_5_port, minus2A_out(4) => 
                           minus2A_s_4_port, minus2A_out(3) => minus2A_s_3_port
                           , minus2A_out(2) => minus2A_s_2_port, minus2A_out(1)
                           => minus2A_s_1_port, minus2A_out(0) => 
                           minus2A_s_0_port, plus4A_out(63) => nextA_63_port, 
                           plus4A_out(62) => nextA_62_port, plus4A_out(61) => 
                           nextA_61_port, plus4A_out(60) => nextA_60_port, 
                           plus4A_out(59) => nextA_59_port, plus4A_out(58) => 
                           nextA_58_port, plus4A_out(57) => n3, plus4A_out(56) 
                           => nextA_56_port, plus4A_out(55) => nextA_55_port, 
                           plus4A_out(54) => nextA_54_port, plus4A_out(53) => 
                           nextA_53_port, plus4A_out(52) => nextA_52_port, 
                           plus4A_out(51) => nextA_51_port, plus4A_out(50) => 
                           nextA_50_port, plus4A_out(49) => nextA_49_port, 
                           plus4A_out(48) => nextA_48_port, plus4A_out(47) => 
                           nextA_47_port, plus4A_out(46) => nextA_46_port, 
                           plus4A_out(45) => nextA_45_port, plus4A_out(44) => 
                           nextA_44_port, plus4A_out(43) => nextA_43_port, 
                           plus4A_out(42) => nextA_42_port, plus4A_out(41) => 
                           nextA_41_port, plus4A_out(40) => nextA_40_port, 
                           plus4A_out(39) => nextA_39_port, plus4A_out(38) => 
                           nextA_38_port, plus4A_out(37) => nextA_37_port, 
                           plus4A_out(36) => nextA_36_port, plus4A_out(35) => 
                           nextA_35_port, plus4A_out(34) => nextA_34_port, 
                           plus4A_out(33) => nextA_33_port, plus4A_out(32) => 
                           nextA_32_port, plus4A_out(31) => nextA_31_port, 
                           plus4A_out(30) => nextA_30_port, plus4A_out(29) => 
                           nextA_29_port, plus4A_out(28) => nextA_28_port, 
                           plus4A_out(27) => nextA_27_port, plus4A_out(26) => 
                           nextA_26_port, plus4A_out(25) => nextA_25_port, 
                           plus4A_out(24) => nextA_24_port, plus4A_out(23) => 
                           nextA_23_port, plus4A_out(22) => nextA_22_port, 
                           plus4A_out(21) => nextA_21_port, plus4A_out(20) => 
                           nextA_20_port, plus4A_out(19) => nextA_19_port, 
                           plus4A_out(18) => nextA_18_port, plus4A_out(17) => 
                           nextA_17_port, plus4A_out(16) => nextA_16_port, 
                           plus4A_out(15) => nextA_15_port, plus4A_out(14) => 
                           nextA_14_port, plus4A_out(13) => nextA_13_port, 
                           plus4A_out(12) => nextA_12_port, plus4A_out(11) => 
                           nextA_11_port, plus4A_out(10) => nextA_10_port, 
                           plus4A_out(9) => nextA_9_port, plus4A_out(8) => 
                           nextA_8_port, plus4A_out(7) => nextA_7_port, 
                           plus4A_out(6) => nextA_6_port, plus4A_out(5) => 
                           nextA_5_port, plus4A_out(4) => nextA_4_port, 
                           plus4A_out(3) => nextA_3_port, plus4A_out(2) => 
                           nextA_2_port, plus4A_out(1) => nextA_1_port, 
                           plus4A_out(0) => n_3212, minus4A_out(63) => 
                           minus4A_s_63_port, minus4A_out(62) => 
                           minus4A_s_62_port, minus4A_out(61) => 
                           minus4A_s_61_port, minus4A_out(60) => 
                           minus4A_s_60_port, minus4A_out(59) => 
                           minus4A_s_59_port, minus4A_out(58) => 
                           minus4A_s_58_port, minus4A_out(57) => 
                           minus4A_s_57_port, minus4A_out(56) => 
                           minus4A_s_56_port, minus4A_out(55) => 
                           minus4A_s_55_port, minus4A_out(54) => 
                           minus4A_s_54_port, minus4A_out(53) => 
                           minus4A_s_53_port, minus4A_out(52) => 
                           minus4A_s_52_port, minus4A_out(51) => 
                           minus4A_s_51_port, minus4A_out(50) => 
                           minus4A_s_50_port, minus4A_out(49) => 
                           minus4A_s_49_port, minus4A_out(48) => 
                           minus4A_s_48_port, minus4A_out(47) => 
                           minus4A_s_47_port, minus4A_out(46) => 
                           minus4A_s_46_port, minus4A_out(45) => 
                           minus4A_s_45_port, minus4A_out(44) => 
                           minus4A_s_44_port, minus4A_out(43) => 
                           minus4A_s_43_port, minus4A_out(42) => 
                           minus4A_s_42_port, minus4A_out(41) => 
                           minus4A_s_41_port, minus4A_out(40) => 
                           minus4A_s_40_port, minus4A_out(39) => 
                           minus4A_s_39_port, minus4A_out(38) => 
                           minus4A_s_38_port, minus4A_out(37) => 
                           minus4A_s_37_port, minus4A_out(36) => 
                           minus4A_s_36_port, minus4A_out(35) => 
                           minus4A_s_35_port, minus4A_out(34) => 
                           minus4A_s_34_port, minus4A_out(33) => 
                           minus4A_s_33_port, minus4A_out(32) => 
                           minus4A_s_32_port, minus4A_out(31) => 
                           minus4A_s_31_port, minus4A_out(30) => 
                           minus4A_s_30_port, minus4A_out(29) => 
                           minus4A_s_29_port, minus4A_out(28) => 
                           minus4A_s_28_port, minus4A_out(27) => 
                           minus4A_s_27_port, minus4A_out(26) => 
                           minus4A_s_26_port, minus4A_out(25) => 
                           minus4A_s_25_port, minus4A_out(24) => 
                           minus4A_s_24_port, minus4A_out(23) => 
                           minus4A_s_23_port, minus4A_out(22) => 
                           minus4A_s_22_port, minus4A_out(21) => 
                           minus4A_s_21_port, minus4A_out(20) => 
                           minus4A_s_20_port, minus4A_out(19) => 
                           minus4A_s_19_port, minus4A_out(18) => 
                           minus4A_s_18_port, minus4A_out(17) => 
                           minus4A_s_17_port, minus4A_out(16) => 
                           minus4A_s_16_port, minus4A_out(15) => 
                           minus4A_s_15_port, minus4A_out(14) => 
                           minus4A_s_14_port, minus4A_out(13) => 
                           minus4A_s_13_port, minus4A_out(12) => 
                           minus4A_s_12_port, minus4A_out(11) => 
                           minus4A_s_11_port, minus4A_out(10) => 
                           minus4A_s_10_port, minus4A_out(9) => 
                           minus4A_s_9_port, minus4A_out(8) => minus4A_s_8_port
                           , minus4A_out(7) => minus4A_s_7_port, minus4A_out(6)
                           => minus4A_s_6_port, minus4A_out(5) => 
                           minus4A_s_5_port, minus4A_out(4) => minus4A_s_4_port
                           , minus4A_out(3) => minus4A_s_3_port, minus4A_out(2)
                           => minus4A_s_2_port, minus4A_out(1) => 
                           minus4A_s_1_port, minus4A_out(0) => minus4A_s_0_port
                           );
   mux_1 : MUX_GENERIC_N64_RADIX3_13 port map( plusA(63) => plus2A_s_63_port, 
                           plusA(62) => plus2A_s_62_port, plusA(61) => 
                           plus2A_s_61_port, plusA(60) => plus2A_s_60_port, 
                           plusA(59) => plus2A_s_59_port, plusA(58) => 
                           plus2A_s_58_port, plusA(57) => plus2A_s_57_port, 
                           plusA(56) => plus2A_s_56_port, plusA(55) => 
                           plus2A_s_55_port, plusA(54) => plus2A_s_54_port, 
                           plusA(53) => plus2A_s_53_port, plusA(52) => 
                           plus2A_s_52_port, plusA(51) => plus2A_s_51_port, 
                           plusA(50) => plus2A_s_50_port, plusA(49) => 
                           plus2A_s_49_port, plusA(48) => plus2A_s_48_port, 
                           plusA(47) => plus2A_s_47_port, plusA(46) => 
                           plus2A_s_46_port, plusA(45) => plus2A_s_45_port, 
                           plusA(44) => plus2A_s_44_port, plusA(43) => 
                           plus2A_s_43_port, plusA(42) => plus2A_s_42_port, 
                           plusA(41) => plus2A_s_41_port, plusA(40) => 
                           plus2A_s_40_port, plusA(39) => plus2A_s_39_port, 
                           plusA(38) => plus2A_s_38_port, plusA(37) => 
                           plus2A_s_37_port, plusA(36) => plus2A_s_36_port, 
                           plusA(35) => plus2A_s_35_port, plusA(34) => 
                           plus2A_s_34_port, plusA(33) => plus2A_s_33_port, 
                           plusA(32) => plus2A_s_32_port, plusA(31) => 
                           plus2A_s_31_port, plusA(30) => plus2A_s_30_port, 
                           plusA(29) => plus2A_s_29_port, plusA(28) => 
                           plus2A_s_28_port, plusA(27) => plus2A_s_27_port, 
                           plusA(26) => plus2A_s_26_port, plusA(25) => 
                           plus2A_s_25_port, plusA(24) => plus2A_s_24_port, 
                           plusA(23) => plus2A_s_23_port, plusA(22) => 
                           plus2A_s_22_port, plusA(21) => plus2A_s_21_port, 
                           plusA(20) => plus2A_s_20_port, plusA(19) => 
                           plus2A_s_19_port, plusA(18) => plus2A_s_18_port, 
                           plusA(17) => plus2A_s_17_port, plusA(16) => 
                           plus2A_s_16_port, plusA(15) => plus2A_s_15_port, 
                           plusA(14) => plus2A_s_14_port, plusA(13) => 
                           plus2A_s_13_port, plusA(12) => plus2A_s_12_port, 
                           plusA(11) => plus2A_s_11_port, plusA(10) => 
                           plus2A_s_10_port, plusA(9) => plus2A_s_9_port, 
                           plusA(8) => plus2A_s_8_port, plusA(7) => 
                           plus2A_s_7_port, plusA(6) => plus2A_s_6_port, 
                           plusA(5) => plus2A_s_5_port, plusA(4) => 
                           plus2A_s_4_port, plusA(3) => plus2A_s_3_port, 
                           plusA(2) => plus2A_s_2_port, plusA(1) => 
                           plus2A_s_1_port, plusA(0) => nextA_0_port, 
                           minusA(63) => minus2A_s_63_port, minusA(62) => 
                           minus2A_s_62_port, minusA(61) => minus2A_s_61_port, 
                           minusA(60) => minus2A_s_60_port, minusA(59) => 
                           minus2A_s_59_port, minusA(58) => minus2A_s_58_port, 
                           minusA(57) => minus2A_s_57_port, minusA(56) => 
                           minus2A_s_56_port, minusA(55) => minus2A_s_55_port, 
                           minusA(54) => minus2A_s_54_port, minusA(53) => 
                           minus2A_s_53_port, minusA(52) => minus2A_s_52_port, 
                           minusA(51) => minus2A_s_51_port, minusA(50) => 
                           minus2A_s_50_port, minusA(49) => minus2A_s_49_port, 
                           minusA(48) => minus2A_s_48_port, minusA(47) => 
                           minus2A_s_47_port, minusA(46) => minus2A_s_46_port, 
                           minusA(45) => minus2A_s_45_port, minusA(44) => 
                           minus2A_s_44_port, minusA(43) => minus2A_s_43_port, 
                           minusA(42) => minus2A_s_42_port, minusA(41) => 
                           minus2A_s_41_port, minusA(40) => minus2A_s_40_port, 
                           minusA(39) => minus2A_s_39_port, minusA(38) => 
                           minus2A_s_38_port, minusA(37) => minus2A_s_37_port, 
                           minusA(36) => minus2A_s_36_port, minusA(35) => 
                           minus2A_s_35_port, minusA(34) => minus2A_s_34_port, 
                           minusA(33) => minus2A_s_33_port, minusA(32) => 
                           minus2A_s_32_port, minusA(31) => minus2A_s_31_port, 
                           minusA(30) => minus2A_s_30_port, minusA(29) => 
                           minus2A_s_29_port, minusA(28) => minus2A_s_28_port, 
                           minusA(27) => minus2A_s_27_port, minusA(26) => 
                           minus2A_s_26_port, minusA(25) => minus2A_s_25_port, 
                           minusA(24) => minus2A_s_24_port, minusA(23) => 
                           minus2A_s_23_port, minusA(22) => minus2A_s_22_port, 
                           minusA(21) => minus2A_s_21_port, minusA(20) => 
                           minus2A_s_20_port, minusA(19) => minus2A_s_19_port, 
                           minusA(18) => minus2A_s_18_port, minusA(17) => 
                           minus2A_s_17_port, minusA(16) => minus2A_s_16_port, 
                           minusA(15) => minus2A_s_15_port, minusA(14) => 
                           minus2A_s_14_port, minusA(13) => minus2A_s_13_port, 
                           minusA(12) => minus2A_s_12_port, minusA(11) => 
                           minus2A_s_11_port, minusA(10) => minus2A_s_10_port, 
                           minusA(9) => minus2A_s_9_port, minusA(8) => 
                           minus2A_s_8_port, minusA(7) => minus2A_s_7_port, 
                           minusA(6) => minus2A_s_6_port, minusA(5) => 
                           minus2A_s_5_port, minusA(4) => minus2A_s_4_port, 
                           minusA(3) => minus2A_s_3_port, minusA(2) => 
                           minus2A_s_2_port, minusA(1) => minus2A_s_1_port, 
                           minusA(0) => minus2A_s_0_port, plus2A(63) => 
                           nextA_63_port, plus2A(62) => nextA_62_port, 
                           plus2A(61) => nextA_61_port, plus2A(60) => 
                           nextA_60_port, plus2A(59) => nextA_59_port, 
                           plus2A(58) => nextA_58_port, plus2A(57) => 
                           nextA_57_port, plus2A(56) => nextA_56_port, 
                           plus2A(55) => nextA_55_port, plus2A(54) => 
                           nextA_54_port, plus2A(53) => nextA_53_port, 
                           plus2A(52) => nextA_52_port, plus2A(51) => 
                           nextA_51_port, plus2A(50) => nextA_50_port, 
                           plus2A(49) => nextA_49_port, plus2A(48) => 
                           nextA_48_port, plus2A(47) => nextA_47_port, 
                           plus2A(46) => nextA_46_port, plus2A(45) => 
                           nextA_45_port, plus2A(44) => nextA_44_port, 
                           plus2A(43) => nextA_43_port, plus2A(42) => 
                           nextA_42_port, plus2A(41) => nextA_41_port, 
                           plus2A(40) => nextA_40_port, plus2A(39) => 
                           nextA_39_port, plus2A(38) => nextA_38_port, 
                           plus2A(37) => nextA_37_port, plus2A(36) => 
                           nextA_36_port, plus2A(35) => nextA_35_port, 
                           plus2A(34) => nextA_34_port, plus2A(33) => 
                           nextA_33_port, plus2A(32) => nextA_32_port, 
                           plus2A(31) => nextA_31_port, plus2A(30) => 
                           nextA_30_port, plus2A(29) => nextA_29_port, 
                           plus2A(28) => nextA_28_port, plus2A(27) => 
                           nextA_27_port, plus2A(26) => nextA_26_port, 
                           plus2A(25) => nextA_25_port, plus2A(24) => 
                           nextA_24_port, plus2A(23) => nextA_23_port, 
                           plus2A(22) => nextA_22_port, plus2A(21) => 
                           nextA_21_port, plus2A(20) => nextA_20_port, 
                           plus2A(19) => nextA_19_port, plus2A(18) => 
                           nextA_18_port, plus2A(17) => nextA_17_port, 
                           plus2A(16) => nextA_16_port, plus2A(15) => 
                           nextA_15_port, plus2A(14) => nextA_14_port, 
                           plus2A(13) => nextA_13_port, plus2A(12) => 
                           nextA_12_port, plus2A(11) => nextA_11_port, 
                           plus2A(10) => nextA_10_port, plus2A(9) => 
                           nextA_9_port, plus2A(8) => nextA_8_port, plus2A(7) 
                           => nextA_7_port, plus2A(6) => nextA_6_port, 
                           plus2A(5) => nextA_5_port, plus2A(4) => nextA_4_port
                           , plus2A(3) => nextA_3_port, plus2A(2) => 
                           nextA_2_port, plus2A(1) => nextA_1_port, plus2A(0) 
                           => nextA_0_port, minus2A(63) => minus4A_s_63_port, 
                           minus2A(62) => minus4A_s_62_port, minus2A(61) => 
                           minus4A_s_61_port, minus2A(60) => minus4A_s_60_port,
                           minus2A(59) => minus4A_s_59_port, minus2A(58) => 
                           minus4A_s_58_port, minus2A(57) => minus4A_s_57_port,
                           minus2A(56) => minus4A_s_56_port, minus2A(55) => 
                           minus4A_s_55_port, minus2A(54) => minus4A_s_54_port,
                           minus2A(53) => minus4A_s_53_port, minus2A(52) => 
                           minus4A_s_52_port, minus2A(51) => minus4A_s_51_port,
                           minus2A(50) => minus4A_s_50_port, minus2A(49) => 
                           minus4A_s_49_port, minus2A(48) => minus4A_s_48_port,
                           minus2A(47) => minus4A_s_47_port, minus2A(46) => 
                           minus4A_s_46_port, minus2A(45) => minus4A_s_45_port,
                           minus2A(44) => minus4A_s_44_port, minus2A(43) => 
                           minus4A_s_43_port, minus2A(42) => minus4A_s_42_port,
                           minus2A(41) => minus4A_s_41_port, minus2A(40) => 
                           minus4A_s_40_port, minus2A(39) => minus4A_s_39_port,
                           minus2A(38) => minus4A_s_38_port, minus2A(37) => 
                           minus4A_s_37_port, minus2A(36) => minus4A_s_36_port,
                           minus2A(35) => minus4A_s_35_port, minus2A(34) => 
                           minus4A_s_34_port, minus2A(33) => minus4A_s_33_port,
                           minus2A(32) => minus4A_s_32_port, minus2A(31) => 
                           minus4A_s_31_port, minus2A(30) => minus4A_s_30_port,
                           minus2A(29) => minus4A_s_29_port, minus2A(28) => 
                           minus4A_s_28_port, minus2A(27) => minus4A_s_27_port,
                           minus2A(26) => minus4A_s_26_port, minus2A(25) => 
                           minus4A_s_25_port, minus2A(24) => minus4A_s_24_port,
                           minus2A(23) => minus4A_s_23_port, minus2A(22) => 
                           minus4A_s_22_port, minus2A(21) => minus4A_s_21_port,
                           minus2A(20) => minus4A_s_20_port, minus2A(19) => 
                           minus4A_s_19_port, minus2A(18) => minus4A_s_18_port,
                           minus2A(17) => minus4A_s_17_port, minus2A(16) => 
                           minus4A_s_16_port, minus2A(15) => minus4A_s_15_port,
                           minus2A(14) => minus4A_s_14_port, minus2A(13) => 
                           minus4A_s_13_port, minus2A(12) => minus4A_s_12_port,
                           minus2A(11) => minus4A_s_11_port, minus2A(10) => 
                           minus4A_s_10_port, minus2A(9) => minus4A_s_9_port, 
                           minus2A(8) => minus4A_s_8_port, minus2A(7) => 
                           minus4A_s_7_port, minus2A(6) => minus4A_s_6_port, 
                           minus2A(5) => minus4A_s_5_port, minus2A(4) => 
                           minus4A_s_4_port, minus2A(3) => minus4A_s_3_port, 
                           minus2A(2) => minus4A_s_2_port, minus2A(1) => 
                           minus4A_s_1_port, minus2A(0) => minus4A_s_0_port, 
                           SEL(2) => encoder_to_mux_2_port, SEL(1) => 
                           encoder_to_mux_1_port, SEL(0) => 
                           encoder_to_mux_0_port, Y(63) => mux_to_adder_63_port
                           , Y(62) => mux_to_adder_62_port, Y(61) => 
                           mux_to_adder_61_port, Y(60) => mux_to_adder_60_port,
                           Y(59) => mux_to_adder_59_port, Y(58) => 
                           mux_to_adder_58_port, Y(57) => mux_to_adder_57_port,
                           Y(56) => mux_to_adder_56_port, Y(55) => 
                           mux_to_adder_55_port, Y(54) => mux_to_adder_54_port,
                           Y(53) => mux_to_adder_53_port, Y(52) => 
                           mux_to_adder_52_port, Y(51) => mux_to_adder_51_port,
                           Y(50) => mux_to_adder_50_port, Y(49) => 
                           mux_to_adder_49_port, Y(48) => mux_to_adder_48_port,
                           Y(47) => mux_to_adder_47_port, Y(46) => 
                           mux_to_adder_46_port, Y(45) => mux_to_adder_45_port,
                           Y(44) => mux_to_adder_44_port, Y(43) => 
                           mux_to_adder_43_port, Y(42) => mux_to_adder_42_port,
                           Y(41) => mux_to_adder_41_port, Y(40) => 
                           mux_to_adder_40_port, Y(39) => mux_to_adder_39_port,
                           Y(38) => mux_to_adder_38_port, Y(37) => 
                           mux_to_adder_37_port, Y(36) => mux_to_adder_36_port,
                           Y(35) => mux_to_adder_35_port, Y(34) => 
                           mux_to_adder_34_port, Y(33) => mux_to_adder_33_port,
                           Y(32) => mux_to_adder_32_port, Y(31) => 
                           mux_to_adder_31_port, Y(30) => mux_to_adder_30_port,
                           Y(29) => mux_to_adder_29_port, Y(28) => 
                           mux_to_adder_28_port, Y(27) => mux_to_adder_27_port,
                           Y(26) => mux_to_adder_26_port, Y(25) => 
                           mux_to_adder_25_port, Y(24) => mux_to_adder_24_port,
                           Y(23) => mux_to_adder_23_port, Y(22) => 
                           mux_to_adder_22_port, Y(21) => mux_to_adder_21_port,
                           Y(20) => mux_to_adder_20_port, Y(19) => 
                           mux_to_adder_19_port, Y(18) => mux_to_adder_18_port,
                           Y(17) => mux_to_adder_17_port, Y(16) => 
                           mux_to_adder_16_port, Y(15) => mux_to_adder_15_port,
                           Y(14) => mux_to_adder_14_port, Y(13) => 
                           mux_to_adder_13_port, Y(12) => mux_to_adder_12_port,
                           Y(11) => mux_to_adder_11_port, Y(10) => 
                           mux_to_adder_10_port, Y(9) => mux_to_adder_9_port, 
                           Y(8) => mux_to_adder_8_port, Y(7) => 
                           mux_to_adder_7_port, Y(6) => mux_to_adder_6_port, 
                           Y(5) => mux_to_adder_5_port, Y(4) => 
                           mux_to_adder_4_port, Y(3) => mux_to_adder_3_port, 
                           Y(2) => mux_to_adder_2_port, Y(1) => 
                           mux_to_adder_1_port, Y(0) => mux_to_adder_0_port);
   rca_1 : RCA_N64_13 port map( A(63) => mux_to_adder_63_port, A(62) => 
                           mux_to_adder_62_port, A(61) => mux_to_adder_61_port,
                           A(60) => mux_to_adder_60_port, A(59) => 
                           mux_to_adder_59_port, A(58) => mux_to_adder_58_port,
                           A(57) => mux_to_adder_57_port, A(56) => 
                           mux_to_adder_56_port, A(55) => mux_to_adder_55_port,
                           A(54) => mux_to_adder_54_port, A(53) => 
                           mux_to_adder_53_port, A(52) => mux_to_adder_52_port,
                           A(51) => mux_to_adder_51_port, A(50) => 
                           mux_to_adder_50_port, A(49) => mux_to_adder_49_port,
                           A(48) => mux_to_adder_48_port, A(47) => 
                           mux_to_adder_47_port, A(46) => mux_to_adder_46_port,
                           A(45) => mux_to_adder_45_port, A(44) => 
                           mux_to_adder_44_port, A(43) => mux_to_adder_43_port,
                           A(42) => mux_to_adder_42_port, A(41) => 
                           mux_to_adder_41_port, A(40) => mux_to_adder_40_port,
                           A(39) => mux_to_adder_39_port, A(38) => 
                           mux_to_adder_38_port, A(37) => mux_to_adder_37_port,
                           A(36) => mux_to_adder_36_port, A(35) => 
                           mux_to_adder_35_port, A(34) => mux_to_adder_34_port,
                           A(33) => mux_to_adder_33_port, A(32) => 
                           mux_to_adder_32_port, A(31) => mux_to_adder_31_port,
                           A(30) => mux_to_adder_30_port, A(29) => 
                           mux_to_adder_29_port, A(28) => mux_to_adder_28_port,
                           A(27) => mux_to_adder_27_port, A(26) => 
                           mux_to_adder_26_port, A(25) => mux_to_adder_25_port,
                           A(24) => mux_to_adder_24_port, A(23) => 
                           mux_to_adder_23_port, A(22) => mux_to_adder_22_port,
                           A(21) => mux_to_adder_21_port, A(20) => 
                           mux_to_adder_20_port, A(19) => mux_to_adder_19_port,
                           A(18) => mux_to_adder_18_port, A(17) => 
                           mux_to_adder_17_port, A(16) => mux_to_adder_16_port,
                           A(15) => mux_to_adder_15_port, A(14) => 
                           mux_to_adder_14_port, A(13) => mux_to_adder_13_port,
                           A(12) => mux_to_adder_12_port, A(11) => 
                           mux_to_adder_11_port, A(10) => mux_to_adder_10_port,
                           A(9) => mux_to_adder_9_port, A(8) => 
                           mux_to_adder_8_port, A(7) => mux_to_adder_7_port, 
                           A(6) => mux_to_adder_6_port, A(5) => 
                           mux_to_adder_5_port, A(4) => mux_to_adder_4_port, 
                           A(3) => mux_to_adder_3_port, A(2) => 
                           mux_to_adder_2_port, A(1) => mux_to_adder_1_port, 
                           A(0) => mux_to_adder_0_port, B(63) => prevSum(63), 
                           B(62) => prevSum(62), B(61) => prevSum(61), B(60) =>
                           prevSum(60), B(59) => prevSum(59), B(58) => 
                           prevSum(58), B(57) => prevSum(57), B(56) => 
                           prevSum(56), B(55) => prevSum(55), B(54) => 
                           prevSum(54), B(53) => prevSum(53), B(52) => 
                           prevSum(52), B(51) => prevSum(51), B(50) => 
                           prevSum(50), B(49) => prevSum(49), B(48) => 
                           prevSum(48), B(47) => prevSum(47), B(46) => 
                           prevSum(46), B(45) => prevSum(45), B(44) => 
                           prevSum(44), B(43) => prevSum(43), B(42) => 
                           prevSum(42), B(41) => prevSum(41), B(40) => 
                           prevSum(40), B(39) => prevSum(39), B(38) => 
                           prevSum(38), B(37) => prevSum(37), B(36) => 
                           prevSum(36), B(35) => prevSum(35), B(34) => 
                           prevSum(34), B(33) => prevSum(33), B(32) => 
                           prevSum(32), B(31) => prevSum(31), B(30) => 
                           prevSum(30), B(29) => prevSum(29), B(28) => 
                           prevSum(28), B(27) => prevSum(27), B(26) => 
                           prevSum(26), B(25) => prevSum(25), B(24) => 
                           prevSum(24), B(23) => prevSum(23), B(22) => 
                           prevSum(22), B(21) => prevSum(21), B(20) => 
                           prevSum(20), B(19) => prevSum(19), B(18) => 
                           prevSum(18), B(17) => prevSum(17), B(16) => 
                           prevSum(16), B(15) => prevSum(15), B(14) => 
                           prevSum(14), B(13) => prevSum(13), B(12) => 
                           prevSum(12), B(11) => prevSum(11), B(10) => 
                           prevSum(10), B(9) => prevSum(9), B(8) => prevSum(8),
                           B(7) => prevSum(7), B(6) => prevSum(6), B(5) => 
                           prevSum(5), B(4) => prevSum(4), B(3) => prevSum(3), 
                           B(2) => prevSum(2), B(1) => prevSum(1), B(0) => 
                           prevSum(0), Ci => X_Logic0_port, S(63) => 
                           nextSum(63), S(62) => nextSum(62), S(61) => 
                           nextSum(61), S(60) => nextSum(60), S(59) => 
                           nextSum(59), S(58) => nextSum(58), S(57) => 
                           nextSum(57), S(56) => nextSum(56), S(55) => 
                           nextSum(55), S(54) => nextSum(54), S(53) => 
                           nextSum(53), S(52) => nextSum(52), S(51) => 
                           nextSum(51), S(50) => nextSum(50), S(49) => 
                           nextSum(49), S(48) => nextSum(48), S(47) => 
                           nextSum(47), S(46) => nextSum(46), S(45) => 
                           nextSum(45), S(44) => nextSum(44), S(43) => 
                           nextSum(43), S(42) => nextSum(42), S(41) => 
                           nextSum(41), S(40) => nextSum(40), S(39) => 
                           nextSum(39), S(38) => nextSum(38), S(37) => 
                           nextSum(37), S(36) => nextSum(36), S(35) => 
                           nextSum(35), S(34) => nextSum(34), S(33) => 
                           nextSum(33), S(32) => nextSum(32), S(31) => 
                           nextSum(31), S(30) => nextSum(30), S(29) => 
                           nextSum(29), S(28) => nextSum(28), S(27) => 
                           nextSum(27), S(26) => nextSum(26), S(25) => 
                           nextSum(25), S(24) => nextSum(24), S(23) => 
                           nextSum(23), S(22) => nextSum(22), S(21) => 
                           nextSum(21), S(20) => nextSum(20), S(19) => 
                           nextSum(19), S(18) => nextSum(18), S(17) => 
                           nextSum(17), S(16) => nextSum(16), S(15) => 
                           nextSum(15), S(14) => nextSum(14), S(13) => 
                           nextSum(13), S(12) => nextSum(12), S(11) => 
                           nextSum(11), S(10) => nextSum(10), S(9) => 
                           nextSum(9), S(8) => nextSum(8), S(7) => nextSum(7), 
                           S(6) => nextSum(6), S(5) => nextSum(5), S(4) => 
                           nextSum(4), S(3) => nextSum(3), S(2) => nextSum(2), 
                           S(1) => nextSum(1), S(0) => nextSum(0), Co => n_3213
                           );
   U3 : BUF_X1 port map( A => n3, Z => nextA_57_port);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity booth_mul_row_N64_RADIX3_14 is

   port( prevA, prevSum : in std_logic_vector (63 downto 0);  encoderIn : in 
         std_logic_vector (2 downto 0);  nextA, nextSum : out std_logic_vector 
         (63 downto 0));

end booth_mul_row_N64_RADIX3_14;

architecture SYN_struct of booth_mul_row_N64_RADIX3_14 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component RCA_N64_14
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component MUX_GENERIC_N64_RADIX3_14
      port( plusA, minusA, plus2A, minus2A : in std_logic_vector (63 downto 0);
            SEL : in std_logic_vector (2 downto 0);  Y : out std_logic_vector 
            (63 downto 0));
   end component;
   
   component ShiftnCompl_N64_14
      port( plusA : in std_logic_vector (63 downto 0);  plus2A_out, minus2A_out
            , plus4A_out, minus4A_out : out std_logic_vector (63 downto 0));
   end component;
   
   component encoder_N64_RADIX3_14
      port( X : in std_logic_vector (2 downto 0);  Z : out std_logic_vector (2 
            downto 0));
   end component;
   
   signal X_Logic0_port, nextA_63_port, nextA_62_port, nextA_61_port, 
      nextA_60_port, nextA_59_port, nextA_58_port, n3, nextA_56_port, 
      nextA_55_port, nextA_54_port, nextA_53_port, nextA_52_port, nextA_51_port
      , nextA_50_port, nextA_49_port, nextA_48_port, nextA_47_port, 
      nextA_46_port, nextA_45_port, nextA_44_port, nextA_43_port, nextA_42_port
      , nextA_41_port, nextA_40_port, nextA_39_port, nextA_38_port, 
      nextA_37_port, nextA_36_port, nextA_35_port, nextA_34_port, nextA_33_port
      , nextA_32_port, nextA_31_port, nextA_30_port, nextA_29_port, 
      nextA_28_port, nextA_27_port, nextA_26_port, nextA_25_port, nextA_24_port
      , nextA_23_port, nextA_22_port, nextA_21_port, nextA_20_port, 
      nextA_19_port, nextA_18_port, nextA_17_port, nextA_16_port, nextA_15_port
      , nextA_14_port, nextA_13_port, nextA_12_port, nextA_11_port, 
      nextA_10_port, nextA_9_port, nextA_8_port, nextA_7_port, nextA_6_port, 
      nextA_5_port, nextA_4_port, nextA_3_port, nextA_2_port, nextA_1_port, 
      encoder_to_mux_2_port, encoder_to_mux_1_port, encoder_to_mux_0_port, 
      plus2A_s_63_port, plus2A_s_62_port, plus2A_s_61_port, plus2A_s_60_port, 
      plus2A_s_59_port, plus2A_s_58_port, plus2A_s_57_port, plus2A_s_56_port, 
      plus2A_s_55_port, plus2A_s_54_port, plus2A_s_53_port, plus2A_s_52_port, 
      plus2A_s_51_port, plus2A_s_50_port, plus2A_s_49_port, plus2A_s_48_port, 
      plus2A_s_47_port, plus2A_s_46_port, plus2A_s_45_port, plus2A_s_44_port, 
      plus2A_s_43_port, plus2A_s_42_port, plus2A_s_41_port, plus2A_s_40_port, 
      plus2A_s_39_port, plus2A_s_38_port, plus2A_s_37_port, plus2A_s_36_port, 
      plus2A_s_35_port, plus2A_s_34_port, plus2A_s_33_port, plus2A_s_32_port, 
      plus2A_s_31_port, plus2A_s_30_port, plus2A_s_29_port, plus2A_s_28_port, 
      plus2A_s_27_port, plus2A_s_26_port, plus2A_s_25_port, plus2A_s_24_port, 
      plus2A_s_23_port, plus2A_s_22_port, plus2A_s_21_port, plus2A_s_20_port, 
      plus2A_s_19_port, plus2A_s_18_port, plus2A_s_17_port, plus2A_s_16_port, 
      plus2A_s_15_port, plus2A_s_14_port, plus2A_s_13_port, plus2A_s_12_port, 
      plus2A_s_11_port, plus2A_s_10_port, plus2A_s_9_port, plus2A_s_8_port, 
      plus2A_s_7_port, plus2A_s_6_port, plus2A_s_5_port, plus2A_s_4_port, 
      plus2A_s_3_port, plus2A_s_2_port, plus2A_s_1_port, minus2A_s_63_port, 
      minus2A_s_62_port, minus2A_s_61_port, minus2A_s_60_port, 
      minus2A_s_59_port, minus2A_s_58_port, minus2A_s_57_port, 
      minus2A_s_56_port, minus2A_s_55_port, minus2A_s_54_port, 
      minus2A_s_53_port, minus2A_s_52_port, minus2A_s_51_port, 
      minus2A_s_50_port, minus2A_s_49_port, minus2A_s_48_port, 
      minus2A_s_47_port, minus2A_s_46_port, minus2A_s_45_port, 
      minus2A_s_44_port, minus2A_s_43_port, minus2A_s_42_port, 
      minus2A_s_41_port, minus2A_s_40_port, minus2A_s_39_port, 
      minus2A_s_38_port, minus2A_s_37_port, minus2A_s_36_port, 
      minus2A_s_35_port, minus2A_s_34_port, minus2A_s_33_port, 
      minus2A_s_32_port, minus2A_s_31_port, minus2A_s_30_port, 
      minus2A_s_29_port, minus2A_s_28_port, minus2A_s_27_port, 
      minus2A_s_26_port, minus2A_s_25_port, minus2A_s_24_port, 
      minus2A_s_23_port, minus2A_s_22_port, minus2A_s_21_port, 
      minus2A_s_20_port, minus2A_s_19_port, minus2A_s_18_port, 
      minus2A_s_17_port, minus2A_s_16_port, minus2A_s_15_port, 
      minus2A_s_14_port, minus2A_s_13_port, minus2A_s_12_port, 
      minus2A_s_11_port, minus2A_s_10_port, minus2A_s_9_port, minus2A_s_8_port,
      minus2A_s_7_port, minus2A_s_6_port, minus2A_s_5_port, minus2A_s_4_port, 
      minus2A_s_3_port, minus2A_s_2_port, minus2A_s_1_port, minus2A_s_0_port, 
      minus4A_s_63_port, minus4A_s_62_port, minus4A_s_61_port, 
      minus4A_s_60_port, minus4A_s_59_port, minus4A_s_58_port, 
      minus4A_s_57_port, minus4A_s_56_port, minus4A_s_55_port, 
      minus4A_s_54_port, minus4A_s_53_port, minus4A_s_52_port, 
      minus4A_s_51_port, minus4A_s_50_port, minus4A_s_49_port, 
      minus4A_s_48_port, minus4A_s_47_port, minus4A_s_46_port, 
      minus4A_s_45_port, minus4A_s_44_port, minus4A_s_43_port, 
      minus4A_s_42_port, minus4A_s_41_port, minus4A_s_40_port, 
      minus4A_s_39_port, minus4A_s_38_port, minus4A_s_37_port, 
      minus4A_s_36_port, minus4A_s_35_port, minus4A_s_34_port, 
      minus4A_s_33_port, minus4A_s_32_port, minus4A_s_31_port, 
      minus4A_s_30_port, minus4A_s_29_port, minus4A_s_28_port, 
      minus4A_s_27_port, minus4A_s_26_port, minus4A_s_25_port, 
      minus4A_s_24_port, minus4A_s_23_port, minus4A_s_22_port, 
      minus4A_s_21_port, minus4A_s_20_port, minus4A_s_19_port, 
      minus4A_s_18_port, minus4A_s_17_port, minus4A_s_16_port, 
      minus4A_s_15_port, minus4A_s_14_port, minus4A_s_13_port, 
      minus4A_s_12_port, minus4A_s_11_port, minus4A_s_10_port, minus4A_s_9_port
      , minus4A_s_8_port, minus4A_s_7_port, minus4A_s_6_port, minus4A_s_5_port,
      minus4A_s_4_port, minus4A_s_3_port, minus4A_s_2_port, minus4A_s_1_port, 
      minus4A_s_0_port, mux_to_adder_63_port, mux_to_adder_62_port, 
      mux_to_adder_61_port, mux_to_adder_60_port, mux_to_adder_59_port, 
      mux_to_adder_58_port, mux_to_adder_57_port, mux_to_adder_56_port, 
      mux_to_adder_55_port, mux_to_adder_54_port, mux_to_adder_53_port, 
      mux_to_adder_52_port, mux_to_adder_51_port, mux_to_adder_50_port, 
      mux_to_adder_49_port, mux_to_adder_48_port, mux_to_adder_47_port, 
      mux_to_adder_46_port, mux_to_adder_45_port, mux_to_adder_44_port, 
      mux_to_adder_43_port, mux_to_adder_42_port, mux_to_adder_41_port, 
      mux_to_adder_40_port, mux_to_adder_39_port, mux_to_adder_38_port, 
      mux_to_adder_37_port, mux_to_adder_36_port, mux_to_adder_35_port, 
      mux_to_adder_34_port, mux_to_adder_33_port, mux_to_adder_32_port, 
      mux_to_adder_31_port, mux_to_adder_30_port, mux_to_adder_29_port, 
      mux_to_adder_28_port, mux_to_adder_27_port, mux_to_adder_26_port, 
      mux_to_adder_25_port, mux_to_adder_24_port, mux_to_adder_23_port, 
      mux_to_adder_22_port, mux_to_adder_21_port, mux_to_adder_20_port, 
      mux_to_adder_19_port, mux_to_adder_18_port, mux_to_adder_17_port, 
      mux_to_adder_16_port, mux_to_adder_15_port, mux_to_adder_14_port, 
      mux_to_adder_13_port, mux_to_adder_12_port, mux_to_adder_11_port, 
      mux_to_adder_10_port, mux_to_adder_9_port, mux_to_adder_8_port, 
      mux_to_adder_7_port, mux_to_adder_6_port, mux_to_adder_5_port, 
      mux_to_adder_4_port, mux_to_adder_3_port, mux_to_adder_2_port, 
      mux_to_adder_1_port, mux_to_adder_0_port, nextA_0_port, nextA_57_port, 
      n_3214, n_3215, n_3216 : std_logic;

begin
   nextA <= ( nextA_63_port, nextA_62_port, nextA_61_port, nextA_60_port, 
      nextA_59_port, nextA_58_port, nextA_57_port, nextA_56_port, nextA_55_port
      , nextA_54_port, nextA_53_port, nextA_52_port, nextA_51_port, 
      nextA_50_port, nextA_49_port, nextA_48_port, nextA_47_port, nextA_46_port
      , nextA_45_port, nextA_44_port, nextA_43_port, nextA_42_port, 
      nextA_41_port, nextA_40_port, nextA_39_port, nextA_38_port, nextA_37_port
      , nextA_36_port, nextA_35_port, nextA_34_port, nextA_33_port, 
      nextA_32_port, nextA_31_port, nextA_30_port, nextA_29_port, nextA_28_port
      , nextA_27_port, nextA_26_port, nextA_25_port, nextA_24_port, 
      nextA_23_port, nextA_22_port, nextA_21_port, nextA_20_port, nextA_19_port
      , nextA_18_port, nextA_17_port, nextA_16_port, nextA_15_port, 
      nextA_14_port, nextA_13_port, nextA_12_port, nextA_11_port, nextA_10_port
      , nextA_9_port, nextA_8_port, nextA_7_port, nextA_6_port, nextA_5_port, 
      nextA_4_port, nextA_3_port, nextA_2_port, nextA_1_port, nextA_0_port );
   
   X_Logic0_port <= '0';
   nextA_0_port <= '0';
   encoder_1 : encoder_N64_RADIX3_14 port map( X(2) => encoderIn(2), X(1) => 
                           encoderIn(1), X(0) => encoderIn(0), Z(2) => 
                           encoder_to_mux_2_port, Z(1) => encoder_to_mux_1_port
                           , Z(0) => encoder_to_mux_0_port);
   ShiftnCompl_1 : ShiftnCompl_N64_14 port map( plusA(63) => prevA(63), 
                           plusA(62) => prevA(62), plusA(61) => prevA(61), 
                           plusA(60) => prevA(60), plusA(59) => prevA(59), 
                           plusA(58) => prevA(58), plusA(57) => prevA(57), 
                           plusA(56) => prevA(56), plusA(55) => prevA(55), 
                           plusA(54) => prevA(54), plusA(53) => prevA(53), 
                           plusA(52) => prevA(52), plusA(51) => prevA(51), 
                           plusA(50) => prevA(50), plusA(49) => prevA(49), 
                           plusA(48) => prevA(48), plusA(47) => prevA(47), 
                           plusA(46) => prevA(46), plusA(45) => prevA(45), 
                           plusA(44) => prevA(44), plusA(43) => prevA(43), 
                           plusA(42) => prevA(42), plusA(41) => prevA(41), 
                           plusA(40) => prevA(40), plusA(39) => prevA(39), 
                           plusA(38) => prevA(38), plusA(37) => prevA(37), 
                           plusA(36) => prevA(36), plusA(35) => prevA(35), 
                           plusA(34) => prevA(34), plusA(33) => prevA(33), 
                           plusA(32) => prevA(32), plusA(31) => prevA(31), 
                           plusA(30) => prevA(30), plusA(29) => prevA(29), 
                           plusA(28) => prevA(28), plusA(27) => prevA(27), 
                           plusA(26) => prevA(26), plusA(25) => prevA(25), 
                           plusA(24) => prevA(24), plusA(23) => prevA(23), 
                           plusA(22) => prevA(22), plusA(21) => prevA(21), 
                           plusA(20) => prevA(20), plusA(19) => prevA(19), 
                           plusA(18) => prevA(18), plusA(17) => prevA(17), 
                           plusA(16) => prevA(16), plusA(15) => prevA(15), 
                           plusA(14) => prevA(14), plusA(13) => prevA(13), 
                           plusA(12) => prevA(12), plusA(11) => prevA(11), 
                           plusA(10) => prevA(10), plusA(9) => prevA(9), 
                           plusA(8) => prevA(8), plusA(7) => prevA(7), plusA(6)
                           => prevA(6), plusA(5) => prevA(5), plusA(4) => 
                           prevA(4), plusA(3) => prevA(3), plusA(2) => prevA(2)
                           , plusA(1) => prevA(1), plusA(0) => prevA(0), 
                           plus2A_out(63) => plus2A_s_63_port, plus2A_out(62) 
                           => plus2A_s_62_port, plus2A_out(61) => 
                           plus2A_s_61_port, plus2A_out(60) => plus2A_s_60_port
                           , plus2A_out(59) => plus2A_s_59_port, plus2A_out(58)
                           => plus2A_s_58_port, plus2A_out(57) => 
                           plus2A_s_57_port, plus2A_out(56) => plus2A_s_56_port
                           , plus2A_out(55) => plus2A_s_55_port, plus2A_out(54)
                           => plus2A_s_54_port, plus2A_out(53) => 
                           plus2A_s_53_port, plus2A_out(52) => plus2A_s_52_port
                           , plus2A_out(51) => plus2A_s_51_port, plus2A_out(50)
                           => plus2A_s_50_port, plus2A_out(49) => 
                           plus2A_s_49_port, plus2A_out(48) => plus2A_s_48_port
                           , plus2A_out(47) => plus2A_s_47_port, plus2A_out(46)
                           => plus2A_s_46_port, plus2A_out(45) => 
                           plus2A_s_45_port, plus2A_out(44) => plus2A_s_44_port
                           , plus2A_out(43) => plus2A_s_43_port, plus2A_out(42)
                           => plus2A_s_42_port, plus2A_out(41) => 
                           plus2A_s_41_port, plus2A_out(40) => plus2A_s_40_port
                           , plus2A_out(39) => plus2A_s_39_port, plus2A_out(38)
                           => plus2A_s_38_port, plus2A_out(37) => 
                           plus2A_s_37_port, plus2A_out(36) => plus2A_s_36_port
                           , plus2A_out(35) => plus2A_s_35_port, plus2A_out(34)
                           => plus2A_s_34_port, plus2A_out(33) => 
                           plus2A_s_33_port, plus2A_out(32) => plus2A_s_32_port
                           , plus2A_out(31) => plus2A_s_31_port, plus2A_out(30)
                           => plus2A_s_30_port, plus2A_out(29) => 
                           plus2A_s_29_port, plus2A_out(28) => plus2A_s_28_port
                           , plus2A_out(27) => plus2A_s_27_port, plus2A_out(26)
                           => plus2A_s_26_port, plus2A_out(25) => 
                           plus2A_s_25_port, plus2A_out(24) => plus2A_s_24_port
                           , plus2A_out(23) => plus2A_s_23_port, plus2A_out(22)
                           => plus2A_s_22_port, plus2A_out(21) => 
                           plus2A_s_21_port, plus2A_out(20) => plus2A_s_20_port
                           , plus2A_out(19) => plus2A_s_19_port, plus2A_out(18)
                           => plus2A_s_18_port, plus2A_out(17) => 
                           plus2A_s_17_port, plus2A_out(16) => plus2A_s_16_port
                           , plus2A_out(15) => plus2A_s_15_port, plus2A_out(14)
                           => plus2A_s_14_port, plus2A_out(13) => 
                           plus2A_s_13_port, plus2A_out(12) => plus2A_s_12_port
                           , plus2A_out(11) => plus2A_s_11_port, plus2A_out(10)
                           => plus2A_s_10_port, plus2A_out(9) => 
                           plus2A_s_9_port, plus2A_out(8) => plus2A_s_8_port, 
                           plus2A_out(7) => plus2A_s_7_port, plus2A_out(6) => 
                           plus2A_s_6_port, plus2A_out(5) => plus2A_s_5_port, 
                           plus2A_out(4) => plus2A_s_4_port, plus2A_out(3) => 
                           plus2A_s_3_port, plus2A_out(2) => plus2A_s_2_port, 
                           plus2A_out(1) => plus2A_s_1_port, plus2A_out(0) => 
                           n_3214, minus2A_out(63) => minus2A_s_63_port, 
                           minus2A_out(62) => minus2A_s_62_port, 
                           minus2A_out(61) => minus2A_s_61_port, 
                           minus2A_out(60) => minus2A_s_60_port, 
                           minus2A_out(59) => minus2A_s_59_port, 
                           minus2A_out(58) => minus2A_s_58_port, 
                           minus2A_out(57) => minus2A_s_57_port, 
                           minus2A_out(56) => minus2A_s_56_port, 
                           minus2A_out(55) => minus2A_s_55_port, 
                           minus2A_out(54) => minus2A_s_54_port, 
                           minus2A_out(53) => minus2A_s_53_port, 
                           minus2A_out(52) => minus2A_s_52_port, 
                           minus2A_out(51) => minus2A_s_51_port, 
                           minus2A_out(50) => minus2A_s_50_port, 
                           minus2A_out(49) => minus2A_s_49_port, 
                           minus2A_out(48) => minus2A_s_48_port, 
                           minus2A_out(47) => minus2A_s_47_port, 
                           minus2A_out(46) => minus2A_s_46_port, 
                           minus2A_out(45) => minus2A_s_45_port, 
                           minus2A_out(44) => minus2A_s_44_port, 
                           minus2A_out(43) => minus2A_s_43_port, 
                           minus2A_out(42) => minus2A_s_42_port, 
                           minus2A_out(41) => minus2A_s_41_port, 
                           minus2A_out(40) => minus2A_s_40_port, 
                           minus2A_out(39) => minus2A_s_39_port, 
                           minus2A_out(38) => minus2A_s_38_port, 
                           minus2A_out(37) => minus2A_s_37_port, 
                           minus2A_out(36) => minus2A_s_36_port, 
                           minus2A_out(35) => minus2A_s_35_port, 
                           minus2A_out(34) => minus2A_s_34_port, 
                           minus2A_out(33) => minus2A_s_33_port, 
                           minus2A_out(32) => minus2A_s_32_port, 
                           minus2A_out(31) => minus2A_s_31_port, 
                           minus2A_out(30) => minus2A_s_30_port, 
                           minus2A_out(29) => minus2A_s_29_port, 
                           minus2A_out(28) => minus2A_s_28_port, 
                           minus2A_out(27) => minus2A_s_27_port, 
                           minus2A_out(26) => minus2A_s_26_port, 
                           minus2A_out(25) => minus2A_s_25_port, 
                           minus2A_out(24) => minus2A_s_24_port, 
                           minus2A_out(23) => minus2A_s_23_port, 
                           minus2A_out(22) => minus2A_s_22_port, 
                           minus2A_out(21) => minus2A_s_21_port, 
                           minus2A_out(20) => minus2A_s_20_port, 
                           minus2A_out(19) => minus2A_s_19_port, 
                           minus2A_out(18) => minus2A_s_18_port, 
                           minus2A_out(17) => minus2A_s_17_port, 
                           minus2A_out(16) => minus2A_s_16_port, 
                           minus2A_out(15) => minus2A_s_15_port, 
                           minus2A_out(14) => minus2A_s_14_port, 
                           minus2A_out(13) => minus2A_s_13_port, 
                           minus2A_out(12) => minus2A_s_12_port, 
                           minus2A_out(11) => minus2A_s_11_port, 
                           minus2A_out(10) => minus2A_s_10_port, minus2A_out(9)
                           => minus2A_s_9_port, minus2A_out(8) => 
                           minus2A_s_8_port, minus2A_out(7) => minus2A_s_7_port
                           , minus2A_out(6) => minus2A_s_6_port, minus2A_out(5)
                           => minus2A_s_5_port, minus2A_out(4) => 
                           minus2A_s_4_port, minus2A_out(3) => minus2A_s_3_port
                           , minus2A_out(2) => minus2A_s_2_port, minus2A_out(1)
                           => minus2A_s_1_port, minus2A_out(0) => 
                           minus2A_s_0_port, plus4A_out(63) => nextA_63_port, 
                           plus4A_out(62) => nextA_62_port, plus4A_out(61) => 
                           nextA_61_port, plus4A_out(60) => nextA_60_port, 
                           plus4A_out(59) => nextA_59_port, plus4A_out(58) => 
                           nextA_58_port, plus4A_out(57) => n3, plus4A_out(56) 
                           => nextA_56_port, plus4A_out(55) => nextA_55_port, 
                           plus4A_out(54) => nextA_54_port, plus4A_out(53) => 
                           nextA_53_port, plus4A_out(52) => nextA_52_port, 
                           plus4A_out(51) => nextA_51_port, plus4A_out(50) => 
                           nextA_50_port, plus4A_out(49) => nextA_49_port, 
                           plus4A_out(48) => nextA_48_port, plus4A_out(47) => 
                           nextA_47_port, plus4A_out(46) => nextA_46_port, 
                           plus4A_out(45) => nextA_45_port, plus4A_out(44) => 
                           nextA_44_port, plus4A_out(43) => nextA_43_port, 
                           plus4A_out(42) => nextA_42_port, plus4A_out(41) => 
                           nextA_41_port, plus4A_out(40) => nextA_40_port, 
                           plus4A_out(39) => nextA_39_port, plus4A_out(38) => 
                           nextA_38_port, plus4A_out(37) => nextA_37_port, 
                           plus4A_out(36) => nextA_36_port, plus4A_out(35) => 
                           nextA_35_port, plus4A_out(34) => nextA_34_port, 
                           plus4A_out(33) => nextA_33_port, plus4A_out(32) => 
                           nextA_32_port, plus4A_out(31) => nextA_31_port, 
                           plus4A_out(30) => nextA_30_port, plus4A_out(29) => 
                           nextA_29_port, plus4A_out(28) => nextA_28_port, 
                           plus4A_out(27) => nextA_27_port, plus4A_out(26) => 
                           nextA_26_port, plus4A_out(25) => nextA_25_port, 
                           plus4A_out(24) => nextA_24_port, plus4A_out(23) => 
                           nextA_23_port, plus4A_out(22) => nextA_22_port, 
                           plus4A_out(21) => nextA_21_port, plus4A_out(20) => 
                           nextA_20_port, plus4A_out(19) => nextA_19_port, 
                           plus4A_out(18) => nextA_18_port, plus4A_out(17) => 
                           nextA_17_port, plus4A_out(16) => nextA_16_port, 
                           plus4A_out(15) => nextA_15_port, plus4A_out(14) => 
                           nextA_14_port, plus4A_out(13) => nextA_13_port, 
                           plus4A_out(12) => nextA_12_port, plus4A_out(11) => 
                           nextA_11_port, plus4A_out(10) => nextA_10_port, 
                           plus4A_out(9) => nextA_9_port, plus4A_out(8) => 
                           nextA_8_port, plus4A_out(7) => nextA_7_port, 
                           plus4A_out(6) => nextA_6_port, plus4A_out(5) => 
                           nextA_5_port, plus4A_out(4) => nextA_4_port, 
                           plus4A_out(3) => nextA_3_port, plus4A_out(2) => 
                           nextA_2_port, plus4A_out(1) => nextA_1_port, 
                           plus4A_out(0) => n_3215, minus4A_out(63) => 
                           minus4A_s_63_port, minus4A_out(62) => 
                           minus4A_s_62_port, minus4A_out(61) => 
                           minus4A_s_61_port, minus4A_out(60) => 
                           minus4A_s_60_port, minus4A_out(59) => 
                           minus4A_s_59_port, minus4A_out(58) => 
                           minus4A_s_58_port, minus4A_out(57) => 
                           minus4A_s_57_port, minus4A_out(56) => 
                           minus4A_s_56_port, minus4A_out(55) => 
                           minus4A_s_55_port, minus4A_out(54) => 
                           minus4A_s_54_port, minus4A_out(53) => 
                           minus4A_s_53_port, minus4A_out(52) => 
                           minus4A_s_52_port, minus4A_out(51) => 
                           minus4A_s_51_port, minus4A_out(50) => 
                           minus4A_s_50_port, minus4A_out(49) => 
                           minus4A_s_49_port, minus4A_out(48) => 
                           minus4A_s_48_port, minus4A_out(47) => 
                           minus4A_s_47_port, minus4A_out(46) => 
                           minus4A_s_46_port, minus4A_out(45) => 
                           minus4A_s_45_port, minus4A_out(44) => 
                           minus4A_s_44_port, minus4A_out(43) => 
                           minus4A_s_43_port, minus4A_out(42) => 
                           minus4A_s_42_port, minus4A_out(41) => 
                           minus4A_s_41_port, minus4A_out(40) => 
                           minus4A_s_40_port, minus4A_out(39) => 
                           minus4A_s_39_port, minus4A_out(38) => 
                           minus4A_s_38_port, minus4A_out(37) => 
                           minus4A_s_37_port, minus4A_out(36) => 
                           minus4A_s_36_port, minus4A_out(35) => 
                           minus4A_s_35_port, minus4A_out(34) => 
                           minus4A_s_34_port, minus4A_out(33) => 
                           minus4A_s_33_port, minus4A_out(32) => 
                           minus4A_s_32_port, minus4A_out(31) => 
                           minus4A_s_31_port, minus4A_out(30) => 
                           minus4A_s_30_port, minus4A_out(29) => 
                           minus4A_s_29_port, minus4A_out(28) => 
                           minus4A_s_28_port, minus4A_out(27) => 
                           minus4A_s_27_port, minus4A_out(26) => 
                           minus4A_s_26_port, minus4A_out(25) => 
                           minus4A_s_25_port, minus4A_out(24) => 
                           minus4A_s_24_port, minus4A_out(23) => 
                           minus4A_s_23_port, minus4A_out(22) => 
                           minus4A_s_22_port, minus4A_out(21) => 
                           minus4A_s_21_port, minus4A_out(20) => 
                           minus4A_s_20_port, minus4A_out(19) => 
                           minus4A_s_19_port, minus4A_out(18) => 
                           minus4A_s_18_port, minus4A_out(17) => 
                           minus4A_s_17_port, minus4A_out(16) => 
                           minus4A_s_16_port, minus4A_out(15) => 
                           minus4A_s_15_port, minus4A_out(14) => 
                           minus4A_s_14_port, minus4A_out(13) => 
                           minus4A_s_13_port, minus4A_out(12) => 
                           minus4A_s_12_port, minus4A_out(11) => 
                           minus4A_s_11_port, minus4A_out(10) => 
                           minus4A_s_10_port, minus4A_out(9) => 
                           minus4A_s_9_port, minus4A_out(8) => minus4A_s_8_port
                           , minus4A_out(7) => minus4A_s_7_port, minus4A_out(6)
                           => minus4A_s_6_port, minus4A_out(5) => 
                           minus4A_s_5_port, minus4A_out(4) => minus4A_s_4_port
                           , minus4A_out(3) => minus4A_s_3_port, minus4A_out(2)
                           => minus4A_s_2_port, minus4A_out(1) => 
                           minus4A_s_1_port, minus4A_out(0) => minus4A_s_0_port
                           );
   mux_1 : MUX_GENERIC_N64_RADIX3_14 port map( plusA(63) => plus2A_s_63_port, 
                           plusA(62) => plus2A_s_62_port, plusA(61) => 
                           plus2A_s_61_port, plusA(60) => plus2A_s_60_port, 
                           plusA(59) => plus2A_s_59_port, plusA(58) => 
                           plus2A_s_58_port, plusA(57) => plus2A_s_57_port, 
                           plusA(56) => plus2A_s_56_port, plusA(55) => 
                           plus2A_s_55_port, plusA(54) => plus2A_s_54_port, 
                           plusA(53) => plus2A_s_53_port, plusA(52) => 
                           plus2A_s_52_port, plusA(51) => plus2A_s_51_port, 
                           plusA(50) => plus2A_s_50_port, plusA(49) => 
                           plus2A_s_49_port, plusA(48) => plus2A_s_48_port, 
                           plusA(47) => plus2A_s_47_port, plusA(46) => 
                           plus2A_s_46_port, plusA(45) => plus2A_s_45_port, 
                           plusA(44) => plus2A_s_44_port, plusA(43) => 
                           plus2A_s_43_port, plusA(42) => plus2A_s_42_port, 
                           plusA(41) => plus2A_s_41_port, plusA(40) => 
                           plus2A_s_40_port, plusA(39) => plus2A_s_39_port, 
                           plusA(38) => plus2A_s_38_port, plusA(37) => 
                           plus2A_s_37_port, plusA(36) => plus2A_s_36_port, 
                           plusA(35) => plus2A_s_35_port, plusA(34) => 
                           plus2A_s_34_port, plusA(33) => plus2A_s_33_port, 
                           plusA(32) => plus2A_s_32_port, plusA(31) => 
                           plus2A_s_31_port, plusA(30) => plus2A_s_30_port, 
                           plusA(29) => plus2A_s_29_port, plusA(28) => 
                           plus2A_s_28_port, plusA(27) => plus2A_s_27_port, 
                           plusA(26) => plus2A_s_26_port, plusA(25) => 
                           plus2A_s_25_port, plusA(24) => plus2A_s_24_port, 
                           plusA(23) => plus2A_s_23_port, plusA(22) => 
                           plus2A_s_22_port, plusA(21) => plus2A_s_21_port, 
                           plusA(20) => plus2A_s_20_port, plusA(19) => 
                           plus2A_s_19_port, plusA(18) => plus2A_s_18_port, 
                           plusA(17) => plus2A_s_17_port, plusA(16) => 
                           plus2A_s_16_port, plusA(15) => plus2A_s_15_port, 
                           plusA(14) => plus2A_s_14_port, plusA(13) => 
                           plus2A_s_13_port, plusA(12) => plus2A_s_12_port, 
                           plusA(11) => plus2A_s_11_port, plusA(10) => 
                           plus2A_s_10_port, plusA(9) => plus2A_s_9_port, 
                           plusA(8) => plus2A_s_8_port, plusA(7) => 
                           plus2A_s_7_port, plusA(6) => plus2A_s_6_port, 
                           plusA(5) => plus2A_s_5_port, plusA(4) => 
                           plus2A_s_4_port, plusA(3) => plus2A_s_3_port, 
                           plusA(2) => plus2A_s_2_port, plusA(1) => 
                           plus2A_s_1_port, plusA(0) => nextA_0_port, 
                           minusA(63) => minus2A_s_63_port, minusA(62) => 
                           minus2A_s_62_port, minusA(61) => minus2A_s_61_port, 
                           minusA(60) => minus2A_s_60_port, minusA(59) => 
                           minus2A_s_59_port, minusA(58) => minus2A_s_58_port, 
                           minusA(57) => minus2A_s_57_port, minusA(56) => 
                           minus2A_s_56_port, minusA(55) => minus2A_s_55_port, 
                           minusA(54) => minus2A_s_54_port, minusA(53) => 
                           minus2A_s_53_port, minusA(52) => minus2A_s_52_port, 
                           minusA(51) => minus2A_s_51_port, minusA(50) => 
                           minus2A_s_50_port, minusA(49) => minus2A_s_49_port, 
                           minusA(48) => minus2A_s_48_port, minusA(47) => 
                           minus2A_s_47_port, minusA(46) => minus2A_s_46_port, 
                           minusA(45) => minus2A_s_45_port, minusA(44) => 
                           minus2A_s_44_port, minusA(43) => minus2A_s_43_port, 
                           minusA(42) => minus2A_s_42_port, minusA(41) => 
                           minus2A_s_41_port, minusA(40) => minus2A_s_40_port, 
                           minusA(39) => minus2A_s_39_port, minusA(38) => 
                           minus2A_s_38_port, minusA(37) => minus2A_s_37_port, 
                           minusA(36) => minus2A_s_36_port, minusA(35) => 
                           minus2A_s_35_port, minusA(34) => minus2A_s_34_port, 
                           minusA(33) => minus2A_s_33_port, minusA(32) => 
                           minus2A_s_32_port, minusA(31) => minus2A_s_31_port, 
                           minusA(30) => minus2A_s_30_port, minusA(29) => 
                           minus2A_s_29_port, minusA(28) => minus2A_s_28_port, 
                           minusA(27) => minus2A_s_27_port, minusA(26) => 
                           minus2A_s_26_port, minusA(25) => minus2A_s_25_port, 
                           minusA(24) => minus2A_s_24_port, minusA(23) => 
                           minus2A_s_23_port, minusA(22) => minus2A_s_22_port, 
                           minusA(21) => minus2A_s_21_port, minusA(20) => 
                           minus2A_s_20_port, minusA(19) => minus2A_s_19_port, 
                           minusA(18) => minus2A_s_18_port, minusA(17) => 
                           minus2A_s_17_port, minusA(16) => minus2A_s_16_port, 
                           minusA(15) => minus2A_s_15_port, minusA(14) => 
                           minus2A_s_14_port, minusA(13) => minus2A_s_13_port, 
                           minusA(12) => minus2A_s_12_port, minusA(11) => 
                           minus2A_s_11_port, minusA(10) => minus2A_s_10_port, 
                           minusA(9) => minus2A_s_9_port, minusA(8) => 
                           minus2A_s_8_port, minusA(7) => minus2A_s_7_port, 
                           minusA(6) => minus2A_s_6_port, minusA(5) => 
                           minus2A_s_5_port, minusA(4) => minus2A_s_4_port, 
                           minusA(3) => minus2A_s_3_port, minusA(2) => 
                           minus2A_s_2_port, minusA(1) => minus2A_s_1_port, 
                           minusA(0) => minus2A_s_0_port, plus2A(63) => 
                           nextA_63_port, plus2A(62) => nextA_62_port, 
                           plus2A(61) => nextA_61_port, plus2A(60) => 
                           nextA_60_port, plus2A(59) => nextA_59_port, 
                           plus2A(58) => nextA_58_port, plus2A(57) => 
                           nextA_57_port, plus2A(56) => nextA_56_port, 
                           plus2A(55) => nextA_55_port, plus2A(54) => 
                           nextA_54_port, plus2A(53) => nextA_53_port, 
                           plus2A(52) => nextA_52_port, plus2A(51) => 
                           nextA_51_port, plus2A(50) => nextA_50_port, 
                           plus2A(49) => nextA_49_port, plus2A(48) => 
                           nextA_48_port, plus2A(47) => nextA_47_port, 
                           plus2A(46) => nextA_46_port, plus2A(45) => 
                           nextA_45_port, plus2A(44) => nextA_44_port, 
                           plus2A(43) => nextA_43_port, plus2A(42) => 
                           nextA_42_port, plus2A(41) => nextA_41_port, 
                           plus2A(40) => nextA_40_port, plus2A(39) => 
                           nextA_39_port, plus2A(38) => nextA_38_port, 
                           plus2A(37) => nextA_37_port, plus2A(36) => 
                           nextA_36_port, plus2A(35) => nextA_35_port, 
                           plus2A(34) => nextA_34_port, plus2A(33) => 
                           nextA_33_port, plus2A(32) => nextA_32_port, 
                           plus2A(31) => nextA_31_port, plus2A(30) => 
                           nextA_30_port, plus2A(29) => nextA_29_port, 
                           plus2A(28) => nextA_28_port, plus2A(27) => 
                           nextA_27_port, plus2A(26) => nextA_26_port, 
                           plus2A(25) => nextA_25_port, plus2A(24) => 
                           nextA_24_port, plus2A(23) => nextA_23_port, 
                           plus2A(22) => nextA_22_port, plus2A(21) => 
                           nextA_21_port, plus2A(20) => nextA_20_port, 
                           plus2A(19) => nextA_19_port, plus2A(18) => 
                           nextA_18_port, plus2A(17) => nextA_17_port, 
                           plus2A(16) => nextA_16_port, plus2A(15) => 
                           nextA_15_port, plus2A(14) => nextA_14_port, 
                           plus2A(13) => nextA_13_port, plus2A(12) => 
                           nextA_12_port, plus2A(11) => nextA_11_port, 
                           plus2A(10) => nextA_10_port, plus2A(9) => 
                           nextA_9_port, plus2A(8) => nextA_8_port, plus2A(7) 
                           => nextA_7_port, plus2A(6) => nextA_6_port, 
                           plus2A(5) => nextA_5_port, plus2A(4) => nextA_4_port
                           , plus2A(3) => nextA_3_port, plus2A(2) => 
                           nextA_2_port, plus2A(1) => nextA_1_port, plus2A(0) 
                           => nextA_0_port, minus2A(63) => minus4A_s_63_port, 
                           minus2A(62) => minus4A_s_62_port, minus2A(61) => 
                           minus4A_s_61_port, minus2A(60) => minus4A_s_60_port,
                           minus2A(59) => minus4A_s_59_port, minus2A(58) => 
                           minus4A_s_58_port, minus2A(57) => minus4A_s_57_port,
                           minus2A(56) => minus4A_s_56_port, minus2A(55) => 
                           minus4A_s_55_port, minus2A(54) => minus4A_s_54_port,
                           minus2A(53) => minus4A_s_53_port, minus2A(52) => 
                           minus4A_s_52_port, minus2A(51) => minus4A_s_51_port,
                           minus2A(50) => minus4A_s_50_port, minus2A(49) => 
                           minus4A_s_49_port, minus2A(48) => minus4A_s_48_port,
                           minus2A(47) => minus4A_s_47_port, minus2A(46) => 
                           minus4A_s_46_port, minus2A(45) => minus4A_s_45_port,
                           minus2A(44) => minus4A_s_44_port, minus2A(43) => 
                           minus4A_s_43_port, minus2A(42) => minus4A_s_42_port,
                           minus2A(41) => minus4A_s_41_port, minus2A(40) => 
                           minus4A_s_40_port, minus2A(39) => minus4A_s_39_port,
                           minus2A(38) => minus4A_s_38_port, minus2A(37) => 
                           minus4A_s_37_port, minus2A(36) => minus4A_s_36_port,
                           minus2A(35) => minus4A_s_35_port, minus2A(34) => 
                           minus4A_s_34_port, minus2A(33) => minus4A_s_33_port,
                           minus2A(32) => minus4A_s_32_port, minus2A(31) => 
                           minus4A_s_31_port, minus2A(30) => minus4A_s_30_port,
                           minus2A(29) => minus4A_s_29_port, minus2A(28) => 
                           minus4A_s_28_port, minus2A(27) => minus4A_s_27_port,
                           minus2A(26) => minus4A_s_26_port, minus2A(25) => 
                           minus4A_s_25_port, minus2A(24) => minus4A_s_24_port,
                           minus2A(23) => minus4A_s_23_port, minus2A(22) => 
                           minus4A_s_22_port, minus2A(21) => minus4A_s_21_port,
                           minus2A(20) => minus4A_s_20_port, minus2A(19) => 
                           minus4A_s_19_port, minus2A(18) => minus4A_s_18_port,
                           minus2A(17) => minus4A_s_17_port, minus2A(16) => 
                           minus4A_s_16_port, minus2A(15) => minus4A_s_15_port,
                           minus2A(14) => minus4A_s_14_port, minus2A(13) => 
                           minus4A_s_13_port, minus2A(12) => minus4A_s_12_port,
                           minus2A(11) => minus4A_s_11_port, minus2A(10) => 
                           minus4A_s_10_port, minus2A(9) => minus4A_s_9_port, 
                           minus2A(8) => minus4A_s_8_port, minus2A(7) => 
                           minus4A_s_7_port, minus2A(6) => minus4A_s_6_port, 
                           minus2A(5) => minus4A_s_5_port, minus2A(4) => 
                           minus4A_s_4_port, minus2A(3) => minus4A_s_3_port, 
                           minus2A(2) => minus4A_s_2_port, minus2A(1) => 
                           minus4A_s_1_port, minus2A(0) => minus4A_s_0_port, 
                           SEL(2) => encoder_to_mux_2_port, SEL(1) => 
                           encoder_to_mux_1_port, SEL(0) => 
                           encoder_to_mux_0_port, Y(63) => mux_to_adder_63_port
                           , Y(62) => mux_to_adder_62_port, Y(61) => 
                           mux_to_adder_61_port, Y(60) => mux_to_adder_60_port,
                           Y(59) => mux_to_adder_59_port, Y(58) => 
                           mux_to_adder_58_port, Y(57) => mux_to_adder_57_port,
                           Y(56) => mux_to_adder_56_port, Y(55) => 
                           mux_to_adder_55_port, Y(54) => mux_to_adder_54_port,
                           Y(53) => mux_to_adder_53_port, Y(52) => 
                           mux_to_adder_52_port, Y(51) => mux_to_adder_51_port,
                           Y(50) => mux_to_adder_50_port, Y(49) => 
                           mux_to_adder_49_port, Y(48) => mux_to_adder_48_port,
                           Y(47) => mux_to_adder_47_port, Y(46) => 
                           mux_to_adder_46_port, Y(45) => mux_to_adder_45_port,
                           Y(44) => mux_to_adder_44_port, Y(43) => 
                           mux_to_adder_43_port, Y(42) => mux_to_adder_42_port,
                           Y(41) => mux_to_adder_41_port, Y(40) => 
                           mux_to_adder_40_port, Y(39) => mux_to_adder_39_port,
                           Y(38) => mux_to_adder_38_port, Y(37) => 
                           mux_to_adder_37_port, Y(36) => mux_to_adder_36_port,
                           Y(35) => mux_to_adder_35_port, Y(34) => 
                           mux_to_adder_34_port, Y(33) => mux_to_adder_33_port,
                           Y(32) => mux_to_adder_32_port, Y(31) => 
                           mux_to_adder_31_port, Y(30) => mux_to_adder_30_port,
                           Y(29) => mux_to_adder_29_port, Y(28) => 
                           mux_to_adder_28_port, Y(27) => mux_to_adder_27_port,
                           Y(26) => mux_to_adder_26_port, Y(25) => 
                           mux_to_adder_25_port, Y(24) => mux_to_adder_24_port,
                           Y(23) => mux_to_adder_23_port, Y(22) => 
                           mux_to_adder_22_port, Y(21) => mux_to_adder_21_port,
                           Y(20) => mux_to_adder_20_port, Y(19) => 
                           mux_to_adder_19_port, Y(18) => mux_to_adder_18_port,
                           Y(17) => mux_to_adder_17_port, Y(16) => 
                           mux_to_adder_16_port, Y(15) => mux_to_adder_15_port,
                           Y(14) => mux_to_adder_14_port, Y(13) => 
                           mux_to_adder_13_port, Y(12) => mux_to_adder_12_port,
                           Y(11) => mux_to_adder_11_port, Y(10) => 
                           mux_to_adder_10_port, Y(9) => mux_to_adder_9_port, 
                           Y(8) => mux_to_adder_8_port, Y(7) => 
                           mux_to_adder_7_port, Y(6) => mux_to_adder_6_port, 
                           Y(5) => mux_to_adder_5_port, Y(4) => 
                           mux_to_adder_4_port, Y(3) => mux_to_adder_3_port, 
                           Y(2) => mux_to_adder_2_port, Y(1) => 
                           mux_to_adder_1_port, Y(0) => mux_to_adder_0_port);
   rca_1 : RCA_N64_14 port map( A(63) => mux_to_adder_63_port, A(62) => 
                           mux_to_adder_62_port, A(61) => mux_to_adder_61_port,
                           A(60) => mux_to_adder_60_port, A(59) => 
                           mux_to_adder_59_port, A(58) => mux_to_adder_58_port,
                           A(57) => mux_to_adder_57_port, A(56) => 
                           mux_to_adder_56_port, A(55) => mux_to_adder_55_port,
                           A(54) => mux_to_adder_54_port, A(53) => 
                           mux_to_adder_53_port, A(52) => mux_to_adder_52_port,
                           A(51) => mux_to_adder_51_port, A(50) => 
                           mux_to_adder_50_port, A(49) => mux_to_adder_49_port,
                           A(48) => mux_to_adder_48_port, A(47) => 
                           mux_to_adder_47_port, A(46) => mux_to_adder_46_port,
                           A(45) => mux_to_adder_45_port, A(44) => 
                           mux_to_adder_44_port, A(43) => mux_to_adder_43_port,
                           A(42) => mux_to_adder_42_port, A(41) => 
                           mux_to_adder_41_port, A(40) => mux_to_adder_40_port,
                           A(39) => mux_to_adder_39_port, A(38) => 
                           mux_to_adder_38_port, A(37) => mux_to_adder_37_port,
                           A(36) => mux_to_adder_36_port, A(35) => 
                           mux_to_adder_35_port, A(34) => mux_to_adder_34_port,
                           A(33) => mux_to_adder_33_port, A(32) => 
                           mux_to_adder_32_port, A(31) => mux_to_adder_31_port,
                           A(30) => mux_to_adder_30_port, A(29) => 
                           mux_to_adder_29_port, A(28) => mux_to_adder_28_port,
                           A(27) => mux_to_adder_27_port, A(26) => 
                           mux_to_adder_26_port, A(25) => mux_to_adder_25_port,
                           A(24) => mux_to_adder_24_port, A(23) => 
                           mux_to_adder_23_port, A(22) => mux_to_adder_22_port,
                           A(21) => mux_to_adder_21_port, A(20) => 
                           mux_to_adder_20_port, A(19) => mux_to_adder_19_port,
                           A(18) => mux_to_adder_18_port, A(17) => 
                           mux_to_adder_17_port, A(16) => mux_to_adder_16_port,
                           A(15) => mux_to_adder_15_port, A(14) => 
                           mux_to_adder_14_port, A(13) => mux_to_adder_13_port,
                           A(12) => mux_to_adder_12_port, A(11) => 
                           mux_to_adder_11_port, A(10) => mux_to_adder_10_port,
                           A(9) => mux_to_adder_9_port, A(8) => 
                           mux_to_adder_8_port, A(7) => mux_to_adder_7_port, 
                           A(6) => mux_to_adder_6_port, A(5) => 
                           mux_to_adder_5_port, A(4) => mux_to_adder_4_port, 
                           A(3) => mux_to_adder_3_port, A(2) => 
                           mux_to_adder_2_port, A(1) => mux_to_adder_1_port, 
                           A(0) => mux_to_adder_0_port, B(63) => prevSum(63), 
                           B(62) => prevSum(62), B(61) => prevSum(61), B(60) =>
                           prevSum(60), B(59) => prevSum(59), B(58) => 
                           prevSum(58), B(57) => prevSum(57), B(56) => 
                           prevSum(56), B(55) => prevSum(55), B(54) => 
                           prevSum(54), B(53) => prevSum(53), B(52) => 
                           prevSum(52), B(51) => prevSum(51), B(50) => 
                           prevSum(50), B(49) => prevSum(49), B(48) => 
                           prevSum(48), B(47) => prevSum(47), B(46) => 
                           prevSum(46), B(45) => prevSum(45), B(44) => 
                           prevSum(44), B(43) => prevSum(43), B(42) => 
                           prevSum(42), B(41) => prevSum(41), B(40) => 
                           prevSum(40), B(39) => prevSum(39), B(38) => 
                           prevSum(38), B(37) => prevSum(37), B(36) => 
                           prevSum(36), B(35) => prevSum(35), B(34) => 
                           prevSum(34), B(33) => prevSum(33), B(32) => 
                           prevSum(32), B(31) => prevSum(31), B(30) => 
                           prevSum(30), B(29) => prevSum(29), B(28) => 
                           prevSum(28), B(27) => prevSum(27), B(26) => 
                           prevSum(26), B(25) => prevSum(25), B(24) => 
                           prevSum(24), B(23) => prevSum(23), B(22) => 
                           prevSum(22), B(21) => prevSum(21), B(20) => 
                           prevSum(20), B(19) => prevSum(19), B(18) => 
                           prevSum(18), B(17) => prevSum(17), B(16) => 
                           prevSum(16), B(15) => prevSum(15), B(14) => 
                           prevSum(14), B(13) => prevSum(13), B(12) => 
                           prevSum(12), B(11) => prevSum(11), B(10) => 
                           prevSum(10), B(9) => prevSum(9), B(8) => prevSum(8),
                           B(7) => prevSum(7), B(6) => prevSum(6), B(5) => 
                           prevSum(5), B(4) => prevSum(4), B(3) => prevSum(3), 
                           B(2) => prevSum(2), B(1) => prevSum(1), B(0) => 
                           prevSum(0), Ci => X_Logic0_port, S(63) => 
                           nextSum(63), S(62) => nextSum(62), S(61) => 
                           nextSum(61), S(60) => nextSum(60), S(59) => 
                           nextSum(59), S(58) => nextSum(58), S(57) => 
                           nextSum(57), S(56) => nextSum(56), S(55) => 
                           nextSum(55), S(54) => nextSum(54), S(53) => 
                           nextSum(53), S(52) => nextSum(52), S(51) => 
                           nextSum(51), S(50) => nextSum(50), S(49) => 
                           nextSum(49), S(48) => nextSum(48), S(47) => 
                           nextSum(47), S(46) => nextSum(46), S(45) => 
                           nextSum(45), S(44) => nextSum(44), S(43) => 
                           nextSum(43), S(42) => nextSum(42), S(41) => 
                           nextSum(41), S(40) => nextSum(40), S(39) => 
                           nextSum(39), S(38) => nextSum(38), S(37) => 
                           nextSum(37), S(36) => nextSum(36), S(35) => 
                           nextSum(35), S(34) => nextSum(34), S(33) => 
                           nextSum(33), S(32) => nextSum(32), S(31) => 
                           nextSum(31), S(30) => nextSum(30), S(29) => 
                           nextSum(29), S(28) => nextSum(28), S(27) => 
                           nextSum(27), S(26) => nextSum(26), S(25) => 
                           nextSum(25), S(24) => nextSum(24), S(23) => 
                           nextSum(23), S(22) => nextSum(22), S(21) => 
                           nextSum(21), S(20) => nextSum(20), S(19) => 
                           nextSum(19), S(18) => nextSum(18), S(17) => 
                           nextSum(17), S(16) => nextSum(16), S(15) => 
                           nextSum(15), S(14) => nextSum(14), S(13) => 
                           nextSum(13), S(12) => nextSum(12), S(11) => 
                           nextSum(11), S(10) => nextSum(10), S(9) => 
                           nextSum(9), S(8) => nextSum(8), S(7) => nextSum(7), 
                           S(6) => nextSum(6), S(5) => nextSum(5), S(4) => 
                           nextSum(4), S(3) => nextSum(3), S(2) => nextSum(2), 
                           S(1) => nextSum(1), S(0) => nextSum(0), Co => n_3216
                           );
   U3 : BUF_X1 port map( A => n3, Z => nextA_57_port);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity booth_mul_row_N64_RADIX3_0 is

   port( prevA, prevSum : in std_logic_vector (63 downto 0);  encoderIn : in 
         std_logic_vector (2 downto 0);  nextA, nextSum : out std_logic_vector 
         (63 downto 0));

end booth_mul_row_N64_RADIX3_0;

architecture SYN_struct of booth_mul_row_N64_RADIX3_0 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component RCA_N64_0
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component MUX_GENERIC_N64_RADIX3_15
      port( plusA, minusA, plus2A, minus2A : in std_logic_vector (63 downto 0);
            SEL : in std_logic_vector (2 downto 0);  Y : out std_logic_vector 
            (63 downto 0));
   end component;
   
   component ShiftnCompl_N64_0
      port( plusA : in std_logic_vector (63 downto 0);  plus2A_out, minus2A_out
            , plus4A_out, minus4A_out : out std_logic_vector (63 downto 0));
   end component;
   
   component encoder_N64_RADIX3_15
      port( X : in std_logic_vector (2 downto 0);  Z : out std_logic_vector (2 
            downto 0));
   end component;
   
   signal X_Logic0_port, nextA_63_port, nextA_62_port, nextA_61_port, 
      nextA_60_port, nextA_59_port, nextA_58_port, n3, nextA_56_port, 
      nextA_55_port, nextA_54_port, nextA_53_port, nextA_52_port, nextA_51_port
      , nextA_50_port, nextA_49_port, nextA_48_port, nextA_47_port, 
      nextA_46_port, nextA_45_port, nextA_44_port, nextA_43_port, nextA_42_port
      , nextA_41_port, nextA_40_port, nextA_39_port, nextA_38_port, 
      nextA_37_port, nextA_36_port, nextA_35_port, nextA_34_port, nextA_33_port
      , nextA_32_port, nextA_31_port, nextA_30_port, nextA_29_port, 
      nextA_28_port, nextA_27_port, nextA_26_port, nextA_25_port, nextA_24_port
      , nextA_23_port, nextA_22_port, nextA_21_port, nextA_20_port, 
      nextA_19_port, nextA_18_port, nextA_17_port, nextA_16_port, nextA_15_port
      , nextA_14_port, nextA_13_port, nextA_12_port, nextA_11_port, 
      nextA_10_port, nextA_9_port, nextA_8_port, nextA_7_port, nextA_6_port, 
      nextA_5_port, nextA_4_port, nextA_3_port, nextA_2_port, nextA_1_port, 
      encoder_to_mux_2_port, encoder_to_mux_1_port, encoder_to_mux_0_port, 
      plus2A_s_63_port, plus2A_s_62_port, plus2A_s_61_port, plus2A_s_60_port, 
      plus2A_s_59_port, plus2A_s_58_port, plus2A_s_57_port, plus2A_s_56_port, 
      plus2A_s_55_port, plus2A_s_54_port, plus2A_s_53_port, plus2A_s_52_port, 
      plus2A_s_51_port, plus2A_s_50_port, plus2A_s_49_port, plus2A_s_48_port, 
      plus2A_s_47_port, plus2A_s_46_port, plus2A_s_45_port, plus2A_s_44_port, 
      plus2A_s_43_port, plus2A_s_42_port, plus2A_s_41_port, plus2A_s_40_port, 
      plus2A_s_39_port, plus2A_s_38_port, plus2A_s_37_port, plus2A_s_36_port, 
      plus2A_s_35_port, plus2A_s_34_port, plus2A_s_33_port, plus2A_s_32_port, 
      plus2A_s_31_port, plus2A_s_30_port, plus2A_s_29_port, plus2A_s_28_port, 
      plus2A_s_27_port, plus2A_s_26_port, plus2A_s_25_port, plus2A_s_24_port, 
      plus2A_s_23_port, plus2A_s_22_port, plus2A_s_21_port, plus2A_s_20_port, 
      plus2A_s_19_port, plus2A_s_18_port, plus2A_s_17_port, plus2A_s_16_port, 
      plus2A_s_15_port, plus2A_s_14_port, plus2A_s_13_port, plus2A_s_12_port, 
      plus2A_s_11_port, plus2A_s_10_port, plus2A_s_9_port, plus2A_s_8_port, 
      plus2A_s_7_port, plus2A_s_6_port, plus2A_s_5_port, plus2A_s_4_port, 
      plus2A_s_3_port, plus2A_s_2_port, plus2A_s_1_port, minus2A_s_63_port, 
      minus2A_s_62_port, minus2A_s_61_port, minus2A_s_60_port, 
      minus2A_s_59_port, minus2A_s_58_port, minus2A_s_57_port, 
      minus2A_s_56_port, minus2A_s_55_port, minus2A_s_54_port, 
      minus2A_s_53_port, minus2A_s_52_port, minus2A_s_51_port, 
      minus2A_s_50_port, minus2A_s_49_port, minus2A_s_48_port, 
      minus2A_s_47_port, minus2A_s_46_port, minus2A_s_45_port, 
      minus2A_s_44_port, minus2A_s_43_port, minus2A_s_42_port, 
      minus2A_s_41_port, minus2A_s_40_port, minus2A_s_39_port, 
      minus2A_s_38_port, minus2A_s_37_port, minus2A_s_36_port, 
      minus2A_s_35_port, minus2A_s_34_port, minus2A_s_33_port, 
      minus2A_s_32_port, minus2A_s_31_port, minus2A_s_30_port, 
      minus2A_s_29_port, minus2A_s_28_port, minus2A_s_27_port, 
      minus2A_s_26_port, minus2A_s_25_port, minus2A_s_24_port, 
      minus2A_s_23_port, minus2A_s_22_port, minus2A_s_21_port, 
      minus2A_s_20_port, minus2A_s_19_port, minus2A_s_18_port, 
      minus2A_s_17_port, minus2A_s_16_port, minus2A_s_15_port, 
      minus2A_s_14_port, minus2A_s_13_port, minus2A_s_12_port, 
      minus2A_s_11_port, minus2A_s_10_port, minus2A_s_9_port, minus2A_s_8_port,
      minus2A_s_7_port, minus2A_s_6_port, minus2A_s_5_port, minus2A_s_4_port, 
      minus2A_s_3_port, minus2A_s_2_port, minus2A_s_1_port, minus2A_s_0_port, 
      minus4A_s_63_port, minus4A_s_62_port, minus4A_s_61_port, 
      minus4A_s_60_port, minus4A_s_59_port, minus4A_s_58_port, 
      minus4A_s_57_port, minus4A_s_56_port, minus4A_s_55_port, 
      minus4A_s_54_port, minus4A_s_53_port, minus4A_s_52_port, 
      minus4A_s_51_port, minus4A_s_50_port, minus4A_s_49_port, 
      minus4A_s_48_port, minus4A_s_47_port, minus4A_s_46_port, 
      minus4A_s_45_port, minus4A_s_44_port, minus4A_s_43_port, 
      minus4A_s_42_port, minus4A_s_41_port, minus4A_s_40_port, 
      minus4A_s_39_port, minus4A_s_38_port, minus4A_s_37_port, 
      minus4A_s_36_port, minus4A_s_35_port, minus4A_s_34_port, 
      minus4A_s_33_port, minus4A_s_32_port, minus4A_s_31_port, 
      minus4A_s_30_port, minus4A_s_29_port, minus4A_s_28_port, 
      minus4A_s_27_port, minus4A_s_26_port, minus4A_s_25_port, 
      minus4A_s_24_port, minus4A_s_23_port, minus4A_s_22_port, 
      minus4A_s_21_port, minus4A_s_20_port, minus4A_s_19_port, 
      minus4A_s_18_port, minus4A_s_17_port, minus4A_s_16_port, 
      minus4A_s_15_port, minus4A_s_14_port, minus4A_s_13_port, 
      minus4A_s_12_port, minus4A_s_11_port, minus4A_s_10_port, minus4A_s_9_port
      , minus4A_s_8_port, minus4A_s_7_port, minus4A_s_6_port, minus4A_s_5_port,
      minus4A_s_4_port, minus4A_s_3_port, minus4A_s_2_port, minus4A_s_1_port, 
      minus4A_s_0_port, mux_to_adder_63_port, mux_to_adder_62_port, 
      mux_to_adder_61_port, mux_to_adder_60_port, mux_to_adder_59_port, 
      mux_to_adder_58_port, mux_to_adder_57_port, mux_to_adder_56_port, 
      mux_to_adder_55_port, mux_to_adder_54_port, mux_to_adder_53_port, 
      mux_to_adder_52_port, mux_to_adder_51_port, mux_to_adder_50_port, 
      mux_to_adder_49_port, mux_to_adder_48_port, mux_to_adder_47_port, 
      mux_to_adder_46_port, mux_to_adder_45_port, mux_to_adder_44_port, 
      mux_to_adder_43_port, mux_to_adder_42_port, mux_to_adder_41_port, 
      mux_to_adder_40_port, mux_to_adder_39_port, mux_to_adder_38_port, 
      mux_to_adder_37_port, mux_to_adder_36_port, mux_to_adder_35_port, 
      mux_to_adder_34_port, mux_to_adder_33_port, mux_to_adder_32_port, 
      mux_to_adder_31_port, mux_to_adder_30_port, mux_to_adder_29_port, 
      mux_to_adder_28_port, mux_to_adder_27_port, mux_to_adder_26_port, 
      mux_to_adder_25_port, mux_to_adder_24_port, mux_to_adder_23_port, 
      mux_to_adder_22_port, mux_to_adder_21_port, mux_to_adder_20_port, 
      mux_to_adder_19_port, mux_to_adder_18_port, mux_to_adder_17_port, 
      mux_to_adder_16_port, mux_to_adder_15_port, mux_to_adder_14_port, 
      mux_to_adder_13_port, mux_to_adder_12_port, mux_to_adder_11_port, 
      mux_to_adder_10_port, mux_to_adder_9_port, mux_to_adder_8_port, 
      mux_to_adder_7_port, mux_to_adder_6_port, mux_to_adder_5_port, 
      mux_to_adder_4_port, mux_to_adder_3_port, mux_to_adder_2_port, 
      mux_to_adder_1_port, mux_to_adder_0_port, nextA_0_port, nextA_57_port, 
      n_3217, n_3218, n_3219 : std_logic;

begin
   nextA <= ( nextA_63_port, nextA_62_port, nextA_61_port, nextA_60_port, 
      nextA_59_port, nextA_58_port, nextA_57_port, nextA_56_port, nextA_55_port
      , nextA_54_port, nextA_53_port, nextA_52_port, nextA_51_port, 
      nextA_50_port, nextA_49_port, nextA_48_port, nextA_47_port, nextA_46_port
      , nextA_45_port, nextA_44_port, nextA_43_port, nextA_42_port, 
      nextA_41_port, nextA_40_port, nextA_39_port, nextA_38_port, nextA_37_port
      , nextA_36_port, nextA_35_port, nextA_34_port, nextA_33_port, 
      nextA_32_port, nextA_31_port, nextA_30_port, nextA_29_port, nextA_28_port
      , nextA_27_port, nextA_26_port, nextA_25_port, nextA_24_port, 
      nextA_23_port, nextA_22_port, nextA_21_port, nextA_20_port, nextA_19_port
      , nextA_18_port, nextA_17_port, nextA_16_port, nextA_15_port, 
      nextA_14_port, nextA_13_port, nextA_12_port, nextA_11_port, nextA_10_port
      , nextA_9_port, nextA_8_port, nextA_7_port, nextA_6_port, nextA_5_port, 
      nextA_4_port, nextA_3_port, nextA_2_port, nextA_1_port, nextA_0_port );
   
   X_Logic0_port <= '0';
   nextA_0_port <= '0';
   encoder_1 : encoder_N64_RADIX3_15 port map( X(2) => encoderIn(2), X(1) => 
                           encoderIn(1), X(0) => encoderIn(0), Z(2) => 
                           encoder_to_mux_2_port, Z(1) => encoder_to_mux_1_port
                           , Z(0) => encoder_to_mux_0_port);
   ShiftnCompl_1 : ShiftnCompl_N64_0 port map( plusA(63) => prevA(63), 
                           plusA(62) => prevA(62), plusA(61) => prevA(61), 
                           plusA(60) => prevA(60), plusA(59) => prevA(59), 
                           plusA(58) => prevA(58), plusA(57) => prevA(57), 
                           plusA(56) => prevA(56), plusA(55) => prevA(55), 
                           plusA(54) => prevA(54), plusA(53) => prevA(53), 
                           plusA(52) => prevA(52), plusA(51) => prevA(51), 
                           plusA(50) => prevA(50), plusA(49) => prevA(49), 
                           plusA(48) => prevA(48), plusA(47) => prevA(47), 
                           plusA(46) => prevA(46), plusA(45) => prevA(45), 
                           plusA(44) => prevA(44), plusA(43) => prevA(43), 
                           plusA(42) => prevA(42), plusA(41) => prevA(41), 
                           plusA(40) => prevA(40), plusA(39) => prevA(39), 
                           plusA(38) => prevA(38), plusA(37) => prevA(37), 
                           plusA(36) => prevA(36), plusA(35) => prevA(35), 
                           plusA(34) => prevA(34), plusA(33) => prevA(33), 
                           plusA(32) => prevA(32), plusA(31) => prevA(31), 
                           plusA(30) => prevA(30), plusA(29) => prevA(29), 
                           plusA(28) => prevA(28), plusA(27) => prevA(27), 
                           plusA(26) => prevA(26), plusA(25) => prevA(25), 
                           plusA(24) => prevA(24), plusA(23) => prevA(23), 
                           plusA(22) => prevA(22), plusA(21) => prevA(21), 
                           plusA(20) => prevA(20), plusA(19) => prevA(19), 
                           plusA(18) => prevA(18), plusA(17) => prevA(17), 
                           plusA(16) => prevA(16), plusA(15) => prevA(15), 
                           plusA(14) => prevA(14), plusA(13) => prevA(13), 
                           plusA(12) => prevA(12), plusA(11) => prevA(11), 
                           plusA(10) => prevA(10), plusA(9) => prevA(9), 
                           plusA(8) => prevA(8), plusA(7) => prevA(7), plusA(6)
                           => prevA(6), plusA(5) => prevA(5), plusA(4) => 
                           prevA(4), plusA(3) => prevA(3), plusA(2) => prevA(2)
                           , plusA(1) => prevA(1), plusA(0) => prevA(0), 
                           plus2A_out(63) => plus2A_s_63_port, plus2A_out(62) 
                           => plus2A_s_62_port, plus2A_out(61) => 
                           plus2A_s_61_port, plus2A_out(60) => plus2A_s_60_port
                           , plus2A_out(59) => plus2A_s_59_port, plus2A_out(58)
                           => plus2A_s_58_port, plus2A_out(57) => 
                           plus2A_s_57_port, plus2A_out(56) => plus2A_s_56_port
                           , plus2A_out(55) => plus2A_s_55_port, plus2A_out(54)
                           => plus2A_s_54_port, plus2A_out(53) => 
                           plus2A_s_53_port, plus2A_out(52) => plus2A_s_52_port
                           , plus2A_out(51) => plus2A_s_51_port, plus2A_out(50)
                           => plus2A_s_50_port, plus2A_out(49) => 
                           plus2A_s_49_port, plus2A_out(48) => plus2A_s_48_port
                           , plus2A_out(47) => plus2A_s_47_port, plus2A_out(46)
                           => plus2A_s_46_port, plus2A_out(45) => 
                           plus2A_s_45_port, plus2A_out(44) => plus2A_s_44_port
                           , plus2A_out(43) => plus2A_s_43_port, plus2A_out(42)
                           => plus2A_s_42_port, plus2A_out(41) => 
                           plus2A_s_41_port, plus2A_out(40) => plus2A_s_40_port
                           , plus2A_out(39) => plus2A_s_39_port, plus2A_out(38)
                           => plus2A_s_38_port, plus2A_out(37) => 
                           plus2A_s_37_port, plus2A_out(36) => plus2A_s_36_port
                           , plus2A_out(35) => plus2A_s_35_port, plus2A_out(34)
                           => plus2A_s_34_port, plus2A_out(33) => 
                           plus2A_s_33_port, plus2A_out(32) => plus2A_s_32_port
                           , plus2A_out(31) => plus2A_s_31_port, plus2A_out(30)
                           => plus2A_s_30_port, plus2A_out(29) => 
                           plus2A_s_29_port, plus2A_out(28) => plus2A_s_28_port
                           , plus2A_out(27) => plus2A_s_27_port, plus2A_out(26)
                           => plus2A_s_26_port, plus2A_out(25) => 
                           plus2A_s_25_port, plus2A_out(24) => plus2A_s_24_port
                           , plus2A_out(23) => plus2A_s_23_port, plus2A_out(22)
                           => plus2A_s_22_port, plus2A_out(21) => 
                           plus2A_s_21_port, plus2A_out(20) => plus2A_s_20_port
                           , plus2A_out(19) => plus2A_s_19_port, plus2A_out(18)
                           => plus2A_s_18_port, plus2A_out(17) => 
                           plus2A_s_17_port, plus2A_out(16) => plus2A_s_16_port
                           , plus2A_out(15) => plus2A_s_15_port, plus2A_out(14)
                           => plus2A_s_14_port, plus2A_out(13) => 
                           plus2A_s_13_port, plus2A_out(12) => plus2A_s_12_port
                           , plus2A_out(11) => plus2A_s_11_port, plus2A_out(10)
                           => plus2A_s_10_port, plus2A_out(9) => 
                           plus2A_s_9_port, plus2A_out(8) => plus2A_s_8_port, 
                           plus2A_out(7) => plus2A_s_7_port, plus2A_out(6) => 
                           plus2A_s_6_port, plus2A_out(5) => plus2A_s_5_port, 
                           plus2A_out(4) => plus2A_s_4_port, plus2A_out(3) => 
                           plus2A_s_3_port, plus2A_out(2) => plus2A_s_2_port, 
                           plus2A_out(1) => plus2A_s_1_port, plus2A_out(0) => 
                           n_3217, minus2A_out(63) => minus2A_s_63_port, 
                           minus2A_out(62) => minus2A_s_62_port, 
                           minus2A_out(61) => minus2A_s_61_port, 
                           minus2A_out(60) => minus2A_s_60_port, 
                           minus2A_out(59) => minus2A_s_59_port, 
                           minus2A_out(58) => minus2A_s_58_port, 
                           minus2A_out(57) => minus2A_s_57_port, 
                           minus2A_out(56) => minus2A_s_56_port, 
                           minus2A_out(55) => minus2A_s_55_port, 
                           minus2A_out(54) => minus2A_s_54_port, 
                           minus2A_out(53) => minus2A_s_53_port, 
                           minus2A_out(52) => minus2A_s_52_port, 
                           minus2A_out(51) => minus2A_s_51_port, 
                           minus2A_out(50) => minus2A_s_50_port, 
                           minus2A_out(49) => minus2A_s_49_port, 
                           minus2A_out(48) => minus2A_s_48_port, 
                           minus2A_out(47) => minus2A_s_47_port, 
                           minus2A_out(46) => minus2A_s_46_port, 
                           minus2A_out(45) => minus2A_s_45_port, 
                           minus2A_out(44) => minus2A_s_44_port, 
                           minus2A_out(43) => minus2A_s_43_port, 
                           minus2A_out(42) => minus2A_s_42_port, 
                           minus2A_out(41) => minus2A_s_41_port, 
                           minus2A_out(40) => minus2A_s_40_port, 
                           minus2A_out(39) => minus2A_s_39_port, 
                           minus2A_out(38) => minus2A_s_38_port, 
                           minus2A_out(37) => minus2A_s_37_port, 
                           minus2A_out(36) => minus2A_s_36_port, 
                           minus2A_out(35) => minus2A_s_35_port, 
                           minus2A_out(34) => minus2A_s_34_port, 
                           minus2A_out(33) => minus2A_s_33_port, 
                           minus2A_out(32) => minus2A_s_32_port, 
                           minus2A_out(31) => minus2A_s_31_port, 
                           minus2A_out(30) => minus2A_s_30_port, 
                           minus2A_out(29) => minus2A_s_29_port, 
                           minus2A_out(28) => minus2A_s_28_port, 
                           minus2A_out(27) => minus2A_s_27_port, 
                           minus2A_out(26) => minus2A_s_26_port, 
                           minus2A_out(25) => minus2A_s_25_port, 
                           minus2A_out(24) => minus2A_s_24_port, 
                           minus2A_out(23) => minus2A_s_23_port, 
                           minus2A_out(22) => minus2A_s_22_port, 
                           minus2A_out(21) => minus2A_s_21_port, 
                           minus2A_out(20) => minus2A_s_20_port, 
                           minus2A_out(19) => minus2A_s_19_port, 
                           minus2A_out(18) => minus2A_s_18_port, 
                           minus2A_out(17) => minus2A_s_17_port, 
                           minus2A_out(16) => minus2A_s_16_port, 
                           minus2A_out(15) => minus2A_s_15_port, 
                           minus2A_out(14) => minus2A_s_14_port, 
                           minus2A_out(13) => minus2A_s_13_port, 
                           minus2A_out(12) => minus2A_s_12_port, 
                           minus2A_out(11) => minus2A_s_11_port, 
                           minus2A_out(10) => minus2A_s_10_port, minus2A_out(9)
                           => minus2A_s_9_port, minus2A_out(8) => 
                           minus2A_s_8_port, minus2A_out(7) => minus2A_s_7_port
                           , minus2A_out(6) => minus2A_s_6_port, minus2A_out(5)
                           => minus2A_s_5_port, minus2A_out(4) => 
                           minus2A_s_4_port, minus2A_out(3) => minus2A_s_3_port
                           , minus2A_out(2) => minus2A_s_2_port, minus2A_out(1)
                           => minus2A_s_1_port, minus2A_out(0) => 
                           minus2A_s_0_port, plus4A_out(63) => nextA_63_port, 
                           plus4A_out(62) => nextA_62_port, plus4A_out(61) => 
                           nextA_61_port, plus4A_out(60) => nextA_60_port, 
                           plus4A_out(59) => nextA_59_port, plus4A_out(58) => 
                           nextA_58_port, plus4A_out(57) => n3, plus4A_out(56) 
                           => nextA_56_port, plus4A_out(55) => nextA_55_port, 
                           plus4A_out(54) => nextA_54_port, plus4A_out(53) => 
                           nextA_53_port, plus4A_out(52) => nextA_52_port, 
                           plus4A_out(51) => nextA_51_port, plus4A_out(50) => 
                           nextA_50_port, plus4A_out(49) => nextA_49_port, 
                           plus4A_out(48) => nextA_48_port, plus4A_out(47) => 
                           nextA_47_port, plus4A_out(46) => nextA_46_port, 
                           plus4A_out(45) => nextA_45_port, plus4A_out(44) => 
                           nextA_44_port, plus4A_out(43) => nextA_43_port, 
                           plus4A_out(42) => nextA_42_port, plus4A_out(41) => 
                           nextA_41_port, plus4A_out(40) => nextA_40_port, 
                           plus4A_out(39) => nextA_39_port, plus4A_out(38) => 
                           nextA_38_port, plus4A_out(37) => nextA_37_port, 
                           plus4A_out(36) => nextA_36_port, plus4A_out(35) => 
                           nextA_35_port, plus4A_out(34) => nextA_34_port, 
                           plus4A_out(33) => nextA_33_port, plus4A_out(32) => 
                           nextA_32_port, plus4A_out(31) => nextA_31_port, 
                           plus4A_out(30) => nextA_30_port, plus4A_out(29) => 
                           nextA_29_port, plus4A_out(28) => nextA_28_port, 
                           plus4A_out(27) => nextA_27_port, plus4A_out(26) => 
                           nextA_26_port, plus4A_out(25) => nextA_25_port, 
                           plus4A_out(24) => nextA_24_port, plus4A_out(23) => 
                           nextA_23_port, plus4A_out(22) => nextA_22_port, 
                           plus4A_out(21) => nextA_21_port, plus4A_out(20) => 
                           nextA_20_port, plus4A_out(19) => nextA_19_port, 
                           plus4A_out(18) => nextA_18_port, plus4A_out(17) => 
                           nextA_17_port, plus4A_out(16) => nextA_16_port, 
                           plus4A_out(15) => nextA_15_port, plus4A_out(14) => 
                           nextA_14_port, plus4A_out(13) => nextA_13_port, 
                           plus4A_out(12) => nextA_12_port, plus4A_out(11) => 
                           nextA_11_port, plus4A_out(10) => nextA_10_port, 
                           plus4A_out(9) => nextA_9_port, plus4A_out(8) => 
                           nextA_8_port, plus4A_out(7) => nextA_7_port, 
                           plus4A_out(6) => nextA_6_port, plus4A_out(5) => 
                           nextA_5_port, plus4A_out(4) => nextA_4_port, 
                           plus4A_out(3) => nextA_3_port, plus4A_out(2) => 
                           nextA_2_port, plus4A_out(1) => nextA_1_port, 
                           plus4A_out(0) => n_3218, minus4A_out(63) => 
                           minus4A_s_63_port, minus4A_out(62) => 
                           minus4A_s_62_port, minus4A_out(61) => 
                           minus4A_s_61_port, minus4A_out(60) => 
                           minus4A_s_60_port, minus4A_out(59) => 
                           minus4A_s_59_port, minus4A_out(58) => 
                           minus4A_s_58_port, minus4A_out(57) => 
                           minus4A_s_57_port, minus4A_out(56) => 
                           minus4A_s_56_port, minus4A_out(55) => 
                           minus4A_s_55_port, minus4A_out(54) => 
                           minus4A_s_54_port, minus4A_out(53) => 
                           minus4A_s_53_port, minus4A_out(52) => 
                           minus4A_s_52_port, minus4A_out(51) => 
                           minus4A_s_51_port, minus4A_out(50) => 
                           minus4A_s_50_port, minus4A_out(49) => 
                           minus4A_s_49_port, minus4A_out(48) => 
                           minus4A_s_48_port, minus4A_out(47) => 
                           minus4A_s_47_port, minus4A_out(46) => 
                           minus4A_s_46_port, minus4A_out(45) => 
                           minus4A_s_45_port, minus4A_out(44) => 
                           minus4A_s_44_port, minus4A_out(43) => 
                           minus4A_s_43_port, minus4A_out(42) => 
                           minus4A_s_42_port, minus4A_out(41) => 
                           minus4A_s_41_port, minus4A_out(40) => 
                           minus4A_s_40_port, minus4A_out(39) => 
                           minus4A_s_39_port, minus4A_out(38) => 
                           minus4A_s_38_port, minus4A_out(37) => 
                           minus4A_s_37_port, minus4A_out(36) => 
                           minus4A_s_36_port, minus4A_out(35) => 
                           minus4A_s_35_port, minus4A_out(34) => 
                           minus4A_s_34_port, minus4A_out(33) => 
                           minus4A_s_33_port, minus4A_out(32) => 
                           minus4A_s_32_port, minus4A_out(31) => 
                           minus4A_s_31_port, minus4A_out(30) => 
                           minus4A_s_30_port, minus4A_out(29) => 
                           minus4A_s_29_port, minus4A_out(28) => 
                           minus4A_s_28_port, minus4A_out(27) => 
                           minus4A_s_27_port, minus4A_out(26) => 
                           minus4A_s_26_port, minus4A_out(25) => 
                           minus4A_s_25_port, minus4A_out(24) => 
                           minus4A_s_24_port, minus4A_out(23) => 
                           minus4A_s_23_port, minus4A_out(22) => 
                           minus4A_s_22_port, minus4A_out(21) => 
                           minus4A_s_21_port, minus4A_out(20) => 
                           minus4A_s_20_port, minus4A_out(19) => 
                           minus4A_s_19_port, minus4A_out(18) => 
                           minus4A_s_18_port, minus4A_out(17) => 
                           minus4A_s_17_port, minus4A_out(16) => 
                           minus4A_s_16_port, minus4A_out(15) => 
                           minus4A_s_15_port, minus4A_out(14) => 
                           minus4A_s_14_port, minus4A_out(13) => 
                           minus4A_s_13_port, minus4A_out(12) => 
                           minus4A_s_12_port, minus4A_out(11) => 
                           minus4A_s_11_port, minus4A_out(10) => 
                           minus4A_s_10_port, minus4A_out(9) => 
                           minus4A_s_9_port, minus4A_out(8) => minus4A_s_8_port
                           , minus4A_out(7) => minus4A_s_7_port, minus4A_out(6)
                           => minus4A_s_6_port, minus4A_out(5) => 
                           minus4A_s_5_port, minus4A_out(4) => minus4A_s_4_port
                           , minus4A_out(3) => minus4A_s_3_port, minus4A_out(2)
                           => minus4A_s_2_port, minus4A_out(1) => 
                           minus4A_s_1_port, minus4A_out(0) => minus4A_s_0_port
                           );
   mux_1 : MUX_GENERIC_N64_RADIX3_15 port map( plusA(63) => plus2A_s_63_port, 
                           plusA(62) => plus2A_s_62_port, plusA(61) => 
                           plus2A_s_61_port, plusA(60) => plus2A_s_60_port, 
                           plusA(59) => plus2A_s_59_port, plusA(58) => 
                           plus2A_s_58_port, plusA(57) => plus2A_s_57_port, 
                           plusA(56) => plus2A_s_56_port, plusA(55) => 
                           plus2A_s_55_port, plusA(54) => plus2A_s_54_port, 
                           plusA(53) => plus2A_s_53_port, plusA(52) => 
                           plus2A_s_52_port, plusA(51) => plus2A_s_51_port, 
                           plusA(50) => plus2A_s_50_port, plusA(49) => 
                           plus2A_s_49_port, plusA(48) => plus2A_s_48_port, 
                           plusA(47) => plus2A_s_47_port, plusA(46) => 
                           plus2A_s_46_port, plusA(45) => plus2A_s_45_port, 
                           plusA(44) => plus2A_s_44_port, plusA(43) => 
                           plus2A_s_43_port, plusA(42) => plus2A_s_42_port, 
                           plusA(41) => plus2A_s_41_port, plusA(40) => 
                           plus2A_s_40_port, plusA(39) => plus2A_s_39_port, 
                           plusA(38) => plus2A_s_38_port, plusA(37) => 
                           plus2A_s_37_port, plusA(36) => plus2A_s_36_port, 
                           plusA(35) => plus2A_s_35_port, plusA(34) => 
                           plus2A_s_34_port, plusA(33) => plus2A_s_33_port, 
                           plusA(32) => plus2A_s_32_port, plusA(31) => 
                           plus2A_s_31_port, plusA(30) => plus2A_s_30_port, 
                           plusA(29) => plus2A_s_29_port, plusA(28) => 
                           plus2A_s_28_port, plusA(27) => plus2A_s_27_port, 
                           plusA(26) => plus2A_s_26_port, plusA(25) => 
                           plus2A_s_25_port, plusA(24) => plus2A_s_24_port, 
                           plusA(23) => plus2A_s_23_port, plusA(22) => 
                           plus2A_s_22_port, plusA(21) => plus2A_s_21_port, 
                           plusA(20) => plus2A_s_20_port, plusA(19) => 
                           plus2A_s_19_port, plusA(18) => plus2A_s_18_port, 
                           plusA(17) => plus2A_s_17_port, plusA(16) => 
                           plus2A_s_16_port, plusA(15) => plus2A_s_15_port, 
                           plusA(14) => plus2A_s_14_port, plusA(13) => 
                           plus2A_s_13_port, plusA(12) => plus2A_s_12_port, 
                           plusA(11) => plus2A_s_11_port, plusA(10) => 
                           plus2A_s_10_port, plusA(9) => plus2A_s_9_port, 
                           plusA(8) => plus2A_s_8_port, plusA(7) => 
                           plus2A_s_7_port, plusA(6) => plus2A_s_6_port, 
                           plusA(5) => plus2A_s_5_port, plusA(4) => 
                           plus2A_s_4_port, plusA(3) => plus2A_s_3_port, 
                           plusA(2) => plus2A_s_2_port, plusA(1) => 
                           plus2A_s_1_port, plusA(0) => nextA_0_port, 
                           minusA(63) => minus2A_s_63_port, minusA(62) => 
                           minus2A_s_62_port, minusA(61) => minus2A_s_61_port, 
                           minusA(60) => minus2A_s_60_port, minusA(59) => 
                           minus2A_s_59_port, minusA(58) => minus2A_s_58_port, 
                           minusA(57) => minus2A_s_57_port, minusA(56) => 
                           minus2A_s_56_port, minusA(55) => minus2A_s_55_port, 
                           minusA(54) => minus2A_s_54_port, minusA(53) => 
                           minus2A_s_53_port, minusA(52) => minus2A_s_52_port, 
                           minusA(51) => minus2A_s_51_port, minusA(50) => 
                           minus2A_s_50_port, minusA(49) => minus2A_s_49_port, 
                           minusA(48) => minus2A_s_48_port, minusA(47) => 
                           minus2A_s_47_port, minusA(46) => minus2A_s_46_port, 
                           minusA(45) => minus2A_s_45_port, minusA(44) => 
                           minus2A_s_44_port, minusA(43) => minus2A_s_43_port, 
                           minusA(42) => minus2A_s_42_port, minusA(41) => 
                           minus2A_s_41_port, minusA(40) => minus2A_s_40_port, 
                           minusA(39) => minus2A_s_39_port, minusA(38) => 
                           minus2A_s_38_port, minusA(37) => minus2A_s_37_port, 
                           minusA(36) => minus2A_s_36_port, minusA(35) => 
                           minus2A_s_35_port, minusA(34) => minus2A_s_34_port, 
                           minusA(33) => minus2A_s_33_port, minusA(32) => 
                           minus2A_s_32_port, minusA(31) => minus2A_s_31_port, 
                           minusA(30) => minus2A_s_30_port, minusA(29) => 
                           minus2A_s_29_port, minusA(28) => minus2A_s_28_port, 
                           minusA(27) => minus2A_s_27_port, minusA(26) => 
                           minus2A_s_26_port, minusA(25) => minus2A_s_25_port, 
                           minusA(24) => minus2A_s_24_port, minusA(23) => 
                           minus2A_s_23_port, minusA(22) => minus2A_s_22_port, 
                           minusA(21) => minus2A_s_21_port, minusA(20) => 
                           minus2A_s_20_port, minusA(19) => minus2A_s_19_port, 
                           minusA(18) => minus2A_s_18_port, minusA(17) => 
                           minus2A_s_17_port, minusA(16) => minus2A_s_16_port, 
                           minusA(15) => minus2A_s_15_port, minusA(14) => 
                           minus2A_s_14_port, minusA(13) => minus2A_s_13_port, 
                           minusA(12) => minus2A_s_12_port, minusA(11) => 
                           minus2A_s_11_port, minusA(10) => minus2A_s_10_port, 
                           minusA(9) => minus2A_s_9_port, minusA(8) => 
                           minus2A_s_8_port, minusA(7) => minus2A_s_7_port, 
                           minusA(6) => minus2A_s_6_port, minusA(5) => 
                           minus2A_s_5_port, minusA(4) => minus2A_s_4_port, 
                           minusA(3) => minus2A_s_3_port, minusA(2) => 
                           minus2A_s_2_port, minusA(1) => minus2A_s_1_port, 
                           minusA(0) => minus2A_s_0_port, plus2A(63) => 
                           nextA_63_port, plus2A(62) => nextA_62_port, 
                           plus2A(61) => nextA_61_port, plus2A(60) => 
                           nextA_60_port, plus2A(59) => nextA_59_port, 
                           plus2A(58) => nextA_58_port, plus2A(57) => 
                           nextA_57_port, plus2A(56) => nextA_56_port, 
                           plus2A(55) => nextA_55_port, plus2A(54) => 
                           nextA_54_port, plus2A(53) => nextA_53_port, 
                           plus2A(52) => nextA_52_port, plus2A(51) => 
                           nextA_51_port, plus2A(50) => nextA_50_port, 
                           plus2A(49) => nextA_49_port, plus2A(48) => 
                           nextA_48_port, plus2A(47) => nextA_47_port, 
                           plus2A(46) => nextA_46_port, plus2A(45) => 
                           nextA_45_port, plus2A(44) => nextA_44_port, 
                           plus2A(43) => nextA_43_port, plus2A(42) => 
                           nextA_42_port, plus2A(41) => nextA_41_port, 
                           plus2A(40) => nextA_40_port, plus2A(39) => 
                           nextA_39_port, plus2A(38) => nextA_38_port, 
                           plus2A(37) => nextA_37_port, plus2A(36) => 
                           nextA_36_port, plus2A(35) => nextA_35_port, 
                           plus2A(34) => nextA_34_port, plus2A(33) => 
                           nextA_33_port, plus2A(32) => nextA_32_port, 
                           plus2A(31) => nextA_31_port, plus2A(30) => 
                           nextA_30_port, plus2A(29) => nextA_29_port, 
                           plus2A(28) => nextA_28_port, plus2A(27) => 
                           nextA_27_port, plus2A(26) => nextA_26_port, 
                           plus2A(25) => nextA_25_port, plus2A(24) => 
                           nextA_24_port, plus2A(23) => nextA_23_port, 
                           plus2A(22) => nextA_22_port, plus2A(21) => 
                           nextA_21_port, plus2A(20) => nextA_20_port, 
                           plus2A(19) => nextA_19_port, plus2A(18) => 
                           nextA_18_port, plus2A(17) => nextA_17_port, 
                           plus2A(16) => nextA_16_port, plus2A(15) => 
                           nextA_15_port, plus2A(14) => nextA_14_port, 
                           plus2A(13) => nextA_13_port, plus2A(12) => 
                           nextA_12_port, plus2A(11) => nextA_11_port, 
                           plus2A(10) => nextA_10_port, plus2A(9) => 
                           nextA_9_port, plus2A(8) => nextA_8_port, plus2A(7) 
                           => nextA_7_port, plus2A(6) => nextA_6_port, 
                           plus2A(5) => nextA_5_port, plus2A(4) => nextA_4_port
                           , plus2A(3) => nextA_3_port, plus2A(2) => 
                           nextA_2_port, plus2A(1) => nextA_1_port, plus2A(0) 
                           => nextA_0_port, minus2A(63) => minus4A_s_63_port, 
                           minus2A(62) => minus4A_s_62_port, minus2A(61) => 
                           minus4A_s_61_port, minus2A(60) => minus4A_s_60_port,
                           minus2A(59) => minus4A_s_59_port, minus2A(58) => 
                           minus4A_s_58_port, minus2A(57) => minus4A_s_57_port,
                           minus2A(56) => minus4A_s_56_port, minus2A(55) => 
                           minus4A_s_55_port, minus2A(54) => minus4A_s_54_port,
                           minus2A(53) => minus4A_s_53_port, minus2A(52) => 
                           minus4A_s_52_port, minus2A(51) => minus4A_s_51_port,
                           minus2A(50) => minus4A_s_50_port, minus2A(49) => 
                           minus4A_s_49_port, minus2A(48) => minus4A_s_48_port,
                           minus2A(47) => minus4A_s_47_port, minus2A(46) => 
                           minus4A_s_46_port, minus2A(45) => minus4A_s_45_port,
                           minus2A(44) => minus4A_s_44_port, minus2A(43) => 
                           minus4A_s_43_port, minus2A(42) => minus4A_s_42_port,
                           minus2A(41) => minus4A_s_41_port, minus2A(40) => 
                           minus4A_s_40_port, minus2A(39) => minus4A_s_39_port,
                           minus2A(38) => minus4A_s_38_port, minus2A(37) => 
                           minus4A_s_37_port, minus2A(36) => minus4A_s_36_port,
                           minus2A(35) => minus4A_s_35_port, minus2A(34) => 
                           minus4A_s_34_port, minus2A(33) => minus4A_s_33_port,
                           minus2A(32) => minus4A_s_32_port, minus2A(31) => 
                           minus4A_s_31_port, minus2A(30) => minus4A_s_30_port,
                           minus2A(29) => minus4A_s_29_port, minus2A(28) => 
                           minus4A_s_28_port, minus2A(27) => minus4A_s_27_port,
                           minus2A(26) => minus4A_s_26_port, minus2A(25) => 
                           minus4A_s_25_port, minus2A(24) => minus4A_s_24_port,
                           minus2A(23) => minus4A_s_23_port, minus2A(22) => 
                           minus4A_s_22_port, minus2A(21) => minus4A_s_21_port,
                           minus2A(20) => minus4A_s_20_port, minus2A(19) => 
                           minus4A_s_19_port, minus2A(18) => minus4A_s_18_port,
                           minus2A(17) => minus4A_s_17_port, minus2A(16) => 
                           minus4A_s_16_port, minus2A(15) => minus4A_s_15_port,
                           minus2A(14) => minus4A_s_14_port, minus2A(13) => 
                           minus4A_s_13_port, minus2A(12) => minus4A_s_12_port,
                           minus2A(11) => minus4A_s_11_port, minus2A(10) => 
                           minus4A_s_10_port, minus2A(9) => minus4A_s_9_port, 
                           minus2A(8) => minus4A_s_8_port, minus2A(7) => 
                           minus4A_s_7_port, minus2A(6) => minus4A_s_6_port, 
                           minus2A(5) => minus4A_s_5_port, minus2A(4) => 
                           minus4A_s_4_port, minus2A(3) => minus4A_s_3_port, 
                           minus2A(2) => minus4A_s_2_port, minus2A(1) => 
                           minus4A_s_1_port, minus2A(0) => minus4A_s_0_port, 
                           SEL(2) => encoder_to_mux_2_port, SEL(1) => 
                           encoder_to_mux_1_port, SEL(0) => 
                           encoder_to_mux_0_port, Y(63) => mux_to_adder_63_port
                           , Y(62) => mux_to_adder_62_port, Y(61) => 
                           mux_to_adder_61_port, Y(60) => mux_to_adder_60_port,
                           Y(59) => mux_to_adder_59_port, Y(58) => 
                           mux_to_adder_58_port, Y(57) => mux_to_adder_57_port,
                           Y(56) => mux_to_adder_56_port, Y(55) => 
                           mux_to_adder_55_port, Y(54) => mux_to_adder_54_port,
                           Y(53) => mux_to_adder_53_port, Y(52) => 
                           mux_to_adder_52_port, Y(51) => mux_to_adder_51_port,
                           Y(50) => mux_to_adder_50_port, Y(49) => 
                           mux_to_adder_49_port, Y(48) => mux_to_adder_48_port,
                           Y(47) => mux_to_adder_47_port, Y(46) => 
                           mux_to_adder_46_port, Y(45) => mux_to_adder_45_port,
                           Y(44) => mux_to_adder_44_port, Y(43) => 
                           mux_to_adder_43_port, Y(42) => mux_to_adder_42_port,
                           Y(41) => mux_to_adder_41_port, Y(40) => 
                           mux_to_adder_40_port, Y(39) => mux_to_adder_39_port,
                           Y(38) => mux_to_adder_38_port, Y(37) => 
                           mux_to_adder_37_port, Y(36) => mux_to_adder_36_port,
                           Y(35) => mux_to_adder_35_port, Y(34) => 
                           mux_to_adder_34_port, Y(33) => mux_to_adder_33_port,
                           Y(32) => mux_to_adder_32_port, Y(31) => 
                           mux_to_adder_31_port, Y(30) => mux_to_adder_30_port,
                           Y(29) => mux_to_adder_29_port, Y(28) => 
                           mux_to_adder_28_port, Y(27) => mux_to_adder_27_port,
                           Y(26) => mux_to_adder_26_port, Y(25) => 
                           mux_to_adder_25_port, Y(24) => mux_to_adder_24_port,
                           Y(23) => mux_to_adder_23_port, Y(22) => 
                           mux_to_adder_22_port, Y(21) => mux_to_adder_21_port,
                           Y(20) => mux_to_adder_20_port, Y(19) => 
                           mux_to_adder_19_port, Y(18) => mux_to_adder_18_port,
                           Y(17) => mux_to_adder_17_port, Y(16) => 
                           mux_to_adder_16_port, Y(15) => mux_to_adder_15_port,
                           Y(14) => mux_to_adder_14_port, Y(13) => 
                           mux_to_adder_13_port, Y(12) => mux_to_adder_12_port,
                           Y(11) => mux_to_adder_11_port, Y(10) => 
                           mux_to_adder_10_port, Y(9) => mux_to_adder_9_port, 
                           Y(8) => mux_to_adder_8_port, Y(7) => 
                           mux_to_adder_7_port, Y(6) => mux_to_adder_6_port, 
                           Y(5) => mux_to_adder_5_port, Y(4) => 
                           mux_to_adder_4_port, Y(3) => mux_to_adder_3_port, 
                           Y(2) => mux_to_adder_2_port, Y(1) => 
                           mux_to_adder_1_port, Y(0) => mux_to_adder_0_port);
   rca_1 : RCA_N64_0 port map( A(63) => mux_to_adder_63_port, A(62) => 
                           mux_to_adder_62_port, A(61) => mux_to_adder_61_port,
                           A(60) => mux_to_adder_60_port, A(59) => 
                           mux_to_adder_59_port, A(58) => mux_to_adder_58_port,
                           A(57) => mux_to_adder_57_port, A(56) => 
                           mux_to_adder_56_port, A(55) => mux_to_adder_55_port,
                           A(54) => mux_to_adder_54_port, A(53) => 
                           mux_to_adder_53_port, A(52) => mux_to_adder_52_port,
                           A(51) => mux_to_adder_51_port, A(50) => 
                           mux_to_adder_50_port, A(49) => mux_to_adder_49_port,
                           A(48) => mux_to_adder_48_port, A(47) => 
                           mux_to_adder_47_port, A(46) => mux_to_adder_46_port,
                           A(45) => mux_to_adder_45_port, A(44) => 
                           mux_to_adder_44_port, A(43) => mux_to_adder_43_port,
                           A(42) => mux_to_adder_42_port, A(41) => 
                           mux_to_adder_41_port, A(40) => mux_to_adder_40_port,
                           A(39) => mux_to_adder_39_port, A(38) => 
                           mux_to_adder_38_port, A(37) => mux_to_adder_37_port,
                           A(36) => mux_to_adder_36_port, A(35) => 
                           mux_to_adder_35_port, A(34) => mux_to_adder_34_port,
                           A(33) => mux_to_adder_33_port, A(32) => 
                           mux_to_adder_32_port, A(31) => mux_to_adder_31_port,
                           A(30) => mux_to_adder_30_port, A(29) => 
                           mux_to_adder_29_port, A(28) => mux_to_adder_28_port,
                           A(27) => mux_to_adder_27_port, A(26) => 
                           mux_to_adder_26_port, A(25) => mux_to_adder_25_port,
                           A(24) => mux_to_adder_24_port, A(23) => 
                           mux_to_adder_23_port, A(22) => mux_to_adder_22_port,
                           A(21) => mux_to_adder_21_port, A(20) => 
                           mux_to_adder_20_port, A(19) => mux_to_adder_19_port,
                           A(18) => mux_to_adder_18_port, A(17) => 
                           mux_to_adder_17_port, A(16) => mux_to_adder_16_port,
                           A(15) => mux_to_adder_15_port, A(14) => 
                           mux_to_adder_14_port, A(13) => mux_to_adder_13_port,
                           A(12) => mux_to_adder_12_port, A(11) => 
                           mux_to_adder_11_port, A(10) => mux_to_adder_10_port,
                           A(9) => mux_to_adder_9_port, A(8) => 
                           mux_to_adder_8_port, A(7) => mux_to_adder_7_port, 
                           A(6) => mux_to_adder_6_port, A(5) => 
                           mux_to_adder_5_port, A(4) => mux_to_adder_4_port, 
                           A(3) => mux_to_adder_3_port, A(2) => 
                           mux_to_adder_2_port, A(1) => mux_to_adder_1_port, 
                           A(0) => mux_to_adder_0_port, B(63) => prevSum(63), 
                           B(62) => prevSum(62), B(61) => prevSum(61), B(60) =>
                           prevSum(60), B(59) => prevSum(59), B(58) => 
                           prevSum(58), B(57) => prevSum(57), B(56) => 
                           prevSum(56), B(55) => prevSum(55), B(54) => 
                           prevSum(54), B(53) => prevSum(53), B(52) => 
                           prevSum(52), B(51) => prevSum(51), B(50) => 
                           prevSum(50), B(49) => prevSum(49), B(48) => 
                           prevSum(48), B(47) => prevSum(47), B(46) => 
                           prevSum(46), B(45) => prevSum(45), B(44) => 
                           prevSum(44), B(43) => prevSum(43), B(42) => 
                           prevSum(42), B(41) => prevSum(41), B(40) => 
                           prevSum(40), B(39) => prevSum(39), B(38) => 
                           prevSum(38), B(37) => prevSum(37), B(36) => 
                           prevSum(36), B(35) => prevSum(35), B(34) => 
                           prevSum(34), B(33) => prevSum(33), B(32) => 
                           prevSum(32), B(31) => prevSum(31), B(30) => 
                           prevSum(30), B(29) => prevSum(29), B(28) => 
                           prevSum(28), B(27) => prevSum(27), B(26) => 
                           prevSum(26), B(25) => prevSum(25), B(24) => 
                           prevSum(24), B(23) => prevSum(23), B(22) => 
                           prevSum(22), B(21) => prevSum(21), B(20) => 
                           prevSum(20), B(19) => prevSum(19), B(18) => 
                           prevSum(18), B(17) => prevSum(17), B(16) => 
                           prevSum(16), B(15) => prevSum(15), B(14) => 
                           prevSum(14), B(13) => prevSum(13), B(12) => 
                           prevSum(12), B(11) => prevSum(11), B(10) => 
                           prevSum(10), B(9) => prevSum(9), B(8) => prevSum(8),
                           B(7) => prevSum(7), B(6) => prevSum(6), B(5) => 
                           prevSum(5), B(4) => prevSum(4), B(3) => prevSum(3), 
                           B(2) => prevSum(2), B(1) => prevSum(1), B(0) => 
                           prevSum(0), Ci => X_Logic0_port, S(63) => 
                           nextSum(63), S(62) => nextSum(62), S(61) => 
                           nextSum(61), S(60) => nextSum(60), S(59) => 
                           nextSum(59), S(58) => nextSum(58), S(57) => 
                           nextSum(57), S(56) => nextSum(56), S(55) => 
                           nextSum(55), S(54) => nextSum(54), S(53) => 
                           nextSum(53), S(52) => nextSum(52), S(51) => 
                           nextSum(51), S(50) => nextSum(50), S(49) => 
                           nextSum(49), S(48) => nextSum(48), S(47) => 
                           nextSum(47), S(46) => nextSum(46), S(45) => 
                           nextSum(45), S(44) => nextSum(44), S(43) => 
                           nextSum(43), S(42) => nextSum(42), S(41) => 
                           nextSum(41), S(40) => nextSum(40), S(39) => 
                           nextSum(39), S(38) => nextSum(38), S(37) => 
                           nextSum(37), S(36) => nextSum(36), S(35) => 
                           nextSum(35), S(34) => nextSum(34), S(33) => 
                           nextSum(33), S(32) => nextSum(32), S(31) => 
                           nextSum(31), S(30) => nextSum(30), S(29) => 
                           nextSum(29), S(28) => nextSum(28), S(27) => 
                           nextSum(27), S(26) => nextSum(26), S(25) => 
                           nextSum(25), S(24) => nextSum(24), S(23) => 
                           nextSum(23), S(22) => nextSum(22), S(21) => 
                           nextSum(21), S(20) => nextSum(20), S(19) => 
                           nextSum(19), S(18) => nextSum(18), S(17) => 
                           nextSum(17), S(16) => nextSum(16), S(15) => 
                           nextSum(15), S(14) => nextSum(14), S(13) => 
                           nextSum(13), S(12) => nextSum(12), S(11) => 
                           nextSum(11), S(10) => nextSum(10), S(9) => 
                           nextSum(9), S(8) => nextSum(8), S(7) => nextSum(7), 
                           S(6) => nextSum(6), S(5) => nextSum(5), S(4) => 
                           nextSum(4), S(3) => nextSum(3), S(2) => nextSum(2), 
                           S(1) => nextSum(1), S(0) => nextSum(0), Co => n_3219
                           );
   U3 : BUF_X1 port map( A => n3, Z => nextA_57_port);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity booth_mul_row_special_N64_RADIX3 is

   port( A : in std_logic_vector (63 downto 0);  encoderIn : in 
         std_logic_vector (2 downto 0);  nextA, nextSum : out std_logic_vector 
         (63 downto 0));

end booth_mul_row_special_N64_RADIX3;

architecture SYN_struct of booth_mul_row_special_N64_RADIX3 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX_GENERIC_N64_RADIX3_0
      port( plusA, minusA, plus2A, minus2A : in std_logic_vector (63 downto 0);
            SEL : in std_logic_vector (2 downto 0);  Y : out std_logic_vector 
            (63 downto 0));
   end component;
   
   component ShiftnCompl_special_N64
      port( plusA : in std_logic_vector (63 downto 0);  plusA_out, minusA_out, 
            plus2A_out, minus2A_out : out std_logic_vector (63 downto 0));
   end component;
   
   component encoder_N64_RADIX3_0
      port( X : in std_logic_vector (2 downto 0);  Z : out std_logic_vector (2 
            downto 0));
   end component;
   
   signal nextA_63_port, nextA_62_port, nextA_61_port, nextA_60_port, 
      nextA_59_port, nextA_58_port, n3, nextA_56_port, nextA_55_port, 
      nextA_54_port, nextA_53_port, nextA_52_port, nextA_51_port, nextA_50_port
      , nextA_49_port, nextA_48_port, nextA_47_port, nextA_46_port, 
      nextA_45_port, nextA_44_port, nextA_43_port, nextA_42_port, nextA_41_port
      , nextA_40_port, nextA_39_port, nextA_38_port, nextA_37_port, 
      nextA_36_port, nextA_35_port, nextA_34_port, nextA_33_port, nextA_32_port
      , nextA_31_port, nextA_30_port, nextA_29_port, nextA_28_port, 
      nextA_27_port, nextA_26_port, nextA_25_port, nextA_24_port, nextA_23_port
      , nextA_22_port, nextA_21_port, nextA_20_port, nextA_19_port, 
      nextA_18_port, nextA_17_port, nextA_16_port, nextA_15_port, nextA_14_port
      , nextA_13_port, nextA_12_port, nextA_11_port, nextA_10_port, 
      nextA_9_port, nextA_8_port, nextA_7_port, nextA_6_port, nextA_5_port, 
      nextA_4_port, nextA_3_port, nextA_2_port, nextA_1_port, 
      encoder_to_mux_2_port, encoder_to_mux_1_port, encoder_to_mux_0_port, 
      plusA_s_63_port, plusA_s_62_port, plusA_s_61_port, plusA_s_60_port, 
      plusA_s_59_port, plusA_s_58_port, plusA_s_57_port, plusA_s_56_port, 
      plusA_s_55_port, plusA_s_54_port, plusA_s_53_port, plusA_s_52_port, 
      plusA_s_51_port, plusA_s_50_port, plusA_s_49_port, plusA_s_48_port, 
      plusA_s_47_port, plusA_s_46_port, plusA_s_45_port, plusA_s_44_port, 
      plusA_s_43_port, plusA_s_42_port, plusA_s_41_port, plusA_s_40_port, 
      plusA_s_39_port, plusA_s_38_port, plusA_s_37_port, plusA_s_36_port, 
      plusA_s_35_port, plusA_s_34_port, plusA_s_33_port, plusA_s_32_port, 
      plusA_s_31_port, plusA_s_30_port, plusA_s_29_port, plusA_s_28_port, 
      plusA_s_27_port, plusA_s_26_port, plusA_s_25_port, plusA_s_24_port, 
      plusA_s_23_port, plusA_s_22_port, plusA_s_21_port, plusA_s_20_port, 
      plusA_s_19_port, plusA_s_18_port, plusA_s_17_port, plusA_s_16_port, 
      plusA_s_15_port, plusA_s_14_port, plusA_s_13_port, plusA_s_12_port, 
      plusA_s_11_port, plusA_s_10_port, plusA_s_9_port, plusA_s_8_port, 
      plusA_s_7_port, plusA_s_6_port, plusA_s_5_port, plusA_s_4_port, 
      plusA_s_3_port, plusA_s_2_port, plusA_s_1_port, plusA_s_0_port, 
      minusA_s_63_port, minusA_s_62_port, minusA_s_61_port, minusA_s_60_port, 
      minusA_s_59_port, minusA_s_58_port, minusA_s_57_port, minusA_s_56_port, 
      minusA_s_55_port, minusA_s_54_port, minusA_s_53_port, minusA_s_52_port, 
      minusA_s_51_port, minusA_s_50_port, minusA_s_49_port, minusA_s_48_port, 
      minusA_s_47_port, minusA_s_46_port, minusA_s_45_port, minusA_s_44_port, 
      minusA_s_43_port, minusA_s_42_port, minusA_s_41_port, minusA_s_40_port, 
      minusA_s_39_port, minusA_s_38_port, minusA_s_37_port, minusA_s_36_port, 
      minusA_s_35_port, minusA_s_34_port, minusA_s_33_port, minusA_s_32_port, 
      minusA_s_31_port, minusA_s_30_port, minusA_s_29_port, minusA_s_28_port, 
      minusA_s_27_port, minusA_s_26_port, minusA_s_25_port, minusA_s_24_port, 
      minusA_s_23_port, minusA_s_22_port, minusA_s_21_port, minusA_s_20_port, 
      minusA_s_19_port, minusA_s_18_port, minusA_s_17_port, minusA_s_16_port, 
      minusA_s_15_port, minusA_s_14_port, minusA_s_13_port, minusA_s_12_port, 
      minusA_s_11_port, minusA_s_10_port, minusA_s_9_port, minusA_s_8_port, 
      minusA_s_7_port, minusA_s_6_port, minusA_s_5_port, minusA_s_4_port, 
      minusA_s_3_port, minusA_s_2_port, minusA_s_1_port, minusA_s_0_port, 
      minus2A_s_63_port, minus2A_s_62_port, minus2A_s_61_port, 
      minus2A_s_60_port, minus2A_s_59_port, minus2A_s_58_port, 
      minus2A_s_57_port, minus2A_s_56_port, minus2A_s_55_port, 
      minus2A_s_54_port, minus2A_s_53_port, minus2A_s_52_port, 
      minus2A_s_51_port, minus2A_s_50_port, minus2A_s_49_port, 
      minus2A_s_48_port, minus2A_s_47_port, minus2A_s_46_port, 
      minus2A_s_45_port, minus2A_s_44_port, minus2A_s_43_port, 
      minus2A_s_42_port, minus2A_s_41_port, minus2A_s_40_port, 
      minus2A_s_39_port, minus2A_s_38_port, minus2A_s_37_port, 
      minus2A_s_36_port, minus2A_s_35_port, minus2A_s_34_port, 
      minus2A_s_33_port, minus2A_s_32_port, minus2A_s_31_port, 
      minus2A_s_30_port, minus2A_s_29_port, minus2A_s_28_port, 
      minus2A_s_27_port, minus2A_s_26_port, minus2A_s_25_port, 
      minus2A_s_24_port, minus2A_s_23_port, minus2A_s_22_port, 
      minus2A_s_21_port, minus2A_s_20_port, minus2A_s_19_port, 
      minus2A_s_18_port, minus2A_s_17_port, minus2A_s_16_port, 
      minus2A_s_15_port, minus2A_s_14_port, minus2A_s_13_port, 
      minus2A_s_12_port, minus2A_s_11_port, minus2A_s_10_port, minus2A_s_9_port
      , minus2A_s_8_port, minus2A_s_7_port, minus2A_s_6_port, minus2A_s_5_port,
      minus2A_s_4_port, minus2A_s_3_port, minus2A_s_2_port, minus2A_s_1_port, 
      minus2A_s_0_port, nextA_0_port, nextA_57_port, n_3220 : std_logic;

begin
   nextA <= ( nextA_63_port, nextA_62_port, nextA_61_port, nextA_60_port, 
      nextA_59_port, nextA_58_port, nextA_57_port, nextA_56_port, nextA_55_port
      , nextA_54_port, nextA_53_port, nextA_52_port, nextA_51_port, 
      nextA_50_port, nextA_49_port, nextA_48_port, nextA_47_port, nextA_46_port
      , nextA_45_port, nextA_44_port, nextA_43_port, nextA_42_port, 
      nextA_41_port, nextA_40_port, nextA_39_port, nextA_38_port, nextA_37_port
      , nextA_36_port, nextA_35_port, nextA_34_port, nextA_33_port, 
      nextA_32_port, nextA_31_port, nextA_30_port, nextA_29_port, nextA_28_port
      , nextA_27_port, nextA_26_port, nextA_25_port, nextA_24_port, 
      nextA_23_port, nextA_22_port, nextA_21_port, nextA_20_port, nextA_19_port
      , nextA_18_port, nextA_17_port, nextA_16_port, nextA_15_port, 
      nextA_14_port, nextA_13_port, nextA_12_port, nextA_11_port, nextA_10_port
      , nextA_9_port, nextA_8_port, nextA_7_port, nextA_6_port, nextA_5_port, 
      nextA_4_port, nextA_3_port, nextA_2_port, nextA_1_port, nextA_0_port );
   
   nextA_0_port <= '0';
   encoder_1 : encoder_N64_RADIX3_0 port map( X(2) => encoderIn(2), X(1) => 
                           encoderIn(1), X(0) => encoderIn(0), Z(2) => 
                           encoder_to_mux_2_port, Z(1) => encoder_to_mux_1_port
                           , Z(0) => encoder_to_mux_0_port);
   ShiftnCompl_special_1 : ShiftnCompl_special_N64 port map( plusA(63) => A(63)
                           , plusA(62) => A(62), plusA(61) => A(61), plusA(60) 
                           => A(60), plusA(59) => A(59), plusA(58) => A(58), 
                           plusA(57) => A(57), plusA(56) => A(56), plusA(55) =>
                           A(55), plusA(54) => A(54), plusA(53) => A(53), 
                           plusA(52) => A(52), plusA(51) => A(51), plusA(50) =>
                           A(50), plusA(49) => A(49), plusA(48) => A(48), 
                           plusA(47) => A(47), plusA(46) => A(46), plusA(45) =>
                           A(45), plusA(44) => A(44), plusA(43) => A(43), 
                           plusA(42) => A(42), plusA(41) => A(41), plusA(40) =>
                           A(40), plusA(39) => A(39), plusA(38) => A(38), 
                           plusA(37) => A(37), plusA(36) => A(36), plusA(35) =>
                           A(35), plusA(34) => A(34), plusA(33) => A(33), 
                           plusA(32) => A(32), plusA(31) => A(31), plusA(30) =>
                           A(30), plusA(29) => A(29), plusA(28) => A(28), 
                           plusA(27) => A(27), plusA(26) => A(26), plusA(25) =>
                           A(25), plusA(24) => A(24), plusA(23) => A(23), 
                           plusA(22) => A(22), plusA(21) => A(21), plusA(20) =>
                           A(20), plusA(19) => A(19), plusA(18) => A(18), 
                           plusA(17) => A(17), plusA(16) => A(16), plusA(15) =>
                           A(15), plusA(14) => A(14), plusA(13) => A(13), 
                           plusA(12) => A(12), plusA(11) => A(11), plusA(10) =>
                           A(10), plusA(9) => A(9), plusA(8) => A(8), plusA(7) 
                           => A(7), plusA(6) => A(6), plusA(5) => A(5), 
                           plusA(4) => A(4), plusA(3) => A(3), plusA(2) => A(2)
                           , plusA(1) => A(1), plusA(0) => A(0), plusA_out(63) 
                           => plusA_s_63_port, plusA_out(62) => plusA_s_62_port
                           , plusA_out(61) => plusA_s_61_port, plusA_out(60) =>
                           plusA_s_60_port, plusA_out(59) => plusA_s_59_port, 
                           plusA_out(58) => plusA_s_58_port, plusA_out(57) => 
                           plusA_s_57_port, plusA_out(56) => plusA_s_56_port, 
                           plusA_out(55) => plusA_s_55_port, plusA_out(54) => 
                           plusA_s_54_port, plusA_out(53) => plusA_s_53_port, 
                           plusA_out(52) => plusA_s_52_port, plusA_out(51) => 
                           plusA_s_51_port, plusA_out(50) => plusA_s_50_port, 
                           plusA_out(49) => plusA_s_49_port, plusA_out(48) => 
                           plusA_s_48_port, plusA_out(47) => plusA_s_47_port, 
                           plusA_out(46) => plusA_s_46_port, plusA_out(45) => 
                           plusA_s_45_port, plusA_out(44) => plusA_s_44_port, 
                           plusA_out(43) => plusA_s_43_port, plusA_out(42) => 
                           plusA_s_42_port, plusA_out(41) => plusA_s_41_port, 
                           plusA_out(40) => plusA_s_40_port, plusA_out(39) => 
                           plusA_s_39_port, plusA_out(38) => plusA_s_38_port, 
                           plusA_out(37) => plusA_s_37_port, plusA_out(36) => 
                           plusA_s_36_port, plusA_out(35) => plusA_s_35_port, 
                           plusA_out(34) => plusA_s_34_port, plusA_out(33) => 
                           plusA_s_33_port, plusA_out(32) => plusA_s_32_port, 
                           plusA_out(31) => plusA_s_31_port, plusA_out(30) => 
                           plusA_s_30_port, plusA_out(29) => plusA_s_29_port, 
                           plusA_out(28) => plusA_s_28_port, plusA_out(27) => 
                           plusA_s_27_port, plusA_out(26) => plusA_s_26_port, 
                           plusA_out(25) => plusA_s_25_port, plusA_out(24) => 
                           plusA_s_24_port, plusA_out(23) => plusA_s_23_port, 
                           plusA_out(22) => plusA_s_22_port, plusA_out(21) => 
                           plusA_s_21_port, plusA_out(20) => plusA_s_20_port, 
                           plusA_out(19) => plusA_s_19_port, plusA_out(18) => 
                           plusA_s_18_port, plusA_out(17) => plusA_s_17_port, 
                           plusA_out(16) => plusA_s_16_port, plusA_out(15) => 
                           plusA_s_15_port, plusA_out(14) => plusA_s_14_port, 
                           plusA_out(13) => plusA_s_13_port, plusA_out(12) => 
                           plusA_s_12_port, plusA_out(11) => plusA_s_11_port, 
                           plusA_out(10) => plusA_s_10_port, plusA_out(9) => 
                           plusA_s_9_port, plusA_out(8) => plusA_s_8_port, 
                           plusA_out(7) => plusA_s_7_port, plusA_out(6) => 
                           plusA_s_6_port, plusA_out(5) => plusA_s_5_port, 
                           plusA_out(4) => plusA_s_4_port, plusA_out(3) => 
                           plusA_s_3_port, plusA_out(2) => plusA_s_2_port, 
                           plusA_out(1) => plusA_s_1_port, plusA_out(0) => 
                           plusA_s_0_port, minusA_out(63) => minusA_s_63_port, 
                           minusA_out(62) => minusA_s_62_port, minusA_out(61) 
                           => minusA_s_61_port, minusA_out(60) => 
                           minusA_s_60_port, minusA_out(59) => minusA_s_59_port
                           , minusA_out(58) => minusA_s_58_port, minusA_out(57)
                           => minusA_s_57_port, minusA_out(56) => 
                           minusA_s_56_port, minusA_out(55) => minusA_s_55_port
                           , minusA_out(54) => minusA_s_54_port, minusA_out(53)
                           => minusA_s_53_port, minusA_out(52) => 
                           minusA_s_52_port, minusA_out(51) => minusA_s_51_port
                           , minusA_out(50) => minusA_s_50_port, minusA_out(49)
                           => minusA_s_49_port, minusA_out(48) => 
                           minusA_s_48_port, minusA_out(47) => minusA_s_47_port
                           , minusA_out(46) => minusA_s_46_port, minusA_out(45)
                           => minusA_s_45_port, minusA_out(44) => 
                           minusA_s_44_port, minusA_out(43) => minusA_s_43_port
                           , minusA_out(42) => minusA_s_42_port, minusA_out(41)
                           => minusA_s_41_port, minusA_out(40) => 
                           minusA_s_40_port, minusA_out(39) => minusA_s_39_port
                           , minusA_out(38) => minusA_s_38_port, minusA_out(37)
                           => minusA_s_37_port, minusA_out(36) => 
                           minusA_s_36_port, minusA_out(35) => minusA_s_35_port
                           , minusA_out(34) => minusA_s_34_port, minusA_out(33)
                           => minusA_s_33_port, minusA_out(32) => 
                           minusA_s_32_port, minusA_out(31) => minusA_s_31_port
                           , minusA_out(30) => minusA_s_30_port, minusA_out(29)
                           => minusA_s_29_port, minusA_out(28) => 
                           minusA_s_28_port, minusA_out(27) => minusA_s_27_port
                           , minusA_out(26) => minusA_s_26_port, minusA_out(25)
                           => minusA_s_25_port, minusA_out(24) => 
                           minusA_s_24_port, minusA_out(23) => minusA_s_23_port
                           , minusA_out(22) => minusA_s_22_port, minusA_out(21)
                           => minusA_s_21_port, minusA_out(20) => 
                           minusA_s_20_port, minusA_out(19) => minusA_s_19_port
                           , minusA_out(18) => minusA_s_18_port, minusA_out(17)
                           => minusA_s_17_port, minusA_out(16) => 
                           minusA_s_16_port, minusA_out(15) => minusA_s_15_port
                           , minusA_out(14) => minusA_s_14_port, minusA_out(13)
                           => minusA_s_13_port, minusA_out(12) => 
                           minusA_s_12_port, minusA_out(11) => minusA_s_11_port
                           , minusA_out(10) => minusA_s_10_port, minusA_out(9) 
                           => minusA_s_9_port, minusA_out(8) => minusA_s_8_port
                           , minusA_out(7) => minusA_s_7_port, minusA_out(6) =>
                           minusA_s_6_port, minusA_out(5) => minusA_s_5_port, 
                           minusA_out(4) => minusA_s_4_port, minusA_out(3) => 
                           minusA_s_3_port, minusA_out(2) => minusA_s_2_port, 
                           minusA_out(1) => minusA_s_1_port, minusA_out(0) => 
                           minusA_s_0_port, plus2A_out(63) => nextA_63_port, 
                           plus2A_out(62) => nextA_62_port, plus2A_out(61) => 
                           nextA_61_port, plus2A_out(60) => nextA_60_port, 
                           plus2A_out(59) => nextA_59_port, plus2A_out(58) => 
                           nextA_58_port, plus2A_out(57) => n3, plus2A_out(56) 
                           => nextA_56_port, plus2A_out(55) => nextA_55_port, 
                           plus2A_out(54) => nextA_54_port, plus2A_out(53) => 
                           nextA_53_port, plus2A_out(52) => nextA_52_port, 
                           plus2A_out(51) => nextA_51_port, plus2A_out(50) => 
                           nextA_50_port, plus2A_out(49) => nextA_49_port, 
                           plus2A_out(48) => nextA_48_port, plus2A_out(47) => 
                           nextA_47_port, plus2A_out(46) => nextA_46_port, 
                           plus2A_out(45) => nextA_45_port, plus2A_out(44) => 
                           nextA_44_port, plus2A_out(43) => nextA_43_port, 
                           plus2A_out(42) => nextA_42_port, plus2A_out(41) => 
                           nextA_41_port, plus2A_out(40) => nextA_40_port, 
                           plus2A_out(39) => nextA_39_port, plus2A_out(38) => 
                           nextA_38_port, plus2A_out(37) => nextA_37_port, 
                           plus2A_out(36) => nextA_36_port, plus2A_out(35) => 
                           nextA_35_port, plus2A_out(34) => nextA_34_port, 
                           plus2A_out(33) => nextA_33_port, plus2A_out(32) => 
                           nextA_32_port, plus2A_out(31) => nextA_31_port, 
                           plus2A_out(30) => nextA_30_port, plus2A_out(29) => 
                           nextA_29_port, plus2A_out(28) => nextA_28_port, 
                           plus2A_out(27) => nextA_27_port, plus2A_out(26) => 
                           nextA_26_port, plus2A_out(25) => nextA_25_port, 
                           plus2A_out(24) => nextA_24_port, plus2A_out(23) => 
                           nextA_23_port, plus2A_out(22) => nextA_22_port, 
                           plus2A_out(21) => nextA_21_port, plus2A_out(20) => 
                           nextA_20_port, plus2A_out(19) => nextA_19_port, 
                           plus2A_out(18) => nextA_18_port, plus2A_out(17) => 
                           nextA_17_port, plus2A_out(16) => nextA_16_port, 
                           plus2A_out(15) => nextA_15_port, plus2A_out(14) => 
                           nextA_14_port, plus2A_out(13) => nextA_13_port, 
                           plus2A_out(12) => nextA_12_port, plus2A_out(11) => 
                           nextA_11_port, plus2A_out(10) => nextA_10_port, 
                           plus2A_out(9) => nextA_9_port, plus2A_out(8) => 
                           nextA_8_port, plus2A_out(7) => nextA_7_port, 
                           plus2A_out(6) => nextA_6_port, plus2A_out(5) => 
                           nextA_5_port, plus2A_out(4) => nextA_4_port, 
                           plus2A_out(3) => nextA_3_port, plus2A_out(2) => 
                           nextA_2_port, plus2A_out(1) => nextA_1_port, 
                           plus2A_out(0) => n_3220, minus2A_out(63) => 
                           minus2A_s_63_port, minus2A_out(62) => 
                           minus2A_s_62_port, minus2A_out(61) => 
                           minus2A_s_61_port, minus2A_out(60) => 
                           minus2A_s_60_port, minus2A_out(59) => 
                           minus2A_s_59_port, minus2A_out(58) => 
                           minus2A_s_58_port, minus2A_out(57) => 
                           minus2A_s_57_port, minus2A_out(56) => 
                           minus2A_s_56_port, minus2A_out(55) => 
                           minus2A_s_55_port, minus2A_out(54) => 
                           minus2A_s_54_port, minus2A_out(53) => 
                           minus2A_s_53_port, minus2A_out(52) => 
                           minus2A_s_52_port, minus2A_out(51) => 
                           minus2A_s_51_port, minus2A_out(50) => 
                           minus2A_s_50_port, minus2A_out(49) => 
                           minus2A_s_49_port, minus2A_out(48) => 
                           minus2A_s_48_port, minus2A_out(47) => 
                           minus2A_s_47_port, minus2A_out(46) => 
                           minus2A_s_46_port, minus2A_out(45) => 
                           minus2A_s_45_port, minus2A_out(44) => 
                           minus2A_s_44_port, minus2A_out(43) => 
                           minus2A_s_43_port, minus2A_out(42) => 
                           minus2A_s_42_port, minus2A_out(41) => 
                           minus2A_s_41_port, minus2A_out(40) => 
                           minus2A_s_40_port, minus2A_out(39) => 
                           minus2A_s_39_port, minus2A_out(38) => 
                           minus2A_s_38_port, minus2A_out(37) => 
                           minus2A_s_37_port, minus2A_out(36) => 
                           minus2A_s_36_port, minus2A_out(35) => 
                           minus2A_s_35_port, minus2A_out(34) => 
                           minus2A_s_34_port, minus2A_out(33) => 
                           minus2A_s_33_port, minus2A_out(32) => 
                           minus2A_s_32_port, minus2A_out(31) => 
                           minus2A_s_31_port, minus2A_out(30) => 
                           minus2A_s_30_port, minus2A_out(29) => 
                           minus2A_s_29_port, minus2A_out(28) => 
                           minus2A_s_28_port, minus2A_out(27) => 
                           minus2A_s_27_port, minus2A_out(26) => 
                           minus2A_s_26_port, minus2A_out(25) => 
                           minus2A_s_25_port, minus2A_out(24) => 
                           minus2A_s_24_port, minus2A_out(23) => 
                           minus2A_s_23_port, minus2A_out(22) => 
                           minus2A_s_22_port, minus2A_out(21) => 
                           minus2A_s_21_port, minus2A_out(20) => 
                           minus2A_s_20_port, minus2A_out(19) => 
                           minus2A_s_19_port, minus2A_out(18) => 
                           minus2A_s_18_port, minus2A_out(17) => 
                           minus2A_s_17_port, minus2A_out(16) => 
                           minus2A_s_16_port, minus2A_out(15) => 
                           minus2A_s_15_port, minus2A_out(14) => 
                           minus2A_s_14_port, minus2A_out(13) => 
                           minus2A_s_13_port, minus2A_out(12) => 
                           minus2A_s_12_port, minus2A_out(11) => 
                           minus2A_s_11_port, minus2A_out(10) => 
                           minus2A_s_10_port, minus2A_out(9) => 
                           minus2A_s_9_port, minus2A_out(8) => minus2A_s_8_port
                           , minus2A_out(7) => minus2A_s_7_port, minus2A_out(6)
                           => minus2A_s_6_port, minus2A_out(5) => 
                           minus2A_s_5_port, minus2A_out(4) => minus2A_s_4_port
                           , minus2A_out(3) => minus2A_s_3_port, minus2A_out(2)
                           => minus2A_s_2_port, minus2A_out(1) => 
                           minus2A_s_1_port, minus2A_out(0) => minus2A_s_0_port
                           );
   mux_1 : MUX_GENERIC_N64_RADIX3_0 port map( plusA(63) => plusA_s_63_port, 
                           plusA(62) => plusA_s_62_port, plusA(61) => 
                           plusA_s_61_port, plusA(60) => plusA_s_60_port, 
                           plusA(59) => plusA_s_59_port, plusA(58) => 
                           plusA_s_58_port, plusA(57) => plusA_s_57_port, 
                           plusA(56) => plusA_s_56_port, plusA(55) => 
                           plusA_s_55_port, plusA(54) => plusA_s_54_port, 
                           plusA(53) => plusA_s_53_port, plusA(52) => 
                           plusA_s_52_port, plusA(51) => plusA_s_51_port, 
                           plusA(50) => plusA_s_50_port, plusA(49) => 
                           plusA_s_49_port, plusA(48) => plusA_s_48_port, 
                           plusA(47) => plusA_s_47_port, plusA(46) => 
                           plusA_s_46_port, plusA(45) => plusA_s_45_port, 
                           plusA(44) => plusA_s_44_port, plusA(43) => 
                           plusA_s_43_port, plusA(42) => plusA_s_42_port, 
                           plusA(41) => plusA_s_41_port, plusA(40) => 
                           plusA_s_40_port, plusA(39) => plusA_s_39_port, 
                           plusA(38) => plusA_s_38_port, plusA(37) => 
                           plusA_s_37_port, plusA(36) => plusA_s_36_port, 
                           plusA(35) => plusA_s_35_port, plusA(34) => 
                           plusA_s_34_port, plusA(33) => plusA_s_33_port, 
                           plusA(32) => plusA_s_32_port, plusA(31) => 
                           plusA_s_31_port, plusA(30) => plusA_s_30_port, 
                           plusA(29) => plusA_s_29_port, plusA(28) => 
                           plusA_s_28_port, plusA(27) => plusA_s_27_port, 
                           plusA(26) => plusA_s_26_port, plusA(25) => 
                           plusA_s_25_port, plusA(24) => plusA_s_24_port, 
                           plusA(23) => plusA_s_23_port, plusA(22) => 
                           plusA_s_22_port, plusA(21) => plusA_s_21_port, 
                           plusA(20) => plusA_s_20_port, plusA(19) => 
                           plusA_s_19_port, plusA(18) => plusA_s_18_port, 
                           plusA(17) => plusA_s_17_port, plusA(16) => 
                           plusA_s_16_port, plusA(15) => plusA_s_15_port, 
                           plusA(14) => plusA_s_14_port, plusA(13) => 
                           plusA_s_13_port, plusA(12) => plusA_s_12_port, 
                           plusA(11) => plusA_s_11_port, plusA(10) => 
                           plusA_s_10_port, plusA(9) => plusA_s_9_port, 
                           plusA(8) => plusA_s_8_port, plusA(7) => 
                           plusA_s_7_port, plusA(6) => plusA_s_6_port, plusA(5)
                           => plusA_s_5_port, plusA(4) => plusA_s_4_port, 
                           plusA(3) => plusA_s_3_port, plusA(2) => 
                           plusA_s_2_port, plusA(1) => plusA_s_1_port, plusA(0)
                           => plusA_s_0_port, minusA(63) => minusA_s_63_port, 
                           minusA(62) => minusA_s_62_port, minusA(61) => 
                           minusA_s_61_port, minusA(60) => minusA_s_60_port, 
                           minusA(59) => minusA_s_59_port, minusA(58) => 
                           minusA_s_58_port, minusA(57) => minusA_s_57_port, 
                           minusA(56) => minusA_s_56_port, minusA(55) => 
                           minusA_s_55_port, minusA(54) => minusA_s_54_port, 
                           minusA(53) => minusA_s_53_port, minusA(52) => 
                           minusA_s_52_port, minusA(51) => minusA_s_51_port, 
                           minusA(50) => minusA_s_50_port, minusA(49) => 
                           minusA_s_49_port, minusA(48) => minusA_s_48_port, 
                           minusA(47) => minusA_s_47_port, minusA(46) => 
                           minusA_s_46_port, minusA(45) => minusA_s_45_port, 
                           minusA(44) => minusA_s_44_port, minusA(43) => 
                           minusA_s_43_port, minusA(42) => minusA_s_42_port, 
                           minusA(41) => minusA_s_41_port, minusA(40) => 
                           minusA_s_40_port, minusA(39) => minusA_s_39_port, 
                           minusA(38) => minusA_s_38_port, minusA(37) => 
                           minusA_s_37_port, minusA(36) => minusA_s_36_port, 
                           minusA(35) => minusA_s_35_port, minusA(34) => 
                           minusA_s_34_port, minusA(33) => minusA_s_33_port, 
                           minusA(32) => minusA_s_32_port, minusA(31) => 
                           minusA_s_31_port, minusA(30) => minusA_s_30_port, 
                           minusA(29) => minusA_s_29_port, minusA(28) => 
                           minusA_s_28_port, minusA(27) => minusA_s_27_port, 
                           minusA(26) => minusA_s_26_port, minusA(25) => 
                           minusA_s_25_port, minusA(24) => minusA_s_24_port, 
                           minusA(23) => minusA_s_23_port, minusA(22) => 
                           minusA_s_22_port, minusA(21) => minusA_s_21_port, 
                           minusA(20) => minusA_s_20_port, minusA(19) => 
                           minusA_s_19_port, minusA(18) => minusA_s_18_port, 
                           minusA(17) => minusA_s_17_port, minusA(16) => 
                           minusA_s_16_port, minusA(15) => minusA_s_15_port, 
                           minusA(14) => minusA_s_14_port, minusA(13) => 
                           minusA_s_13_port, minusA(12) => minusA_s_12_port, 
                           minusA(11) => minusA_s_11_port, minusA(10) => 
                           minusA_s_10_port, minusA(9) => minusA_s_9_port, 
                           minusA(8) => minusA_s_8_port, minusA(7) => 
                           minusA_s_7_port, minusA(6) => minusA_s_6_port, 
                           minusA(5) => minusA_s_5_port, minusA(4) => 
                           minusA_s_4_port, minusA(3) => minusA_s_3_port, 
                           minusA(2) => minusA_s_2_port, minusA(1) => 
                           minusA_s_1_port, minusA(0) => minusA_s_0_port, 
                           plus2A(63) => nextA_63_port, plus2A(62) => 
                           nextA_62_port, plus2A(61) => nextA_61_port, 
                           plus2A(60) => nextA_60_port, plus2A(59) => 
                           nextA_59_port, plus2A(58) => nextA_58_port, 
                           plus2A(57) => nextA_57_port, plus2A(56) => 
                           nextA_56_port, plus2A(55) => nextA_55_port, 
                           plus2A(54) => nextA_54_port, plus2A(53) => 
                           nextA_53_port, plus2A(52) => nextA_52_port, 
                           plus2A(51) => nextA_51_port, plus2A(50) => 
                           nextA_50_port, plus2A(49) => nextA_49_port, 
                           plus2A(48) => nextA_48_port, plus2A(47) => 
                           nextA_47_port, plus2A(46) => nextA_46_port, 
                           plus2A(45) => nextA_45_port, plus2A(44) => 
                           nextA_44_port, plus2A(43) => nextA_43_port, 
                           plus2A(42) => nextA_42_port, plus2A(41) => 
                           nextA_41_port, plus2A(40) => nextA_40_port, 
                           plus2A(39) => nextA_39_port, plus2A(38) => 
                           nextA_38_port, plus2A(37) => nextA_37_port, 
                           plus2A(36) => nextA_36_port, plus2A(35) => 
                           nextA_35_port, plus2A(34) => nextA_34_port, 
                           plus2A(33) => nextA_33_port, plus2A(32) => 
                           nextA_32_port, plus2A(31) => nextA_31_port, 
                           plus2A(30) => nextA_30_port, plus2A(29) => 
                           nextA_29_port, plus2A(28) => nextA_28_port, 
                           plus2A(27) => nextA_27_port, plus2A(26) => 
                           nextA_26_port, plus2A(25) => nextA_25_port, 
                           plus2A(24) => nextA_24_port, plus2A(23) => 
                           nextA_23_port, plus2A(22) => nextA_22_port, 
                           plus2A(21) => nextA_21_port, plus2A(20) => 
                           nextA_20_port, plus2A(19) => nextA_19_port, 
                           plus2A(18) => nextA_18_port, plus2A(17) => 
                           nextA_17_port, plus2A(16) => nextA_16_port, 
                           plus2A(15) => nextA_15_port, plus2A(14) => 
                           nextA_14_port, plus2A(13) => nextA_13_port, 
                           plus2A(12) => nextA_12_port, plus2A(11) => 
                           nextA_11_port, plus2A(10) => nextA_10_port, 
                           plus2A(9) => nextA_9_port, plus2A(8) => nextA_8_port
                           , plus2A(7) => nextA_7_port, plus2A(6) => 
                           nextA_6_port, plus2A(5) => nextA_5_port, plus2A(4) 
                           => nextA_4_port, plus2A(3) => nextA_3_port, 
                           plus2A(2) => nextA_2_port, plus2A(1) => nextA_1_port
                           , plus2A(0) => nextA_0_port, minus2A(63) => 
                           minus2A_s_63_port, minus2A(62) => minus2A_s_62_port,
                           minus2A(61) => minus2A_s_61_port, minus2A(60) => 
                           minus2A_s_60_port, minus2A(59) => minus2A_s_59_port,
                           minus2A(58) => minus2A_s_58_port, minus2A(57) => 
                           minus2A_s_57_port, minus2A(56) => minus2A_s_56_port,
                           minus2A(55) => minus2A_s_55_port, minus2A(54) => 
                           minus2A_s_54_port, minus2A(53) => minus2A_s_53_port,
                           minus2A(52) => minus2A_s_52_port, minus2A(51) => 
                           minus2A_s_51_port, minus2A(50) => minus2A_s_50_port,
                           minus2A(49) => minus2A_s_49_port, minus2A(48) => 
                           minus2A_s_48_port, minus2A(47) => minus2A_s_47_port,
                           minus2A(46) => minus2A_s_46_port, minus2A(45) => 
                           minus2A_s_45_port, minus2A(44) => minus2A_s_44_port,
                           minus2A(43) => minus2A_s_43_port, minus2A(42) => 
                           minus2A_s_42_port, minus2A(41) => minus2A_s_41_port,
                           minus2A(40) => minus2A_s_40_port, minus2A(39) => 
                           minus2A_s_39_port, minus2A(38) => minus2A_s_38_port,
                           minus2A(37) => minus2A_s_37_port, minus2A(36) => 
                           minus2A_s_36_port, minus2A(35) => minus2A_s_35_port,
                           minus2A(34) => minus2A_s_34_port, minus2A(33) => 
                           minus2A_s_33_port, minus2A(32) => minus2A_s_32_port,
                           minus2A(31) => minus2A_s_31_port, minus2A(30) => 
                           minus2A_s_30_port, minus2A(29) => minus2A_s_29_port,
                           minus2A(28) => minus2A_s_28_port, minus2A(27) => 
                           minus2A_s_27_port, minus2A(26) => minus2A_s_26_port,
                           minus2A(25) => minus2A_s_25_port, minus2A(24) => 
                           minus2A_s_24_port, minus2A(23) => minus2A_s_23_port,
                           minus2A(22) => minus2A_s_22_port, minus2A(21) => 
                           minus2A_s_21_port, minus2A(20) => minus2A_s_20_port,
                           minus2A(19) => minus2A_s_19_port, minus2A(18) => 
                           minus2A_s_18_port, minus2A(17) => minus2A_s_17_port,
                           minus2A(16) => minus2A_s_16_port, minus2A(15) => 
                           minus2A_s_15_port, minus2A(14) => minus2A_s_14_port,
                           minus2A(13) => minus2A_s_13_port, minus2A(12) => 
                           minus2A_s_12_port, minus2A(11) => minus2A_s_11_port,
                           minus2A(10) => minus2A_s_10_port, minus2A(9) => 
                           minus2A_s_9_port, minus2A(8) => minus2A_s_8_port, 
                           minus2A(7) => minus2A_s_7_port, minus2A(6) => 
                           minus2A_s_6_port, minus2A(5) => minus2A_s_5_port, 
                           minus2A(4) => minus2A_s_4_port, minus2A(3) => 
                           minus2A_s_3_port, minus2A(2) => minus2A_s_2_port, 
                           minus2A(1) => minus2A_s_1_port, minus2A(0) => 
                           minus2A_s_0_port, SEL(2) => encoder_to_mux_2_port, 
                           SEL(1) => encoder_to_mux_1_port, SEL(0) => 
                           encoder_to_mux_0_port, Y(63) => nextSum(63), Y(62) 
                           => nextSum(62), Y(61) => nextSum(61), Y(60) => 
                           nextSum(60), Y(59) => nextSum(59), Y(58) => 
                           nextSum(58), Y(57) => nextSum(57), Y(56) => 
                           nextSum(56), Y(55) => nextSum(55), Y(54) => 
                           nextSum(54), Y(53) => nextSum(53), Y(52) => 
                           nextSum(52), Y(51) => nextSum(51), Y(50) => 
                           nextSum(50), Y(49) => nextSum(49), Y(48) => 
                           nextSum(48), Y(47) => nextSum(47), Y(46) => 
                           nextSum(46), Y(45) => nextSum(45), Y(44) => 
                           nextSum(44), Y(43) => nextSum(43), Y(42) => 
                           nextSum(42), Y(41) => nextSum(41), Y(40) => 
                           nextSum(40), Y(39) => nextSum(39), Y(38) => 
                           nextSum(38), Y(37) => nextSum(37), Y(36) => 
                           nextSum(36), Y(35) => nextSum(35), Y(34) => 
                           nextSum(34), Y(33) => nextSum(33), Y(32) => 
                           nextSum(32), Y(31) => nextSum(31), Y(30) => 
                           nextSum(30), Y(29) => nextSum(29), Y(28) => 
                           nextSum(28), Y(27) => nextSum(27), Y(26) => 
                           nextSum(26), Y(25) => nextSum(25), Y(24) => 
                           nextSum(24), Y(23) => nextSum(23), Y(22) => 
                           nextSum(22), Y(21) => nextSum(21), Y(20) => 
                           nextSum(20), Y(19) => nextSum(19), Y(18) => 
                           nextSum(18), Y(17) => nextSum(17), Y(16) => 
                           nextSum(16), Y(15) => nextSum(15), Y(14) => 
                           nextSum(14), Y(13) => nextSum(13), Y(12) => 
                           nextSum(12), Y(11) => nextSum(11), Y(10) => 
                           nextSum(10), Y(9) => nextSum(9), Y(8) => nextSum(8),
                           Y(7) => nextSum(7), Y(6) => nextSum(6), Y(5) => 
                           nextSum(5), Y(4) => nextSum(4), Y(3) => nextSum(3), 
                           Y(2) => nextSum(2), Y(1) => nextSum(1), Y(0) => 
                           nextSum(0));
   U2 : BUF_X1 port map( A => n3, Z => nextA_57_port);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Booth.all;

entity Booth is

   port( A, B : in std_logic_vector (31 downto 0);  P : out std_logic_vector 
         (63 downto 0));

end Booth;

architecture SYN_booth_struct of Booth is

   component booth_mul_row_N64_RADIX3_1
      port( prevA, prevSum : in std_logic_vector (63 downto 0);  encoderIn : in
            std_logic_vector (2 downto 0);  nextA, nextSum : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component booth_mul_row_N64_RADIX3_2
      port( prevA, prevSum : in std_logic_vector (63 downto 0);  encoderIn : in
            std_logic_vector (2 downto 0);  nextA, nextSum : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component booth_mul_row_N64_RADIX3_3
      port( prevA, prevSum : in std_logic_vector (63 downto 0);  encoderIn : in
            std_logic_vector (2 downto 0);  nextA, nextSum : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component booth_mul_row_N64_RADIX3_4
      port( prevA, prevSum : in std_logic_vector (63 downto 0);  encoderIn : in
            std_logic_vector (2 downto 0);  nextA, nextSum : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component booth_mul_row_N64_RADIX3_5
      port( prevA, prevSum : in std_logic_vector (63 downto 0);  encoderIn : in
            std_logic_vector (2 downto 0);  nextA, nextSum : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component booth_mul_row_N64_RADIX3_6
      port( prevA, prevSum : in std_logic_vector (63 downto 0);  encoderIn : in
            std_logic_vector (2 downto 0);  nextA, nextSum : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component booth_mul_row_N64_RADIX3_7
      port( prevA, prevSum : in std_logic_vector (63 downto 0);  encoderIn : in
            std_logic_vector (2 downto 0);  nextA, nextSum : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component booth_mul_row_N64_RADIX3_8
      port( prevA, prevSum : in std_logic_vector (63 downto 0);  encoderIn : in
            std_logic_vector (2 downto 0);  nextA, nextSum : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component booth_mul_row_N64_RADIX3_9
      port( prevA, prevSum : in std_logic_vector (63 downto 0);  encoderIn : in
            std_logic_vector (2 downto 0);  nextA, nextSum : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component booth_mul_row_N64_RADIX3_10
      port( prevA, prevSum : in std_logic_vector (63 downto 0);  encoderIn : in
            std_logic_vector (2 downto 0);  nextA, nextSum : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component booth_mul_row_N64_RADIX3_11
      port( prevA, prevSum : in std_logic_vector (63 downto 0);  encoderIn : in
            std_logic_vector (2 downto 0);  nextA, nextSum : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component booth_mul_row_N64_RADIX3_12
      port( prevA, prevSum : in std_logic_vector (63 downto 0);  encoderIn : in
            std_logic_vector (2 downto 0);  nextA, nextSum : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component booth_mul_row_N64_RADIX3_13
      port( prevA, prevSum : in std_logic_vector (63 downto 0);  encoderIn : in
            std_logic_vector (2 downto 0);  nextA, nextSum : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component booth_mul_row_N64_RADIX3_14
      port( prevA, prevSum : in std_logic_vector (63 downto 0);  encoderIn : in
            std_logic_vector (2 downto 0);  nextA, nextSum : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component booth_mul_row_N64_RADIX3_0
      port( prevA, prevSum : in std_logic_vector (63 downto 0);  encoderIn : in
            std_logic_vector (2 downto 0);  nextA, nextSum : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component booth_mul_row_special_N64_RADIX3
      port( A : in std_logic_vector (63 downto 0);  encoderIn : in 
            std_logic_vector (2 downto 0);  nextA, nextSum : out 
            std_logic_vector (63 downto 0));
   end component;
   
   signal X_Logic0_port, sigMatrix_0_127_port, sigMatrix_0_126_port, 
      sigMatrix_0_125_port, sigMatrix_0_124_port, sigMatrix_0_123_port, 
      sigMatrix_0_122_port, sigMatrix_0_121_port, sigMatrix_0_120_port, 
      sigMatrix_0_119_port, sigMatrix_0_118_port, sigMatrix_0_117_port, 
      sigMatrix_0_116_port, sigMatrix_0_115_port, sigMatrix_0_114_port, 
      sigMatrix_0_113_port, sigMatrix_0_112_port, sigMatrix_0_111_port, 
      sigMatrix_0_110_port, sigMatrix_0_109_port, sigMatrix_0_108_port, 
      sigMatrix_0_107_port, sigMatrix_0_106_port, sigMatrix_0_105_port, 
      sigMatrix_0_104_port, sigMatrix_0_103_port, sigMatrix_0_102_port, 
      sigMatrix_0_101_port, sigMatrix_0_100_port, sigMatrix_0_99_port, 
      sigMatrix_0_98_port, sigMatrix_0_97_port, sigMatrix_0_96_port, 
      sigMatrix_0_95_port, sigMatrix_0_94_port, sigMatrix_0_93_port, 
      sigMatrix_0_92_port, sigMatrix_0_91_port, sigMatrix_0_90_port, 
      sigMatrix_0_89_port, sigMatrix_0_88_port, sigMatrix_0_87_port, 
      sigMatrix_0_86_port, sigMatrix_0_85_port, sigMatrix_0_84_port, 
      sigMatrix_0_83_port, sigMatrix_0_82_port, sigMatrix_0_81_port, 
      sigMatrix_0_80_port, sigMatrix_0_79_port, sigMatrix_0_78_port, 
      sigMatrix_0_77_port, sigMatrix_0_76_port, sigMatrix_0_75_port, 
      sigMatrix_0_74_port, sigMatrix_0_73_port, sigMatrix_0_72_port, 
      sigMatrix_0_71_port, sigMatrix_0_70_port, sigMatrix_0_69_port, 
      sigMatrix_0_68_port, sigMatrix_0_67_port, sigMatrix_0_66_port, 
      sigMatrix_0_65_port, sigMatrix_0_63_port, sigMatrix_0_62_port, 
      sigMatrix_0_61_port, sigMatrix_0_60_port, sigMatrix_0_59_port, 
      sigMatrix_0_58_port, sigMatrix_0_57_port, sigMatrix_0_56_port, 
      sigMatrix_0_55_port, sigMatrix_0_54_port, sigMatrix_0_53_port, 
      sigMatrix_0_52_port, sigMatrix_0_51_port, sigMatrix_0_50_port, 
      sigMatrix_0_49_port, sigMatrix_0_48_port, sigMatrix_0_47_port, 
      sigMatrix_0_46_port, sigMatrix_0_45_port, sigMatrix_0_44_port, 
      sigMatrix_0_43_port, sigMatrix_0_42_port, sigMatrix_0_41_port, 
      sigMatrix_0_40_port, sigMatrix_0_39_port, sigMatrix_0_38_port, 
      sigMatrix_0_37_port, sigMatrix_0_36_port, sigMatrix_0_35_port, 
      sigMatrix_0_34_port, sigMatrix_0_33_port, sigMatrix_0_32_port, 
      sigMatrix_0_31_port, sigMatrix_0_30_port, sigMatrix_0_29_port, 
      sigMatrix_0_28_port, sigMatrix_0_27_port, sigMatrix_0_26_port, 
      sigMatrix_0_25_port, sigMatrix_0_24_port, sigMatrix_0_23_port, 
      sigMatrix_0_22_port, sigMatrix_0_21_port, sigMatrix_0_20_port, 
      sigMatrix_0_19_port, sigMatrix_0_18_port, sigMatrix_0_17_port, 
      sigMatrix_0_16_port, sigMatrix_0_15_port, sigMatrix_0_14_port, 
      sigMatrix_0_13_port, sigMatrix_0_12_port, sigMatrix_0_11_port, 
      sigMatrix_0_10_port, sigMatrix_0_9_port, sigMatrix_0_8_port, 
      sigMatrix_0_7_port, sigMatrix_0_6_port, sigMatrix_0_5_port, 
      sigMatrix_0_4_port, sigMatrix_0_3_port, sigMatrix_0_2_port, 
      sigMatrix_0_1_port, sigMatrix_0_0_port, sigMatrix_1_127_port, 
      sigMatrix_1_126_port, sigMatrix_1_125_port, sigMatrix_1_124_port, 
      sigMatrix_1_123_port, sigMatrix_1_122_port, sigMatrix_1_121_port, 
      sigMatrix_1_120_port, sigMatrix_1_119_port, sigMatrix_1_118_port, 
      sigMatrix_1_117_port, sigMatrix_1_116_port, sigMatrix_1_115_port, 
      sigMatrix_1_114_port, sigMatrix_1_113_port, sigMatrix_1_112_port, 
      sigMatrix_1_111_port, sigMatrix_1_110_port, sigMatrix_1_109_port, 
      sigMatrix_1_108_port, sigMatrix_1_107_port, sigMatrix_1_106_port, 
      sigMatrix_1_105_port, sigMatrix_1_104_port, sigMatrix_1_103_port, 
      sigMatrix_1_102_port, sigMatrix_1_101_port, sigMatrix_1_100_port, 
      sigMatrix_1_99_port, sigMatrix_1_98_port, sigMatrix_1_97_port, 
      sigMatrix_1_96_port, sigMatrix_1_95_port, sigMatrix_1_94_port, 
      sigMatrix_1_93_port, sigMatrix_1_92_port, sigMatrix_1_91_port, 
      sigMatrix_1_90_port, sigMatrix_1_89_port, sigMatrix_1_88_port, 
      sigMatrix_1_87_port, sigMatrix_1_86_port, sigMatrix_1_85_port, 
      sigMatrix_1_84_port, sigMatrix_1_83_port, sigMatrix_1_82_port, 
      sigMatrix_1_81_port, sigMatrix_1_80_port, sigMatrix_1_79_port, 
      sigMatrix_1_78_port, sigMatrix_1_77_port, sigMatrix_1_76_port, 
      sigMatrix_1_75_port, sigMatrix_1_74_port, sigMatrix_1_73_port, 
      sigMatrix_1_72_port, sigMatrix_1_71_port, sigMatrix_1_70_port, 
      sigMatrix_1_69_port, sigMatrix_1_68_port, sigMatrix_1_67_port, 
      sigMatrix_1_66_port, sigMatrix_1_65_port, sigMatrix_1_63_port, 
      sigMatrix_1_62_port, sigMatrix_1_61_port, sigMatrix_1_60_port, 
      sigMatrix_1_59_port, sigMatrix_1_58_port, sigMatrix_1_57_port, 
      sigMatrix_1_56_port, sigMatrix_1_55_port, sigMatrix_1_54_port, 
      sigMatrix_1_53_port, sigMatrix_1_52_port, sigMatrix_1_51_port, 
      sigMatrix_1_50_port, sigMatrix_1_49_port, sigMatrix_1_48_port, 
      sigMatrix_1_47_port, sigMatrix_1_46_port, sigMatrix_1_45_port, 
      sigMatrix_1_44_port, sigMatrix_1_43_port, sigMatrix_1_42_port, 
      sigMatrix_1_41_port, sigMatrix_1_40_port, sigMatrix_1_39_port, 
      sigMatrix_1_38_port, sigMatrix_1_37_port, sigMatrix_1_36_port, 
      sigMatrix_1_35_port, sigMatrix_1_34_port, sigMatrix_1_33_port, 
      sigMatrix_1_32_port, sigMatrix_1_31_port, sigMatrix_1_30_port, 
      sigMatrix_1_29_port, sigMatrix_1_28_port, sigMatrix_1_27_port, 
      sigMatrix_1_26_port, sigMatrix_1_25_port, sigMatrix_1_24_port, 
      sigMatrix_1_23_port, sigMatrix_1_22_port, sigMatrix_1_21_port, 
      sigMatrix_1_20_port, sigMatrix_1_19_port, sigMatrix_1_18_port, 
      sigMatrix_1_17_port, sigMatrix_1_16_port, sigMatrix_1_15_port, 
      sigMatrix_1_14_port, sigMatrix_1_13_port, sigMatrix_1_12_port, 
      sigMatrix_1_11_port, sigMatrix_1_10_port, sigMatrix_1_9_port, 
      sigMatrix_1_8_port, sigMatrix_1_7_port, sigMatrix_1_6_port, 
      sigMatrix_1_5_port, sigMatrix_1_4_port, sigMatrix_1_3_port, 
      sigMatrix_1_2_port, sigMatrix_1_1_port, sigMatrix_1_0_port, 
      sigMatrix_2_127_port, sigMatrix_2_126_port, sigMatrix_2_125_port, 
      sigMatrix_2_124_port, sigMatrix_2_123_port, sigMatrix_2_122_port, 
      sigMatrix_2_121_port, sigMatrix_2_120_port, sigMatrix_2_119_port, 
      sigMatrix_2_118_port, sigMatrix_2_117_port, sigMatrix_2_116_port, 
      sigMatrix_2_115_port, sigMatrix_2_114_port, sigMatrix_2_113_port, 
      sigMatrix_2_112_port, sigMatrix_2_111_port, sigMatrix_2_110_port, 
      sigMatrix_2_109_port, sigMatrix_2_108_port, sigMatrix_2_107_port, 
      sigMatrix_2_106_port, sigMatrix_2_105_port, sigMatrix_2_104_port, 
      sigMatrix_2_103_port, sigMatrix_2_102_port, sigMatrix_2_101_port, 
      sigMatrix_2_100_port, sigMatrix_2_99_port, sigMatrix_2_98_port, 
      sigMatrix_2_97_port, sigMatrix_2_96_port, sigMatrix_2_95_port, 
      sigMatrix_2_94_port, sigMatrix_2_93_port, sigMatrix_2_92_port, 
      sigMatrix_2_91_port, sigMatrix_2_90_port, sigMatrix_2_89_port, 
      sigMatrix_2_88_port, sigMatrix_2_87_port, sigMatrix_2_86_port, 
      sigMatrix_2_85_port, sigMatrix_2_84_port, sigMatrix_2_83_port, 
      sigMatrix_2_82_port, sigMatrix_2_81_port, sigMatrix_2_80_port, 
      sigMatrix_2_79_port, sigMatrix_2_78_port, sigMatrix_2_77_port, 
      sigMatrix_2_76_port, sigMatrix_2_75_port, sigMatrix_2_74_port, 
      sigMatrix_2_73_port, sigMatrix_2_72_port, sigMatrix_2_71_port, 
      sigMatrix_2_70_port, sigMatrix_2_69_port, sigMatrix_2_68_port, 
      sigMatrix_2_67_port, sigMatrix_2_66_port, sigMatrix_2_65_port, 
      sigMatrix_2_63_port, sigMatrix_2_62_port, sigMatrix_2_61_port, 
      sigMatrix_2_60_port, sigMatrix_2_59_port, sigMatrix_2_58_port, 
      sigMatrix_2_57_port, sigMatrix_2_56_port, sigMatrix_2_55_port, 
      sigMatrix_2_54_port, sigMatrix_2_53_port, sigMatrix_2_52_port, 
      sigMatrix_2_51_port, sigMatrix_2_50_port, sigMatrix_2_49_port, 
      sigMatrix_2_48_port, sigMatrix_2_47_port, sigMatrix_2_46_port, 
      sigMatrix_2_45_port, sigMatrix_2_44_port, sigMatrix_2_43_port, 
      sigMatrix_2_42_port, sigMatrix_2_41_port, sigMatrix_2_40_port, 
      sigMatrix_2_39_port, sigMatrix_2_38_port, sigMatrix_2_37_port, 
      sigMatrix_2_36_port, sigMatrix_2_35_port, sigMatrix_2_34_port, 
      sigMatrix_2_33_port, sigMatrix_2_32_port, sigMatrix_2_31_port, 
      sigMatrix_2_30_port, sigMatrix_2_29_port, sigMatrix_2_28_port, 
      sigMatrix_2_27_port, sigMatrix_2_26_port, sigMatrix_2_25_port, 
      sigMatrix_2_24_port, sigMatrix_2_23_port, sigMatrix_2_22_port, 
      sigMatrix_2_21_port, sigMatrix_2_20_port, sigMatrix_2_19_port, 
      sigMatrix_2_18_port, sigMatrix_2_17_port, sigMatrix_2_16_port, 
      sigMatrix_2_15_port, sigMatrix_2_14_port, sigMatrix_2_13_port, 
      sigMatrix_2_12_port, sigMatrix_2_11_port, sigMatrix_2_10_port, 
      sigMatrix_2_9_port, sigMatrix_2_8_port, sigMatrix_2_7_port, 
      sigMatrix_2_6_port, sigMatrix_2_5_port, sigMatrix_2_4_port, 
      sigMatrix_2_3_port, sigMatrix_2_2_port, sigMatrix_2_1_port, 
      sigMatrix_2_0_port, sigMatrix_3_127_port, sigMatrix_3_126_port, 
      sigMatrix_3_125_port, sigMatrix_3_124_port, sigMatrix_3_123_port, 
      sigMatrix_3_122_port, sigMatrix_3_121_port, sigMatrix_3_120_port, 
      sigMatrix_3_119_port, sigMatrix_3_118_port, sigMatrix_3_117_port, 
      sigMatrix_3_116_port, sigMatrix_3_115_port, sigMatrix_3_114_port, 
      sigMatrix_3_113_port, sigMatrix_3_112_port, sigMatrix_3_111_port, 
      sigMatrix_3_110_port, sigMatrix_3_109_port, sigMatrix_3_108_port, 
      sigMatrix_3_107_port, sigMatrix_3_106_port, sigMatrix_3_105_port, 
      sigMatrix_3_104_port, sigMatrix_3_103_port, sigMatrix_3_102_port, 
      sigMatrix_3_101_port, sigMatrix_3_100_port, sigMatrix_3_99_port, 
      sigMatrix_3_98_port, sigMatrix_3_97_port, sigMatrix_3_96_port, 
      sigMatrix_3_95_port, sigMatrix_3_94_port, sigMatrix_3_93_port, 
      sigMatrix_3_92_port, sigMatrix_3_91_port, sigMatrix_3_90_port, 
      sigMatrix_3_89_port, sigMatrix_3_88_port, sigMatrix_3_87_port, 
      sigMatrix_3_86_port, sigMatrix_3_85_port, sigMatrix_3_84_port, 
      sigMatrix_3_83_port, sigMatrix_3_82_port, sigMatrix_3_81_port, 
      sigMatrix_3_80_port, sigMatrix_3_79_port, sigMatrix_3_78_port, 
      sigMatrix_3_77_port, sigMatrix_3_76_port, sigMatrix_3_75_port, 
      sigMatrix_3_74_port, sigMatrix_3_73_port, sigMatrix_3_72_port, 
      sigMatrix_3_71_port, sigMatrix_3_70_port, sigMatrix_3_69_port, 
      sigMatrix_3_68_port, sigMatrix_3_67_port, sigMatrix_3_66_port, 
      sigMatrix_3_65_port, sigMatrix_3_63_port, sigMatrix_3_62_port, 
      sigMatrix_3_61_port, sigMatrix_3_60_port, sigMatrix_3_59_port, 
      sigMatrix_3_58_port, sigMatrix_3_57_port, sigMatrix_3_56_port, 
      sigMatrix_3_55_port, sigMatrix_3_54_port, sigMatrix_3_53_port, 
      sigMatrix_3_52_port, sigMatrix_3_51_port, sigMatrix_3_50_port, 
      sigMatrix_3_49_port, sigMatrix_3_48_port, sigMatrix_3_47_port, 
      sigMatrix_3_46_port, sigMatrix_3_45_port, sigMatrix_3_44_port, 
      sigMatrix_3_43_port, sigMatrix_3_42_port, sigMatrix_3_41_port, 
      sigMatrix_3_40_port, sigMatrix_3_39_port, sigMatrix_3_38_port, 
      sigMatrix_3_37_port, sigMatrix_3_36_port, sigMatrix_3_35_port, 
      sigMatrix_3_34_port, sigMatrix_3_33_port, sigMatrix_3_32_port, 
      sigMatrix_3_31_port, sigMatrix_3_30_port, sigMatrix_3_29_port, 
      sigMatrix_3_28_port, sigMatrix_3_27_port, sigMatrix_3_26_port, 
      sigMatrix_3_25_port, sigMatrix_3_24_port, sigMatrix_3_23_port, 
      sigMatrix_3_22_port, sigMatrix_3_21_port, sigMatrix_3_20_port, 
      sigMatrix_3_19_port, sigMatrix_3_18_port, sigMatrix_3_17_port, 
      sigMatrix_3_16_port, sigMatrix_3_15_port, sigMatrix_3_14_port, 
      sigMatrix_3_13_port, sigMatrix_3_12_port, sigMatrix_3_11_port, 
      sigMatrix_3_10_port, sigMatrix_3_9_port, sigMatrix_3_8_port, 
      sigMatrix_3_7_port, sigMatrix_3_6_port, sigMatrix_3_5_port, 
      sigMatrix_3_4_port, sigMatrix_3_3_port, sigMatrix_3_2_port, 
      sigMatrix_3_1_port, sigMatrix_3_0_port, sigMatrix_4_127_port, 
      sigMatrix_4_126_port, sigMatrix_4_125_port, sigMatrix_4_124_port, 
      sigMatrix_4_123_port, sigMatrix_4_122_port, sigMatrix_4_121_port, 
      sigMatrix_4_120_port, sigMatrix_4_119_port, sigMatrix_4_118_port, 
      sigMatrix_4_117_port, sigMatrix_4_116_port, sigMatrix_4_115_port, 
      sigMatrix_4_114_port, sigMatrix_4_113_port, sigMatrix_4_112_port, 
      sigMatrix_4_111_port, sigMatrix_4_110_port, sigMatrix_4_109_port, 
      sigMatrix_4_108_port, sigMatrix_4_107_port, sigMatrix_4_106_port, 
      sigMatrix_4_105_port, sigMatrix_4_104_port, sigMatrix_4_103_port, 
      sigMatrix_4_102_port, sigMatrix_4_101_port, sigMatrix_4_100_port, 
      sigMatrix_4_99_port, sigMatrix_4_98_port, sigMatrix_4_97_port, 
      sigMatrix_4_96_port, sigMatrix_4_95_port, sigMatrix_4_94_port, 
      sigMatrix_4_93_port, sigMatrix_4_92_port, sigMatrix_4_91_port, 
      sigMatrix_4_90_port, sigMatrix_4_89_port, sigMatrix_4_88_port, 
      sigMatrix_4_87_port, sigMatrix_4_86_port, sigMatrix_4_85_port, 
      sigMatrix_4_84_port, sigMatrix_4_83_port, sigMatrix_4_82_port, 
      sigMatrix_4_81_port, sigMatrix_4_80_port, sigMatrix_4_79_port, 
      sigMatrix_4_78_port, sigMatrix_4_77_port, sigMatrix_4_76_port, 
      sigMatrix_4_75_port, sigMatrix_4_74_port, sigMatrix_4_73_port, 
      sigMatrix_4_72_port, sigMatrix_4_71_port, sigMatrix_4_70_port, 
      sigMatrix_4_69_port, sigMatrix_4_68_port, sigMatrix_4_67_port, 
      sigMatrix_4_66_port, sigMatrix_4_65_port, sigMatrix_4_63_port, 
      sigMatrix_4_62_port, sigMatrix_4_61_port, sigMatrix_4_60_port, 
      sigMatrix_4_59_port, sigMatrix_4_58_port, sigMatrix_4_57_port, 
      sigMatrix_4_56_port, sigMatrix_4_55_port, sigMatrix_4_54_port, 
      sigMatrix_4_53_port, sigMatrix_4_52_port, sigMatrix_4_51_port, 
      sigMatrix_4_50_port, sigMatrix_4_49_port, sigMatrix_4_48_port, 
      sigMatrix_4_47_port, sigMatrix_4_46_port, sigMatrix_4_45_port, 
      sigMatrix_4_44_port, sigMatrix_4_43_port, sigMatrix_4_42_port, 
      sigMatrix_4_41_port, sigMatrix_4_40_port, sigMatrix_4_39_port, 
      sigMatrix_4_38_port, sigMatrix_4_37_port, sigMatrix_4_36_port, 
      sigMatrix_4_35_port, sigMatrix_4_34_port, sigMatrix_4_33_port, 
      sigMatrix_4_32_port, sigMatrix_4_31_port, sigMatrix_4_30_port, 
      sigMatrix_4_29_port, sigMatrix_4_28_port, sigMatrix_4_27_port, 
      sigMatrix_4_26_port, sigMatrix_4_25_port, sigMatrix_4_24_port, 
      sigMatrix_4_23_port, sigMatrix_4_22_port, sigMatrix_4_21_port, 
      sigMatrix_4_20_port, sigMatrix_4_19_port, sigMatrix_4_18_port, 
      sigMatrix_4_17_port, sigMatrix_4_16_port, sigMatrix_4_15_port, 
      sigMatrix_4_14_port, sigMatrix_4_13_port, sigMatrix_4_12_port, 
      sigMatrix_4_11_port, sigMatrix_4_10_port, sigMatrix_4_9_port, 
      sigMatrix_4_8_port, sigMatrix_4_7_port, sigMatrix_4_6_port, 
      sigMatrix_4_5_port, sigMatrix_4_4_port, sigMatrix_4_3_port, 
      sigMatrix_4_2_port, sigMatrix_4_1_port, sigMatrix_4_0_port, 
      sigMatrix_5_127_port, sigMatrix_5_126_port, sigMatrix_5_125_port, 
      sigMatrix_5_124_port, sigMatrix_5_123_port, sigMatrix_5_122_port, 
      sigMatrix_5_121_port, sigMatrix_5_120_port, sigMatrix_5_119_port, 
      sigMatrix_5_118_port, sigMatrix_5_117_port, sigMatrix_5_116_port, 
      sigMatrix_5_115_port, sigMatrix_5_114_port, sigMatrix_5_113_port, 
      sigMatrix_5_112_port, sigMatrix_5_111_port, sigMatrix_5_110_port, 
      sigMatrix_5_109_port, sigMatrix_5_108_port, sigMatrix_5_107_port, 
      sigMatrix_5_106_port, sigMatrix_5_105_port, sigMatrix_5_104_port, 
      sigMatrix_5_103_port, sigMatrix_5_102_port, sigMatrix_5_101_port, 
      sigMatrix_5_100_port, sigMatrix_5_99_port, sigMatrix_5_98_port, 
      sigMatrix_5_97_port, sigMatrix_5_96_port, sigMatrix_5_95_port, 
      sigMatrix_5_94_port, sigMatrix_5_93_port, sigMatrix_5_92_port, 
      sigMatrix_5_91_port, sigMatrix_5_90_port, sigMatrix_5_89_port, 
      sigMatrix_5_88_port, sigMatrix_5_87_port, sigMatrix_5_86_port, 
      sigMatrix_5_85_port, sigMatrix_5_84_port, sigMatrix_5_83_port, 
      sigMatrix_5_82_port, sigMatrix_5_81_port, sigMatrix_5_80_port, 
      sigMatrix_5_79_port, sigMatrix_5_78_port, sigMatrix_5_77_port, 
      sigMatrix_5_76_port, sigMatrix_5_75_port, sigMatrix_5_74_port, 
      sigMatrix_5_73_port, sigMatrix_5_72_port, sigMatrix_5_71_port, 
      sigMatrix_5_70_port, sigMatrix_5_69_port, sigMatrix_5_68_port, 
      sigMatrix_5_67_port, sigMatrix_5_66_port, sigMatrix_5_65_port, 
      sigMatrix_5_63_port, sigMatrix_5_62_port, sigMatrix_5_61_port, 
      sigMatrix_5_60_port, sigMatrix_5_59_port, sigMatrix_5_58_port, 
      sigMatrix_5_57_port, sigMatrix_5_56_port, sigMatrix_5_55_port, 
      sigMatrix_5_54_port, sigMatrix_5_53_port, sigMatrix_5_52_port, 
      sigMatrix_5_51_port, sigMatrix_5_50_port, sigMatrix_5_49_port, 
      sigMatrix_5_48_port, sigMatrix_5_47_port, sigMatrix_5_46_port, 
      sigMatrix_5_45_port, sigMatrix_5_44_port, sigMatrix_5_43_port, 
      sigMatrix_5_42_port, sigMatrix_5_41_port, sigMatrix_5_40_port, 
      sigMatrix_5_39_port, sigMatrix_5_38_port, sigMatrix_5_37_port, 
      sigMatrix_5_36_port, sigMatrix_5_35_port, sigMatrix_5_34_port, 
      sigMatrix_5_33_port, sigMatrix_5_32_port, sigMatrix_5_31_port, 
      sigMatrix_5_30_port, sigMatrix_5_29_port, sigMatrix_5_28_port, 
      sigMatrix_5_27_port, sigMatrix_5_26_port, sigMatrix_5_25_port, 
      sigMatrix_5_24_port, sigMatrix_5_23_port, sigMatrix_5_22_port, 
      sigMatrix_5_21_port, sigMatrix_5_20_port, sigMatrix_5_19_port, 
      sigMatrix_5_18_port, sigMatrix_5_17_port, sigMatrix_5_16_port, 
      sigMatrix_5_15_port, sigMatrix_5_14_port, sigMatrix_5_13_port, 
      sigMatrix_5_12_port, sigMatrix_5_11_port, sigMatrix_5_10_port, 
      sigMatrix_5_9_port, sigMatrix_5_8_port, sigMatrix_5_7_port, 
      sigMatrix_5_6_port, sigMatrix_5_5_port, sigMatrix_5_4_port, 
      sigMatrix_5_3_port, sigMatrix_5_2_port, sigMatrix_5_1_port, 
      sigMatrix_5_0_port, sigMatrix_6_127_port, sigMatrix_6_126_port, 
      sigMatrix_6_125_port, sigMatrix_6_124_port, sigMatrix_6_123_port, 
      sigMatrix_6_122_port, sigMatrix_6_121_port, sigMatrix_6_120_port, 
      sigMatrix_6_119_port, sigMatrix_6_118_port, sigMatrix_6_117_port, 
      sigMatrix_6_116_port, sigMatrix_6_115_port, sigMatrix_6_114_port, 
      sigMatrix_6_113_port, sigMatrix_6_112_port, sigMatrix_6_111_port, 
      sigMatrix_6_110_port, sigMatrix_6_109_port, sigMatrix_6_108_port, 
      sigMatrix_6_107_port, sigMatrix_6_106_port, sigMatrix_6_105_port, 
      sigMatrix_6_104_port, sigMatrix_6_103_port, sigMatrix_6_102_port, 
      sigMatrix_6_101_port, sigMatrix_6_100_port, sigMatrix_6_99_port, 
      sigMatrix_6_98_port, sigMatrix_6_97_port, sigMatrix_6_96_port, 
      sigMatrix_6_95_port, sigMatrix_6_94_port, sigMatrix_6_93_port, 
      sigMatrix_6_92_port, sigMatrix_6_91_port, sigMatrix_6_90_port, 
      sigMatrix_6_89_port, sigMatrix_6_88_port, sigMatrix_6_87_port, 
      sigMatrix_6_86_port, sigMatrix_6_85_port, sigMatrix_6_84_port, 
      sigMatrix_6_83_port, sigMatrix_6_82_port, sigMatrix_6_81_port, 
      sigMatrix_6_80_port, sigMatrix_6_79_port, sigMatrix_6_78_port, 
      sigMatrix_6_77_port, sigMatrix_6_76_port, sigMatrix_6_75_port, 
      sigMatrix_6_74_port, sigMatrix_6_73_port, sigMatrix_6_72_port, 
      sigMatrix_6_71_port, sigMatrix_6_70_port, sigMatrix_6_69_port, 
      sigMatrix_6_68_port, sigMatrix_6_67_port, sigMatrix_6_66_port, 
      sigMatrix_6_65_port, sigMatrix_6_63_port, sigMatrix_6_62_port, 
      sigMatrix_6_61_port, sigMatrix_6_60_port, sigMatrix_6_59_port, 
      sigMatrix_6_58_port, sigMatrix_6_57_port, sigMatrix_6_56_port, 
      sigMatrix_6_55_port, sigMatrix_6_54_port, sigMatrix_6_53_port, 
      sigMatrix_6_52_port, sigMatrix_6_51_port, sigMatrix_6_50_port, 
      sigMatrix_6_49_port, sigMatrix_6_48_port, sigMatrix_6_47_port, 
      sigMatrix_6_46_port, sigMatrix_6_45_port, sigMatrix_6_44_port, 
      sigMatrix_6_43_port, sigMatrix_6_42_port, sigMatrix_6_41_port, 
      sigMatrix_6_40_port, sigMatrix_6_39_port, sigMatrix_6_38_port, 
      sigMatrix_6_37_port, sigMatrix_6_36_port, sigMatrix_6_35_port, 
      sigMatrix_6_34_port, sigMatrix_6_33_port, sigMatrix_6_32_port, 
      sigMatrix_6_31_port, sigMatrix_6_30_port, sigMatrix_6_29_port, 
      sigMatrix_6_28_port, sigMatrix_6_27_port, sigMatrix_6_26_port, 
      sigMatrix_6_25_port, sigMatrix_6_24_port, sigMatrix_6_23_port, 
      sigMatrix_6_22_port, sigMatrix_6_21_port, sigMatrix_6_20_port, 
      sigMatrix_6_19_port, sigMatrix_6_18_port, sigMatrix_6_17_port, 
      sigMatrix_6_16_port, sigMatrix_6_15_port, sigMatrix_6_14_port, 
      sigMatrix_6_13_port, sigMatrix_6_12_port, sigMatrix_6_11_port, 
      sigMatrix_6_10_port, sigMatrix_6_9_port, sigMatrix_6_8_port, 
      sigMatrix_6_7_port, sigMatrix_6_6_port, sigMatrix_6_5_port, 
      sigMatrix_6_4_port, sigMatrix_6_3_port, sigMatrix_6_2_port, 
      sigMatrix_6_1_port, sigMatrix_6_0_port, sigMatrix_7_127_port, 
      sigMatrix_7_126_port, sigMatrix_7_125_port, sigMatrix_7_124_port, 
      sigMatrix_7_123_port, sigMatrix_7_122_port, sigMatrix_7_121_port, 
      sigMatrix_7_120_port, sigMatrix_7_119_port, sigMatrix_7_118_port, 
      sigMatrix_7_117_port, sigMatrix_7_116_port, sigMatrix_7_115_port, 
      sigMatrix_7_114_port, sigMatrix_7_113_port, sigMatrix_7_112_port, 
      sigMatrix_7_111_port, sigMatrix_7_110_port, sigMatrix_7_109_port, 
      sigMatrix_7_108_port, sigMatrix_7_107_port, sigMatrix_7_106_port, 
      sigMatrix_7_105_port, sigMatrix_7_104_port, sigMatrix_7_103_port, 
      sigMatrix_7_102_port, sigMatrix_7_101_port, sigMatrix_7_100_port, 
      sigMatrix_7_99_port, sigMatrix_7_98_port, sigMatrix_7_97_port, 
      sigMatrix_7_96_port, sigMatrix_7_95_port, sigMatrix_7_94_port, 
      sigMatrix_7_93_port, sigMatrix_7_92_port, sigMatrix_7_91_port, 
      sigMatrix_7_90_port, sigMatrix_7_89_port, sigMatrix_7_88_port, 
      sigMatrix_7_87_port, sigMatrix_7_86_port, sigMatrix_7_85_port, 
      sigMatrix_7_84_port, sigMatrix_7_83_port, sigMatrix_7_82_port, 
      sigMatrix_7_81_port, sigMatrix_7_80_port, sigMatrix_7_79_port, 
      sigMatrix_7_78_port, sigMatrix_7_77_port, sigMatrix_7_76_port, 
      sigMatrix_7_75_port, sigMatrix_7_74_port, sigMatrix_7_73_port, 
      sigMatrix_7_72_port, sigMatrix_7_71_port, sigMatrix_7_70_port, 
      sigMatrix_7_69_port, sigMatrix_7_68_port, sigMatrix_7_67_port, 
      sigMatrix_7_66_port, sigMatrix_7_65_port, sigMatrix_7_63_port, 
      sigMatrix_7_62_port, sigMatrix_7_61_port, sigMatrix_7_60_port, 
      sigMatrix_7_59_port, sigMatrix_7_58_port, sigMatrix_7_57_port, 
      sigMatrix_7_56_port, sigMatrix_7_55_port, sigMatrix_7_54_port, 
      sigMatrix_7_53_port, sigMatrix_7_52_port, sigMatrix_7_51_port, 
      sigMatrix_7_50_port, sigMatrix_7_49_port, sigMatrix_7_48_port, 
      sigMatrix_7_47_port, sigMatrix_7_46_port, sigMatrix_7_45_port, 
      sigMatrix_7_44_port, sigMatrix_7_43_port, sigMatrix_7_42_port, 
      sigMatrix_7_41_port, sigMatrix_7_40_port, sigMatrix_7_39_port, 
      sigMatrix_7_38_port, sigMatrix_7_37_port, sigMatrix_7_36_port, 
      sigMatrix_7_35_port, sigMatrix_7_34_port, sigMatrix_7_33_port, 
      sigMatrix_7_32_port, sigMatrix_7_31_port, sigMatrix_7_30_port, 
      sigMatrix_7_29_port, sigMatrix_7_28_port, sigMatrix_7_27_port, 
      sigMatrix_7_26_port, sigMatrix_7_25_port, sigMatrix_7_24_port, 
      sigMatrix_7_23_port, sigMatrix_7_22_port, sigMatrix_7_21_port, 
      sigMatrix_7_20_port, sigMatrix_7_19_port, sigMatrix_7_18_port, 
      sigMatrix_7_17_port, sigMatrix_7_16_port, sigMatrix_7_15_port, 
      sigMatrix_7_14_port, sigMatrix_7_13_port, sigMatrix_7_12_port, 
      sigMatrix_7_11_port, sigMatrix_7_10_port, sigMatrix_7_9_port, 
      sigMatrix_7_8_port, sigMatrix_7_7_port, sigMatrix_7_6_port, 
      sigMatrix_7_5_port, sigMatrix_7_4_port, sigMatrix_7_3_port, 
      sigMatrix_7_2_port, sigMatrix_7_1_port, sigMatrix_7_0_port, 
      sigMatrix_8_127_port, sigMatrix_8_126_port, sigMatrix_8_125_port, 
      sigMatrix_8_124_port, sigMatrix_8_123_port, sigMatrix_8_122_port, 
      sigMatrix_8_121_port, sigMatrix_8_120_port, sigMatrix_8_119_port, 
      sigMatrix_8_118_port, sigMatrix_8_117_port, sigMatrix_8_116_port, 
      sigMatrix_8_115_port, sigMatrix_8_114_port, sigMatrix_8_113_port, 
      sigMatrix_8_112_port, sigMatrix_8_111_port, sigMatrix_8_110_port, 
      sigMatrix_8_109_port, sigMatrix_8_108_port, sigMatrix_8_107_port, 
      sigMatrix_8_106_port, sigMatrix_8_105_port, sigMatrix_8_104_port, 
      sigMatrix_8_103_port, sigMatrix_8_102_port, sigMatrix_8_101_port, 
      sigMatrix_8_100_port, sigMatrix_8_99_port, sigMatrix_8_98_port, 
      sigMatrix_8_97_port, sigMatrix_8_96_port, sigMatrix_8_95_port, 
      sigMatrix_8_94_port, sigMatrix_8_93_port, sigMatrix_8_92_port, 
      sigMatrix_8_91_port, sigMatrix_8_90_port, sigMatrix_8_89_port, 
      sigMatrix_8_88_port, sigMatrix_8_87_port, sigMatrix_8_86_port, 
      sigMatrix_8_85_port, sigMatrix_8_84_port, sigMatrix_8_83_port, 
      sigMatrix_8_82_port, sigMatrix_8_81_port, sigMatrix_8_80_port, 
      sigMatrix_8_79_port, sigMatrix_8_78_port, sigMatrix_8_77_port, 
      sigMatrix_8_76_port, sigMatrix_8_75_port, sigMatrix_8_74_port, 
      sigMatrix_8_73_port, sigMatrix_8_72_port, sigMatrix_8_71_port, 
      sigMatrix_8_70_port, sigMatrix_8_69_port, sigMatrix_8_68_port, 
      sigMatrix_8_67_port, sigMatrix_8_66_port, sigMatrix_8_65_port, 
      sigMatrix_8_63_port, sigMatrix_8_62_port, sigMatrix_8_61_port, 
      sigMatrix_8_60_port, sigMatrix_8_59_port, sigMatrix_8_58_port, 
      sigMatrix_8_57_port, sigMatrix_8_56_port, sigMatrix_8_55_port, 
      sigMatrix_8_54_port, sigMatrix_8_53_port, sigMatrix_8_52_port, 
      sigMatrix_8_51_port, sigMatrix_8_50_port, sigMatrix_8_49_port, 
      sigMatrix_8_48_port, sigMatrix_8_47_port, sigMatrix_8_46_port, 
      sigMatrix_8_45_port, sigMatrix_8_44_port, sigMatrix_8_43_port, 
      sigMatrix_8_42_port, sigMatrix_8_41_port, sigMatrix_8_40_port, 
      sigMatrix_8_39_port, sigMatrix_8_38_port, sigMatrix_8_37_port, 
      sigMatrix_8_36_port, sigMatrix_8_35_port, sigMatrix_8_34_port, 
      sigMatrix_8_33_port, sigMatrix_8_32_port, sigMatrix_8_31_port, 
      sigMatrix_8_30_port, sigMatrix_8_29_port, sigMatrix_8_28_port, 
      sigMatrix_8_27_port, sigMatrix_8_26_port, sigMatrix_8_25_port, 
      sigMatrix_8_24_port, sigMatrix_8_23_port, sigMatrix_8_22_port, 
      sigMatrix_8_21_port, sigMatrix_8_20_port, sigMatrix_8_19_port, 
      sigMatrix_8_18_port, sigMatrix_8_17_port, sigMatrix_8_16_port, 
      sigMatrix_8_15_port, sigMatrix_8_14_port, sigMatrix_8_13_port, 
      sigMatrix_8_12_port, sigMatrix_8_11_port, sigMatrix_8_10_port, 
      sigMatrix_8_9_port, sigMatrix_8_8_port, sigMatrix_8_7_port, 
      sigMatrix_8_6_port, sigMatrix_8_5_port, sigMatrix_8_4_port, 
      sigMatrix_8_3_port, sigMatrix_8_2_port, sigMatrix_8_1_port, 
      sigMatrix_8_0_port, sigMatrix_9_127_port, sigMatrix_9_126_port, 
      sigMatrix_9_125_port, sigMatrix_9_124_port, sigMatrix_9_123_port, 
      sigMatrix_9_122_port, sigMatrix_9_121_port, sigMatrix_9_120_port, 
      sigMatrix_9_119_port, sigMatrix_9_118_port, sigMatrix_9_117_port, 
      sigMatrix_9_116_port, sigMatrix_9_115_port, sigMatrix_9_114_port, 
      sigMatrix_9_113_port, sigMatrix_9_112_port, sigMatrix_9_111_port, 
      sigMatrix_9_110_port, sigMatrix_9_109_port, sigMatrix_9_108_port, 
      sigMatrix_9_107_port, sigMatrix_9_106_port, sigMatrix_9_105_port, 
      sigMatrix_9_104_port, sigMatrix_9_103_port, sigMatrix_9_102_port, 
      sigMatrix_9_101_port, sigMatrix_9_100_port, sigMatrix_9_99_port, 
      sigMatrix_9_98_port, sigMatrix_9_97_port, sigMatrix_9_96_port, 
      sigMatrix_9_95_port, sigMatrix_9_94_port, sigMatrix_9_93_port, 
      sigMatrix_9_92_port, sigMatrix_9_91_port, sigMatrix_9_90_port, 
      sigMatrix_9_89_port, sigMatrix_9_88_port, sigMatrix_9_87_port, 
      sigMatrix_9_86_port, sigMatrix_9_85_port, sigMatrix_9_84_port, 
      sigMatrix_9_83_port, sigMatrix_9_82_port, sigMatrix_9_81_port, 
      sigMatrix_9_80_port, sigMatrix_9_79_port, sigMatrix_9_78_port, 
      sigMatrix_9_77_port, sigMatrix_9_76_port, sigMatrix_9_75_port, 
      sigMatrix_9_74_port, sigMatrix_9_73_port, sigMatrix_9_72_port, 
      sigMatrix_9_71_port, sigMatrix_9_70_port, sigMatrix_9_69_port, 
      sigMatrix_9_68_port, sigMatrix_9_67_port, sigMatrix_9_66_port, 
      sigMatrix_9_65_port, sigMatrix_9_63_port, sigMatrix_9_62_port, 
      sigMatrix_9_61_port, sigMatrix_9_60_port, sigMatrix_9_59_port, 
      sigMatrix_9_58_port, sigMatrix_9_57_port, sigMatrix_9_56_port, 
      sigMatrix_9_55_port, sigMatrix_9_54_port, sigMatrix_9_53_port, 
      sigMatrix_9_52_port, sigMatrix_9_51_port, sigMatrix_9_50_port, 
      sigMatrix_9_49_port, sigMatrix_9_48_port, sigMatrix_9_47_port, 
      sigMatrix_9_46_port, sigMatrix_9_45_port, sigMatrix_9_44_port, 
      sigMatrix_9_43_port, sigMatrix_9_42_port, sigMatrix_9_41_port, 
      sigMatrix_9_40_port, sigMatrix_9_39_port, sigMatrix_9_38_port, 
      sigMatrix_9_37_port, sigMatrix_9_36_port, sigMatrix_9_35_port, 
      sigMatrix_9_34_port, sigMatrix_9_33_port, sigMatrix_9_32_port, 
      sigMatrix_9_31_port, sigMatrix_9_30_port, sigMatrix_9_29_port, 
      sigMatrix_9_28_port, sigMatrix_9_27_port, sigMatrix_9_26_port, 
      sigMatrix_9_25_port, sigMatrix_9_24_port, sigMatrix_9_23_port, 
      sigMatrix_9_22_port, sigMatrix_9_21_port, sigMatrix_9_20_port, 
      sigMatrix_9_19_port, sigMatrix_9_18_port, sigMatrix_9_17_port, 
      sigMatrix_9_16_port, sigMatrix_9_15_port, sigMatrix_9_14_port, 
      sigMatrix_9_13_port, sigMatrix_9_12_port, sigMatrix_9_11_port, 
      sigMatrix_9_10_port, sigMatrix_9_9_port, sigMatrix_9_8_port, 
      sigMatrix_9_7_port, sigMatrix_9_6_port, sigMatrix_9_5_port, 
      sigMatrix_9_4_port, sigMatrix_9_3_port, sigMatrix_9_2_port, 
      sigMatrix_9_1_port, sigMatrix_9_0_port, sigMatrix_10_127_port, 
      sigMatrix_10_126_port, sigMatrix_10_125_port, sigMatrix_10_124_port, 
      sigMatrix_10_123_port, sigMatrix_10_122_port, sigMatrix_10_121_port, 
      sigMatrix_10_120_port, sigMatrix_10_119_port, sigMatrix_10_118_port, 
      sigMatrix_10_117_port, sigMatrix_10_116_port, sigMatrix_10_115_port, 
      sigMatrix_10_114_port, sigMatrix_10_113_port, sigMatrix_10_112_port, 
      sigMatrix_10_111_port, sigMatrix_10_110_port, sigMatrix_10_109_port, 
      sigMatrix_10_108_port, sigMatrix_10_107_port, sigMatrix_10_106_port, 
      sigMatrix_10_105_port, sigMatrix_10_104_port, sigMatrix_10_103_port, 
      sigMatrix_10_102_port, sigMatrix_10_101_port, sigMatrix_10_100_port, 
      sigMatrix_10_99_port, sigMatrix_10_98_port, sigMatrix_10_97_port, 
      sigMatrix_10_96_port, sigMatrix_10_95_port, sigMatrix_10_94_port, 
      sigMatrix_10_93_port, sigMatrix_10_92_port, sigMatrix_10_91_port, 
      sigMatrix_10_90_port, sigMatrix_10_89_port, sigMatrix_10_88_port, 
      sigMatrix_10_87_port, sigMatrix_10_86_port, sigMatrix_10_85_port, 
      sigMatrix_10_84_port, sigMatrix_10_83_port, sigMatrix_10_82_port, 
      sigMatrix_10_81_port, sigMatrix_10_80_port, sigMatrix_10_79_port, 
      sigMatrix_10_78_port, sigMatrix_10_77_port, sigMatrix_10_76_port, 
      sigMatrix_10_75_port, sigMatrix_10_74_port, sigMatrix_10_73_port, 
      sigMatrix_10_72_port, sigMatrix_10_71_port, sigMatrix_10_70_port, 
      sigMatrix_10_69_port, sigMatrix_10_68_port, sigMatrix_10_67_port, 
      sigMatrix_10_66_port, sigMatrix_10_65_port, sigMatrix_10_63_port, 
      sigMatrix_10_62_port, sigMatrix_10_61_port, sigMatrix_10_60_port, 
      sigMatrix_10_59_port, sigMatrix_10_58_port, sigMatrix_10_57_port, 
      sigMatrix_10_56_port, sigMatrix_10_55_port, sigMatrix_10_54_port, 
      sigMatrix_10_53_port, sigMatrix_10_52_port, sigMatrix_10_51_port, 
      sigMatrix_10_50_port, sigMatrix_10_49_port, sigMatrix_10_48_port, 
      sigMatrix_10_47_port, sigMatrix_10_46_port, sigMatrix_10_45_port, 
      sigMatrix_10_44_port, sigMatrix_10_43_port, sigMatrix_10_42_port, 
      sigMatrix_10_41_port, sigMatrix_10_40_port, sigMatrix_10_39_port, 
      sigMatrix_10_38_port, sigMatrix_10_37_port, sigMatrix_10_36_port, 
      sigMatrix_10_35_port, sigMatrix_10_34_port, sigMatrix_10_33_port, 
      sigMatrix_10_32_port, sigMatrix_10_31_port, sigMatrix_10_30_port, 
      sigMatrix_10_29_port, sigMatrix_10_28_port, sigMatrix_10_27_port, 
      sigMatrix_10_26_port, sigMatrix_10_25_port, sigMatrix_10_24_port, 
      sigMatrix_10_23_port, sigMatrix_10_22_port, sigMatrix_10_21_port, 
      sigMatrix_10_20_port, sigMatrix_10_19_port, sigMatrix_10_18_port, 
      sigMatrix_10_17_port, sigMatrix_10_16_port, sigMatrix_10_15_port, 
      sigMatrix_10_14_port, sigMatrix_10_13_port, sigMatrix_10_12_port, 
      sigMatrix_10_11_port, sigMatrix_10_10_port, sigMatrix_10_9_port, 
      sigMatrix_10_8_port, sigMatrix_10_7_port, sigMatrix_10_6_port, 
      sigMatrix_10_5_port, sigMatrix_10_4_port, sigMatrix_10_3_port, 
      sigMatrix_10_2_port, sigMatrix_10_1_port, sigMatrix_10_0_port, 
      sigMatrix_11_127_port, sigMatrix_11_126_port, sigMatrix_11_125_port, 
      sigMatrix_11_124_port, sigMatrix_11_123_port, sigMatrix_11_122_port, 
      sigMatrix_11_121_port, sigMatrix_11_120_port, sigMatrix_11_119_port, 
      sigMatrix_11_118_port, sigMatrix_11_117_port, sigMatrix_11_116_port, 
      sigMatrix_11_115_port, sigMatrix_11_114_port, sigMatrix_11_113_port, 
      sigMatrix_11_112_port, sigMatrix_11_111_port, sigMatrix_11_110_port, 
      sigMatrix_11_109_port, sigMatrix_11_108_port, sigMatrix_11_107_port, 
      sigMatrix_11_106_port, sigMatrix_11_105_port, sigMatrix_11_104_port, 
      sigMatrix_11_103_port, sigMatrix_11_102_port, sigMatrix_11_101_port, 
      sigMatrix_11_100_port, sigMatrix_11_99_port, sigMatrix_11_98_port, 
      sigMatrix_11_97_port, sigMatrix_11_96_port, sigMatrix_11_95_port, 
      sigMatrix_11_94_port, sigMatrix_11_93_port, sigMatrix_11_92_port, 
      sigMatrix_11_91_port, sigMatrix_11_90_port, sigMatrix_11_89_port, 
      sigMatrix_11_88_port, sigMatrix_11_87_port, sigMatrix_11_86_port, 
      sigMatrix_11_85_port, sigMatrix_11_84_port, sigMatrix_11_83_port, 
      sigMatrix_11_82_port, sigMatrix_11_81_port, sigMatrix_11_80_port, 
      sigMatrix_11_79_port, sigMatrix_11_78_port, sigMatrix_11_77_port, 
      sigMatrix_11_76_port, sigMatrix_11_75_port, sigMatrix_11_74_port, 
      sigMatrix_11_73_port, sigMatrix_11_72_port, sigMatrix_11_71_port, 
      sigMatrix_11_70_port, sigMatrix_11_69_port, sigMatrix_11_68_port, 
      sigMatrix_11_67_port, sigMatrix_11_66_port, sigMatrix_11_65_port, 
      sigMatrix_11_63_port, sigMatrix_11_62_port, sigMatrix_11_61_port, 
      sigMatrix_11_60_port, sigMatrix_11_59_port, sigMatrix_11_58_port, 
      sigMatrix_11_57_port, sigMatrix_11_56_port, sigMatrix_11_55_port, 
      sigMatrix_11_54_port, sigMatrix_11_53_port, sigMatrix_11_52_port, 
      sigMatrix_11_51_port, sigMatrix_11_50_port, sigMatrix_11_49_port, 
      sigMatrix_11_48_port, sigMatrix_11_47_port, sigMatrix_11_46_port, 
      sigMatrix_11_45_port, sigMatrix_11_44_port, sigMatrix_11_43_port, 
      sigMatrix_11_42_port, sigMatrix_11_41_port, sigMatrix_11_40_port, 
      sigMatrix_11_39_port, sigMatrix_11_38_port, sigMatrix_11_37_port, 
      sigMatrix_11_36_port, sigMatrix_11_35_port, sigMatrix_11_34_port, 
      sigMatrix_11_33_port, sigMatrix_11_32_port, sigMatrix_11_31_port, 
      sigMatrix_11_30_port, sigMatrix_11_29_port, sigMatrix_11_28_port, 
      sigMatrix_11_27_port, sigMatrix_11_26_port, sigMatrix_11_25_port, 
      sigMatrix_11_24_port, sigMatrix_11_23_port, sigMatrix_11_22_port, 
      sigMatrix_11_21_port, sigMatrix_11_20_port, sigMatrix_11_19_port, 
      sigMatrix_11_18_port, sigMatrix_11_17_port, sigMatrix_11_16_port, 
      sigMatrix_11_15_port, sigMatrix_11_14_port, sigMatrix_11_13_port, 
      sigMatrix_11_12_port, sigMatrix_11_11_port, sigMatrix_11_10_port, 
      sigMatrix_11_9_port, sigMatrix_11_8_port, sigMatrix_11_7_port, 
      sigMatrix_11_6_port, sigMatrix_11_5_port, sigMatrix_11_4_port, 
      sigMatrix_11_3_port, sigMatrix_11_2_port, sigMatrix_11_1_port, 
      sigMatrix_11_0_port, sigMatrix_12_127_port, sigMatrix_12_126_port, 
      sigMatrix_12_125_port, sigMatrix_12_124_port, sigMatrix_12_123_port, 
      sigMatrix_12_122_port, sigMatrix_12_121_port, sigMatrix_12_120_port, 
      sigMatrix_12_119_port, sigMatrix_12_118_port, sigMatrix_12_117_port, 
      sigMatrix_12_116_port, sigMatrix_12_115_port, sigMatrix_12_114_port, 
      sigMatrix_12_113_port, sigMatrix_12_112_port, sigMatrix_12_111_port, 
      sigMatrix_12_110_port, sigMatrix_12_109_port, sigMatrix_12_108_port, 
      sigMatrix_12_107_port, sigMatrix_12_106_port, sigMatrix_12_105_port, 
      sigMatrix_12_104_port, sigMatrix_12_103_port, sigMatrix_12_102_port, 
      sigMatrix_12_101_port, sigMatrix_12_100_port, sigMatrix_12_99_port, 
      sigMatrix_12_98_port, sigMatrix_12_97_port, sigMatrix_12_96_port, 
      sigMatrix_12_95_port, sigMatrix_12_94_port, sigMatrix_12_93_port, 
      sigMatrix_12_92_port, sigMatrix_12_91_port, sigMatrix_12_90_port, 
      sigMatrix_12_89_port, sigMatrix_12_88_port, sigMatrix_12_87_port, 
      sigMatrix_12_86_port, sigMatrix_12_85_port, sigMatrix_12_84_port, 
      sigMatrix_12_83_port, sigMatrix_12_82_port, sigMatrix_12_81_port, 
      sigMatrix_12_80_port, sigMatrix_12_79_port, sigMatrix_12_78_port, 
      sigMatrix_12_77_port, sigMatrix_12_76_port, sigMatrix_12_75_port, 
      sigMatrix_12_74_port, sigMatrix_12_73_port, sigMatrix_12_72_port, 
      sigMatrix_12_71_port, sigMatrix_12_70_port, sigMatrix_12_69_port, 
      sigMatrix_12_68_port, sigMatrix_12_67_port, sigMatrix_12_66_port, 
      sigMatrix_12_65_port, sigMatrix_12_63_port, sigMatrix_12_62_port, 
      sigMatrix_12_61_port, sigMatrix_12_60_port, sigMatrix_12_59_port, 
      sigMatrix_12_58_port, sigMatrix_12_57_port, sigMatrix_12_56_port, 
      sigMatrix_12_55_port, sigMatrix_12_54_port, sigMatrix_12_53_port, 
      sigMatrix_12_52_port, sigMatrix_12_51_port, sigMatrix_12_50_port, 
      sigMatrix_12_49_port, sigMatrix_12_48_port, sigMatrix_12_47_port, 
      sigMatrix_12_46_port, sigMatrix_12_45_port, sigMatrix_12_44_port, 
      sigMatrix_12_43_port, sigMatrix_12_42_port, sigMatrix_12_41_port, 
      sigMatrix_12_40_port, sigMatrix_12_39_port, sigMatrix_12_38_port, 
      sigMatrix_12_37_port, sigMatrix_12_36_port, sigMatrix_12_35_port, 
      sigMatrix_12_34_port, sigMatrix_12_33_port, sigMatrix_12_32_port, 
      sigMatrix_12_31_port, sigMatrix_12_30_port, sigMatrix_12_29_port, 
      sigMatrix_12_28_port, sigMatrix_12_27_port, sigMatrix_12_26_port, 
      sigMatrix_12_25_port, sigMatrix_12_24_port, sigMatrix_12_23_port, 
      sigMatrix_12_22_port, sigMatrix_12_21_port, sigMatrix_12_20_port, 
      sigMatrix_12_19_port, sigMatrix_12_18_port, sigMatrix_12_17_port, 
      sigMatrix_12_16_port, sigMatrix_12_15_port, sigMatrix_12_14_port, 
      sigMatrix_12_13_port, sigMatrix_12_12_port, sigMatrix_12_11_port, 
      sigMatrix_12_10_port, sigMatrix_12_9_port, sigMatrix_12_8_port, 
      sigMatrix_12_7_port, sigMatrix_12_6_port, sigMatrix_12_5_port, 
      sigMatrix_12_4_port, sigMatrix_12_3_port, sigMatrix_12_2_port, 
      sigMatrix_12_1_port, sigMatrix_12_0_port, sigMatrix_13_127_port, 
      sigMatrix_13_126_port, sigMatrix_13_125_port, sigMatrix_13_124_port, 
      sigMatrix_13_123_port, sigMatrix_13_122_port, sigMatrix_13_121_port, 
      sigMatrix_13_120_port, sigMatrix_13_119_port, sigMatrix_13_118_port, 
      sigMatrix_13_117_port, sigMatrix_13_116_port, sigMatrix_13_115_port, 
      sigMatrix_13_114_port, sigMatrix_13_113_port, sigMatrix_13_112_port, 
      sigMatrix_13_111_port, sigMatrix_13_110_port, sigMatrix_13_109_port, 
      sigMatrix_13_108_port, sigMatrix_13_107_port, sigMatrix_13_106_port, 
      sigMatrix_13_105_port, sigMatrix_13_104_port, sigMatrix_13_103_port, 
      sigMatrix_13_102_port, sigMatrix_13_101_port, sigMatrix_13_100_port, 
      sigMatrix_13_99_port, sigMatrix_13_98_port, sigMatrix_13_97_port, 
      sigMatrix_13_96_port, sigMatrix_13_95_port, sigMatrix_13_94_port, 
      sigMatrix_13_93_port, sigMatrix_13_92_port, sigMatrix_13_91_port, 
      sigMatrix_13_90_port, sigMatrix_13_89_port, sigMatrix_13_88_port, 
      sigMatrix_13_87_port, sigMatrix_13_86_port, sigMatrix_13_85_port, 
      sigMatrix_13_84_port, sigMatrix_13_83_port, sigMatrix_13_82_port, 
      sigMatrix_13_81_port, sigMatrix_13_80_port, sigMatrix_13_79_port, 
      sigMatrix_13_78_port, sigMatrix_13_77_port, sigMatrix_13_76_port, 
      sigMatrix_13_75_port, sigMatrix_13_74_port, sigMatrix_13_73_port, 
      sigMatrix_13_72_port, sigMatrix_13_71_port, sigMatrix_13_70_port, 
      sigMatrix_13_69_port, sigMatrix_13_68_port, sigMatrix_13_67_port, 
      sigMatrix_13_66_port, sigMatrix_13_65_port, sigMatrix_13_63_port, 
      sigMatrix_13_62_port, sigMatrix_13_61_port, sigMatrix_13_60_port, 
      sigMatrix_13_59_port, sigMatrix_13_58_port, sigMatrix_13_57_port, 
      sigMatrix_13_56_port, sigMatrix_13_55_port, sigMatrix_13_54_port, 
      sigMatrix_13_53_port, sigMatrix_13_52_port, sigMatrix_13_51_port, 
      sigMatrix_13_50_port, sigMatrix_13_49_port, sigMatrix_13_48_port, 
      sigMatrix_13_47_port, sigMatrix_13_46_port, sigMatrix_13_45_port, 
      sigMatrix_13_44_port, sigMatrix_13_43_port, sigMatrix_13_42_port, 
      sigMatrix_13_41_port, sigMatrix_13_40_port, sigMatrix_13_39_port, 
      sigMatrix_13_38_port, sigMatrix_13_37_port, sigMatrix_13_36_port, 
      sigMatrix_13_35_port, sigMatrix_13_34_port, sigMatrix_13_33_port, 
      sigMatrix_13_32_port, sigMatrix_13_31_port, sigMatrix_13_30_port, 
      sigMatrix_13_29_port, sigMatrix_13_28_port, sigMatrix_13_27_port, 
      sigMatrix_13_26_port, sigMatrix_13_25_port, sigMatrix_13_24_port, 
      sigMatrix_13_23_port, sigMatrix_13_22_port, sigMatrix_13_21_port, 
      sigMatrix_13_20_port, sigMatrix_13_19_port, sigMatrix_13_18_port, 
      sigMatrix_13_17_port, sigMatrix_13_16_port, sigMatrix_13_15_port, 
      sigMatrix_13_14_port, sigMatrix_13_13_port, sigMatrix_13_12_port, 
      sigMatrix_13_11_port, sigMatrix_13_10_port, sigMatrix_13_9_port, 
      sigMatrix_13_8_port, sigMatrix_13_7_port, sigMatrix_13_6_port, 
      sigMatrix_13_5_port, sigMatrix_13_4_port, sigMatrix_13_3_port, 
      sigMatrix_13_2_port, sigMatrix_13_1_port, sigMatrix_13_0_port, 
      sigMatrix_14_127_port, sigMatrix_14_126_port, sigMatrix_14_125_port, 
      sigMatrix_14_124_port, sigMatrix_14_123_port, sigMatrix_14_122_port, 
      sigMatrix_14_121_port, sigMatrix_14_120_port, sigMatrix_14_119_port, 
      sigMatrix_14_118_port, sigMatrix_14_117_port, sigMatrix_14_116_port, 
      sigMatrix_14_115_port, sigMatrix_14_114_port, sigMatrix_14_113_port, 
      sigMatrix_14_112_port, sigMatrix_14_111_port, sigMatrix_14_110_port, 
      sigMatrix_14_109_port, sigMatrix_14_108_port, sigMatrix_14_107_port, 
      sigMatrix_14_106_port, sigMatrix_14_105_port, sigMatrix_14_104_port, 
      sigMatrix_14_103_port, sigMatrix_14_102_port, sigMatrix_14_101_port, 
      sigMatrix_14_100_port, sigMatrix_14_99_port, sigMatrix_14_98_port, 
      sigMatrix_14_97_port, sigMatrix_14_96_port, sigMatrix_14_95_port, 
      sigMatrix_14_94_port, sigMatrix_14_93_port, sigMatrix_14_92_port, 
      sigMatrix_14_91_port, sigMatrix_14_90_port, sigMatrix_14_89_port, 
      sigMatrix_14_88_port, sigMatrix_14_87_port, sigMatrix_14_86_port, 
      sigMatrix_14_85_port, sigMatrix_14_84_port, sigMatrix_14_83_port, 
      sigMatrix_14_82_port, sigMatrix_14_81_port, sigMatrix_14_80_port, 
      sigMatrix_14_79_port, sigMatrix_14_78_port, sigMatrix_14_77_port, 
      sigMatrix_14_76_port, sigMatrix_14_75_port, sigMatrix_14_74_port, 
      sigMatrix_14_73_port, sigMatrix_14_72_port, sigMatrix_14_71_port, 
      sigMatrix_14_70_port, sigMatrix_14_69_port, sigMatrix_14_68_port, 
      sigMatrix_14_67_port, sigMatrix_14_66_port, sigMatrix_14_65_port, 
      sigMatrix_14_63_port, sigMatrix_14_62_port, sigMatrix_14_61_port, 
      sigMatrix_14_60_port, sigMatrix_14_59_port, sigMatrix_14_58_port, 
      sigMatrix_14_57_port, sigMatrix_14_56_port, sigMatrix_14_55_port, 
      sigMatrix_14_54_port, sigMatrix_14_53_port, sigMatrix_14_52_port, 
      sigMatrix_14_51_port, sigMatrix_14_50_port, sigMatrix_14_49_port, 
      sigMatrix_14_48_port, sigMatrix_14_47_port, sigMatrix_14_46_port, 
      sigMatrix_14_45_port, sigMatrix_14_44_port, sigMatrix_14_43_port, 
      sigMatrix_14_42_port, sigMatrix_14_41_port, sigMatrix_14_40_port, 
      sigMatrix_14_39_port, sigMatrix_14_38_port, sigMatrix_14_37_port, 
      sigMatrix_14_36_port, sigMatrix_14_35_port, sigMatrix_14_34_port, 
      sigMatrix_14_33_port, sigMatrix_14_32_port, sigMatrix_14_31_port, 
      sigMatrix_14_30_port, sigMatrix_14_29_port, sigMatrix_14_28_port, 
      sigMatrix_14_27_port, sigMatrix_14_26_port, sigMatrix_14_25_port, 
      sigMatrix_14_24_port, sigMatrix_14_23_port, sigMatrix_14_22_port, 
      sigMatrix_14_21_port, sigMatrix_14_20_port, sigMatrix_14_19_port, 
      sigMatrix_14_18_port, sigMatrix_14_17_port, sigMatrix_14_16_port, 
      sigMatrix_14_15_port, sigMatrix_14_14_port, sigMatrix_14_13_port, 
      sigMatrix_14_12_port, sigMatrix_14_11_port, sigMatrix_14_10_port, 
      sigMatrix_14_9_port, sigMatrix_14_8_port, sigMatrix_14_7_port, 
      sigMatrix_14_6_port, sigMatrix_14_5_port, sigMatrix_14_4_port, 
      sigMatrix_14_3_port, sigMatrix_14_2_port, sigMatrix_14_1_port, 
      sigMatrix_14_0_port, n1, n_3221, n_3222, n_3223, n_3224, n_3225, n_3226, 
      n_3227, n_3228, n_3229, n_3230, n_3231, n_3232, n_3233, n_3234, n_3235, 
      n_3236, n_3237, n_3238, n_3239, n_3240, n_3241, n_3242, n_3243, n_3244, 
      n_3245, n_3246, n_3247, n_3248, n_3249, n_3250, n_3251, n_3252, n_3253, 
      n_3254, n_3255, n_3256, n_3257, n_3258, n_3259, n_3260, n_3261, n_3262, 
      n_3263, n_3264, n_3265, n_3266, n_3267, n_3268, n_3269, n_3270, n_3271, 
      n_3272, n_3273, n_3274, n_3275, n_3276, n_3277, n_3278, n_3279, n_3280, 
      n_3281, n_3282, n_3283, n_3284, n_3285, n_3286, n_3287, n_3288, n_3289, 
      n_3290, n_3291, n_3292, n_3293, n_3294, n_3295, n_3296, n_3297, n_3298, 
      n_3299 : std_logic;

begin
   
   X_Logic0_port <= '0';
   n1 <= '0';
   booth_mul_row_special_1_0 : booth_mul_row_special_N64_RADIX3 port map( A(63)
                           => A(31), A(62) => A(31), A(61) => A(31), A(60) => 
                           A(31), A(59) => A(31), A(58) => A(31), A(57) => 
                           A(31), A(56) => A(31), A(55) => A(31), A(54) => 
                           A(31), A(53) => A(31), A(52) => A(31), A(51) => 
                           A(31), A(50) => A(31), A(49) => A(31), A(48) => 
                           A(31), A(47) => A(31), A(46) => A(31), A(45) => 
                           A(31), A(44) => A(31), A(43) => A(31), A(42) => 
                           A(31), A(41) => A(31), A(40) => A(31), A(39) => 
                           A(31), A(38) => A(31), A(37) => A(31), A(36) => 
                           A(31), A(35) => A(31), A(34) => A(31), A(33) => 
                           A(31), A(32) => A(31), A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), encoderIn(2) => B(1), 
                           encoderIn(1) => B(0), encoderIn(0) => X_Logic0_port,
                           nextA(63) => sigMatrix_0_127_port, nextA(62) => 
                           sigMatrix_0_126_port, nextA(61) => 
                           sigMatrix_0_125_port, nextA(60) => 
                           sigMatrix_0_124_port, nextA(59) => 
                           sigMatrix_0_123_port, nextA(58) => 
                           sigMatrix_0_122_port, nextA(57) => 
                           sigMatrix_0_121_port, nextA(56) => 
                           sigMatrix_0_120_port, nextA(55) => 
                           sigMatrix_0_119_port, nextA(54) => 
                           sigMatrix_0_118_port, nextA(53) => 
                           sigMatrix_0_117_port, nextA(52) => 
                           sigMatrix_0_116_port, nextA(51) => 
                           sigMatrix_0_115_port, nextA(50) => 
                           sigMatrix_0_114_port, nextA(49) => 
                           sigMatrix_0_113_port, nextA(48) => 
                           sigMatrix_0_112_port, nextA(47) => 
                           sigMatrix_0_111_port, nextA(46) => 
                           sigMatrix_0_110_port, nextA(45) => 
                           sigMatrix_0_109_port, nextA(44) => 
                           sigMatrix_0_108_port, nextA(43) => 
                           sigMatrix_0_107_port, nextA(42) => 
                           sigMatrix_0_106_port, nextA(41) => 
                           sigMatrix_0_105_port, nextA(40) => 
                           sigMatrix_0_104_port, nextA(39) => 
                           sigMatrix_0_103_port, nextA(38) => 
                           sigMatrix_0_102_port, nextA(37) => 
                           sigMatrix_0_101_port, nextA(36) => 
                           sigMatrix_0_100_port, nextA(35) => 
                           sigMatrix_0_99_port, nextA(34) => 
                           sigMatrix_0_98_port, nextA(33) => 
                           sigMatrix_0_97_port, nextA(32) => 
                           sigMatrix_0_96_port, nextA(31) => 
                           sigMatrix_0_95_port, nextA(30) => 
                           sigMatrix_0_94_port, nextA(29) => 
                           sigMatrix_0_93_port, nextA(28) => 
                           sigMatrix_0_92_port, nextA(27) => 
                           sigMatrix_0_91_port, nextA(26) => 
                           sigMatrix_0_90_port, nextA(25) => 
                           sigMatrix_0_89_port, nextA(24) => 
                           sigMatrix_0_88_port, nextA(23) => 
                           sigMatrix_0_87_port, nextA(22) => 
                           sigMatrix_0_86_port, nextA(21) => 
                           sigMatrix_0_85_port, nextA(20) => 
                           sigMatrix_0_84_port, nextA(19) => 
                           sigMatrix_0_83_port, nextA(18) => 
                           sigMatrix_0_82_port, nextA(17) => 
                           sigMatrix_0_81_port, nextA(16) => 
                           sigMatrix_0_80_port, nextA(15) => 
                           sigMatrix_0_79_port, nextA(14) => 
                           sigMatrix_0_78_port, nextA(13) => 
                           sigMatrix_0_77_port, nextA(12) => 
                           sigMatrix_0_76_port, nextA(11) => 
                           sigMatrix_0_75_port, nextA(10) => 
                           sigMatrix_0_74_port, nextA(9) => sigMatrix_0_73_port
                           , nextA(8) => sigMatrix_0_72_port, nextA(7) => 
                           sigMatrix_0_71_port, nextA(6) => sigMatrix_0_70_port
                           , nextA(5) => sigMatrix_0_69_port, nextA(4) => 
                           sigMatrix_0_68_port, nextA(3) => sigMatrix_0_67_port
                           , nextA(2) => sigMatrix_0_66_port, nextA(1) => 
                           sigMatrix_0_65_port, nextA(0) => n_3221, nextSum(63)
                           => sigMatrix_0_63_port, nextSum(62) => 
                           sigMatrix_0_62_port, nextSum(61) => 
                           sigMatrix_0_61_port, nextSum(60) => 
                           sigMatrix_0_60_port, nextSum(59) => 
                           sigMatrix_0_59_port, nextSum(58) => 
                           sigMatrix_0_58_port, nextSum(57) => 
                           sigMatrix_0_57_port, nextSum(56) => 
                           sigMatrix_0_56_port, nextSum(55) => 
                           sigMatrix_0_55_port, nextSum(54) => 
                           sigMatrix_0_54_port, nextSum(53) => 
                           sigMatrix_0_53_port, nextSum(52) => 
                           sigMatrix_0_52_port, nextSum(51) => 
                           sigMatrix_0_51_port, nextSum(50) => 
                           sigMatrix_0_50_port, nextSum(49) => 
                           sigMatrix_0_49_port, nextSum(48) => 
                           sigMatrix_0_48_port, nextSum(47) => 
                           sigMatrix_0_47_port, nextSum(46) => 
                           sigMatrix_0_46_port, nextSum(45) => 
                           sigMatrix_0_45_port, nextSum(44) => 
                           sigMatrix_0_44_port, nextSum(43) => 
                           sigMatrix_0_43_port, nextSum(42) => 
                           sigMatrix_0_42_port, nextSum(41) => 
                           sigMatrix_0_41_port, nextSum(40) => 
                           sigMatrix_0_40_port, nextSum(39) => 
                           sigMatrix_0_39_port, nextSum(38) => 
                           sigMatrix_0_38_port, nextSum(37) => 
                           sigMatrix_0_37_port, nextSum(36) => 
                           sigMatrix_0_36_port, nextSum(35) => 
                           sigMatrix_0_35_port, nextSum(34) => 
                           sigMatrix_0_34_port, nextSum(33) => 
                           sigMatrix_0_33_port, nextSum(32) => 
                           sigMatrix_0_32_port, nextSum(31) => 
                           sigMatrix_0_31_port, nextSum(30) => 
                           sigMatrix_0_30_port, nextSum(29) => 
                           sigMatrix_0_29_port, nextSum(28) => 
                           sigMatrix_0_28_port, nextSum(27) => 
                           sigMatrix_0_27_port, nextSum(26) => 
                           sigMatrix_0_26_port, nextSum(25) => 
                           sigMatrix_0_25_port, nextSum(24) => 
                           sigMatrix_0_24_port, nextSum(23) => 
                           sigMatrix_0_23_port, nextSum(22) => 
                           sigMatrix_0_22_port, nextSum(21) => 
                           sigMatrix_0_21_port, nextSum(20) => 
                           sigMatrix_0_20_port, nextSum(19) => 
                           sigMatrix_0_19_port, nextSum(18) => 
                           sigMatrix_0_18_port, nextSum(17) => 
                           sigMatrix_0_17_port, nextSum(16) => 
                           sigMatrix_0_16_port, nextSum(15) => 
                           sigMatrix_0_15_port, nextSum(14) => 
                           sigMatrix_0_14_port, nextSum(13) => 
                           sigMatrix_0_13_port, nextSum(12) => 
                           sigMatrix_0_12_port, nextSum(11) => 
                           sigMatrix_0_11_port, nextSum(10) => 
                           sigMatrix_0_10_port, nextSum(9) => 
                           sigMatrix_0_9_port, nextSum(8) => sigMatrix_0_8_port
                           , nextSum(7) => sigMatrix_0_7_port, nextSum(6) => 
                           sigMatrix_0_6_port, nextSum(5) => sigMatrix_0_5_port
                           , nextSum(4) => sigMatrix_0_4_port, nextSum(3) => 
                           sigMatrix_0_3_port, nextSum(2) => sigMatrix_0_2_port
                           , nextSum(1) => sigMatrix_0_1_port, nextSum(0) => 
                           sigMatrix_0_0_port);
   booth_mul_row_1_1 : booth_mul_row_N64_RADIX3_0 port map( prevA(63) => 
                           sigMatrix_0_127_port, prevA(62) => 
                           sigMatrix_0_126_port, prevA(61) => 
                           sigMatrix_0_125_port, prevA(60) => 
                           sigMatrix_0_124_port, prevA(59) => 
                           sigMatrix_0_123_port, prevA(58) => 
                           sigMatrix_0_122_port, prevA(57) => 
                           sigMatrix_0_121_port, prevA(56) => 
                           sigMatrix_0_120_port, prevA(55) => 
                           sigMatrix_0_119_port, prevA(54) => 
                           sigMatrix_0_118_port, prevA(53) => 
                           sigMatrix_0_117_port, prevA(52) => 
                           sigMatrix_0_116_port, prevA(51) => 
                           sigMatrix_0_115_port, prevA(50) => 
                           sigMatrix_0_114_port, prevA(49) => 
                           sigMatrix_0_113_port, prevA(48) => 
                           sigMatrix_0_112_port, prevA(47) => 
                           sigMatrix_0_111_port, prevA(46) => 
                           sigMatrix_0_110_port, prevA(45) => 
                           sigMatrix_0_109_port, prevA(44) => 
                           sigMatrix_0_108_port, prevA(43) => 
                           sigMatrix_0_107_port, prevA(42) => 
                           sigMatrix_0_106_port, prevA(41) => 
                           sigMatrix_0_105_port, prevA(40) => 
                           sigMatrix_0_104_port, prevA(39) => 
                           sigMatrix_0_103_port, prevA(38) => 
                           sigMatrix_0_102_port, prevA(37) => 
                           sigMatrix_0_101_port, prevA(36) => 
                           sigMatrix_0_100_port, prevA(35) => 
                           sigMatrix_0_99_port, prevA(34) => 
                           sigMatrix_0_98_port, prevA(33) => 
                           sigMatrix_0_97_port, prevA(32) => 
                           sigMatrix_0_96_port, prevA(31) => 
                           sigMatrix_0_95_port, prevA(30) => 
                           sigMatrix_0_94_port, prevA(29) => 
                           sigMatrix_0_93_port, prevA(28) => 
                           sigMatrix_0_92_port, prevA(27) => 
                           sigMatrix_0_91_port, prevA(26) => 
                           sigMatrix_0_90_port, prevA(25) => 
                           sigMatrix_0_89_port, prevA(24) => 
                           sigMatrix_0_88_port, prevA(23) => 
                           sigMatrix_0_87_port, prevA(22) => 
                           sigMatrix_0_86_port, prevA(21) => 
                           sigMatrix_0_85_port, prevA(20) => 
                           sigMatrix_0_84_port, prevA(19) => 
                           sigMatrix_0_83_port, prevA(18) => 
                           sigMatrix_0_82_port, prevA(17) => 
                           sigMatrix_0_81_port, prevA(16) => 
                           sigMatrix_0_80_port, prevA(15) => 
                           sigMatrix_0_79_port, prevA(14) => 
                           sigMatrix_0_78_port, prevA(13) => 
                           sigMatrix_0_77_port, prevA(12) => 
                           sigMatrix_0_76_port, prevA(11) => 
                           sigMatrix_0_75_port, prevA(10) => 
                           sigMatrix_0_74_port, prevA(9) => sigMatrix_0_73_port
                           , prevA(8) => sigMatrix_0_72_port, prevA(7) => 
                           sigMatrix_0_71_port, prevA(6) => sigMatrix_0_70_port
                           , prevA(5) => sigMatrix_0_69_port, prevA(4) => 
                           sigMatrix_0_68_port, prevA(3) => sigMatrix_0_67_port
                           , prevA(2) => sigMatrix_0_66_port, prevA(1) => 
                           sigMatrix_0_65_port, prevA(0) => n1, prevSum(63) => 
                           sigMatrix_0_63_port, prevSum(62) => 
                           sigMatrix_0_62_port, prevSum(61) => 
                           sigMatrix_0_61_port, prevSum(60) => 
                           sigMatrix_0_60_port, prevSum(59) => 
                           sigMatrix_0_59_port, prevSum(58) => 
                           sigMatrix_0_58_port, prevSum(57) => 
                           sigMatrix_0_57_port, prevSum(56) => 
                           sigMatrix_0_56_port, prevSum(55) => 
                           sigMatrix_0_55_port, prevSum(54) => 
                           sigMatrix_0_54_port, prevSum(53) => 
                           sigMatrix_0_53_port, prevSum(52) => 
                           sigMatrix_0_52_port, prevSum(51) => 
                           sigMatrix_0_51_port, prevSum(50) => 
                           sigMatrix_0_50_port, prevSum(49) => 
                           sigMatrix_0_49_port, prevSum(48) => 
                           sigMatrix_0_48_port, prevSum(47) => 
                           sigMatrix_0_47_port, prevSum(46) => 
                           sigMatrix_0_46_port, prevSum(45) => 
                           sigMatrix_0_45_port, prevSum(44) => 
                           sigMatrix_0_44_port, prevSum(43) => 
                           sigMatrix_0_43_port, prevSum(42) => 
                           sigMatrix_0_42_port, prevSum(41) => 
                           sigMatrix_0_41_port, prevSum(40) => 
                           sigMatrix_0_40_port, prevSum(39) => 
                           sigMatrix_0_39_port, prevSum(38) => 
                           sigMatrix_0_38_port, prevSum(37) => 
                           sigMatrix_0_37_port, prevSum(36) => 
                           sigMatrix_0_36_port, prevSum(35) => 
                           sigMatrix_0_35_port, prevSum(34) => 
                           sigMatrix_0_34_port, prevSum(33) => 
                           sigMatrix_0_33_port, prevSum(32) => 
                           sigMatrix_0_32_port, prevSum(31) => 
                           sigMatrix_0_31_port, prevSum(30) => 
                           sigMatrix_0_30_port, prevSum(29) => 
                           sigMatrix_0_29_port, prevSum(28) => 
                           sigMatrix_0_28_port, prevSum(27) => 
                           sigMatrix_0_27_port, prevSum(26) => 
                           sigMatrix_0_26_port, prevSum(25) => 
                           sigMatrix_0_25_port, prevSum(24) => 
                           sigMatrix_0_24_port, prevSum(23) => 
                           sigMatrix_0_23_port, prevSum(22) => 
                           sigMatrix_0_22_port, prevSum(21) => 
                           sigMatrix_0_21_port, prevSum(20) => 
                           sigMatrix_0_20_port, prevSum(19) => 
                           sigMatrix_0_19_port, prevSum(18) => 
                           sigMatrix_0_18_port, prevSum(17) => 
                           sigMatrix_0_17_port, prevSum(16) => 
                           sigMatrix_0_16_port, prevSum(15) => 
                           sigMatrix_0_15_port, prevSum(14) => 
                           sigMatrix_0_14_port, prevSum(13) => 
                           sigMatrix_0_13_port, prevSum(12) => 
                           sigMatrix_0_12_port, prevSum(11) => 
                           sigMatrix_0_11_port, prevSum(10) => 
                           sigMatrix_0_10_port, prevSum(9) => 
                           sigMatrix_0_9_port, prevSum(8) => sigMatrix_0_8_port
                           , prevSum(7) => sigMatrix_0_7_port, prevSum(6) => 
                           sigMatrix_0_6_port, prevSum(5) => sigMatrix_0_5_port
                           , prevSum(4) => sigMatrix_0_4_port, prevSum(3) => 
                           sigMatrix_0_3_port, prevSum(2) => sigMatrix_0_2_port
                           , prevSum(1) => sigMatrix_0_1_port, prevSum(0) => 
                           sigMatrix_0_0_port, encoderIn(2) => B(3), 
                           encoderIn(1) => B(2), encoderIn(0) => B(1), 
                           nextA(63) => sigMatrix_1_127_port, nextA(62) => 
                           sigMatrix_1_126_port, nextA(61) => 
                           sigMatrix_1_125_port, nextA(60) => 
                           sigMatrix_1_124_port, nextA(59) => 
                           sigMatrix_1_123_port, nextA(58) => 
                           sigMatrix_1_122_port, nextA(57) => 
                           sigMatrix_1_121_port, nextA(56) => 
                           sigMatrix_1_120_port, nextA(55) => 
                           sigMatrix_1_119_port, nextA(54) => 
                           sigMatrix_1_118_port, nextA(53) => 
                           sigMatrix_1_117_port, nextA(52) => 
                           sigMatrix_1_116_port, nextA(51) => 
                           sigMatrix_1_115_port, nextA(50) => 
                           sigMatrix_1_114_port, nextA(49) => 
                           sigMatrix_1_113_port, nextA(48) => 
                           sigMatrix_1_112_port, nextA(47) => 
                           sigMatrix_1_111_port, nextA(46) => 
                           sigMatrix_1_110_port, nextA(45) => 
                           sigMatrix_1_109_port, nextA(44) => 
                           sigMatrix_1_108_port, nextA(43) => 
                           sigMatrix_1_107_port, nextA(42) => 
                           sigMatrix_1_106_port, nextA(41) => 
                           sigMatrix_1_105_port, nextA(40) => 
                           sigMatrix_1_104_port, nextA(39) => 
                           sigMatrix_1_103_port, nextA(38) => 
                           sigMatrix_1_102_port, nextA(37) => 
                           sigMatrix_1_101_port, nextA(36) => 
                           sigMatrix_1_100_port, nextA(35) => 
                           sigMatrix_1_99_port, nextA(34) => 
                           sigMatrix_1_98_port, nextA(33) => 
                           sigMatrix_1_97_port, nextA(32) => 
                           sigMatrix_1_96_port, nextA(31) => 
                           sigMatrix_1_95_port, nextA(30) => 
                           sigMatrix_1_94_port, nextA(29) => 
                           sigMatrix_1_93_port, nextA(28) => 
                           sigMatrix_1_92_port, nextA(27) => 
                           sigMatrix_1_91_port, nextA(26) => 
                           sigMatrix_1_90_port, nextA(25) => 
                           sigMatrix_1_89_port, nextA(24) => 
                           sigMatrix_1_88_port, nextA(23) => 
                           sigMatrix_1_87_port, nextA(22) => 
                           sigMatrix_1_86_port, nextA(21) => 
                           sigMatrix_1_85_port, nextA(20) => 
                           sigMatrix_1_84_port, nextA(19) => 
                           sigMatrix_1_83_port, nextA(18) => 
                           sigMatrix_1_82_port, nextA(17) => 
                           sigMatrix_1_81_port, nextA(16) => 
                           sigMatrix_1_80_port, nextA(15) => 
                           sigMatrix_1_79_port, nextA(14) => 
                           sigMatrix_1_78_port, nextA(13) => 
                           sigMatrix_1_77_port, nextA(12) => 
                           sigMatrix_1_76_port, nextA(11) => 
                           sigMatrix_1_75_port, nextA(10) => 
                           sigMatrix_1_74_port, nextA(9) => sigMatrix_1_73_port
                           , nextA(8) => sigMatrix_1_72_port, nextA(7) => 
                           sigMatrix_1_71_port, nextA(6) => sigMatrix_1_70_port
                           , nextA(5) => sigMatrix_1_69_port, nextA(4) => 
                           sigMatrix_1_68_port, nextA(3) => sigMatrix_1_67_port
                           , nextA(2) => sigMatrix_1_66_port, nextA(1) => 
                           sigMatrix_1_65_port, nextA(0) => n_3222, nextSum(63)
                           => sigMatrix_1_63_port, nextSum(62) => 
                           sigMatrix_1_62_port, nextSum(61) => 
                           sigMatrix_1_61_port, nextSum(60) => 
                           sigMatrix_1_60_port, nextSum(59) => 
                           sigMatrix_1_59_port, nextSum(58) => 
                           sigMatrix_1_58_port, nextSum(57) => 
                           sigMatrix_1_57_port, nextSum(56) => 
                           sigMatrix_1_56_port, nextSum(55) => 
                           sigMatrix_1_55_port, nextSum(54) => 
                           sigMatrix_1_54_port, nextSum(53) => 
                           sigMatrix_1_53_port, nextSum(52) => 
                           sigMatrix_1_52_port, nextSum(51) => 
                           sigMatrix_1_51_port, nextSum(50) => 
                           sigMatrix_1_50_port, nextSum(49) => 
                           sigMatrix_1_49_port, nextSum(48) => 
                           sigMatrix_1_48_port, nextSum(47) => 
                           sigMatrix_1_47_port, nextSum(46) => 
                           sigMatrix_1_46_port, nextSum(45) => 
                           sigMatrix_1_45_port, nextSum(44) => 
                           sigMatrix_1_44_port, nextSum(43) => 
                           sigMatrix_1_43_port, nextSum(42) => 
                           sigMatrix_1_42_port, nextSum(41) => 
                           sigMatrix_1_41_port, nextSum(40) => 
                           sigMatrix_1_40_port, nextSum(39) => 
                           sigMatrix_1_39_port, nextSum(38) => 
                           sigMatrix_1_38_port, nextSum(37) => 
                           sigMatrix_1_37_port, nextSum(36) => 
                           sigMatrix_1_36_port, nextSum(35) => 
                           sigMatrix_1_35_port, nextSum(34) => 
                           sigMatrix_1_34_port, nextSum(33) => 
                           sigMatrix_1_33_port, nextSum(32) => 
                           sigMatrix_1_32_port, nextSum(31) => 
                           sigMatrix_1_31_port, nextSum(30) => 
                           sigMatrix_1_30_port, nextSum(29) => 
                           sigMatrix_1_29_port, nextSum(28) => 
                           sigMatrix_1_28_port, nextSum(27) => 
                           sigMatrix_1_27_port, nextSum(26) => 
                           sigMatrix_1_26_port, nextSum(25) => 
                           sigMatrix_1_25_port, nextSum(24) => 
                           sigMatrix_1_24_port, nextSum(23) => 
                           sigMatrix_1_23_port, nextSum(22) => 
                           sigMatrix_1_22_port, nextSum(21) => 
                           sigMatrix_1_21_port, nextSum(20) => 
                           sigMatrix_1_20_port, nextSum(19) => 
                           sigMatrix_1_19_port, nextSum(18) => 
                           sigMatrix_1_18_port, nextSum(17) => 
                           sigMatrix_1_17_port, nextSum(16) => 
                           sigMatrix_1_16_port, nextSum(15) => 
                           sigMatrix_1_15_port, nextSum(14) => 
                           sigMatrix_1_14_port, nextSum(13) => 
                           sigMatrix_1_13_port, nextSum(12) => 
                           sigMatrix_1_12_port, nextSum(11) => 
                           sigMatrix_1_11_port, nextSum(10) => 
                           sigMatrix_1_10_port, nextSum(9) => 
                           sigMatrix_1_9_port, nextSum(8) => sigMatrix_1_8_port
                           , nextSum(7) => sigMatrix_1_7_port, nextSum(6) => 
                           sigMatrix_1_6_port, nextSum(5) => sigMatrix_1_5_port
                           , nextSum(4) => sigMatrix_1_4_port, nextSum(3) => 
                           sigMatrix_1_3_port, nextSum(2) => sigMatrix_1_2_port
                           , nextSum(1) => sigMatrix_1_1_port, nextSum(0) => 
                           sigMatrix_1_0_port);
   booth_mul_row_1_2 : booth_mul_row_N64_RADIX3_14 port map( prevA(63) => 
                           sigMatrix_1_127_port, prevA(62) => 
                           sigMatrix_1_126_port, prevA(61) => 
                           sigMatrix_1_125_port, prevA(60) => 
                           sigMatrix_1_124_port, prevA(59) => 
                           sigMatrix_1_123_port, prevA(58) => 
                           sigMatrix_1_122_port, prevA(57) => 
                           sigMatrix_1_121_port, prevA(56) => 
                           sigMatrix_1_120_port, prevA(55) => 
                           sigMatrix_1_119_port, prevA(54) => 
                           sigMatrix_1_118_port, prevA(53) => 
                           sigMatrix_1_117_port, prevA(52) => 
                           sigMatrix_1_116_port, prevA(51) => 
                           sigMatrix_1_115_port, prevA(50) => 
                           sigMatrix_1_114_port, prevA(49) => 
                           sigMatrix_1_113_port, prevA(48) => 
                           sigMatrix_1_112_port, prevA(47) => 
                           sigMatrix_1_111_port, prevA(46) => 
                           sigMatrix_1_110_port, prevA(45) => 
                           sigMatrix_1_109_port, prevA(44) => 
                           sigMatrix_1_108_port, prevA(43) => 
                           sigMatrix_1_107_port, prevA(42) => 
                           sigMatrix_1_106_port, prevA(41) => 
                           sigMatrix_1_105_port, prevA(40) => 
                           sigMatrix_1_104_port, prevA(39) => 
                           sigMatrix_1_103_port, prevA(38) => 
                           sigMatrix_1_102_port, prevA(37) => 
                           sigMatrix_1_101_port, prevA(36) => 
                           sigMatrix_1_100_port, prevA(35) => 
                           sigMatrix_1_99_port, prevA(34) => 
                           sigMatrix_1_98_port, prevA(33) => 
                           sigMatrix_1_97_port, prevA(32) => 
                           sigMatrix_1_96_port, prevA(31) => 
                           sigMatrix_1_95_port, prevA(30) => 
                           sigMatrix_1_94_port, prevA(29) => 
                           sigMatrix_1_93_port, prevA(28) => 
                           sigMatrix_1_92_port, prevA(27) => 
                           sigMatrix_1_91_port, prevA(26) => 
                           sigMatrix_1_90_port, prevA(25) => 
                           sigMatrix_1_89_port, prevA(24) => 
                           sigMatrix_1_88_port, prevA(23) => 
                           sigMatrix_1_87_port, prevA(22) => 
                           sigMatrix_1_86_port, prevA(21) => 
                           sigMatrix_1_85_port, prevA(20) => 
                           sigMatrix_1_84_port, prevA(19) => 
                           sigMatrix_1_83_port, prevA(18) => 
                           sigMatrix_1_82_port, prevA(17) => 
                           sigMatrix_1_81_port, prevA(16) => 
                           sigMatrix_1_80_port, prevA(15) => 
                           sigMatrix_1_79_port, prevA(14) => 
                           sigMatrix_1_78_port, prevA(13) => 
                           sigMatrix_1_77_port, prevA(12) => 
                           sigMatrix_1_76_port, prevA(11) => 
                           sigMatrix_1_75_port, prevA(10) => 
                           sigMatrix_1_74_port, prevA(9) => sigMatrix_1_73_port
                           , prevA(8) => sigMatrix_1_72_port, prevA(7) => 
                           sigMatrix_1_71_port, prevA(6) => sigMatrix_1_70_port
                           , prevA(5) => sigMatrix_1_69_port, prevA(4) => 
                           sigMatrix_1_68_port, prevA(3) => sigMatrix_1_67_port
                           , prevA(2) => sigMatrix_1_66_port, prevA(1) => 
                           sigMatrix_1_65_port, prevA(0) => n1, prevSum(63) => 
                           sigMatrix_1_63_port, prevSum(62) => 
                           sigMatrix_1_62_port, prevSum(61) => 
                           sigMatrix_1_61_port, prevSum(60) => 
                           sigMatrix_1_60_port, prevSum(59) => 
                           sigMatrix_1_59_port, prevSum(58) => 
                           sigMatrix_1_58_port, prevSum(57) => 
                           sigMatrix_1_57_port, prevSum(56) => 
                           sigMatrix_1_56_port, prevSum(55) => 
                           sigMatrix_1_55_port, prevSum(54) => 
                           sigMatrix_1_54_port, prevSum(53) => 
                           sigMatrix_1_53_port, prevSum(52) => 
                           sigMatrix_1_52_port, prevSum(51) => 
                           sigMatrix_1_51_port, prevSum(50) => 
                           sigMatrix_1_50_port, prevSum(49) => 
                           sigMatrix_1_49_port, prevSum(48) => 
                           sigMatrix_1_48_port, prevSum(47) => 
                           sigMatrix_1_47_port, prevSum(46) => 
                           sigMatrix_1_46_port, prevSum(45) => 
                           sigMatrix_1_45_port, prevSum(44) => 
                           sigMatrix_1_44_port, prevSum(43) => 
                           sigMatrix_1_43_port, prevSum(42) => 
                           sigMatrix_1_42_port, prevSum(41) => 
                           sigMatrix_1_41_port, prevSum(40) => 
                           sigMatrix_1_40_port, prevSum(39) => 
                           sigMatrix_1_39_port, prevSum(38) => 
                           sigMatrix_1_38_port, prevSum(37) => 
                           sigMatrix_1_37_port, prevSum(36) => 
                           sigMatrix_1_36_port, prevSum(35) => 
                           sigMatrix_1_35_port, prevSum(34) => 
                           sigMatrix_1_34_port, prevSum(33) => 
                           sigMatrix_1_33_port, prevSum(32) => 
                           sigMatrix_1_32_port, prevSum(31) => 
                           sigMatrix_1_31_port, prevSum(30) => 
                           sigMatrix_1_30_port, prevSum(29) => 
                           sigMatrix_1_29_port, prevSum(28) => 
                           sigMatrix_1_28_port, prevSum(27) => 
                           sigMatrix_1_27_port, prevSum(26) => 
                           sigMatrix_1_26_port, prevSum(25) => 
                           sigMatrix_1_25_port, prevSum(24) => 
                           sigMatrix_1_24_port, prevSum(23) => 
                           sigMatrix_1_23_port, prevSum(22) => 
                           sigMatrix_1_22_port, prevSum(21) => 
                           sigMatrix_1_21_port, prevSum(20) => 
                           sigMatrix_1_20_port, prevSum(19) => 
                           sigMatrix_1_19_port, prevSum(18) => 
                           sigMatrix_1_18_port, prevSum(17) => 
                           sigMatrix_1_17_port, prevSum(16) => 
                           sigMatrix_1_16_port, prevSum(15) => 
                           sigMatrix_1_15_port, prevSum(14) => 
                           sigMatrix_1_14_port, prevSum(13) => 
                           sigMatrix_1_13_port, prevSum(12) => 
                           sigMatrix_1_12_port, prevSum(11) => 
                           sigMatrix_1_11_port, prevSum(10) => 
                           sigMatrix_1_10_port, prevSum(9) => 
                           sigMatrix_1_9_port, prevSum(8) => sigMatrix_1_8_port
                           , prevSum(7) => sigMatrix_1_7_port, prevSum(6) => 
                           sigMatrix_1_6_port, prevSum(5) => sigMatrix_1_5_port
                           , prevSum(4) => sigMatrix_1_4_port, prevSum(3) => 
                           sigMatrix_1_3_port, prevSum(2) => sigMatrix_1_2_port
                           , prevSum(1) => sigMatrix_1_1_port, prevSum(0) => 
                           sigMatrix_1_0_port, encoderIn(2) => B(5), 
                           encoderIn(1) => B(4), encoderIn(0) => B(3), 
                           nextA(63) => sigMatrix_2_127_port, nextA(62) => 
                           sigMatrix_2_126_port, nextA(61) => 
                           sigMatrix_2_125_port, nextA(60) => 
                           sigMatrix_2_124_port, nextA(59) => 
                           sigMatrix_2_123_port, nextA(58) => 
                           sigMatrix_2_122_port, nextA(57) => 
                           sigMatrix_2_121_port, nextA(56) => 
                           sigMatrix_2_120_port, nextA(55) => 
                           sigMatrix_2_119_port, nextA(54) => 
                           sigMatrix_2_118_port, nextA(53) => 
                           sigMatrix_2_117_port, nextA(52) => 
                           sigMatrix_2_116_port, nextA(51) => 
                           sigMatrix_2_115_port, nextA(50) => 
                           sigMatrix_2_114_port, nextA(49) => 
                           sigMatrix_2_113_port, nextA(48) => 
                           sigMatrix_2_112_port, nextA(47) => 
                           sigMatrix_2_111_port, nextA(46) => 
                           sigMatrix_2_110_port, nextA(45) => 
                           sigMatrix_2_109_port, nextA(44) => 
                           sigMatrix_2_108_port, nextA(43) => 
                           sigMatrix_2_107_port, nextA(42) => 
                           sigMatrix_2_106_port, nextA(41) => 
                           sigMatrix_2_105_port, nextA(40) => 
                           sigMatrix_2_104_port, nextA(39) => 
                           sigMatrix_2_103_port, nextA(38) => 
                           sigMatrix_2_102_port, nextA(37) => 
                           sigMatrix_2_101_port, nextA(36) => 
                           sigMatrix_2_100_port, nextA(35) => 
                           sigMatrix_2_99_port, nextA(34) => 
                           sigMatrix_2_98_port, nextA(33) => 
                           sigMatrix_2_97_port, nextA(32) => 
                           sigMatrix_2_96_port, nextA(31) => 
                           sigMatrix_2_95_port, nextA(30) => 
                           sigMatrix_2_94_port, nextA(29) => 
                           sigMatrix_2_93_port, nextA(28) => 
                           sigMatrix_2_92_port, nextA(27) => 
                           sigMatrix_2_91_port, nextA(26) => 
                           sigMatrix_2_90_port, nextA(25) => 
                           sigMatrix_2_89_port, nextA(24) => 
                           sigMatrix_2_88_port, nextA(23) => 
                           sigMatrix_2_87_port, nextA(22) => 
                           sigMatrix_2_86_port, nextA(21) => 
                           sigMatrix_2_85_port, nextA(20) => 
                           sigMatrix_2_84_port, nextA(19) => 
                           sigMatrix_2_83_port, nextA(18) => 
                           sigMatrix_2_82_port, nextA(17) => 
                           sigMatrix_2_81_port, nextA(16) => 
                           sigMatrix_2_80_port, nextA(15) => 
                           sigMatrix_2_79_port, nextA(14) => 
                           sigMatrix_2_78_port, nextA(13) => 
                           sigMatrix_2_77_port, nextA(12) => 
                           sigMatrix_2_76_port, nextA(11) => 
                           sigMatrix_2_75_port, nextA(10) => 
                           sigMatrix_2_74_port, nextA(9) => sigMatrix_2_73_port
                           , nextA(8) => sigMatrix_2_72_port, nextA(7) => 
                           sigMatrix_2_71_port, nextA(6) => sigMatrix_2_70_port
                           , nextA(5) => sigMatrix_2_69_port, nextA(4) => 
                           sigMatrix_2_68_port, nextA(3) => sigMatrix_2_67_port
                           , nextA(2) => sigMatrix_2_66_port, nextA(1) => 
                           sigMatrix_2_65_port, nextA(0) => n_3223, nextSum(63)
                           => sigMatrix_2_63_port, nextSum(62) => 
                           sigMatrix_2_62_port, nextSum(61) => 
                           sigMatrix_2_61_port, nextSum(60) => 
                           sigMatrix_2_60_port, nextSum(59) => 
                           sigMatrix_2_59_port, nextSum(58) => 
                           sigMatrix_2_58_port, nextSum(57) => 
                           sigMatrix_2_57_port, nextSum(56) => 
                           sigMatrix_2_56_port, nextSum(55) => 
                           sigMatrix_2_55_port, nextSum(54) => 
                           sigMatrix_2_54_port, nextSum(53) => 
                           sigMatrix_2_53_port, nextSum(52) => 
                           sigMatrix_2_52_port, nextSum(51) => 
                           sigMatrix_2_51_port, nextSum(50) => 
                           sigMatrix_2_50_port, nextSum(49) => 
                           sigMatrix_2_49_port, nextSum(48) => 
                           sigMatrix_2_48_port, nextSum(47) => 
                           sigMatrix_2_47_port, nextSum(46) => 
                           sigMatrix_2_46_port, nextSum(45) => 
                           sigMatrix_2_45_port, nextSum(44) => 
                           sigMatrix_2_44_port, nextSum(43) => 
                           sigMatrix_2_43_port, nextSum(42) => 
                           sigMatrix_2_42_port, nextSum(41) => 
                           sigMatrix_2_41_port, nextSum(40) => 
                           sigMatrix_2_40_port, nextSum(39) => 
                           sigMatrix_2_39_port, nextSum(38) => 
                           sigMatrix_2_38_port, nextSum(37) => 
                           sigMatrix_2_37_port, nextSum(36) => 
                           sigMatrix_2_36_port, nextSum(35) => 
                           sigMatrix_2_35_port, nextSum(34) => 
                           sigMatrix_2_34_port, nextSum(33) => 
                           sigMatrix_2_33_port, nextSum(32) => 
                           sigMatrix_2_32_port, nextSum(31) => 
                           sigMatrix_2_31_port, nextSum(30) => 
                           sigMatrix_2_30_port, nextSum(29) => 
                           sigMatrix_2_29_port, nextSum(28) => 
                           sigMatrix_2_28_port, nextSum(27) => 
                           sigMatrix_2_27_port, nextSum(26) => 
                           sigMatrix_2_26_port, nextSum(25) => 
                           sigMatrix_2_25_port, nextSum(24) => 
                           sigMatrix_2_24_port, nextSum(23) => 
                           sigMatrix_2_23_port, nextSum(22) => 
                           sigMatrix_2_22_port, nextSum(21) => 
                           sigMatrix_2_21_port, nextSum(20) => 
                           sigMatrix_2_20_port, nextSum(19) => 
                           sigMatrix_2_19_port, nextSum(18) => 
                           sigMatrix_2_18_port, nextSum(17) => 
                           sigMatrix_2_17_port, nextSum(16) => 
                           sigMatrix_2_16_port, nextSum(15) => 
                           sigMatrix_2_15_port, nextSum(14) => 
                           sigMatrix_2_14_port, nextSum(13) => 
                           sigMatrix_2_13_port, nextSum(12) => 
                           sigMatrix_2_12_port, nextSum(11) => 
                           sigMatrix_2_11_port, nextSum(10) => 
                           sigMatrix_2_10_port, nextSum(9) => 
                           sigMatrix_2_9_port, nextSum(8) => sigMatrix_2_8_port
                           , nextSum(7) => sigMatrix_2_7_port, nextSum(6) => 
                           sigMatrix_2_6_port, nextSum(5) => sigMatrix_2_5_port
                           , nextSum(4) => sigMatrix_2_4_port, nextSum(3) => 
                           sigMatrix_2_3_port, nextSum(2) => sigMatrix_2_2_port
                           , nextSum(1) => sigMatrix_2_1_port, nextSum(0) => 
                           sigMatrix_2_0_port);
   booth_mul_row_1_3 : booth_mul_row_N64_RADIX3_13 port map( prevA(63) => 
                           sigMatrix_2_127_port, prevA(62) => 
                           sigMatrix_2_126_port, prevA(61) => 
                           sigMatrix_2_125_port, prevA(60) => 
                           sigMatrix_2_124_port, prevA(59) => 
                           sigMatrix_2_123_port, prevA(58) => 
                           sigMatrix_2_122_port, prevA(57) => 
                           sigMatrix_2_121_port, prevA(56) => 
                           sigMatrix_2_120_port, prevA(55) => 
                           sigMatrix_2_119_port, prevA(54) => 
                           sigMatrix_2_118_port, prevA(53) => 
                           sigMatrix_2_117_port, prevA(52) => 
                           sigMatrix_2_116_port, prevA(51) => 
                           sigMatrix_2_115_port, prevA(50) => 
                           sigMatrix_2_114_port, prevA(49) => 
                           sigMatrix_2_113_port, prevA(48) => 
                           sigMatrix_2_112_port, prevA(47) => 
                           sigMatrix_2_111_port, prevA(46) => 
                           sigMatrix_2_110_port, prevA(45) => 
                           sigMatrix_2_109_port, prevA(44) => 
                           sigMatrix_2_108_port, prevA(43) => 
                           sigMatrix_2_107_port, prevA(42) => 
                           sigMatrix_2_106_port, prevA(41) => 
                           sigMatrix_2_105_port, prevA(40) => 
                           sigMatrix_2_104_port, prevA(39) => 
                           sigMatrix_2_103_port, prevA(38) => 
                           sigMatrix_2_102_port, prevA(37) => 
                           sigMatrix_2_101_port, prevA(36) => 
                           sigMatrix_2_100_port, prevA(35) => 
                           sigMatrix_2_99_port, prevA(34) => 
                           sigMatrix_2_98_port, prevA(33) => 
                           sigMatrix_2_97_port, prevA(32) => 
                           sigMatrix_2_96_port, prevA(31) => 
                           sigMatrix_2_95_port, prevA(30) => 
                           sigMatrix_2_94_port, prevA(29) => 
                           sigMatrix_2_93_port, prevA(28) => 
                           sigMatrix_2_92_port, prevA(27) => 
                           sigMatrix_2_91_port, prevA(26) => 
                           sigMatrix_2_90_port, prevA(25) => 
                           sigMatrix_2_89_port, prevA(24) => 
                           sigMatrix_2_88_port, prevA(23) => 
                           sigMatrix_2_87_port, prevA(22) => 
                           sigMatrix_2_86_port, prevA(21) => 
                           sigMatrix_2_85_port, prevA(20) => 
                           sigMatrix_2_84_port, prevA(19) => 
                           sigMatrix_2_83_port, prevA(18) => 
                           sigMatrix_2_82_port, prevA(17) => 
                           sigMatrix_2_81_port, prevA(16) => 
                           sigMatrix_2_80_port, prevA(15) => 
                           sigMatrix_2_79_port, prevA(14) => 
                           sigMatrix_2_78_port, prevA(13) => 
                           sigMatrix_2_77_port, prevA(12) => 
                           sigMatrix_2_76_port, prevA(11) => 
                           sigMatrix_2_75_port, prevA(10) => 
                           sigMatrix_2_74_port, prevA(9) => sigMatrix_2_73_port
                           , prevA(8) => sigMatrix_2_72_port, prevA(7) => 
                           sigMatrix_2_71_port, prevA(6) => sigMatrix_2_70_port
                           , prevA(5) => sigMatrix_2_69_port, prevA(4) => 
                           sigMatrix_2_68_port, prevA(3) => sigMatrix_2_67_port
                           , prevA(2) => sigMatrix_2_66_port, prevA(1) => 
                           sigMatrix_2_65_port, prevA(0) => n1, prevSum(63) => 
                           sigMatrix_2_63_port, prevSum(62) => 
                           sigMatrix_2_62_port, prevSum(61) => 
                           sigMatrix_2_61_port, prevSum(60) => 
                           sigMatrix_2_60_port, prevSum(59) => 
                           sigMatrix_2_59_port, prevSum(58) => 
                           sigMatrix_2_58_port, prevSum(57) => 
                           sigMatrix_2_57_port, prevSum(56) => 
                           sigMatrix_2_56_port, prevSum(55) => 
                           sigMatrix_2_55_port, prevSum(54) => 
                           sigMatrix_2_54_port, prevSum(53) => 
                           sigMatrix_2_53_port, prevSum(52) => 
                           sigMatrix_2_52_port, prevSum(51) => 
                           sigMatrix_2_51_port, prevSum(50) => 
                           sigMatrix_2_50_port, prevSum(49) => 
                           sigMatrix_2_49_port, prevSum(48) => 
                           sigMatrix_2_48_port, prevSum(47) => 
                           sigMatrix_2_47_port, prevSum(46) => 
                           sigMatrix_2_46_port, prevSum(45) => 
                           sigMatrix_2_45_port, prevSum(44) => 
                           sigMatrix_2_44_port, prevSum(43) => 
                           sigMatrix_2_43_port, prevSum(42) => 
                           sigMatrix_2_42_port, prevSum(41) => 
                           sigMatrix_2_41_port, prevSum(40) => 
                           sigMatrix_2_40_port, prevSum(39) => 
                           sigMatrix_2_39_port, prevSum(38) => 
                           sigMatrix_2_38_port, prevSum(37) => 
                           sigMatrix_2_37_port, prevSum(36) => 
                           sigMatrix_2_36_port, prevSum(35) => 
                           sigMatrix_2_35_port, prevSum(34) => 
                           sigMatrix_2_34_port, prevSum(33) => 
                           sigMatrix_2_33_port, prevSum(32) => 
                           sigMatrix_2_32_port, prevSum(31) => 
                           sigMatrix_2_31_port, prevSum(30) => 
                           sigMatrix_2_30_port, prevSum(29) => 
                           sigMatrix_2_29_port, prevSum(28) => 
                           sigMatrix_2_28_port, prevSum(27) => 
                           sigMatrix_2_27_port, prevSum(26) => 
                           sigMatrix_2_26_port, prevSum(25) => 
                           sigMatrix_2_25_port, prevSum(24) => 
                           sigMatrix_2_24_port, prevSum(23) => 
                           sigMatrix_2_23_port, prevSum(22) => 
                           sigMatrix_2_22_port, prevSum(21) => 
                           sigMatrix_2_21_port, prevSum(20) => 
                           sigMatrix_2_20_port, prevSum(19) => 
                           sigMatrix_2_19_port, prevSum(18) => 
                           sigMatrix_2_18_port, prevSum(17) => 
                           sigMatrix_2_17_port, prevSum(16) => 
                           sigMatrix_2_16_port, prevSum(15) => 
                           sigMatrix_2_15_port, prevSum(14) => 
                           sigMatrix_2_14_port, prevSum(13) => 
                           sigMatrix_2_13_port, prevSum(12) => 
                           sigMatrix_2_12_port, prevSum(11) => 
                           sigMatrix_2_11_port, prevSum(10) => 
                           sigMatrix_2_10_port, prevSum(9) => 
                           sigMatrix_2_9_port, prevSum(8) => sigMatrix_2_8_port
                           , prevSum(7) => sigMatrix_2_7_port, prevSum(6) => 
                           sigMatrix_2_6_port, prevSum(5) => sigMatrix_2_5_port
                           , prevSum(4) => sigMatrix_2_4_port, prevSum(3) => 
                           sigMatrix_2_3_port, prevSum(2) => sigMatrix_2_2_port
                           , prevSum(1) => sigMatrix_2_1_port, prevSum(0) => 
                           sigMatrix_2_0_port, encoderIn(2) => B(7), 
                           encoderIn(1) => B(6), encoderIn(0) => B(5), 
                           nextA(63) => sigMatrix_3_127_port, nextA(62) => 
                           sigMatrix_3_126_port, nextA(61) => 
                           sigMatrix_3_125_port, nextA(60) => 
                           sigMatrix_3_124_port, nextA(59) => 
                           sigMatrix_3_123_port, nextA(58) => 
                           sigMatrix_3_122_port, nextA(57) => 
                           sigMatrix_3_121_port, nextA(56) => 
                           sigMatrix_3_120_port, nextA(55) => 
                           sigMatrix_3_119_port, nextA(54) => 
                           sigMatrix_3_118_port, nextA(53) => 
                           sigMatrix_3_117_port, nextA(52) => 
                           sigMatrix_3_116_port, nextA(51) => 
                           sigMatrix_3_115_port, nextA(50) => 
                           sigMatrix_3_114_port, nextA(49) => 
                           sigMatrix_3_113_port, nextA(48) => 
                           sigMatrix_3_112_port, nextA(47) => 
                           sigMatrix_3_111_port, nextA(46) => 
                           sigMatrix_3_110_port, nextA(45) => 
                           sigMatrix_3_109_port, nextA(44) => 
                           sigMatrix_3_108_port, nextA(43) => 
                           sigMatrix_3_107_port, nextA(42) => 
                           sigMatrix_3_106_port, nextA(41) => 
                           sigMatrix_3_105_port, nextA(40) => 
                           sigMatrix_3_104_port, nextA(39) => 
                           sigMatrix_3_103_port, nextA(38) => 
                           sigMatrix_3_102_port, nextA(37) => 
                           sigMatrix_3_101_port, nextA(36) => 
                           sigMatrix_3_100_port, nextA(35) => 
                           sigMatrix_3_99_port, nextA(34) => 
                           sigMatrix_3_98_port, nextA(33) => 
                           sigMatrix_3_97_port, nextA(32) => 
                           sigMatrix_3_96_port, nextA(31) => 
                           sigMatrix_3_95_port, nextA(30) => 
                           sigMatrix_3_94_port, nextA(29) => 
                           sigMatrix_3_93_port, nextA(28) => 
                           sigMatrix_3_92_port, nextA(27) => 
                           sigMatrix_3_91_port, nextA(26) => 
                           sigMatrix_3_90_port, nextA(25) => 
                           sigMatrix_3_89_port, nextA(24) => 
                           sigMatrix_3_88_port, nextA(23) => 
                           sigMatrix_3_87_port, nextA(22) => 
                           sigMatrix_3_86_port, nextA(21) => 
                           sigMatrix_3_85_port, nextA(20) => 
                           sigMatrix_3_84_port, nextA(19) => 
                           sigMatrix_3_83_port, nextA(18) => 
                           sigMatrix_3_82_port, nextA(17) => 
                           sigMatrix_3_81_port, nextA(16) => 
                           sigMatrix_3_80_port, nextA(15) => 
                           sigMatrix_3_79_port, nextA(14) => 
                           sigMatrix_3_78_port, nextA(13) => 
                           sigMatrix_3_77_port, nextA(12) => 
                           sigMatrix_3_76_port, nextA(11) => 
                           sigMatrix_3_75_port, nextA(10) => 
                           sigMatrix_3_74_port, nextA(9) => sigMatrix_3_73_port
                           , nextA(8) => sigMatrix_3_72_port, nextA(7) => 
                           sigMatrix_3_71_port, nextA(6) => sigMatrix_3_70_port
                           , nextA(5) => sigMatrix_3_69_port, nextA(4) => 
                           sigMatrix_3_68_port, nextA(3) => sigMatrix_3_67_port
                           , nextA(2) => sigMatrix_3_66_port, nextA(1) => 
                           sigMatrix_3_65_port, nextA(0) => n_3224, nextSum(63)
                           => sigMatrix_3_63_port, nextSum(62) => 
                           sigMatrix_3_62_port, nextSum(61) => 
                           sigMatrix_3_61_port, nextSum(60) => 
                           sigMatrix_3_60_port, nextSum(59) => 
                           sigMatrix_3_59_port, nextSum(58) => 
                           sigMatrix_3_58_port, nextSum(57) => 
                           sigMatrix_3_57_port, nextSum(56) => 
                           sigMatrix_3_56_port, nextSum(55) => 
                           sigMatrix_3_55_port, nextSum(54) => 
                           sigMatrix_3_54_port, nextSum(53) => 
                           sigMatrix_3_53_port, nextSum(52) => 
                           sigMatrix_3_52_port, nextSum(51) => 
                           sigMatrix_3_51_port, nextSum(50) => 
                           sigMatrix_3_50_port, nextSum(49) => 
                           sigMatrix_3_49_port, nextSum(48) => 
                           sigMatrix_3_48_port, nextSum(47) => 
                           sigMatrix_3_47_port, nextSum(46) => 
                           sigMatrix_3_46_port, nextSum(45) => 
                           sigMatrix_3_45_port, nextSum(44) => 
                           sigMatrix_3_44_port, nextSum(43) => 
                           sigMatrix_3_43_port, nextSum(42) => 
                           sigMatrix_3_42_port, nextSum(41) => 
                           sigMatrix_3_41_port, nextSum(40) => 
                           sigMatrix_3_40_port, nextSum(39) => 
                           sigMatrix_3_39_port, nextSum(38) => 
                           sigMatrix_3_38_port, nextSum(37) => 
                           sigMatrix_3_37_port, nextSum(36) => 
                           sigMatrix_3_36_port, nextSum(35) => 
                           sigMatrix_3_35_port, nextSum(34) => 
                           sigMatrix_3_34_port, nextSum(33) => 
                           sigMatrix_3_33_port, nextSum(32) => 
                           sigMatrix_3_32_port, nextSum(31) => 
                           sigMatrix_3_31_port, nextSum(30) => 
                           sigMatrix_3_30_port, nextSum(29) => 
                           sigMatrix_3_29_port, nextSum(28) => 
                           sigMatrix_3_28_port, nextSum(27) => 
                           sigMatrix_3_27_port, nextSum(26) => 
                           sigMatrix_3_26_port, nextSum(25) => 
                           sigMatrix_3_25_port, nextSum(24) => 
                           sigMatrix_3_24_port, nextSum(23) => 
                           sigMatrix_3_23_port, nextSum(22) => 
                           sigMatrix_3_22_port, nextSum(21) => 
                           sigMatrix_3_21_port, nextSum(20) => 
                           sigMatrix_3_20_port, nextSum(19) => 
                           sigMatrix_3_19_port, nextSum(18) => 
                           sigMatrix_3_18_port, nextSum(17) => 
                           sigMatrix_3_17_port, nextSum(16) => 
                           sigMatrix_3_16_port, nextSum(15) => 
                           sigMatrix_3_15_port, nextSum(14) => 
                           sigMatrix_3_14_port, nextSum(13) => 
                           sigMatrix_3_13_port, nextSum(12) => 
                           sigMatrix_3_12_port, nextSum(11) => 
                           sigMatrix_3_11_port, nextSum(10) => 
                           sigMatrix_3_10_port, nextSum(9) => 
                           sigMatrix_3_9_port, nextSum(8) => sigMatrix_3_8_port
                           , nextSum(7) => sigMatrix_3_7_port, nextSum(6) => 
                           sigMatrix_3_6_port, nextSum(5) => sigMatrix_3_5_port
                           , nextSum(4) => sigMatrix_3_4_port, nextSum(3) => 
                           sigMatrix_3_3_port, nextSum(2) => sigMatrix_3_2_port
                           , nextSum(1) => sigMatrix_3_1_port, nextSum(0) => 
                           sigMatrix_3_0_port);
   booth_mul_row_1_4 : booth_mul_row_N64_RADIX3_12 port map( prevA(63) => 
                           sigMatrix_3_127_port, prevA(62) => 
                           sigMatrix_3_126_port, prevA(61) => 
                           sigMatrix_3_125_port, prevA(60) => 
                           sigMatrix_3_124_port, prevA(59) => 
                           sigMatrix_3_123_port, prevA(58) => 
                           sigMatrix_3_122_port, prevA(57) => 
                           sigMatrix_3_121_port, prevA(56) => 
                           sigMatrix_3_120_port, prevA(55) => 
                           sigMatrix_3_119_port, prevA(54) => 
                           sigMatrix_3_118_port, prevA(53) => 
                           sigMatrix_3_117_port, prevA(52) => 
                           sigMatrix_3_116_port, prevA(51) => 
                           sigMatrix_3_115_port, prevA(50) => 
                           sigMatrix_3_114_port, prevA(49) => 
                           sigMatrix_3_113_port, prevA(48) => 
                           sigMatrix_3_112_port, prevA(47) => 
                           sigMatrix_3_111_port, prevA(46) => 
                           sigMatrix_3_110_port, prevA(45) => 
                           sigMatrix_3_109_port, prevA(44) => 
                           sigMatrix_3_108_port, prevA(43) => 
                           sigMatrix_3_107_port, prevA(42) => 
                           sigMatrix_3_106_port, prevA(41) => 
                           sigMatrix_3_105_port, prevA(40) => 
                           sigMatrix_3_104_port, prevA(39) => 
                           sigMatrix_3_103_port, prevA(38) => 
                           sigMatrix_3_102_port, prevA(37) => 
                           sigMatrix_3_101_port, prevA(36) => 
                           sigMatrix_3_100_port, prevA(35) => 
                           sigMatrix_3_99_port, prevA(34) => 
                           sigMatrix_3_98_port, prevA(33) => 
                           sigMatrix_3_97_port, prevA(32) => 
                           sigMatrix_3_96_port, prevA(31) => 
                           sigMatrix_3_95_port, prevA(30) => 
                           sigMatrix_3_94_port, prevA(29) => 
                           sigMatrix_3_93_port, prevA(28) => 
                           sigMatrix_3_92_port, prevA(27) => 
                           sigMatrix_3_91_port, prevA(26) => 
                           sigMatrix_3_90_port, prevA(25) => 
                           sigMatrix_3_89_port, prevA(24) => 
                           sigMatrix_3_88_port, prevA(23) => 
                           sigMatrix_3_87_port, prevA(22) => 
                           sigMatrix_3_86_port, prevA(21) => 
                           sigMatrix_3_85_port, prevA(20) => 
                           sigMatrix_3_84_port, prevA(19) => 
                           sigMatrix_3_83_port, prevA(18) => 
                           sigMatrix_3_82_port, prevA(17) => 
                           sigMatrix_3_81_port, prevA(16) => 
                           sigMatrix_3_80_port, prevA(15) => 
                           sigMatrix_3_79_port, prevA(14) => 
                           sigMatrix_3_78_port, prevA(13) => 
                           sigMatrix_3_77_port, prevA(12) => 
                           sigMatrix_3_76_port, prevA(11) => 
                           sigMatrix_3_75_port, prevA(10) => 
                           sigMatrix_3_74_port, prevA(9) => sigMatrix_3_73_port
                           , prevA(8) => sigMatrix_3_72_port, prevA(7) => 
                           sigMatrix_3_71_port, prevA(6) => sigMatrix_3_70_port
                           , prevA(5) => sigMatrix_3_69_port, prevA(4) => 
                           sigMatrix_3_68_port, prevA(3) => sigMatrix_3_67_port
                           , prevA(2) => sigMatrix_3_66_port, prevA(1) => 
                           sigMatrix_3_65_port, prevA(0) => n1, prevSum(63) => 
                           sigMatrix_3_63_port, prevSum(62) => 
                           sigMatrix_3_62_port, prevSum(61) => 
                           sigMatrix_3_61_port, prevSum(60) => 
                           sigMatrix_3_60_port, prevSum(59) => 
                           sigMatrix_3_59_port, prevSum(58) => 
                           sigMatrix_3_58_port, prevSum(57) => 
                           sigMatrix_3_57_port, prevSum(56) => 
                           sigMatrix_3_56_port, prevSum(55) => 
                           sigMatrix_3_55_port, prevSum(54) => 
                           sigMatrix_3_54_port, prevSum(53) => 
                           sigMatrix_3_53_port, prevSum(52) => 
                           sigMatrix_3_52_port, prevSum(51) => 
                           sigMatrix_3_51_port, prevSum(50) => 
                           sigMatrix_3_50_port, prevSum(49) => 
                           sigMatrix_3_49_port, prevSum(48) => 
                           sigMatrix_3_48_port, prevSum(47) => 
                           sigMatrix_3_47_port, prevSum(46) => 
                           sigMatrix_3_46_port, prevSum(45) => 
                           sigMatrix_3_45_port, prevSum(44) => 
                           sigMatrix_3_44_port, prevSum(43) => 
                           sigMatrix_3_43_port, prevSum(42) => 
                           sigMatrix_3_42_port, prevSum(41) => 
                           sigMatrix_3_41_port, prevSum(40) => 
                           sigMatrix_3_40_port, prevSum(39) => 
                           sigMatrix_3_39_port, prevSum(38) => 
                           sigMatrix_3_38_port, prevSum(37) => 
                           sigMatrix_3_37_port, prevSum(36) => 
                           sigMatrix_3_36_port, prevSum(35) => 
                           sigMatrix_3_35_port, prevSum(34) => 
                           sigMatrix_3_34_port, prevSum(33) => 
                           sigMatrix_3_33_port, prevSum(32) => 
                           sigMatrix_3_32_port, prevSum(31) => 
                           sigMatrix_3_31_port, prevSum(30) => 
                           sigMatrix_3_30_port, prevSum(29) => 
                           sigMatrix_3_29_port, prevSum(28) => 
                           sigMatrix_3_28_port, prevSum(27) => 
                           sigMatrix_3_27_port, prevSum(26) => 
                           sigMatrix_3_26_port, prevSum(25) => 
                           sigMatrix_3_25_port, prevSum(24) => 
                           sigMatrix_3_24_port, prevSum(23) => 
                           sigMatrix_3_23_port, prevSum(22) => 
                           sigMatrix_3_22_port, prevSum(21) => 
                           sigMatrix_3_21_port, prevSum(20) => 
                           sigMatrix_3_20_port, prevSum(19) => 
                           sigMatrix_3_19_port, prevSum(18) => 
                           sigMatrix_3_18_port, prevSum(17) => 
                           sigMatrix_3_17_port, prevSum(16) => 
                           sigMatrix_3_16_port, prevSum(15) => 
                           sigMatrix_3_15_port, prevSum(14) => 
                           sigMatrix_3_14_port, prevSum(13) => 
                           sigMatrix_3_13_port, prevSum(12) => 
                           sigMatrix_3_12_port, prevSum(11) => 
                           sigMatrix_3_11_port, prevSum(10) => 
                           sigMatrix_3_10_port, prevSum(9) => 
                           sigMatrix_3_9_port, prevSum(8) => sigMatrix_3_8_port
                           , prevSum(7) => sigMatrix_3_7_port, prevSum(6) => 
                           sigMatrix_3_6_port, prevSum(5) => sigMatrix_3_5_port
                           , prevSum(4) => sigMatrix_3_4_port, prevSum(3) => 
                           sigMatrix_3_3_port, prevSum(2) => sigMatrix_3_2_port
                           , prevSum(1) => sigMatrix_3_1_port, prevSum(0) => 
                           sigMatrix_3_0_port, encoderIn(2) => B(9), 
                           encoderIn(1) => B(8), encoderIn(0) => B(7), 
                           nextA(63) => sigMatrix_4_127_port, nextA(62) => 
                           sigMatrix_4_126_port, nextA(61) => 
                           sigMatrix_4_125_port, nextA(60) => 
                           sigMatrix_4_124_port, nextA(59) => 
                           sigMatrix_4_123_port, nextA(58) => 
                           sigMatrix_4_122_port, nextA(57) => 
                           sigMatrix_4_121_port, nextA(56) => 
                           sigMatrix_4_120_port, nextA(55) => 
                           sigMatrix_4_119_port, nextA(54) => 
                           sigMatrix_4_118_port, nextA(53) => 
                           sigMatrix_4_117_port, nextA(52) => 
                           sigMatrix_4_116_port, nextA(51) => 
                           sigMatrix_4_115_port, nextA(50) => 
                           sigMatrix_4_114_port, nextA(49) => 
                           sigMatrix_4_113_port, nextA(48) => 
                           sigMatrix_4_112_port, nextA(47) => 
                           sigMatrix_4_111_port, nextA(46) => 
                           sigMatrix_4_110_port, nextA(45) => 
                           sigMatrix_4_109_port, nextA(44) => 
                           sigMatrix_4_108_port, nextA(43) => 
                           sigMatrix_4_107_port, nextA(42) => 
                           sigMatrix_4_106_port, nextA(41) => 
                           sigMatrix_4_105_port, nextA(40) => 
                           sigMatrix_4_104_port, nextA(39) => 
                           sigMatrix_4_103_port, nextA(38) => 
                           sigMatrix_4_102_port, nextA(37) => 
                           sigMatrix_4_101_port, nextA(36) => 
                           sigMatrix_4_100_port, nextA(35) => 
                           sigMatrix_4_99_port, nextA(34) => 
                           sigMatrix_4_98_port, nextA(33) => 
                           sigMatrix_4_97_port, nextA(32) => 
                           sigMatrix_4_96_port, nextA(31) => 
                           sigMatrix_4_95_port, nextA(30) => 
                           sigMatrix_4_94_port, nextA(29) => 
                           sigMatrix_4_93_port, nextA(28) => 
                           sigMatrix_4_92_port, nextA(27) => 
                           sigMatrix_4_91_port, nextA(26) => 
                           sigMatrix_4_90_port, nextA(25) => 
                           sigMatrix_4_89_port, nextA(24) => 
                           sigMatrix_4_88_port, nextA(23) => 
                           sigMatrix_4_87_port, nextA(22) => 
                           sigMatrix_4_86_port, nextA(21) => 
                           sigMatrix_4_85_port, nextA(20) => 
                           sigMatrix_4_84_port, nextA(19) => 
                           sigMatrix_4_83_port, nextA(18) => 
                           sigMatrix_4_82_port, nextA(17) => 
                           sigMatrix_4_81_port, nextA(16) => 
                           sigMatrix_4_80_port, nextA(15) => 
                           sigMatrix_4_79_port, nextA(14) => 
                           sigMatrix_4_78_port, nextA(13) => 
                           sigMatrix_4_77_port, nextA(12) => 
                           sigMatrix_4_76_port, nextA(11) => 
                           sigMatrix_4_75_port, nextA(10) => 
                           sigMatrix_4_74_port, nextA(9) => sigMatrix_4_73_port
                           , nextA(8) => sigMatrix_4_72_port, nextA(7) => 
                           sigMatrix_4_71_port, nextA(6) => sigMatrix_4_70_port
                           , nextA(5) => sigMatrix_4_69_port, nextA(4) => 
                           sigMatrix_4_68_port, nextA(3) => sigMatrix_4_67_port
                           , nextA(2) => sigMatrix_4_66_port, nextA(1) => 
                           sigMatrix_4_65_port, nextA(0) => n_3225, nextSum(63)
                           => sigMatrix_4_63_port, nextSum(62) => 
                           sigMatrix_4_62_port, nextSum(61) => 
                           sigMatrix_4_61_port, nextSum(60) => 
                           sigMatrix_4_60_port, nextSum(59) => 
                           sigMatrix_4_59_port, nextSum(58) => 
                           sigMatrix_4_58_port, nextSum(57) => 
                           sigMatrix_4_57_port, nextSum(56) => 
                           sigMatrix_4_56_port, nextSum(55) => 
                           sigMatrix_4_55_port, nextSum(54) => 
                           sigMatrix_4_54_port, nextSum(53) => 
                           sigMatrix_4_53_port, nextSum(52) => 
                           sigMatrix_4_52_port, nextSum(51) => 
                           sigMatrix_4_51_port, nextSum(50) => 
                           sigMatrix_4_50_port, nextSum(49) => 
                           sigMatrix_4_49_port, nextSum(48) => 
                           sigMatrix_4_48_port, nextSum(47) => 
                           sigMatrix_4_47_port, nextSum(46) => 
                           sigMatrix_4_46_port, nextSum(45) => 
                           sigMatrix_4_45_port, nextSum(44) => 
                           sigMatrix_4_44_port, nextSum(43) => 
                           sigMatrix_4_43_port, nextSum(42) => 
                           sigMatrix_4_42_port, nextSum(41) => 
                           sigMatrix_4_41_port, nextSum(40) => 
                           sigMatrix_4_40_port, nextSum(39) => 
                           sigMatrix_4_39_port, nextSum(38) => 
                           sigMatrix_4_38_port, nextSum(37) => 
                           sigMatrix_4_37_port, nextSum(36) => 
                           sigMatrix_4_36_port, nextSum(35) => 
                           sigMatrix_4_35_port, nextSum(34) => 
                           sigMatrix_4_34_port, nextSum(33) => 
                           sigMatrix_4_33_port, nextSum(32) => 
                           sigMatrix_4_32_port, nextSum(31) => 
                           sigMatrix_4_31_port, nextSum(30) => 
                           sigMatrix_4_30_port, nextSum(29) => 
                           sigMatrix_4_29_port, nextSum(28) => 
                           sigMatrix_4_28_port, nextSum(27) => 
                           sigMatrix_4_27_port, nextSum(26) => 
                           sigMatrix_4_26_port, nextSum(25) => 
                           sigMatrix_4_25_port, nextSum(24) => 
                           sigMatrix_4_24_port, nextSum(23) => 
                           sigMatrix_4_23_port, nextSum(22) => 
                           sigMatrix_4_22_port, nextSum(21) => 
                           sigMatrix_4_21_port, nextSum(20) => 
                           sigMatrix_4_20_port, nextSum(19) => 
                           sigMatrix_4_19_port, nextSum(18) => 
                           sigMatrix_4_18_port, nextSum(17) => 
                           sigMatrix_4_17_port, nextSum(16) => 
                           sigMatrix_4_16_port, nextSum(15) => 
                           sigMatrix_4_15_port, nextSum(14) => 
                           sigMatrix_4_14_port, nextSum(13) => 
                           sigMatrix_4_13_port, nextSum(12) => 
                           sigMatrix_4_12_port, nextSum(11) => 
                           sigMatrix_4_11_port, nextSum(10) => 
                           sigMatrix_4_10_port, nextSum(9) => 
                           sigMatrix_4_9_port, nextSum(8) => sigMatrix_4_8_port
                           , nextSum(7) => sigMatrix_4_7_port, nextSum(6) => 
                           sigMatrix_4_6_port, nextSum(5) => sigMatrix_4_5_port
                           , nextSum(4) => sigMatrix_4_4_port, nextSum(3) => 
                           sigMatrix_4_3_port, nextSum(2) => sigMatrix_4_2_port
                           , nextSum(1) => sigMatrix_4_1_port, nextSum(0) => 
                           sigMatrix_4_0_port);
   booth_mul_row_1_5 : booth_mul_row_N64_RADIX3_11 port map( prevA(63) => 
                           sigMatrix_4_127_port, prevA(62) => 
                           sigMatrix_4_126_port, prevA(61) => 
                           sigMatrix_4_125_port, prevA(60) => 
                           sigMatrix_4_124_port, prevA(59) => 
                           sigMatrix_4_123_port, prevA(58) => 
                           sigMatrix_4_122_port, prevA(57) => 
                           sigMatrix_4_121_port, prevA(56) => 
                           sigMatrix_4_120_port, prevA(55) => 
                           sigMatrix_4_119_port, prevA(54) => 
                           sigMatrix_4_118_port, prevA(53) => 
                           sigMatrix_4_117_port, prevA(52) => 
                           sigMatrix_4_116_port, prevA(51) => 
                           sigMatrix_4_115_port, prevA(50) => 
                           sigMatrix_4_114_port, prevA(49) => 
                           sigMatrix_4_113_port, prevA(48) => 
                           sigMatrix_4_112_port, prevA(47) => 
                           sigMatrix_4_111_port, prevA(46) => 
                           sigMatrix_4_110_port, prevA(45) => 
                           sigMatrix_4_109_port, prevA(44) => 
                           sigMatrix_4_108_port, prevA(43) => 
                           sigMatrix_4_107_port, prevA(42) => 
                           sigMatrix_4_106_port, prevA(41) => 
                           sigMatrix_4_105_port, prevA(40) => 
                           sigMatrix_4_104_port, prevA(39) => 
                           sigMatrix_4_103_port, prevA(38) => 
                           sigMatrix_4_102_port, prevA(37) => 
                           sigMatrix_4_101_port, prevA(36) => 
                           sigMatrix_4_100_port, prevA(35) => 
                           sigMatrix_4_99_port, prevA(34) => 
                           sigMatrix_4_98_port, prevA(33) => 
                           sigMatrix_4_97_port, prevA(32) => 
                           sigMatrix_4_96_port, prevA(31) => 
                           sigMatrix_4_95_port, prevA(30) => 
                           sigMatrix_4_94_port, prevA(29) => 
                           sigMatrix_4_93_port, prevA(28) => 
                           sigMatrix_4_92_port, prevA(27) => 
                           sigMatrix_4_91_port, prevA(26) => 
                           sigMatrix_4_90_port, prevA(25) => 
                           sigMatrix_4_89_port, prevA(24) => 
                           sigMatrix_4_88_port, prevA(23) => 
                           sigMatrix_4_87_port, prevA(22) => 
                           sigMatrix_4_86_port, prevA(21) => 
                           sigMatrix_4_85_port, prevA(20) => 
                           sigMatrix_4_84_port, prevA(19) => 
                           sigMatrix_4_83_port, prevA(18) => 
                           sigMatrix_4_82_port, prevA(17) => 
                           sigMatrix_4_81_port, prevA(16) => 
                           sigMatrix_4_80_port, prevA(15) => 
                           sigMatrix_4_79_port, prevA(14) => 
                           sigMatrix_4_78_port, prevA(13) => 
                           sigMatrix_4_77_port, prevA(12) => 
                           sigMatrix_4_76_port, prevA(11) => 
                           sigMatrix_4_75_port, prevA(10) => 
                           sigMatrix_4_74_port, prevA(9) => sigMatrix_4_73_port
                           , prevA(8) => sigMatrix_4_72_port, prevA(7) => 
                           sigMatrix_4_71_port, prevA(6) => sigMatrix_4_70_port
                           , prevA(5) => sigMatrix_4_69_port, prevA(4) => 
                           sigMatrix_4_68_port, prevA(3) => sigMatrix_4_67_port
                           , prevA(2) => sigMatrix_4_66_port, prevA(1) => 
                           sigMatrix_4_65_port, prevA(0) => n1, prevSum(63) => 
                           sigMatrix_4_63_port, prevSum(62) => 
                           sigMatrix_4_62_port, prevSum(61) => 
                           sigMatrix_4_61_port, prevSum(60) => 
                           sigMatrix_4_60_port, prevSum(59) => 
                           sigMatrix_4_59_port, prevSum(58) => 
                           sigMatrix_4_58_port, prevSum(57) => 
                           sigMatrix_4_57_port, prevSum(56) => 
                           sigMatrix_4_56_port, prevSum(55) => 
                           sigMatrix_4_55_port, prevSum(54) => 
                           sigMatrix_4_54_port, prevSum(53) => 
                           sigMatrix_4_53_port, prevSum(52) => 
                           sigMatrix_4_52_port, prevSum(51) => 
                           sigMatrix_4_51_port, prevSum(50) => 
                           sigMatrix_4_50_port, prevSum(49) => 
                           sigMatrix_4_49_port, prevSum(48) => 
                           sigMatrix_4_48_port, prevSum(47) => 
                           sigMatrix_4_47_port, prevSum(46) => 
                           sigMatrix_4_46_port, prevSum(45) => 
                           sigMatrix_4_45_port, prevSum(44) => 
                           sigMatrix_4_44_port, prevSum(43) => 
                           sigMatrix_4_43_port, prevSum(42) => 
                           sigMatrix_4_42_port, prevSum(41) => 
                           sigMatrix_4_41_port, prevSum(40) => 
                           sigMatrix_4_40_port, prevSum(39) => 
                           sigMatrix_4_39_port, prevSum(38) => 
                           sigMatrix_4_38_port, prevSum(37) => 
                           sigMatrix_4_37_port, prevSum(36) => 
                           sigMatrix_4_36_port, prevSum(35) => 
                           sigMatrix_4_35_port, prevSum(34) => 
                           sigMatrix_4_34_port, prevSum(33) => 
                           sigMatrix_4_33_port, prevSum(32) => 
                           sigMatrix_4_32_port, prevSum(31) => 
                           sigMatrix_4_31_port, prevSum(30) => 
                           sigMatrix_4_30_port, prevSum(29) => 
                           sigMatrix_4_29_port, prevSum(28) => 
                           sigMatrix_4_28_port, prevSum(27) => 
                           sigMatrix_4_27_port, prevSum(26) => 
                           sigMatrix_4_26_port, prevSum(25) => 
                           sigMatrix_4_25_port, prevSum(24) => 
                           sigMatrix_4_24_port, prevSum(23) => 
                           sigMatrix_4_23_port, prevSum(22) => 
                           sigMatrix_4_22_port, prevSum(21) => 
                           sigMatrix_4_21_port, prevSum(20) => 
                           sigMatrix_4_20_port, prevSum(19) => 
                           sigMatrix_4_19_port, prevSum(18) => 
                           sigMatrix_4_18_port, prevSum(17) => 
                           sigMatrix_4_17_port, prevSum(16) => 
                           sigMatrix_4_16_port, prevSum(15) => 
                           sigMatrix_4_15_port, prevSum(14) => 
                           sigMatrix_4_14_port, prevSum(13) => 
                           sigMatrix_4_13_port, prevSum(12) => 
                           sigMatrix_4_12_port, prevSum(11) => 
                           sigMatrix_4_11_port, prevSum(10) => 
                           sigMatrix_4_10_port, prevSum(9) => 
                           sigMatrix_4_9_port, prevSum(8) => sigMatrix_4_8_port
                           , prevSum(7) => sigMatrix_4_7_port, prevSum(6) => 
                           sigMatrix_4_6_port, prevSum(5) => sigMatrix_4_5_port
                           , prevSum(4) => sigMatrix_4_4_port, prevSum(3) => 
                           sigMatrix_4_3_port, prevSum(2) => sigMatrix_4_2_port
                           , prevSum(1) => sigMatrix_4_1_port, prevSum(0) => 
                           sigMatrix_4_0_port, encoderIn(2) => B(11), 
                           encoderIn(1) => B(10), encoderIn(0) => B(9), 
                           nextA(63) => sigMatrix_5_127_port, nextA(62) => 
                           sigMatrix_5_126_port, nextA(61) => 
                           sigMatrix_5_125_port, nextA(60) => 
                           sigMatrix_5_124_port, nextA(59) => 
                           sigMatrix_5_123_port, nextA(58) => 
                           sigMatrix_5_122_port, nextA(57) => 
                           sigMatrix_5_121_port, nextA(56) => 
                           sigMatrix_5_120_port, nextA(55) => 
                           sigMatrix_5_119_port, nextA(54) => 
                           sigMatrix_5_118_port, nextA(53) => 
                           sigMatrix_5_117_port, nextA(52) => 
                           sigMatrix_5_116_port, nextA(51) => 
                           sigMatrix_5_115_port, nextA(50) => 
                           sigMatrix_5_114_port, nextA(49) => 
                           sigMatrix_5_113_port, nextA(48) => 
                           sigMatrix_5_112_port, nextA(47) => 
                           sigMatrix_5_111_port, nextA(46) => 
                           sigMatrix_5_110_port, nextA(45) => 
                           sigMatrix_5_109_port, nextA(44) => 
                           sigMatrix_5_108_port, nextA(43) => 
                           sigMatrix_5_107_port, nextA(42) => 
                           sigMatrix_5_106_port, nextA(41) => 
                           sigMatrix_5_105_port, nextA(40) => 
                           sigMatrix_5_104_port, nextA(39) => 
                           sigMatrix_5_103_port, nextA(38) => 
                           sigMatrix_5_102_port, nextA(37) => 
                           sigMatrix_5_101_port, nextA(36) => 
                           sigMatrix_5_100_port, nextA(35) => 
                           sigMatrix_5_99_port, nextA(34) => 
                           sigMatrix_5_98_port, nextA(33) => 
                           sigMatrix_5_97_port, nextA(32) => 
                           sigMatrix_5_96_port, nextA(31) => 
                           sigMatrix_5_95_port, nextA(30) => 
                           sigMatrix_5_94_port, nextA(29) => 
                           sigMatrix_5_93_port, nextA(28) => 
                           sigMatrix_5_92_port, nextA(27) => 
                           sigMatrix_5_91_port, nextA(26) => 
                           sigMatrix_5_90_port, nextA(25) => 
                           sigMatrix_5_89_port, nextA(24) => 
                           sigMatrix_5_88_port, nextA(23) => 
                           sigMatrix_5_87_port, nextA(22) => 
                           sigMatrix_5_86_port, nextA(21) => 
                           sigMatrix_5_85_port, nextA(20) => 
                           sigMatrix_5_84_port, nextA(19) => 
                           sigMatrix_5_83_port, nextA(18) => 
                           sigMatrix_5_82_port, nextA(17) => 
                           sigMatrix_5_81_port, nextA(16) => 
                           sigMatrix_5_80_port, nextA(15) => 
                           sigMatrix_5_79_port, nextA(14) => 
                           sigMatrix_5_78_port, nextA(13) => 
                           sigMatrix_5_77_port, nextA(12) => 
                           sigMatrix_5_76_port, nextA(11) => 
                           sigMatrix_5_75_port, nextA(10) => 
                           sigMatrix_5_74_port, nextA(9) => sigMatrix_5_73_port
                           , nextA(8) => sigMatrix_5_72_port, nextA(7) => 
                           sigMatrix_5_71_port, nextA(6) => sigMatrix_5_70_port
                           , nextA(5) => sigMatrix_5_69_port, nextA(4) => 
                           sigMatrix_5_68_port, nextA(3) => sigMatrix_5_67_port
                           , nextA(2) => sigMatrix_5_66_port, nextA(1) => 
                           sigMatrix_5_65_port, nextA(0) => n_3226, nextSum(63)
                           => sigMatrix_5_63_port, nextSum(62) => 
                           sigMatrix_5_62_port, nextSum(61) => 
                           sigMatrix_5_61_port, nextSum(60) => 
                           sigMatrix_5_60_port, nextSum(59) => 
                           sigMatrix_5_59_port, nextSum(58) => 
                           sigMatrix_5_58_port, nextSum(57) => 
                           sigMatrix_5_57_port, nextSum(56) => 
                           sigMatrix_5_56_port, nextSum(55) => 
                           sigMatrix_5_55_port, nextSum(54) => 
                           sigMatrix_5_54_port, nextSum(53) => 
                           sigMatrix_5_53_port, nextSum(52) => 
                           sigMatrix_5_52_port, nextSum(51) => 
                           sigMatrix_5_51_port, nextSum(50) => 
                           sigMatrix_5_50_port, nextSum(49) => 
                           sigMatrix_5_49_port, nextSum(48) => 
                           sigMatrix_5_48_port, nextSum(47) => 
                           sigMatrix_5_47_port, nextSum(46) => 
                           sigMatrix_5_46_port, nextSum(45) => 
                           sigMatrix_5_45_port, nextSum(44) => 
                           sigMatrix_5_44_port, nextSum(43) => 
                           sigMatrix_5_43_port, nextSum(42) => 
                           sigMatrix_5_42_port, nextSum(41) => 
                           sigMatrix_5_41_port, nextSum(40) => 
                           sigMatrix_5_40_port, nextSum(39) => 
                           sigMatrix_5_39_port, nextSum(38) => 
                           sigMatrix_5_38_port, nextSum(37) => 
                           sigMatrix_5_37_port, nextSum(36) => 
                           sigMatrix_5_36_port, nextSum(35) => 
                           sigMatrix_5_35_port, nextSum(34) => 
                           sigMatrix_5_34_port, nextSum(33) => 
                           sigMatrix_5_33_port, nextSum(32) => 
                           sigMatrix_5_32_port, nextSum(31) => 
                           sigMatrix_5_31_port, nextSum(30) => 
                           sigMatrix_5_30_port, nextSum(29) => 
                           sigMatrix_5_29_port, nextSum(28) => 
                           sigMatrix_5_28_port, nextSum(27) => 
                           sigMatrix_5_27_port, nextSum(26) => 
                           sigMatrix_5_26_port, nextSum(25) => 
                           sigMatrix_5_25_port, nextSum(24) => 
                           sigMatrix_5_24_port, nextSum(23) => 
                           sigMatrix_5_23_port, nextSum(22) => 
                           sigMatrix_5_22_port, nextSum(21) => 
                           sigMatrix_5_21_port, nextSum(20) => 
                           sigMatrix_5_20_port, nextSum(19) => 
                           sigMatrix_5_19_port, nextSum(18) => 
                           sigMatrix_5_18_port, nextSum(17) => 
                           sigMatrix_5_17_port, nextSum(16) => 
                           sigMatrix_5_16_port, nextSum(15) => 
                           sigMatrix_5_15_port, nextSum(14) => 
                           sigMatrix_5_14_port, nextSum(13) => 
                           sigMatrix_5_13_port, nextSum(12) => 
                           sigMatrix_5_12_port, nextSum(11) => 
                           sigMatrix_5_11_port, nextSum(10) => 
                           sigMatrix_5_10_port, nextSum(9) => 
                           sigMatrix_5_9_port, nextSum(8) => sigMatrix_5_8_port
                           , nextSum(7) => sigMatrix_5_7_port, nextSum(6) => 
                           sigMatrix_5_6_port, nextSum(5) => sigMatrix_5_5_port
                           , nextSum(4) => sigMatrix_5_4_port, nextSum(3) => 
                           sigMatrix_5_3_port, nextSum(2) => sigMatrix_5_2_port
                           , nextSum(1) => sigMatrix_5_1_port, nextSum(0) => 
                           sigMatrix_5_0_port);
   booth_mul_row_1_6 : booth_mul_row_N64_RADIX3_10 port map( prevA(63) => 
                           sigMatrix_5_127_port, prevA(62) => 
                           sigMatrix_5_126_port, prevA(61) => 
                           sigMatrix_5_125_port, prevA(60) => 
                           sigMatrix_5_124_port, prevA(59) => 
                           sigMatrix_5_123_port, prevA(58) => 
                           sigMatrix_5_122_port, prevA(57) => 
                           sigMatrix_5_121_port, prevA(56) => 
                           sigMatrix_5_120_port, prevA(55) => 
                           sigMatrix_5_119_port, prevA(54) => 
                           sigMatrix_5_118_port, prevA(53) => 
                           sigMatrix_5_117_port, prevA(52) => 
                           sigMatrix_5_116_port, prevA(51) => 
                           sigMatrix_5_115_port, prevA(50) => 
                           sigMatrix_5_114_port, prevA(49) => 
                           sigMatrix_5_113_port, prevA(48) => 
                           sigMatrix_5_112_port, prevA(47) => 
                           sigMatrix_5_111_port, prevA(46) => 
                           sigMatrix_5_110_port, prevA(45) => 
                           sigMatrix_5_109_port, prevA(44) => 
                           sigMatrix_5_108_port, prevA(43) => 
                           sigMatrix_5_107_port, prevA(42) => 
                           sigMatrix_5_106_port, prevA(41) => 
                           sigMatrix_5_105_port, prevA(40) => 
                           sigMatrix_5_104_port, prevA(39) => 
                           sigMatrix_5_103_port, prevA(38) => 
                           sigMatrix_5_102_port, prevA(37) => 
                           sigMatrix_5_101_port, prevA(36) => 
                           sigMatrix_5_100_port, prevA(35) => 
                           sigMatrix_5_99_port, prevA(34) => 
                           sigMatrix_5_98_port, prevA(33) => 
                           sigMatrix_5_97_port, prevA(32) => 
                           sigMatrix_5_96_port, prevA(31) => 
                           sigMatrix_5_95_port, prevA(30) => 
                           sigMatrix_5_94_port, prevA(29) => 
                           sigMatrix_5_93_port, prevA(28) => 
                           sigMatrix_5_92_port, prevA(27) => 
                           sigMatrix_5_91_port, prevA(26) => 
                           sigMatrix_5_90_port, prevA(25) => 
                           sigMatrix_5_89_port, prevA(24) => 
                           sigMatrix_5_88_port, prevA(23) => 
                           sigMatrix_5_87_port, prevA(22) => 
                           sigMatrix_5_86_port, prevA(21) => 
                           sigMatrix_5_85_port, prevA(20) => 
                           sigMatrix_5_84_port, prevA(19) => 
                           sigMatrix_5_83_port, prevA(18) => 
                           sigMatrix_5_82_port, prevA(17) => 
                           sigMatrix_5_81_port, prevA(16) => 
                           sigMatrix_5_80_port, prevA(15) => 
                           sigMatrix_5_79_port, prevA(14) => 
                           sigMatrix_5_78_port, prevA(13) => 
                           sigMatrix_5_77_port, prevA(12) => 
                           sigMatrix_5_76_port, prevA(11) => 
                           sigMatrix_5_75_port, prevA(10) => 
                           sigMatrix_5_74_port, prevA(9) => sigMatrix_5_73_port
                           , prevA(8) => sigMatrix_5_72_port, prevA(7) => 
                           sigMatrix_5_71_port, prevA(6) => sigMatrix_5_70_port
                           , prevA(5) => sigMatrix_5_69_port, prevA(4) => 
                           sigMatrix_5_68_port, prevA(3) => sigMatrix_5_67_port
                           , prevA(2) => sigMatrix_5_66_port, prevA(1) => 
                           sigMatrix_5_65_port, prevA(0) => n1, prevSum(63) => 
                           sigMatrix_5_63_port, prevSum(62) => 
                           sigMatrix_5_62_port, prevSum(61) => 
                           sigMatrix_5_61_port, prevSum(60) => 
                           sigMatrix_5_60_port, prevSum(59) => 
                           sigMatrix_5_59_port, prevSum(58) => 
                           sigMatrix_5_58_port, prevSum(57) => 
                           sigMatrix_5_57_port, prevSum(56) => 
                           sigMatrix_5_56_port, prevSum(55) => 
                           sigMatrix_5_55_port, prevSum(54) => 
                           sigMatrix_5_54_port, prevSum(53) => 
                           sigMatrix_5_53_port, prevSum(52) => 
                           sigMatrix_5_52_port, prevSum(51) => 
                           sigMatrix_5_51_port, prevSum(50) => 
                           sigMatrix_5_50_port, prevSum(49) => 
                           sigMatrix_5_49_port, prevSum(48) => 
                           sigMatrix_5_48_port, prevSum(47) => 
                           sigMatrix_5_47_port, prevSum(46) => 
                           sigMatrix_5_46_port, prevSum(45) => 
                           sigMatrix_5_45_port, prevSum(44) => 
                           sigMatrix_5_44_port, prevSum(43) => 
                           sigMatrix_5_43_port, prevSum(42) => 
                           sigMatrix_5_42_port, prevSum(41) => 
                           sigMatrix_5_41_port, prevSum(40) => 
                           sigMatrix_5_40_port, prevSum(39) => 
                           sigMatrix_5_39_port, prevSum(38) => 
                           sigMatrix_5_38_port, prevSum(37) => 
                           sigMatrix_5_37_port, prevSum(36) => 
                           sigMatrix_5_36_port, prevSum(35) => 
                           sigMatrix_5_35_port, prevSum(34) => 
                           sigMatrix_5_34_port, prevSum(33) => 
                           sigMatrix_5_33_port, prevSum(32) => 
                           sigMatrix_5_32_port, prevSum(31) => 
                           sigMatrix_5_31_port, prevSum(30) => 
                           sigMatrix_5_30_port, prevSum(29) => 
                           sigMatrix_5_29_port, prevSum(28) => 
                           sigMatrix_5_28_port, prevSum(27) => 
                           sigMatrix_5_27_port, prevSum(26) => 
                           sigMatrix_5_26_port, prevSum(25) => 
                           sigMatrix_5_25_port, prevSum(24) => 
                           sigMatrix_5_24_port, prevSum(23) => 
                           sigMatrix_5_23_port, prevSum(22) => 
                           sigMatrix_5_22_port, prevSum(21) => 
                           sigMatrix_5_21_port, prevSum(20) => 
                           sigMatrix_5_20_port, prevSum(19) => 
                           sigMatrix_5_19_port, prevSum(18) => 
                           sigMatrix_5_18_port, prevSum(17) => 
                           sigMatrix_5_17_port, prevSum(16) => 
                           sigMatrix_5_16_port, prevSum(15) => 
                           sigMatrix_5_15_port, prevSum(14) => 
                           sigMatrix_5_14_port, prevSum(13) => 
                           sigMatrix_5_13_port, prevSum(12) => 
                           sigMatrix_5_12_port, prevSum(11) => 
                           sigMatrix_5_11_port, prevSum(10) => 
                           sigMatrix_5_10_port, prevSum(9) => 
                           sigMatrix_5_9_port, prevSum(8) => sigMatrix_5_8_port
                           , prevSum(7) => sigMatrix_5_7_port, prevSum(6) => 
                           sigMatrix_5_6_port, prevSum(5) => sigMatrix_5_5_port
                           , prevSum(4) => sigMatrix_5_4_port, prevSum(3) => 
                           sigMatrix_5_3_port, prevSum(2) => sigMatrix_5_2_port
                           , prevSum(1) => sigMatrix_5_1_port, prevSum(0) => 
                           sigMatrix_5_0_port, encoderIn(2) => B(13), 
                           encoderIn(1) => B(12), encoderIn(0) => B(11), 
                           nextA(63) => sigMatrix_6_127_port, nextA(62) => 
                           sigMatrix_6_126_port, nextA(61) => 
                           sigMatrix_6_125_port, nextA(60) => 
                           sigMatrix_6_124_port, nextA(59) => 
                           sigMatrix_6_123_port, nextA(58) => 
                           sigMatrix_6_122_port, nextA(57) => 
                           sigMatrix_6_121_port, nextA(56) => 
                           sigMatrix_6_120_port, nextA(55) => 
                           sigMatrix_6_119_port, nextA(54) => 
                           sigMatrix_6_118_port, nextA(53) => 
                           sigMatrix_6_117_port, nextA(52) => 
                           sigMatrix_6_116_port, nextA(51) => 
                           sigMatrix_6_115_port, nextA(50) => 
                           sigMatrix_6_114_port, nextA(49) => 
                           sigMatrix_6_113_port, nextA(48) => 
                           sigMatrix_6_112_port, nextA(47) => 
                           sigMatrix_6_111_port, nextA(46) => 
                           sigMatrix_6_110_port, nextA(45) => 
                           sigMatrix_6_109_port, nextA(44) => 
                           sigMatrix_6_108_port, nextA(43) => 
                           sigMatrix_6_107_port, nextA(42) => 
                           sigMatrix_6_106_port, nextA(41) => 
                           sigMatrix_6_105_port, nextA(40) => 
                           sigMatrix_6_104_port, nextA(39) => 
                           sigMatrix_6_103_port, nextA(38) => 
                           sigMatrix_6_102_port, nextA(37) => 
                           sigMatrix_6_101_port, nextA(36) => 
                           sigMatrix_6_100_port, nextA(35) => 
                           sigMatrix_6_99_port, nextA(34) => 
                           sigMatrix_6_98_port, nextA(33) => 
                           sigMatrix_6_97_port, nextA(32) => 
                           sigMatrix_6_96_port, nextA(31) => 
                           sigMatrix_6_95_port, nextA(30) => 
                           sigMatrix_6_94_port, nextA(29) => 
                           sigMatrix_6_93_port, nextA(28) => 
                           sigMatrix_6_92_port, nextA(27) => 
                           sigMatrix_6_91_port, nextA(26) => 
                           sigMatrix_6_90_port, nextA(25) => 
                           sigMatrix_6_89_port, nextA(24) => 
                           sigMatrix_6_88_port, nextA(23) => 
                           sigMatrix_6_87_port, nextA(22) => 
                           sigMatrix_6_86_port, nextA(21) => 
                           sigMatrix_6_85_port, nextA(20) => 
                           sigMatrix_6_84_port, nextA(19) => 
                           sigMatrix_6_83_port, nextA(18) => 
                           sigMatrix_6_82_port, nextA(17) => 
                           sigMatrix_6_81_port, nextA(16) => 
                           sigMatrix_6_80_port, nextA(15) => 
                           sigMatrix_6_79_port, nextA(14) => 
                           sigMatrix_6_78_port, nextA(13) => 
                           sigMatrix_6_77_port, nextA(12) => 
                           sigMatrix_6_76_port, nextA(11) => 
                           sigMatrix_6_75_port, nextA(10) => 
                           sigMatrix_6_74_port, nextA(9) => sigMatrix_6_73_port
                           , nextA(8) => sigMatrix_6_72_port, nextA(7) => 
                           sigMatrix_6_71_port, nextA(6) => sigMatrix_6_70_port
                           , nextA(5) => sigMatrix_6_69_port, nextA(4) => 
                           sigMatrix_6_68_port, nextA(3) => sigMatrix_6_67_port
                           , nextA(2) => sigMatrix_6_66_port, nextA(1) => 
                           sigMatrix_6_65_port, nextA(0) => n_3227, nextSum(63)
                           => sigMatrix_6_63_port, nextSum(62) => 
                           sigMatrix_6_62_port, nextSum(61) => 
                           sigMatrix_6_61_port, nextSum(60) => 
                           sigMatrix_6_60_port, nextSum(59) => 
                           sigMatrix_6_59_port, nextSum(58) => 
                           sigMatrix_6_58_port, nextSum(57) => 
                           sigMatrix_6_57_port, nextSum(56) => 
                           sigMatrix_6_56_port, nextSum(55) => 
                           sigMatrix_6_55_port, nextSum(54) => 
                           sigMatrix_6_54_port, nextSum(53) => 
                           sigMatrix_6_53_port, nextSum(52) => 
                           sigMatrix_6_52_port, nextSum(51) => 
                           sigMatrix_6_51_port, nextSum(50) => 
                           sigMatrix_6_50_port, nextSum(49) => 
                           sigMatrix_6_49_port, nextSum(48) => 
                           sigMatrix_6_48_port, nextSum(47) => 
                           sigMatrix_6_47_port, nextSum(46) => 
                           sigMatrix_6_46_port, nextSum(45) => 
                           sigMatrix_6_45_port, nextSum(44) => 
                           sigMatrix_6_44_port, nextSum(43) => 
                           sigMatrix_6_43_port, nextSum(42) => 
                           sigMatrix_6_42_port, nextSum(41) => 
                           sigMatrix_6_41_port, nextSum(40) => 
                           sigMatrix_6_40_port, nextSum(39) => 
                           sigMatrix_6_39_port, nextSum(38) => 
                           sigMatrix_6_38_port, nextSum(37) => 
                           sigMatrix_6_37_port, nextSum(36) => 
                           sigMatrix_6_36_port, nextSum(35) => 
                           sigMatrix_6_35_port, nextSum(34) => 
                           sigMatrix_6_34_port, nextSum(33) => 
                           sigMatrix_6_33_port, nextSum(32) => 
                           sigMatrix_6_32_port, nextSum(31) => 
                           sigMatrix_6_31_port, nextSum(30) => 
                           sigMatrix_6_30_port, nextSum(29) => 
                           sigMatrix_6_29_port, nextSum(28) => 
                           sigMatrix_6_28_port, nextSum(27) => 
                           sigMatrix_6_27_port, nextSum(26) => 
                           sigMatrix_6_26_port, nextSum(25) => 
                           sigMatrix_6_25_port, nextSum(24) => 
                           sigMatrix_6_24_port, nextSum(23) => 
                           sigMatrix_6_23_port, nextSum(22) => 
                           sigMatrix_6_22_port, nextSum(21) => 
                           sigMatrix_6_21_port, nextSum(20) => 
                           sigMatrix_6_20_port, nextSum(19) => 
                           sigMatrix_6_19_port, nextSum(18) => 
                           sigMatrix_6_18_port, nextSum(17) => 
                           sigMatrix_6_17_port, nextSum(16) => 
                           sigMatrix_6_16_port, nextSum(15) => 
                           sigMatrix_6_15_port, nextSum(14) => 
                           sigMatrix_6_14_port, nextSum(13) => 
                           sigMatrix_6_13_port, nextSum(12) => 
                           sigMatrix_6_12_port, nextSum(11) => 
                           sigMatrix_6_11_port, nextSum(10) => 
                           sigMatrix_6_10_port, nextSum(9) => 
                           sigMatrix_6_9_port, nextSum(8) => sigMatrix_6_8_port
                           , nextSum(7) => sigMatrix_6_7_port, nextSum(6) => 
                           sigMatrix_6_6_port, nextSum(5) => sigMatrix_6_5_port
                           , nextSum(4) => sigMatrix_6_4_port, nextSum(3) => 
                           sigMatrix_6_3_port, nextSum(2) => sigMatrix_6_2_port
                           , nextSum(1) => sigMatrix_6_1_port, nextSum(0) => 
                           sigMatrix_6_0_port);
   booth_mul_row_1_7 : booth_mul_row_N64_RADIX3_9 port map( prevA(63) => 
                           sigMatrix_6_127_port, prevA(62) => 
                           sigMatrix_6_126_port, prevA(61) => 
                           sigMatrix_6_125_port, prevA(60) => 
                           sigMatrix_6_124_port, prevA(59) => 
                           sigMatrix_6_123_port, prevA(58) => 
                           sigMatrix_6_122_port, prevA(57) => 
                           sigMatrix_6_121_port, prevA(56) => 
                           sigMatrix_6_120_port, prevA(55) => 
                           sigMatrix_6_119_port, prevA(54) => 
                           sigMatrix_6_118_port, prevA(53) => 
                           sigMatrix_6_117_port, prevA(52) => 
                           sigMatrix_6_116_port, prevA(51) => 
                           sigMatrix_6_115_port, prevA(50) => 
                           sigMatrix_6_114_port, prevA(49) => 
                           sigMatrix_6_113_port, prevA(48) => 
                           sigMatrix_6_112_port, prevA(47) => 
                           sigMatrix_6_111_port, prevA(46) => 
                           sigMatrix_6_110_port, prevA(45) => 
                           sigMatrix_6_109_port, prevA(44) => 
                           sigMatrix_6_108_port, prevA(43) => 
                           sigMatrix_6_107_port, prevA(42) => 
                           sigMatrix_6_106_port, prevA(41) => 
                           sigMatrix_6_105_port, prevA(40) => 
                           sigMatrix_6_104_port, prevA(39) => 
                           sigMatrix_6_103_port, prevA(38) => 
                           sigMatrix_6_102_port, prevA(37) => 
                           sigMatrix_6_101_port, prevA(36) => 
                           sigMatrix_6_100_port, prevA(35) => 
                           sigMatrix_6_99_port, prevA(34) => 
                           sigMatrix_6_98_port, prevA(33) => 
                           sigMatrix_6_97_port, prevA(32) => 
                           sigMatrix_6_96_port, prevA(31) => 
                           sigMatrix_6_95_port, prevA(30) => 
                           sigMatrix_6_94_port, prevA(29) => 
                           sigMatrix_6_93_port, prevA(28) => 
                           sigMatrix_6_92_port, prevA(27) => 
                           sigMatrix_6_91_port, prevA(26) => 
                           sigMatrix_6_90_port, prevA(25) => 
                           sigMatrix_6_89_port, prevA(24) => 
                           sigMatrix_6_88_port, prevA(23) => 
                           sigMatrix_6_87_port, prevA(22) => 
                           sigMatrix_6_86_port, prevA(21) => 
                           sigMatrix_6_85_port, prevA(20) => 
                           sigMatrix_6_84_port, prevA(19) => 
                           sigMatrix_6_83_port, prevA(18) => 
                           sigMatrix_6_82_port, prevA(17) => 
                           sigMatrix_6_81_port, prevA(16) => 
                           sigMatrix_6_80_port, prevA(15) => 
                           sigMatrix_6_79_port, prevA(14) => 
                           sigMatrix_6_78_port, prevA(13) => 
                           sigMatrix_6_77_port, prevA(12) => 
                           sigMatrix_6_76_port, prevA(11) => 
                           sigMatrix_6_75_port, prevA(10) => 
                           sigMatrix_6_74_port, prevA(9) => sigMatrix_6_73_port
                           , prevA(8) => sigMatrix_6_72_port, prevA(7) => 
                           sigMatrix_6_71_port, prevA(6) => sigMatrix_6_70_port
                           , prevA(5) => sigMatrix_6_69_port, prevA(4) => 
                           sigMatrix_6_68_port, prevA(3) => sigMatrix_6_67_port
                           , prevA(2) => sigMatrix_6_66_port, prevA(1) => 
                           sigMatrix_6_65_port, prevA(0) => n1, prevSum(63) => 
                           sigMatrix_6_63_port, prevSum(62) => 
                           sigMatrix_6_62_port, prevSum(61) => 
                           sigMatrix_6_61_port, prevSum(60) => 
                           sigMatrix_6_60_port, prevSum(59) => 
                           sigMatrix_6_59_port, prevSum(58) => 
                           sigMatrix_6_58_port, prevSum(57) => 
                           sigMatrix_6_57_port, prevSum(56) => 
                           sigMatrix_6_56_port, prevSum(55) => 
                           sigMatrix_6_55_port, prevSum(54) => 
                           sigMatrix_6_54_port, prevSum(53) => 
                           sigMatrix_6_53_port, prevSum(52) => 
                           sigMatrix_6_52_port, prevSum(51) => 
                           sigMatrix_6_51_port, prevSum(50) => 
                           sigMatrix_6_50_port, prevSum(49) => 
                           sigMatrix_6_49_port, prevSum(48) => 
                           sigMatrix_6_48_port, prevSum(47) => 
                           sigMatrix_6_47_port, prevSum(46) => 
                           sigMatrix_6_46_port, prevSum(45) => 
                           sigMatrix_6_45_port, prevSum(44) => 
                           sigMatrix_6_44_port, prevSum(43) => 
                           sigMatrix_6_43_port, prevSum(42) => 
                           sigMatrix_6_42_port, prevSum(41) => 
                           sigMatrix_6_41_port, prevSum(40) => 
                           sigMatrix_6_40_port, prevSum(39) => 
                           sigMatrix_6_39_port, prevSum(38) => 
                           sigMatrix_6_38_port, prevSum(37) => 
                           sigMatrix_6_37_port, prevSum(36) => 
                           sigMatrix_6_36_port, prevSum(35) => 
                           sigMatrix_6_35_port, prevSum(34) => 
                           sigMatrix_6_34_port, prevSum(33) => 
                           sigMatrix_6_33_port, prevSum(32) => 
                           sigMatrix_6_32_port, prevSum(31) => 
                           sigMatrix_6_31_port, prevSum(30) => 
                           sigMatrix_6_30_port, prevSum(29) => 
                           sigMatrix_6_29_port, prevSum(28) => 
                           sigMatrix_6_28_port, prevSum(27) => 
                           sigMatrix_6_27_port, prevSum(26) => 
                           sigMatrix_6_26_port, prevSum(25) => 
                           sigMatrix_6_25_port, prevSum(24) => 
                           sigMatrix_6_24_port, prevSum(23) => 
                           sigMatrix_6_23_port, prevSum(22) => 
                           sigMatrix_6_22_port, prevSum(21) => 
                           sigMatrix_6_21_port, prevSum(20) => 
                           sigMatrix_6_20_port, prevSum(19) => 
                           sigMatrix_6_19_port, prevSum(18) => 
                           sigMatrix_6_18_port, prevSum(17) => 
                           sigMatrix_6_17_port, prevSum(16) => 
                           sigMatrix_6_16_port, prevSum(15) => 
                           sigMatrix_6_15_port, prevSum(14) => 
                           sigMatrix_6_14_port, prevSum(13) => 
                           sigMatrix_6_13_port, prevSum(12) => 
                           sigMatrix_6_12_port, prevSum(11) => 
                           sigMatrix_6_11_port, prevSum(10) => 
                           sigMatrix_6_10_port, prevSum(9) => 
                           sigMatrix_6_9_port, prevSum(8) => sigMatrix_6_8_port
                           , prevSum(7) => sigMatrix_6_7_port, prevSum(6) => 
                           sigMatrix_6_6_port, prevSum(5) => sigMatrix_6_5_port
                           , prevSum(4) => sigMatrix_6_4_port, prevSum(3) => 
                           sigMatrix_6_3_port, prevSum(2) => sigMatrix_6_2_port
                           , prevSum(1) => sigMatrix_6_1_port, prevSum(0) => 
                           sigMatrix_6_0_port, encoderIn(2) => B(15), 
                           encoderIn(1) => B(14), encoderIn(0) => B(13), 
                           nextA(63) => sigMatrix_7_127_port, nextA(62) => 
                           sigMatrix_7_126_port, nextA(61) => 
                           sigMatrix_7_125_port, nextA(60) => 
                           sigMatrix_7_124_port, nextA(59) => 
                           sigMatrix_7_123_port, nextA(58) => 
                           sigMatrix_7_122_port, nextA(57) => 
                           sigMatrix_7_121_port, nextA(56) => 
                           sigMatrix_7_120_port, nextA(55) => 
                           sigMatrix_7_119_port, nextA(54) => 
                           sigMatrix_7_118_port, nextA(53) => 
                           sigMatrix_7_117_port, nextA(52) => 
                           sigMatrix_7_116_port, nextA(51) => 
                           sigMatrix_7_115_port, nextA(50) => 
                           sigMatrix_7_114_port, nextA(49) => 
                           sigMatrix_7_113_port, nextA(48) => 
                           sigMatrix_7_112_port, nextA(47) => 
                           sigMatrix_7_111_port, nextA(46) => 
                           sigMatrix_7_110_port, nextA(45) => 
                           sigMatrix_7_109_port, nextA(44) => 
                           sigMatrix_7_108_port, nextA(43) => 
                           sigMatrix_7_107_port, nextA(42) => 
                           sigMatrix_7_106_port, nextA(41) => 
                           sigMatrix_7_105_port, nextA(40) => 
                           sigMatrix_7_104_port, nextA(39) => 
                           sigMatrix_7_103_port, nextA(38) => 
                           sigMatrix_7_102_port, nextA(37) => 
                           sigMatrix_7_101_port, nextA(36) => 
                           sigMatrix_7_100_port, nextA(35) => 
                           sigMatrix_7_99_port, nextA(34) => 
                           sigMatrix_7_98_port, nextA(33) => 
                           sigMatrix_7_97_port, nextA(32) => 
                           sigMatrix_7_96_port, nextA(31) => 
                           sigMatrix_7_95_port, nextA(30) => 
                           sigMatrix_7_94_port, nextA(29) => 
                           sigMatrix_7_93_port, nextA(28) => 
                           sigMatrix_7_92_port, nextA(27) => 
                           sigMatrix_7_91_port, nextA(26) => 
                           sigMatrix_7_90_port, nextA(25) => 
                           sigMatrix_7_89_port, nextA(24) => 
                           sigMatrix_7_88_port, nextA(23) => 
                           sigMatrix_7_87_port, nextA(22) => 
                           sigMatrix_7_86_port, nextA(21) => 
                           sigMatrix_7_85_port, nextA(20) => 
                           sigMatrix_7_84_port, nextA(19) => 
                           sigMatrix_7_83_port, nextA(18) => 
                           sigMatrix_7_82_port, nextA(17) => 
                           sigMatrix_7_81_port, nextA(16) => 
                           sigMatrix_7_80_port, nextA(15) => 
                           sigMatrix_7_79_port, nextA(14) => 
                           sigMatrix_7_78_port, nextA(13) => 
                           sigMatrix_7_77_port, nextA(12) => 
                           sigMatrix_7_76_port, nextA(11) => 
                           sigMatrix_7_75_port, nextA(10) => 
                           sigMatrix_7_74_port, nextA(9) => sigMatrix_7_73_port
                           , nextA(8) => sigMatrix_7_72_port, nextA(7) => 
                           sigMatrix_7_71_port, nextA(6) => sigMatrix_7_70_port
                           , nextA(5) => sigMatrix_7_69_port, nextA(4) => 
                           sigMatrix_7_68_port, nextA(3) => sigMatrix_7_67_port
                           , nextA(2) => sigMatrix_7_66_port, nextA(1) => 
                           sigMatrix_7_65_port, nextA(0) => n_3228, nextSum(63)
                           => sigMatrix_7_63_port, nextSum(62) => 
                           sigMatrix_7_62_port, nextSum(61) => 
                           sigMatrix_7_61_port, nextSum(60) => 
                           sigMatrix_7_60_port, nextSum(59) => 
                           sigMatrix_7_59_port, nextSum(58) => 
                           sigMatrix_7_58_port, nextSum(57) => 
                           sigMatrix_7_57_port, nextSum(56) => 
                           sigMatrix_7_56_port, nextSum(55) => 
                           sigMatrix_7_55_port, nextSum(54) => 
                           sigMatrix_7_54_port, nextSum(53) => 
                           sigMatrix_7_53_port, nextSum(52) => 
                           sigMatrix_7_52_port, nextSum(51) => 
                           sigMatrix_7_51_port, nextSum(50) => 
                           sigMatrix_7_50_port, nextSum(49) => 
                           sigMatrix_7_49_port, nextSum(48) => 
                           sigMatrix_7_48_port, nextSum(47) => 
                           sigMatrix_7_47_port, nextSum(46) => 
                           sigMatrix_7_46_port, nextSum(45) => 
                           sigMatrix_7_45_port, nextSum(44) => 
                           sigMatrix_7_44_port, nextSum(43) => 
                           sigMatrix_7_43_port, nextSum(42) => 
                           sigMatrix_7_42_port, nextSum(41) => 
                           sigMatrix_7_41_port, nextSum(40) => 
                           sigMatrix_7_40_port, nextSum(39) => 
                           sigMatrix_7_39_port, nextSum(38) => 
                           sigMatrix_7_38_port, nextSum(37) => 
                           sigMatrix_7_37_port, nextSum(36) => 
                           sigMatrix_7_36_port, nextSum(35) => 
                           sigMatrix_7_35_port, nextSum(34) => 
                           sigMatrix_7_34_port, nextSum(33) => 
                           sigMatrix_7_33_port, nextSum(32) => 
                           sigMatrix_7_32_port, nextSum(31) => 
                           sigMatrix_7_31_port, nextSum(30) => 
                           sigMatrix_7_30_port, nextSum(29) => 
                           sigMatrix_7_29_port, nextSum(28) => 
                           sigMatrix_7_28_port, nextSum(27) => 
                           sigMatrix_7_27_port, nextSum(26) => 
                           sigMatrix_7_26_port, nextSum(25) => 
                           sigMatrix_7_25_port, nextSum(24) => 
                           sigMatrix_7_24_port, nextSum(23) => 
                           sigMatrix_7_23_port, nextSum(22) => 
                           sigMatrix_7_22_port, nextSum(21) => 
                           sigMatrix_7_21_port, nextSum(20) => 
                           sigMatrix_7_20_port, nextSum(19) => 
                           sigMatrix_7_19_port, nextSum(18) => 
                           sigMatrix_7_18_port, nextSum(17) => 
                           sigMatrix_7_17_port, nextSum(16) => 
                           sigMatrix_7_16_port, nextSum(15) => 
                           sigMatrix_7_15_port, nextSum(14) => 
                           sigMatrix_7_14_port, nextSum(13) => 
                           sigMatrix_7_13_port, nextSum(12) => 
                           sigMatrix_7_12_port, nextSum(11) => 
                           sigMatrix_7_11_port, nextSum(10) => 
                           sigMatrix_7_10_port, nextSum(9) => 
                           sigMatrix_7_9_port, nextSum(8) => sigMatrix_7_8_port
                           , nextSum(7) => sigMatrix_7_7_port, nextSum(6) => 
                           sigMatrix_7_6_port, nextSum(5) => sigMatrix_7_5_port
                           , nextSum(4) => sigMatrix_7_4_port, nextSum(3) => 
                           sigMatrix_7_3_port, nextSum(2) => sigMatrix_7_2_port
                           , nextSum(1) => sigMatrix_7_1_port, nextSum(0) => 
                           sigMatrix_7_0_port);
   booth_mul_row_1_8 : booth_mul_row_N64_RADIX3_8 port map( prevA(63) => 
                           sigMatrix_7_127_port, prevA(62) => 
                           sigMatrix_7_126_port, prevA(61) => 
                           sigMatrix_7_125_port, prevA(60) => 
                           sigMatrix_7_124_port, prevA(59) => 
                           sigMatrix_7_123_port, prevA(58) => 
                           sigMatrix_7_122_port, prevA(57) => 
                           sigMatrix_7_121_port, prevA(56) => 
                           sigMatrix_7_120_port, prevA(55) => 
                           sigMatrix_7_119_port, prevA(54) => 
                           sigMatrix_7_118_port, prevA(53) => 
                           sigMatrix_7_117_port, prevA(52) => 
                           sigMatrix_7_116_port, prevA(51) => 
                           sigMatrix_7_115_port, prevA(50) => 
                           sigMatrix_7_114_port, prevA(49) => 
                           sigMatrix_7_113_port, prevA(48) => 
                           sigMatrix_7_112_port, prevA(47) => 
                           sigMatrix_7_111_port, prevA(46) => 
                           sigMatrix_7_110_port, prevA(45) => 
                           sigMatrix_7_109_port, prevA(44) => 
                           sigMatrix_7_108_port, prevA(43) => 
                           sigMatrix_7_107_port, prevA(42) => 
                           sigMatrix_7_106_port, prevA(41) => 
                           sigMatrix_7_105_port, prevA(40) => 
                           sigMatrix_7_104_port, prevA(39) => 
                           sigMatrix_7_103_port, prevA(38) => 
                           sigMatrix_7_102_port, prevA(37) => 
                           sigMatrix_7_101_port, prevA(36) => 
                           sigMatrix_7_100_port, prevA(35) => 
                           sigMatrix_7_99_port, prevA(34) => 
                           sigMatrix_7_98_port, prevA(33) => 
                           sigMatrix_7_97_port, prevA(32) => 
                           sigMatrix_7_96_port, prevA(31) => 
                           sigMatrix_7_95_port, prevA(30) => 
                           sigMatrix_7_94_port, prevA(29) => 
                           sigMatrix_7_93_port, prevA(28) => 
                           sigMatrix_7_92_port, prevA(27) => 
                           sigMatrix_7_91_port, prevA(26) => 
                           sigMatrix_7_90_port, prevA(25) => 
                           sigMatrix_7_89_port, prevA(24) => 
                           sigMatrix_7_88_port, prevA(23) => 
                           sigMatrix_7_87_port, prevA(22) => 
                           sigMatrix_7_86_port, prevA(21) => 
                           sigMatrix_7_85_port, prevA(20) => 
                           sigMatrix_7_84_port, prevA(19) => 
                           sigMatrix_7_83_port, prevA(18) => 
                           sigMatrix_7_82_port, prevA(17) => 
                           sigMatrix_7_81_port, prevA(16) => 
                           sigMatrix_7_80_port, prevA(15) => 
                           sigMatrix_7_79_port, prevA(14) => 
                           sigMatrix_7_78_port, prevA(13) => 
                           sigMatrix_7_77_port, prevA(12) => 
                           sigMatrix_7_76_port, prevA(11) => 
                           sigMatrix_7_75_port, prevA(10) => 
                           sigMatrix_7_74_port, prevA(9) => sigMatrix_7_73_port
                           , prevA(8) => sigMatrix_7_72_port, prevA(7) => 
                           sigMatrix_7_71_port, prevA(6) => sigMatrix_7_70_port
                           , prevA(5) => sigMatrix_7_69_port, prevA(4) => 
                           sigMatrix_7_68_port, prevA(3) => sigMatrix_7_67_port
                           , prevA(2) => sigMatrix_7_66_port, prevA(1) => 
                           sigMatrix_7_65_port, prevA(0) => n1, prevSum(63) => 
                           sigMatrix_7_63_port, prevSum(62) => 
                           sigMatrix_7_62_port, prevSum(61) => 
                           sigMatrix_7_61_port, prevSum(60) => 
                           sigMatrix_7_60_port, prevSum(59) => 
                           sigMatrix_7_59_port, prevSum(58) => 
                           sigMatrix_7_58_port, prevSum(57) => 
                           sigMatrix_7_57_port, prevSum(56) => 
                           sigMatrix_7_56_port, prevSum(55) => 
                           sigMatrix_7_55_port, prevSum(54) => 
                           sigMatrix_7_54_port, prevSum(53) => 
                           sigMatrix_7_53_port, prevSum(52) => 
                           sigMatrix_7_52_port, prevSum(51) => 
                           sigMatrix_7_51_port, prevSum(50) => 
                           sigMatrix_7_50_port, prevSum(49) => 
                           sigMatrix_7_49_port, prevSum(48) => 
                           sigMatrix_7_48_port, prevSum(47) => 
                           sigMatrix_7_47_port, prevSum(46) => 
                           sigMatrix_7_46_port, prevSum(45) => 
                           sigMatrix_7_45_port, prevSum(44) => 
                           sigMatrix_7_44_port, prevSum(43) => 
                           sigMatrix_7_43_port, prevSum(42) => 
                           sigMatrix_7_42_port, prevSum(41) => 
                           sigMatrix_7_41_port, prevSum(40) => 
                           sigMatrix_7_40_port, prevSum(39) => 
                           sigMatrix_7_39_port, prevSum(38) => 
                           sigMatrix_7_38_port, prevSum(37) => 
                           sigMatrix_7_37_port, prevSum(36) => 
                           sigMatrix_7_36_port, prevSum(35) => 
                           sigMatrix_7_35_port, prevSum(34) => 
                           sigMatrix_7_34_port, prevSum(33) => 
                           sigMatrix_7_33_port, prevSum(32) => 
                           sigMatrix_7_32_port, prevSum(31) => 
                           sigMatrix_7_31_port, prevSum(30) => 
                           sigMatrix_7_30_port, prevSum(29) => 
                           sigMatrix_7_29_port, prevSum(28) => 
                           sigMatrix_7_28_port, prevSum(27) => 
                           sigMatrix_7_27_port, prevSum(26) => 
                           sigMatrix_7_26_port, prevSum(25) => 
                           sigMatrix_7_25_port, prevSum(24) => 
                           sigMatrix_7_24_port, prevSum(23) => 
                           sigMatrix_7_23_port, prevSum(22) => 
                           sigMatrix_7_22_port, prevSum(21) => 
                           sigMatrix_7_21_port, prevSum(20) => 
                           sigMatrix_7_20_port, prevSum(19) => 
                           sigMatrix_7_19_port, prevSum(18) => 
                           sigMatrix_7_18_port, prevSum(17) => 
                           sigMatrix_7_17_port, prevSum(16) => 
                           sigMatrix_7_16_port, prevSum(15) => 
                           sigMatrix_7_15_port, prevSum(14) => 
                           sigMatrix_7_14_port, prevSum(13) => 
                           sigMatrix_7_13_port, prevSum(12) => 
                           sigMatrix_7_12_port, prevSum(11) => 
                           sigMatrix_7_11_port, prevSum(10) => 
                           sigMatrix_7_10_port, prevSum(9) => 
                           sigMatrix_7_9_port, prevSum(8) => sigMatrix_7_8_port
                           , prevSum(7) => sigMatrix_7_7_port, prevSum(6) => 
                           sigMatrix_7_6_port, prevSum(5) => sigMatrix_7_5_port
                           , prevSum(4) => sigMatrix_7_4_port, prevSum(3) => 
                           sigMatrix_7_3_port, prevSum(2) => sigMatrix_7_2_port
                           , prevSum(1) => sigMatrix_7_1_port, prevSum(0) => 
                           sigMatrix_7_0_port, encoderIn(2) => B(17), 
                           encoderIn(1) => B(16), encoderIn(0) => B(15), 
                           nextA(63) => sigMatrix_8_127_port, nextA(62) => 
                           sigMatrix_8_126_port, nextA(61) => 
                           sigMatrix_8_125_port, nextA(60) => 
                           sigMatrix_8_124_port, nextA(59) => 
                           sigMatrix_8_123_port, nextA(58) => 
                           sigMatrix_8_122_port, nextA(57) => 
                           sigMatrix_8_121_port, nextA(56) => 
                           sigMatrix_8_120_port, nextA(55) => 
                           sigMatrix_8_119_port, nextA(54) => 
                           sigMatrix_8_118_port, nextA(53) => 
                           sigMatrix_8_117_port, nextA(52) => 
                           sigMatrix_8_116_port, nextA(51) => 
                           sigMatrix_8_115_port, nextA(50) => 
                           sigMatrix_8_114_port, nextA(49) => 
                           sigMatrix_8_113_port, nextA(48) => 
                           sigMatrix_8_112_port, nextA(47) => 
                           sigMatrix_8_111_port, nextA(46) => 
                           sigMatrix_8_110_port, nextA(45) => 
                           sigMatrix_8_109_port, nextA(44) => 
                           sigMatrix_8_108_port, nextA(43) => 
                           sigMatrix_8_107_port, nextA(42) => 
                           sigMatrix_8_106_port, nextA(41) => 
                           sigMatrix_8_105_port, nextA(40) => 
                           sigMatrix_8_104_port, nextA(39) => 
                           sigMatrix_8_103_port, nextA(38) => 
                           sigMatrix_8_102_port, nextA(37) => 
                           sigMatrix_8_101_port, nextA(36) => 
                           sigMatrix_8_100_port, nextA(35) => 
                           sigMatrix_8_99_port, nextA(34) => 
                           sigMatrix_8_98_port, nextA(33) => 
                           sigMatrix_8_97_port, nextA(32) => 
                           sigMatrix_8_96_port, nextA(31) => 
                           sigMatrix_8_95_port, nextA(30) => 
                           sigMatrix_8_94_port, nextA(29) => 
                           sigMatrix_8_93_port, nextA(28) => 
                           sigMatrix_8_92_port, nextA(27) => 
                           sigMatrix_8_91_port, nextA(26) => 
                           sigMatrix_8_90_port, nextA(25) => 
                           sigMatrix_8_89_port, nextA(24) => 
                           sigMatrix_8_88_port, nextA(23) => 
                           sigMatrix_8_87_port, nextA(22) => 
                           sigMatrix_8_86_port, nextA(21) => 
                           sigMatrix_8_85_port, nextA(20) => 
                           sigMatrix_8_84_port, nextA(19) => 
                           sigMatrix_8_83_port, nextA(18) => 
                           sigMatrix_8_82_port, nextA(17) => 
                           sigMatrix_8_81_port, nextA(16) => 
                           sigMatrix_8_80_port, nextA(15) => 
                           sigMatrix_8_79_port, nextA(14) => 
                           sigMatrix_8_78_port, nextA(13) => 
                           sigMatrix_8_77_port, nextA(12) => 
                           sigMatrix_8_76_port, nextA(11) => 
                           sigMatrix_8_75_port, nextA(10) => 
                           sigMatrix_8_74_port, nextA(9) => sigMatrix_8_73_port
                           , nextA(8) => sigMatrix_8_72_port, nextA(7) => 
                           sigMatrix_8_71_port, nextA(6) => sigMatrix_8_70_port
                           , nextA(5) => sigMatrix_8_69_port, nextA(4) => 
                           sigMatrix_8_68_port, nextA(3) => sigMatrix_8_67_port
                           , nextA(2) => sigMatrix_8_66_port, nextA(1) => 
                           sigMatrix_8_65_port, nextA(0) => n_3229, nextSum(63)
                           => sigMatrix_8_63_port, nextSum(62) => 
                           sigMatrix_8_62_port, nextSum(61) => 
                           sigMatrix_8_61_port, nextSum(60) => 
                           sigMatrix_8_60_port, nextSum(59) => 
                           sigMatrix_8_59_port, nextSum(58) => 
                           sigMatrix_8_58_port, nextSum(57) => 
                           sigMatrix_8_57_port, nextSum(56) => 
                           sigMatrix_8_56_port, nextSum(55) => 
                           sigMatrix_8_55_port, nextSum(54) => 
                           sigMatrix_8_54_port, nextSum(53) => 
                           sigMatrix_8_53_port, nextSum(52) => 
                           sigMatrix_8_52_port, nextSum(51) => 
                           sigMatrix_8_51_port, nextSum(50) => 
                           sigMatrix_8_50_port, nextSum(49) => 
                           sigMatrix_8_49_port, nextSum(48) => 
                           sigMatrix_8_48_port, nextSum(47) => 
                           sigMatrix_8_47_port, nextSum(46) => 
                           sigMatrix_8_46_port, nextSum(45) => 
                           sigMatrix_8_45_port, nextSum(44) => 
                           sigMatrix_8_44_port, nextSum(43) => 
                           sigMatrix_8_43_port, nextSum(42) => 
                           sigMatrix_8_42_port, nextSum(41) => 
                           sigMatrix_8_41_port, nextSum(40) => 
                           sigMatrix_8_40_port, nextSum(39) => 
                           sigMatrix_8_39_port, nextSum(38) => 
                           sigMatrix_8_38_port, nextSum(37) => 
                           sigMatrix_8_37_port, nextSum(36) => 
                           sigMatrix_8_36_port, nextSum(35) => 
                           sigMatrix_8_35_port, nextSum(34) => 
                           sigMatrix_8_34_port, nextSum(33) => 
                           sigMatrix_8_33_port, nextSum(32) => 
                           sigMatrix_8_32_port, nextSum(31) => 
                           sigMatrix_8_31_port, nextSum(30) => 
                           sigMatrix_8_30_port, nextSum(29) => 
                           sigMatrix_8_29_port, nextSum(28) => 
                           sigMatrix_8_28_port, nextSum(27) => 
                           sigMatrix_8_27_port, nextSum(26) => 
                           sigMatrix_8_26_port, nextSum(25) => 
                           sigMatrix_8_25_port, nextSum(24) => 
                           sigMatrix_8_24_port, nextSum(23) => 
                           sigMatrix_8_23_port, nextSum(22) => 
                           sigMatrix_8_22_port, nextSum(21) => 
                           sigMatrix_8_21_port, nextSum(20) => 
                           sigMatrix_8_20_port, nextSum(19) => 
                           sigMatrix_8_19_port, nextSum(18) => 
                           sigMatrix_8_18_port, nextSum(17) => 
                           sigMatrix_8_17_port, nextSum(16) => 
                           sigMatrix_8_16_port, nextSum(15) => 
                           sigMatrix_8_15_port, nextSum(14) => 
                           sigMatrix_8_14_port, nextSum(13) => 
                           sigMatrix_8_13_port, nextSum(12) => 
                           sigMatrix_8_12_port, nextSum(11) => 
                           sigMatrix_8_11_port, nextSum(10) => 
                           sigMatrix_8_10_port, nextSum(9) => 
                           sigMatrix_8_9_port, nextSum(8) => sigMatrix_8_8_port
                           , nextSum(7) => sigMatrix_8_7_port, nextSum(6) => 
                           sigMatrix_8_6_port, nextSum(5) => sigMatrix_8_5_port
                           , nextSum(4) => sigMatrix_8_4_port, nextSum(3) => 
                           sigMatrix_8_3_port, nextSum(2) => sigMatrix_8_2_port
                           , nextSum(1) => sigMatrix_8_1_port, nextSum(0) => 
                           sigMatrix_8_0_port);
   booth_mul_row_1_9 : booth_mul_row_N64_RADIX3_7 port map( prevA(63) => 
                           sigMatrix_8_127_port, prevA(62) => 
                           sigMatrix_8_126_port, prevA(61) => 
                           sigMatrix_8_125_port, prevA(60) => 
                           sigMatrix_8_124_port, prevA(59) => 
                           sigMatrix_8_123_port, prevA(58) => 
                           sigMatrix_8_122_port, prevA(57) => 
                           sigMatrix_8_121_port, prevA(56) => 
                           sigMatrix_8_120_port, prevA(55) => 
                           sigMatrix_8_119_port, prevA(54) => 
                           sigMatrix_8_118_port, prevA(53) => 
                           sigMatrix_8_117_port, prevA(52) => 
                           sigMatrix_8_116_port, prevA(51) => 
                           sigMatrix_8_115_port, prevA(50) => 
                           sigMatrix_8_114_port, prevA(49) => 
                           sigMatrix_8_113_port, prevA(48) => 
                           sigMatrix_8_112_port, prevA(47) => 
                           sigMatrix_8_111_port, prevA(46) => 
                           sigMatrix_8_110_port, prevA(45) => 
                           sigMatrix_8_109_port, prevA(44) => 
                           sigMatrix_8_108_port, prevA(43) => 
                           sigMatrix_8_107_port, prevA(42) => 
                           sigMatrix_8_106_port, prevA(41) => 
                           sigMatrix_8_105_port, prevA(40) => 
                           sigMatrix_8_104_port, prevA(39) => 
                           sigMatrix_8_103_port, prevA(38) => 
                           sigMatrix_8_102_port, prevA(37) => 
                           sigMatrix_8_101_port, prevA(36) => 
                           sigMatrix_8_100_port, prevA(35) => 
                           sigMatrix_8_99_port, prevA(34) => 
                           sigMatrix_8_98_port, prevA(33) => 
                           sigMatrix_8_97_port, prevA(32) => 
                           sigMatrix_8_96_port, prevA(31) => 
                           sigMatrix_8_95_port, prevA(30) => 
                           sigMatrix_8_94_port, prevA(29) => 
                           sigMatrix_8_93_port, prevA(28) => 
                           sigMatrix_8_92_port, prevA(27) => 
                           sigMatrix_8_91_port, prevA(26) => 
                           sigMatrix_8_90_port, prevA(25) => 
                           sigMatrix_8_89_port, prevA(24) => 
                           sigMatrix_8_88_port, prevA(23) => 
                           sigMatrix_8_87_port, prevA(22) => 
                           sigMatrix_8_86_port, prevA(21) => 
                           sigMatrix_8_85_port, prevA(20) => 
                           sigMatrix_8_84_port, prevA(19) => 
                           sigMatrix_8_83_port, prevA(18) => 
                           sigMatrix_8_82_port, prevA(17) => 
                           sigMatrix_8_81_port, prevA(16) => 
                           sigMatrix_8_80_port, prevA(15) => 
                           sigMatrix_8_79_port, prevA(14) => 
                           sigMatrix_8_78_port, prevA(13) => 
                           sigMatrix_8_77_port, prevA(12) => 
                           sigMatrix_8_76_port, prevA(11) => 
                           sigMatrix_8_75_port, prevA(10) => 
                           sigMatrix_8_74_port, prevA(9) => sigMatrix_8_73_port
                           , prevA(8) => sigMatrix_8_72_port, prevA(7) => 
                           sigMatrix_8_71_port, prevA(6) => sigMatrix_8_70_port
                           , prevA(5) => sigMatrix_8_69_port, prevA(4) => 
                           sigMatrix_8_68_port, prevA(3) => sigMatrix_8_67_port
                           , prevA(2) => sigMatrix_8_66_port, prevA(1) => 
                           sigMatrix_8_65_port, prevA(0) => n1, prevSum(63) => 
                           sigMatrix_8_63_port, prevSum(62) => 
                           sigMatrix_8_62_port, prevSum(61) => 
                           sigMatrix_8_61_port, prevSum(60) => 
                           sigMatrix_8_60_port, prevSum(59) => 
                           sigMatrix_8_59_port, prevSum(58) => 
                           sigMatrix_8_58_port, prevSum(57) => 
                           sigMatrix_8_57_port, prevSum(56) => 
                           sigMatrix_8_56_port, prevSum(55) => 
                           sigMatrix_8_55_port, prevSum(54) => 
                           sigMatrix_8_54_port, prevSum(53) => 
                           sigMatrix_8_53_port, prevSum(52) => 
                           sigMatrix_8_52_port, prevSum(51) => 
                           sigMatrix_8_51_port, prevSum(50) => 
                           sigMatrix_8_50_port, prevSum(49) => 
                           sigMatrix_8_49_port, prevSum(48) => 
                           sigMatrix_8_48_port, prevSum(47) => 
                           sigMatrix_8_47_port, prevSum(46) => 
                           sigMatrix_8_46_port, prevSum(45) => 
                           sigMatrix_8_45_port, prevSum(44) => 
                           sigMatrix_8_44_port, prevSum(43) => 
                           sigMatrix_8_43_port, prevSum(42) => 
                           sigMatrix_8_42_port, prevSum(41) => 
                           sigMatrix_8_41_port, prevSum(40) => 
                           sigMatrix_8_40_port, prevSum(39) => 
                           sigMatrix_8_39_port, prevSum(38) => 
                           sigMatrix_8_38_port, prevSum(37) => 
                           sigMatrix_8_37_port, prevSum(36) => 
                           sigMatrix_8_36_port, prevSum(35) => 
                           sigMatrix_8_35_port, prevSum(34) => 
                           sigMatrix_8_34_port, prevSum(33) => 
                           sigMatrix_8_33_port, prevSum(32) => 
                           sigMatrix_8_32_port, prevSum(31) => 
                           sigMatrix_8_31_port, prevSum(30) => 
                           sigMatrix_8_30_port, prevSum(29) => 
                           sigMatrix_8_29_port, prevSum(28) => 
                           sigMatrix_8_28_port, prevSum(27) => 
                           sigMatrix_8_27_port, prevSum(26) => 
                           sigMatrix_8_26_port, prevSum(25) => 
                           sigMatrix_8_25_port, prevSum(24) => 
                           sigMatrix_8_24_port, prevSum(23) => 
                           sigMatrix_8_23_port, prevSum(22) => 
                           sigMatrix_8_22_port, prevSum(21) => 
                           sigMatrix_8_21_port, prevSum(20) => 
                           sigMatrix_8_20_port, prevSum(19) => 
                           sigMatrix_8_19_port, prevSum(18) => 
                           sigMatrix_8_18_port, prevSum(17) => 
                           sigMatrix_8_17_port, prevSum(16) => 
                           sigMatrix_8_16_port, prevSum(15) => 
                           sigMatrix_8_15_port, prevSum(14) => 
                           sigMatrix_8_14_port, prevSum(13) => 
                           sigMatrix_8_13_port, prevSum(12) => 
                           sigMatrix_8_12_port, prevSum(11) => 
                           sigMatrix_8_11_port, prevSum(10) => 
                           sigMatrix_8_10_port, prevSum(9) => 
                           sigMatrix_8_9_port, prevSum(8) => sigMatrix_8_8_port
                           , prevSum(7) => sigMatrix_8_7_port, prevSum(6) => 
                           sigMatrix_8_6_port, prevSum(5) => sigMatrix_8_5_port
                           , prevSum(4) => sigMatrix_8_4_port, prevSum(3) => 
                           sigMatrix_8_3_port, prevSum(2) => sigMatrix_8_2_port
                           , prevSum(1) => sigMatrix_8_1_port, prevSum(0) => 
                           sigMatrix_8_0_port, encoderIn(2) => B(19), 
                           encoderIn(1) => B(18), encoderIn(0) => B(17), 
                           nextA(63) => sigMatrix_9_127_port, nextA(62) => 
                           sigMatrix_9_126_port, nextA(61) => 
                           sigMatrix_9_125_port, nextA(60) => 
                           sigMatrix_9_124_port, nextA(59) => 
                           sigMatrix_9_123_port, nextA(58) => 
                           sigMatrix_9_122_port, nextA(57) => 
                           sigMatrix_9_121_port, nextA(56) => 
                           sigMatrix_9_120_port, nextA(55) => 
                           sigMatrix_9_119_port, nextA(54) => 
                           sigMatrix_9_118_port, nextA(53) => 
                           sigMatrix_9_117_port, nextA(52) => 
                           sigMatrix_9_116_port, nextA(51) => 
                           sigMatrix_9_115_port, nextA(50) => 
                           sigMatrix_9_114_port, nextA(49) => 
                           sigMatrix_9_113_port, nextA(48) => 
                           sigMatrix_9_112_port, nextA(47) => 
                           sigMatrix_9_111_port, nextA(46) => 
                           sigMatrix_9_110_port, nextA(45) => 
                           sigMatrix_9_109_port, nextA(44) => 
                           sigMatrix_9_108_port, nextA(43) => 
                           sigMatrix_9_107_port, nextA(42) => 
                           sigMatrix_9_106_port, nextA(41) => 
                           sigMatrix_9_105_port, nextA(40) => 
                           sigMatrix_9_104_port, nextA(39) => 
                           sigMatrix_9_103_port, nextA(38) => 
                           sigMatrix_9_102_port, nextA(37) => 
                           sigMatrix_9_101_port, nextA(36) => 
                           sigMatrix_9_100_port, nextA(35) => 
                           sigMatrix_9_99_port, nextA(34) => 
                           sigMatrix_9_98_port, nextA(33) => 
                           sigMatrix_9_97_port, nextA(32) => 
                           sigMatrix_9_96_port, nextA(31) => 
                           sigMatrix_9_95_port, nextA(30) => 
                           sigMatrix_9_94_port, nextA(29) => 
                           sigMatrix_9_93_port, nextA(28) => 
                           sigMatrix_9_92_port, nextA(27) => 
                           sigMatrix_9_91_port, nextA(26) => 
                           sigMatrix_9_90_port, nextA(25) => 
                           sigMatrix_9_89_port, nextA(24) => 
                           sigMatrix_9_88_port, nextA(23) => 
                           sigMatrix_9_87_port, nextA(22) => 
                           sigMatrix_9_86_port, nextA(21) => 
                           sigMatrix_9_85_port, nextA(20) => 
                           sigMatrix_9_84_port, nextA(19) => 
                           sigMatrix_9_83_port, nextA(18) => 
                           sigMatrix_9_82_port, nextA(17) => 
                           sigMatrix_9_81_port, nextA(16) => 
                           sigMatrix_9_80_port, nextA(15) => 
                           sigMatrix_9_79_port, nextA(14) => 
                           sigMatrix_9_78_port, nextA(13) => 
                           sigMatrix_9_77_port, nextA(12) => 
                           sigMatrix_9_76_port, nextA(11) => 
                           sigMatrix_9_75_port, nextA(10) => 
                           sigMatrix_9_74_port, nextA(9) => sigMatrix_9_73_port
                           , nextA(8) => sigMatrix_9_72_port, nextA(7) => 
                           sigMatrix_9_71_port, nextA(6) => sigMatrix_9_70_port
                           , nextA(5) => sigMatrix_9_69_port, nextA(4) => 
                           sigMatrix_9_68_port, nextA(3) => sigMatrix_9_67_port
                           , nextA(2) => sigMatrix_9_66_port, nextA(1) => 
                           sigMatrix_9_65_port, nextA(0) => n_3230, nextSum(63)
                           => sigMatrix_9_63_port, nextSum(62) => 
                           sigMatrix_9_62_port, nextSum(61) => 
                           sigMatrix_9_61_port, nextSum(60) => 
                           sigMatrix_9_60_port, nextSum(59) => 
                           sigMatrix_9_59_port, nextSum(58) => 
                           sigMatrix_9_58_port, nextSum(57) => 
                           sigMatrix_9_57_port, nextSum(56) => 
                           sigMatrix_9_56_port, nextSum(55) => 
                           sigMatrix_9_55_port, nextSum(54) => 
                           sigMatrix_9_54_port, nextSum(53) => 
                           sigMatrix_9_53_port, nextSum(52) => 
                           sigMatrix_9_52_port, nextSum(51) => 
                           sigMatrix_9_51_port, nextSum(50) => 
                           sigMatrix_9_50_port, nextSum(49) => 
                           sigMatrix_9_49_port, nextSum(48) => 
                           sigMatrix_9_48_port, nextSum(47) => 
                           sigMatrix_9_47_port, nextSum(46) => 
                           sigMatrix_9_46_port, nextSum(45) => 
                           sigMatrix_9_45_port, nextSum(44) => 
                           sigMatrix_9_44_port, nextSum(43) => 
                           sigMatrix_9_43_port, nextSum(42) => 
                           sigMatrix_9_42_port, nextSum(41) => 
                           sigMatrix_9_41_port, nextSum(40) => 
                           sigMatrix_9_40_port, nextSum(39) => 
                           sigMatrix_9_39_port, nextSum(38) => 
                           sigMatrix_9_38_port, nextSum(37) => 
                           sigMatrix_9_37_port, nextSum(36) => 
                           sigMatrix_9_36_port, nextSum(35) => 
                           sigMatrix_9_35_port, nextSum(34) => 
                           sigMatrix_9_34_port, nextSum(33) => 
                           sigMatrix_9_33_port, nextSum(32) => 
                           sigMatrix_9_32_port, nextSum(31) => 
                           sigMatrix_9_31_port, nextSum(30) => 
                           sigMatrix_9_30_port, nextSum(29) => 
                           sigMatrix_9_29_port, nextSum(28) => 
                           sigMatrix_9_28_port, nextSum(27) => 
                           sigMatrix_9_27_port, nextSum(26) => 
                           sigMatrix_9_26_port, nextSum(25) => 
                           sigMatrix_9_25_port, nextSum(24) => 
                           sigMatrix_9_24_port, nextSum(23) => 
                           sigMatrix_9_23_port, nextSum(22) => 
                           sigMatrix_9_22_port, nextSum(21) => 
                           sigMatrix_9_21_port, nextSum(20) => 
                           sigMatrix_9_20_port, nextSum(19) => 
                           sigMatrix_9_19_port, nextSum(18) => 
                           sigMatrix_9_18_port, nextSum(17) => 
                           sigMatrix_9_17_port, nextSum(16) => 
                           sigMatrix_9_16_port, nextSum(15) => 
                           sigMatrix_9_15_port, nextSum(14) => 
                           sigMatrix_9_14_port, nextSum(13) => 
                           sigMatrix_9_13_port, nextSum(12) => 
                           sigMatrix_9_12_port, nextSum(11) => 
                           sigMatrix_9_11_port, nextSum(10) => 
                           sigMatrix_9_10_port, nextSum(9) => 
                           sigMatrix_9_9_port, nextSum(8) => sigMatrix_9_8_port
                           , nextSum(7) => sigMatrix_9_7_port, nextSum(6) => 
                           sigMatrix_9_6_port, nextSum(5) => sigMatrix_9_5_port
                           , nextSum(4) => sigMatrix_9_4_port, nextSum(3) => 
                           sigMatrix_9_3_port, nextSum(2) => sigMatrix_9_2_port
                           , nextSum(1) => sigMatrix_9_1_port, nextSum(0) => 
                           sigMatrix_9_0_port);
   booth_mul_row_1_10 : booth_mul_row_N64_RADIX3_6 port map( prevA(63) => 
                           sigMatrix_9_127_port, prevA(62) => 
                           sigMatrix_9_126_port, prevA(61) => 
                           sigMatrix_9_125_port, prevA(60) => 
                           sigMatrix_9_124_port, prevA(59) => 
                           sigMatrix_9_123_port, prevA(58) => 
                           sigMatrix_9_122_port, prevA(57) => 
                           sigMatrix_9_121_port, prevA(56) => 
                           sigMatrix_9_120_port, prevA(55) => 
                           sigMatrix_9_119_port, prevA(54) => 
                           sigMatrix_9_118_port, prevA(53) => 
                           sigMatrix_9_117_port, prevA(52) => 
                           sigMatrix_9_116_port, prevA(51) => 
                           sigMatrix_9_115_port, prevA(50) => 
                           sigMatrix_9_114_port, prevA(49) => 
                           sigMatrix_9_113_port, prevA(48) => 
                           sigMatrix_9_112_port, prevA(47) => 
                           sigMatrix_9_111_port, prevA(46) => 
                           sigMatrix_9_110_port, prevA(45) => 
                           sigMatrix_9_109_port, prevA(44) => 
                           sigMatrix_9_108_port, prevA(43) => 
                           sigMatrix_9_107_port, prevA(42) => 
                           sigMatrix_9_106_port, prevA(41) => 
                           sigMatrix_9_105_port, prevA(40) => 
                           sigMatrix_9_104_port, prevA(39) => 
                           sigMatrix_9_103_port, prevA(38) => 
                           sigMatrix_9_102_port, prevA(37) => 
                           sigMatrix_9_101_port, prevA(36) => 
                           sigMatrix_9_100_port, prevA(35) => 
                           sigMatrix_9_99_port, prevA(34) => 
                           sigMatrix_9_98_port, prevA(33) => 
                           sigMatrix_9_97_port, prevA(32) => 
                           sigMatrix_9_96_port, prevA(31) => 
                           sigMatrix_9_95_port, prevA(30) => 
                           sigMatrix_9_94_port, prevA(29) => 
                           sigMatrix_9_93_port, prevA(28) => 
                           sigMatrix_9_92_port, prevA(27) => 
                           sigMatrix_9_91_port, prevA(26) => 
                           sigMatrix_9_90_port, prevA(25) => 
                           sigMatrix_9_89_port, prevA(24) => 
                           sigMatrix_9_88_port, prevA(23) => 
                           sigMatrix_9_87_port, prevA(22) => 
                           sigMatrix_9_86_port, prevA(21) => 
                           sigMatrix_9_85_port, prevA(20) => 
                           sigMatrix_9_84_port, prevA(19) => 
                           sigMatrix_9_83_port, prevA(18) => 
                           sigMatrix_9_82_port, prevA(17) => 
                           sigMatrix_9_81_port, prevA(16) => 
                           sigMatrix_9_80_port, prevA(15) => 
                           sigMatrix_9_79_port, prevA(14) => 
                           sigMatrix_9_78_port, prevA(13) => 
                           sigMatrix_9_77_port, prevA(12) => 
                           sigMatrix_9_76_port, prevA(11) => 
                           sigMatrix_9_75_port, prevA(10) => 
                           sigMatrix_9_74_port, prevA(9) => sigMatrix_9_73_port
                           , prevA(8) => sigMatrix_9_72_port, prevA(7) => 
                           sigMatrix_9_71_port, prevA(6) => sigMatrix_9_70_port
                           , prevA(5) => sigMatrix_9_69_port, prevA(4) => 
                           sigMatrix_9_68_port, prevA(3) => sigMatrix_9_67_port
                           , prevA(2) => sigMatrix_9_66_port, prevA(1) => 
                           sigMatrix_9_65_port, prevA(0) => n1, prevSum(63) => 
                           sigMatrix_9_63_port, prevSum(62) => 
                           sigMatrix_9_62_port, prevSum(61) => 
                           sigMatrix_9_61_port, prevSum(60) => 
                           sigMatrix_9_60_port, prevSum(59) => 
                           sigMatrix_9_59_port, prevSum(58) => 
                           sigMatrix_9_58_port, prevSum(57) => 
                           sigMatrix_9_57_port, prevSum(56) => 
                           sigMatrix_9_56_port, prevSum(55) => 
                           sigMatrix_9_55_port, prevSum(54) => 
                           sigMatrix_9_54_port, prevSum(53) => 
                           sigMatrix_9_53_port, prevSum(52) => 
                           sigMatrix_9_52_port, prevSum(51) => 
                           sigMatrix_9_51_port, prevSum(50) => 
                           sigMatrix_9_50_port, prevSum(49) => 
                           sigMatrix_9_49_port, prevSum(48) => 
                           sigMatrix_9_48_port, prevSum(47) => 
                           sigMatrix_9_47_port, prevSum(46) => 
                           sigMatrix_9_46_port, prevSum(45) => 
                           sigMatrix_9_45_port, prevSum(44) => 
                           sigMatrix_9_44_port, prevSum(43) => 
                           sigMatrix_9_43_port, prevSum(42) => 
                           sigMatrix_9_42_port, prevSum(41) => 
                           sigMatrix_9_41_port, prevSum(40) => 
                           sigMatrix_9_40_port, prevSum(39) => 
                           sigMatrix_9_39_port, prevSum(38) => 
                           sigMatrix_9_38_port, prevSum(37) => 
                           sigMatrix_9_37_port, prevSum(36) => 
                           sigMatrix_9_36_port, prevSum(35) => 
                           sigMatrix_9_35_port, prevSum(34) => 
                           sigMatrix_9_34_port, prevSum(33) => 
                           sigMatrix_9_33_port, prevSum(32) => 
                           sigMatrix_9_32_port, prevSum(31) => 
                           sigMatrix_9_31_port, prevSum(30) => 
                           sigMatrix_9_30_port, prevSum(29) => 
                           sigMatrix_9_29_port, prevSum(28) => 
                           sigMatrix_9_28_port, prevSum(27) => 
                           sigMatrix_9_27_port, prevSum(26) => 
                           sigMatrix_9_26_port, prevSum(25) => 
                           sigMatrix_9_25_port, prevSum(24) => 
                           sigMatrix_9_24_port, prevSum(23) => 
                           sigMatrix_9_23_port, prevSum(22) => 
                           sigMatrix_9_22_port, prevSum(21) => 
                           sigMatrix_9_21_port, prevSum(20) => 
                           sigMatrix_9_20_port, prevSum(19) => 
                           sigMatrix_9_19_port, prevSum(18) => 
                           sigMatrix_9_18_port, prevSum(17) => 
                           sigMatrix_9_17_port, prevSum(16) => 
                           sigMatrix_9_16_port, prevSum(15) => 
                           sigMatrix_9_15_port, prevSum(14) => 
                           sigMatrix_9_14_port, prevSum(13) => 
                           sigMatrix_9_13_port, prevSum(12) => 
                           sigMatrix_9_12_port, prevSum(11) => 
                           sigMatrix_9_11_port, prevSum(10) => 
                           sigMatrix_9_10_port, prevSum(9) => 
                           sigMatrix_9_9_port, prevSum(8) => sigMatrix_9_8_port
                           , prevSum(7) => sigMatrix_9_7_port, prevSum(6) => 
                           sigMatrix_9_6_port, prevSum(5) => sigMatrix_9_5_port
                           , prevSum(4) => sigMatrix_9_4_port, prevSum(3) => 
                           sigMatrix_9_3_port, prevSum(2) => sigMatrix_9_2_port
                           , prevSum(1) => sigMatrix_9_1_port, prevSum(0) => 
                           sigMatrix_9_0_port, encoderIn(2) => B(21), 
                           encoderIn(1) => B(20), encoderIn(0) => B(19), 
                           nextA(63) => sigMatrix_10_127_port, nextA(62) => 
                           sigMatrix_10_126_port, nextA(61) => 
                           sigMatrix_10_125_port, nextA(60) => 
                           sigMatrix_10_124_port, nextA(59) => 
                           sigMatrix_10_123_port, nextA(58) => 
                           sigMatrix_10_122_port, nextA(57) => 
                           sigMatrix_10_121_port, nextA(56) => 
                           sigMatrix_10_120_port, nextA(55) => 
                           sigMatrix_10_119_port, nextA(54) => 
                           sigMatrix_10_118_port, nextA(53) => 
                           sigMatrix_10_117_port, nextA(52) => 
                           sigMatrix_10_116_port, nextA(51) => 
                           sigMatrix_10_115_port, nextA(50) => 
                           sigMatrix_10_114_port, nextA(49) => 
                           sigMatrix_10_113_port, nextA(48) => 
                           sigMatrix_10_112_port, nextA(47) => 
                           sigMatrix_10_111_port, nextA(46) => 
                           sigMatrix_10_110_port, nextA(45) => 
                           sigMatrix_10_109_port, nextA(44) => 
                           sigMatrix_10_108_port, nextA(43) => 
                           sigMatrix_10_107_port, nextA(42) => 
                           sigMatrix_10_106_port, nextA(41) => 
                           sigMatrix_10_105_port, nextA(40) => 
                           sigMatrix_10_104_port, nextA(39) => 
                           sigMatrix_10_103_port, nextA(38) => 
                           sigMatrix_10_102_port, nextA(37) => 
                           sigMatrix_10_101_port, nextA(36) => 
                           sigMatrix_10_100_port, nextA(35) => 
                           sigMatrix_10_99_port, nextA(34) => 
                           sigMatrix_10_98_port, nextA(33) => 
                           sigMatrix_10_97_port, nextA(32) => 
                           sigMatrix_10_96_port, nextA(31) => 
                           sigMatrix_10_95_port, nextA(30) => 
                           sigMatrix_10_94_port, nextA(29) => 
                           sigMatrix_10_93_port, nextA(28) => 
                           sigMatrix_10_92_port, nextA(27) => 
                           sigMatrix_10_91_port, nextA(26) => 
                           sigMatrix_10_90_port, nextA(25) => 
                           sigMatrix_10_89_port, nextA(24) => 
                           sigMatrix_10_88_port, nextA(23) => 
                           sigMatrix_10_87_port, nextA(22) => 
                           sigMatrix_10_86_port, nextA(21) => 
                           sigMatrix_10_85_port, nextA(20) => 
                           sigMatrix_10_84_port, nextA(19) => 
                           sigMatrix_10_83_port, nextA(18) => 
                           sigMatrix_10_82_port, nextA(17) => 
                           sigMatrix_10_81_port, nextA(16) => 
                           sigMatrix_10_80_port, nextA(15) => 
                           sigMatrix_10_79_port, nextA(14) => 
                           sigMatrix_10_78_port, nextA(13) => 
                           sigMatrix_10_77_port, nextA(12) => 
                           sigMatrix_10_76_port, nextA(11) => 
                           sigMatrix_10_75_port, nextA(10) => 
                           sigMatrix_10_74_port, nextA(9) => 
                           sigMatrix_10_73_port, nextA(8) => 
                           sigMatrix_10_72_port, nextA(7) => 
                           sigMatrix_10_71_port, nextA(6) => 
                           sigMatrix_10_70_port, nextA(5) => 
                           sigMatrix_10_69_port, nextA(4) => 
                           sigMatrix_10_68_port, nextA(3) => 
                           sigMatrix_10_67_port, nextA(2) => 
                           sigMatrix_10_66_port, nextA(1) => 
                           sigMatrix_10_65_port, nextA(0) => n_3231, 
                           nextSum(63) => sigMatrix_10_63_port, nextSum(62) => 
                           sigMatrix_10_62_port, nextSum(61) => 
                           sigMatrix_10_61_port, nextSum(60) => 
                           sigMatrix_10_60_port, nextSum(59) => 
                           sigMatrix_10_59_port, nextSum(58) => 
                           sigMatrix_10_58_port, nextSum(57) => 
                           sigMatrix_10_57_port, nextSum(56) => 
                           sigMatrix_10_56_port, nextSum(55) => 
                           sigMatrix_10_55_port, nextSum(54) => 
                           sigMatrix_10_54_port, nextSum(53) => 
                           sigMatrix_10_53_port, nextSum(52) => 
                           sigMatrix_10_52_port, nextSum(51) => 
                           sigMatrix_10_51_port, nextSum(50) => 
                           sigMatrix_10_50_port, nextSum(49) => 
                           sigMatrix_10_49_port, nextSum(48) => 
                           sigMatrix_10_48_port, nextSum(47) => 
                           sigMatrix_10_47_port, nextSum(46) => 
                           sigMatrix_10_46_port, nextSum(45) => 
                           sigMatrix_10_45_port, nextSum(44) => 
                           sigMatrix_10_44_port, nextSum(43) => 
                           sigMatrix_10_43_port, nextSum(42) => 
                           sigMatrix_10_42_port, nextSum(41) => 
                           sigMatrix_10_41_port, nextSum(40) => 
                           sigMatrix_10_40_port, nextSum(39) => 
                           sigMatrix_10_39_port, nextSum(38) => 
                           sigMatrix_10_38_port, nextSum(37) => 
                           sigMatrix_10_37_port, nextSum(36) => 
                           sigMatrix_10_36_port, nextSum(35) => 
                           sigMatrix_10_35_port, nextSum(34) => 
                           sigMatrix_10_34_port, nextSum(33) => 
                           sigMatrix_10_33_port, nextSum(32) => 
                           sigMatrix_10_32_port, nextSum(31) => 
                           sigMatrix_10_31_port, nextSum(30) => 
                           sigMatrix_10_30_port, nextSum(29) => 
                           sigMatrix_10_29_port, nextSum(28) => 
                           sigMatrix_10_28_port, nextSum(27) => 
                           sigMatrix_10_27_port, nextSum(26) => 
                           sigMatrix_10_26_port, nextSum(25) => 
                           sigMatrix_10_25_port, nextSum(24) => 
                           sigMatrix_10_24_port, nextSum(23) => 
                           sigMatrix_10_23_port, nextSum(22) => 
                           sigMatrix_10_22_port, nextSum(21) => 
                           sigMatrix_10_21_port, nextSum(20) => 
                           sigMatrix_10_20_port, nextSum(19) => 
                           sigMatrix_10_19_port, nextSum(18) => 
                           sigMatrix_10_18_port, nextSum(17) => 
                           sigMatrix_10_17_port, nextSum(16) => 
                           sigMatrix_10_16_port, nextSum(15) => 
                           sigMatrix_10_15_port, nextSum(14) => 
                           sigMatrix_10_14_port, nextSum(13) => 
                           sigMatrix_10_13_port, nextSum(12) => 
                           sigMatrix_10_12_port, nextSum(11) => 
                           sigMatrix_10_11_port, nextSum(10) => 
                           sigMatrix_10_10_port, nextSum(9) => 
                           sigMatrix_10_9_port, nextSum(8) => 
                           sigMatrix_10_8_port, nextSum(7) => 
                           sigMatrix_10_7_port, nextSum(6) => 
                           sigMatrix_10_6_port, nextSum(5) => 
                           sigMatrix_10_5_port, nextSum(4) => 
                           sigMatrix_10_4_port, nextSum(3) => 
                           sigMatrix_10_3_port, nextSum(2) => 
                           sigMatrix_10_2_port, nextSum(1) => 
                           sigMatrix_10_1_port, nextSum(0) => 
                           sigMatrix_10_0_port);
   booth_mul_row_1_11 : booth_mul_row_N64_RADIX3_5 port map( prevA(63) => 
                           sigMatrix_10_127_port, prevA(62) => 
                           sigMatrix_10_126_port, prevA(61) => 
                           sigMatrix_10_125_port, prevA(60) => 
                           sigMatrix_10_124_port, prevA(59) => 
                           sigMatrix_10_123_port, prevA(58) => 
                           sigMatrix_10_122_port, prevA(57) => 
                           sigMatrix_10_121_port, prevA(56) => 
                           sigMatrix_10_120_port, prevA(55) => 
                           sigMatrix_10_119_port, prevA(54) => 
                           sigMatrix_10_118_port, prevA(53) => 
                           sigMatrix_10_117_port, prevA(52) => 
                           sigMatrix_10_116_port, prevA(51) => 
                           sigMatrix_10_115_port, prevA(50) => 
                           sigMatrix_10_114_port, prevA(49) => 
                           sigMatrix_10_113_port, prevA(48) => 
                           sigMatrix_10_112_port, prevA(47) => 
                           sigMatrix_10_111_port, prevA(46) => 
                           sigMatrix_10_110_port, prevA(45) => 
                           sigMatrix_10_109_port, prevA(44) => 
                           sigMatrix_10_108_port, prevA(43) => 
                           sigMatrix_10_107_port, prevA(42) => 
                           sigMatrix_10_106_port, prevA(41) => 
                           sigMatrix_10_105_port, prevA(40) => 
                           sigMatrix_10_104_port, prevA(39) => 
                           sigMatrix_10_103_port, prevA(38) => 
                           sigMatrix_10_102_port, prevA(37) => 
                           sigMatrix_10_101_port, prevA(36) => 
                           sigMatrix_10_100_port, prevA(35) => 
                           sigMatrix_10_99_port, prevA(34) => 
                           sigMatrix_10_98_port, prevA(33) => 
                           sigMatrix_10_97_port, prevA(32) => 
                           sigMatrix_10_96_port, prevA(31) => 
                           sigMatrix_10_95_port, prevA(30) => 
                           sigMatrix_10_94_port, prevA(29) => 
                           sigMatrix_10_93_port, prevA(28) => 
                           sigMatrix_10_92_port, prevA(27) => 
                           sigMatrix_10_91_port, prevA(26) => 
                           sigMatrix_10_90_port, prevA(25) => 
                           sigMatrix_10_89_port, prevA(24) => 
                           sigMatrix_10_88_port, prevA(23) => 
                           sigMatrix_10_87_port, prevA(22) => 
                           sigMatrix_10_86_port, prevA(21) => 
                           sigMatrix_10_85_port, prevA(20) => 
                           sigMatrix_10_84_port, prevA(19) => 
                           sigMatrix_10_83_port, prevA(18) => 
                           sigMatrix_10_82_port, prevA(17) => 
                           sigMatrix_10_81_port, prevA(16) => 
                           sigMatrix_10_80_port, prevA(15) => 
                           sigMatrix_10_79_port, prevA(14) => 
                           sigMatrix_10_78_port, prevA(13) => 
                           sigMatrix_10_77_port, prevA(12) => 
                           sigMatrix_10_76_port, prevA(11) => 
                           sigMatrix_10_75_port, prevA(10) => 
                           sigMatrix_10_74_port, prevA(9) => 
                           sigMatrix_10_73_port, prevA(8) => 
                           sigMatrix_10_72_port, prevA(7) => 
                           sigMatrix_10_71_port, prevA(6) => 
                           sigMatrix_10_70_port, prevA(5) => 
                           sigMatrix_10_69_port, prevA(4) => 
                           sigMatrix_10_68_port, prevA(3) => 
                           sigMatrix_10_67_port, prevA(2) => 
                           sigMatrix_10_66_port, prevA(1) => 
                           sigMatrix_10_65_port, prevA(0) => n1, prevSum(63) =>
                           sigMatrix_10_63_port, prevSum(62) => 
                           sigMatrix_10_62_port, prevSum(61) => 
                           sigMatrix_10_61_port, prevSum(60) => 
                           sigMatrix_10_60_port, prevSum(59) => 
                           sigMatrix_10_59_port, prevSum(58) => 
                           sigMatrix_10_58_port, prevSum(57) => 
                           sigMatrix_10_57_port, prevSum(56) => 
                           sigMatrix_10_56_port, prevSum(55) => 
                           sigMatrix_10_55_port, prevSum(54) => 
                           sigMatrix_10_54_port, prevSum(53) => 
                           sigMatrix_10_53_port, prevSum(52) => 
                           sigMatrix_10_52_port, prevSum(51) => 
                           sigMatrix_10_51_port, prevSum(50) => 
                           sigMatrix_10_50_port, prevSum(49) => 
                           sigMatrix_10_49_port, prevSum(48) => 
                           sigMatrix_10_48_port, prevSum(47) => 
                           sigMatrix_10_47_port, prevSum(46) => 
                           sigMatrix_10_46_port, prevSum(45) => 
                           sigMatrix_10_45_port, prevSum(44) => 
                           sigMatrix_10_44_port, prevSum(43) => 
                           sigMatrix_10_43_port, prevSum(42) => 
                           sigMatrix_10_42_port, prevSum(41) => 
                           sigMatrix_10_41_port, prevSum(40) => 
                           sigMatrix_10_40_port, prevSum(39) => 
                           sigMatrix_10_39_port, prevSum(38) => 
                           sigMatrix_10_38_port, prevSum(37) => 
                           sigMatrix_10_37_port, prevSum(36) => 
                           sigMatrix_10_36_port, prevSum(35) => 
                           sigMatrix_10_35_port, prevSum(34) => 
                           sigMatrix_10_34_port, prevSum(33) => 
                           sigMatrix_10_33_port, prevSum(32) => 
                           sigMatrix_10_32_port, prevSum(31) => 
                           sigMatrix_10_31_port, prevSum(30) => 
                           sigMatrix_10_30_port, prevSum(29) => 
                           sigMatrix_10_29_port, prevSum(28) => 
                           sigMatrix_10_28_port, prevSum(27) => 
                           sigMatrix_10_27_port, prevSum(26) => 
                           sigMatrix_10_26_port, prevSum(25) => 
                           sigMatrix_10_25_port, prevSum(24) => 
                           sigMatrix_10_24_port, prevSum(23) => 
                           sigMatrix_10_23_port, prevSum(22) => 
                           sigMatrix_10_22_port, prevSum(21) => 
                           sigMatrix_10_21_port, prevSum(20) => 
                           sigMatrix_10_20_port, prevSum(19) => 
                           sigMatrix_10_19_port, prevSum(18) => 
                           sigMatrix_10_18_port, prevSum(17) => 
                           sigMatrix_10_17_port, prevSum(16) => 
                           sigMatrix_10_16_port, prevSum(15) => 
                           sigMatrix_10_15_port, prevSum(14) => 
                           sigMatrix_10_14_port, prevSum(13) => 
                           sigMatrix_10_13_port, prevSum(12) => 
                           sigMatrix_10_12_port, prevSum(11) => 
                           sigMatrix_10_11_port, prevSum(10) => 
                           sigMatrix_10_10_port, prevSum(9) => 
                           sigMatrix_10_9_port, prevSum(8) => 
                           sigMatrix_10_8_port, prevSum(7) => 
                           sigMatrix_10_7_port, prevSum(6) => 
                           sigMatrix_10_6_port, prevSum(5) => 
                           sigMatrix_10_5_port, prevSum(4) => 
                           sigMatrix_10_4_port, prevSum(3) => 
                           sigMatrix_10_3_port, prevSum(2) => 
                           sigMatrix_10_2_port, prevSum(1) => 
                           sigMatrix_10_1_port, prevSum(0) => 
                           sigMatrix_10_0_port, encoderIn(2) => B(23), 
                           encoderIn(1) => B(22), encoderIn(0) => B(21), 
                           nextA(63) => sigMatrix_11_127_port, nextA(62) => 
                           sigMatrix_11_126_port, nextA(61) => 
                           sigMatrix_11_125_port, nextA(60) => 
                           sigMatrix_11_124_port, nextA(59) => 
                           sigMatrix_11_123_port, nextA(58) => 
                           sigMatrix_11_122_port, nextA(57) => 
                           sigMatrix_11_121_port, nextA(56) => 
                           sigMatrix_11_120_port, nextA(55) => 
                           sigMatrix_11_119_port, nextA(54) => 
                           sigMatrix_11_118_port, nextA(53) => 
                           sigMatrix_11_117_port, nextA(52) => 
                           sigMatrix_11_116_port, nextA(51) => 
                           sigMatrix_11_115_port, nextA(50) => 
                           sigMatrix_11_114_port, nextA(49) => 
                           sigMatrix_11_113_port, nextA(48) => 
                           sigMatrix_11_112_port, nextA(47) => 
                           sigMatrix_11_111_port, nextA(46) => 
                           sigMatrix_11_110_port, nextA(45) => 
                           sigMatrix_11_109_port, nextA(44) => 
                           sigMatrix_11_108_port, nextA(43) => 
                           sigMatrix_11_107_port, nextA(42) => 
                           sigMatrix_11_106_port, nextA(41) => 
                           sigMatrix_11_105_port, nextA(40) => 
                           sigMatrix_11_104_port, nextA(39) => 
                           sigMatrix_11_103_port, nextA(38) => 
                           sigMatrix_11_102_port, nextA(37) => 
                           sigMatrix_11_101_port, nextA(36) => 
                           sigMatrix_11_100_port, nextA(35) => 
                           sigMatrix_11_99_port, nextA(34) => 
                           sigMatrix_11_98_port, nextA(33) => 
                           sigMatrix_11_97_port, nextA(32) => 
                           sigMatrix_11_96_port, nextA(31) => 
                           sigMatrix_11_95_port, nextA(30) => 
                           sigMatrix_11_94_port, nextA(29) => 
                           sigMatrix_11_93_port, nextA(28) => 
                           sigMatrix_11_92_port, nextA(27) => 
                           sigMatrix_11_91_port, nextA(26) => 
                           sigMatrix_11_90_port, nextA(25) => 
                           sigMatrix_11_89_port, nextA(24) => 
                           sigMatrix_11_88_port, nextA(23) => 
                           sigMatrix_11_87_port, nextA(22) => 
                           sigMatrix_11_86_port, nextA(21) => 
                           sigMatrix_11_85_port, nextA(20) => 
                           sigMatrix_11_84_port, nextA(19) => 
                           sigMatrix_11_83_port, nextA(18) => 
                           sigMatrix_11_82_port, nextA(17) => 
                           sigMatrix_11_81_port, nextA(16) => 
                           sigMatrix_11_80_port, nextA(15) => 
                           sigMatrix_11_79_port, nextA(14) => 
                           sigMatrix_11_78_port, nextA(13) => 
                           sigMatrix_11_77_port, nextA(12) => 
                           sigMatrix_11_76_port, nextA(11) => 
                           sigMatrix_11_75_port, nextA(10) => 
                           sigMatrix_11_74_port, nextA(9) => 
                           sigMatrix_11_73_port, nextA(8) => 
                           sigMatrix_11_72_port, nextA(7) => 
                           sigMatrix_11_71_port, nextA(6) => 
                           sigMatrix_11_70_port, nextA(5) => 
                           sigMatrix_11_69_port, nextA(4) => 
                           sigMatrix_11_68_port, nextA(3) => 
                           sigMatrix_11_67_port, nextA(2) => 
                           sigMatrix_11_66_port, nextA(1) => 
                           sigMatrix_11_65_port, nextA(0) => n_3232, 
                           nextSum(63) => sigMatrix_11_63_port, nextSum(62) => 
                           sigMatrix_11_62_port, nextSum(61) => 
                           sigMatrix_11_61_port, nextSum(60) => 
                           sigMatrix_11_60_port, nextSum(59) => 
                           sigMatrix_11_59_port, nextSum(58) => 
                           sigMatrix_11_58_port, nextSum(57) => 
                           sigMatrix_11_57_port, nextSum(56) => 
                           sigMatrix_11_56_port, nextSum(55) => 
                           sigMatrix_11_55_port, nextSum(54) => 
                           sigMatrix_11_54_port, nextSum(53) => 
                           sigMatrix_11_53_port, nextSum(52) => 
                           sigMatrix_11_52_port, nextSum(51) => 
                           sigMatrix_11_51_port, nextSum(50) => 
                           sigMatrix_11_50_port, nextSum(49) => 
                           sigMatrix_11_49_port, nextSum(48) => 
                           sigMatrix_11_48_port, nextSum(47) => 
                           sigMatrix_11_47_port, nextSum(46) => 
                           sigMatrix_11_46_port, nextSum(45) => 
                           sigMatrix_11_45_port, nextSum(44) => 
                           sigMatrix_11_44_port, nextSum(43) => 
                           sigMatrix_11_43_port, nextSum(42) => 
                           sigMatrix_11_42_port, nextSum(41) => 
                           sigMatrix_11_41_port, nextSum(40) => 
                           sigMatrix_11_40_port, nextSum(39) => 
                           sigMatrix_11_39_port, nextSum(38) => 
                           sigMatrix_11_38_port, nextSum(37) => 
                           sigMatrix_11_37_port, nextSum(36) => 
                           sigMatrix_11_36_port, nextSum(35) => 
                           sigMatrix_11_35_port, nextSum(34) => 
                           sigMatrix_11_34_port, nextSum(33) => 
                           sigMatrix_11_33_port, nextSum(32) => 
                           sigMatrix_11_32_port, nextSum(31) => 
                           sigMatrix_11_31_port, nextSum(30) => 
                           sigMatrix_11_30_port, nextSum(29) => 
                           sigMatrix_11_29_port, nextSum(28) => 
                           sigMatrix_11_28_port, nextSum(27) => 
                           sigMatrix_11_27_port, nextSum(26) => 
                           sigMatrix_11_26_port, nextSum(25) => 
                           sigMatrix_11_25_port, nextSum(24) => 
                           sigMatrix_11_24_port, nextSum(23) => 
                           sigMatrix_11_23_port, nextSum(22) => 
                           sigMatrix_11_22_port, nextSum(21) => 
                           sigMatrix_11_21_port, nextSum(20) => 
                           sigMatrix_11_20_port, nextSum(19) => 
                           sigMatrix_11_19_port, nextSum(18) => 
                           sigMatrix_11_18_port, nextSum(17) => 
                           sigMatrix_11_17_port, nextSum(16) => 
                           sigMatrix_11_16_port, nextSum(15) => 
                           sigMatrix_11_15_port, nextSum(14) => 
                           sigMatrix_11_14_port, nextSum(13) => 
                           sigMatrix_11_13_port, nextSum(12) => 
                           sigMatrix_11_12_port, nextSum(11) => 
                           sigMatrix_11_11_port, nextSum(10) => 
                           sigMatrix_11_10_port, nextSum(9) => 
                           sigMatrix_11_9_port, nextSum(8) => 
                           sigMatrix_11_8_port, nextSum(7) => 
                           sigMatrix_11_7_port, nextSum(6) => 
                           sigMatrix_11_6_port, nextSum(5) => 
                           sigMatrix_11_5_port, nextSum(4) => 
                           sigMatrix_11_4_port, nextSum(3) => 
                           sigMatrix_11_3_port, nextSum(2) => 
                           sigMatrix_11_2_port, nextSum(1) => 
                           sigMatrix_11_1_port, nextSum(0) => 
                           sigMatrix_11_0_port);
   booth_mul_row_1_12 : booth_mul_row_N64_RADIX3_4 port map( prevA(63) => 
                           sigMatrix_11_127_port, prevA(62) => 
                           sigMatrix_11_126_port, prevA(61) => 
                           sigMatrix_11_125_port, prevA(60) => 
                           sigMatrix_11_124_port, prevA(59) => 
                           sigMatrix_11_123_port, prevA(58) => 
                           sigMatrix_11_122_port, prevA(57) => 
                           sigMatrix_11_121_port, prevA(56) => 
                           sigMatrix_11_120_port, prevA(55) => 
                           sigMatrix_11_119_port, prevA(54) => 
                           sigMatrix_11_118_port, prevA(53) => 
                           sigMatrix_11_117_port, prevA(52) => 
                           sigMatrix_11_116_port, prevA(51) => 
                           sigMatrix_11_115_port, prevA(50) => 
                           sigMatrix_11_114_port, prevA(49) => 
                           sigMatrix_11_113_port, prevA(48) => 
                           sigMatrix_11_112_port, prevA(47) => 
                           sigMatrix_11_111_port, prevA(46) => 
                           sigMatrix_11_110_port, prevA(45) => 
                           sigMatrix_11_109_port, prevA(44) => 
                           sigMatrix_11_108_port, prevA(43) => 
                           sigMatrix_11_107_port, prevA(42) => 
                           sigMatrix_11_106_port, prevA(41) => 
                           sigMatrix_11_105_port, prevA(40) => 
                           sigMatrix_11_104_port, prevA(39) => 
                           sigMatrix_11_103_port, prevA(38) => 
                           sigMatrix_11_102_port, prevA(37) => 
                           sigMatrix_11_101_port, prevA(36) => 
                           sigMatrix_11_100_port, prevA(35) => 
                           sigMatrix_11_99_port, prevA(34) => 
                           sigMatrix_11_98_port, prevA(33) => 
                           sigMatrix_11_97_port, prevA(32) => 
                           sigMatrix_11_96_port, prevA(31) => 
                           sigMatrix_11_95_port, prevA(30) => 
                           sigMatrix_11_94_port, prevA(29) => 
                           sigMatrix_11_93_port, prevA(28) => 
                           sigMatrix_11_92_port, prevA(27) => 
                           sigMatrix_11_91_port, prevA(26) => 
                           sigMatrix_11_90_port, prevA(25) => 
                           sigMatrix_11_89_port, prevA(24) => 
                           sigMatrix_11_88_port, prevA(23) => 
                           sigMatrix_11_87_port, prevA(22) => 
                           sigMatrix_11_86_port, prevA(21) => 
                           sigMatrix_11_85_port, prevA(20) => 
                           sigMatrix_11_84_port, prevA(19) => 
                           sigMatrix_11_83_port, prevA(18) => 
                           sigMatrix_11_82_port, prevA(17) => 
                           sigMatrix_11_81_port, prevA(16) => 
                           sigMatrix_11_80_port, prevA(15) => 
                           sigMatrix_11_79_port, prevA(14) => 
                           sigMatrix_11_78_port, prevA(13) => 
                           sigMatrix_11_77_port, prevA(12) => 
                           sigMatrix_11_76_port, prevA(11) => 
                           sigMatrix_11_75_port, prevA(10) => 
                           sigMatrix_11_74_port, prevA(9) => 
                           sigMatrix_11_73_port, prevA(8) => 
                           sigMatrix_11_72_port, prevA(7) => 
                           sigMatrix_11_71_port, prevA(6) => 
                           sigMatrix_11_70_port, prevA(5) => 
                           sigMatrix_11_69_port, prevA(4) => 
                           sigMatrix_11_68_port, prevA(3) => 
                           sigMatrix_11_67_port, prevA(2) => 
                           sigMatrix_11_66_port, prevA(1) => 
                           sigMatrix_11_65_port, prevA(0) => n1, prevSum(63) =>
                           sigMatrix_11_63_port, prevSum(62) => 
                           sigMatrix_11_62_port, prevSum(61) => 
                           sigMatrix_11_61_port, prevSum(60) => 
                           sigMatrix_11_60_port, prevSum(59) => 
                           sigMatrix_11_59_port, prevSum(58) => 
                           sigMatrix_11_58_port, prevSum(57) => 
                           sigMatrix_11_57_port, prevSum(56) => 
                           sigMatrix_11_56_port, prevSum(55) => 
                           sigMatrix_11_55_port, prevSum(54) => 
                           sigMatrix_11_54_port, prevSum(53) => 
                           sigMatrix_11_53_port, prevSum(52) => 
                           sigMatrix_11_52_port, prevSum(51) => 
                           sigMatrix_11_51_port, prevSum(50) => 
                           sigMatrix_11_50_port, prevSum(49) => 
                           sigMatrix_11_49_port, prevSum(48) => 
                           sigMatrix_11_48_port, prevSum(47) => 
                           sigMatrix_11_47_port, prevSum(46) => 
                           sigMatrix_11_46_port, prevSum(45) => 
                           sigMatrix_11_45_port, prevSum(44) => 
                           sigMatrix_11_44_port, prevSum(43) => 
                           sigMatrix_11_43_port, prevSum(42) => 
                           sigMatrix_11_42_port, prevSum(41) => 
                           sigMatrix_11_41_port, prevSum(40) => 
                           sigMatrix_11_40_port, prevSum(39) => 
                           sigMatrix_11_39_port, prevSum(38) => 
                           sigMatrix_11_38_port, prevSum(37) => 
                           sigMatrix_11_37_port, prevSum(36) => 
                           sigMatrix_11_36_port, prevSum(35) => 
                           sigMatrix_11_35_port, prevSum(34) => 
                           sigMatrix_11_34_port, prevSum(33) => 
                           sigMatrix_11_33_port, prevSum(32) => 
                           sigMatrix_11_32_port, prevSum(31) => 
                           sigMatrix_11_31_port, prevSum(30) => 
                           sigMatrix_11_30_port, prevSum(29) => 
                           sigMatrix_11_29_port, prevSum(28) => 
                           sigMatrix_11_28_port, prevSum(27) => 
                           sigMatrix_11_27_port, prevSum(26) => 
                           sigMatrix_11_26_port, prevSum(25) => 
                           sigMatrix_11_25_port, prevSum(24) => 
                           sigMatrix_11_24_port, prevSum(23) => 
                           sigMatrix_11_23_port, prevSum(22) => 
                           sigMatrix_11_22_port, prevSum(21) => 
                           sigMatrix_11_21_port, prevSum(20) => 
                           sigMatrix_11_20_port, prevSum(19) => 
                           sigMatrix_11_19_port, prevSum(18) => 
                           sigMatrix_11_18_port, prevSum(17) => 
                           sigMatrix_11_17_port, prevSum(16) => 
                           sigMatrix_11_16_port, prevSum(15) => 
                           sigMatrix_11_15_port, prevSum(14) => 
                           sigMatrix_11_14_port, prevSum(13) => 
                           sigMatrix_11_13_port, prevSum(12) => 
                           sigMatrix_11_12_port, prevSum(11) => 
                           sigMatrix_11_11_port, prevSum(10) => 
                           sigMatrix_11_10_port, prevSum(9) => 
                           sigMatrix_11_9_port, prevSum(8) => 
                           sigMatrix_11_8_port, prevSum(7) => 
                           sigMatrix_11_7_port, prevSum(6) => 
                           sigMatrix_11_6_port, prevSum(5) => 
                           sigMatrix_11_5_port, prevSum(4) => 
                           sigMatrix_11_4_port, prevSum(3) => 
                           sigMatrix_11_3_port, prevSum(2) => 
                           sigMatrix_11_2_port, prevSum(1) => 
                           sigMatrix_11_1_port, prevSum(0) => 
                           sigMatrix_11_0_port, encoderIn(2) => B(25), 
                           encoderIn(1) => B(24), encoderIn(0) => B(23), 
                           nextA(63) => sigMatrix_12_127_port, nextA(62) => 
                           sigMatrix_12_126_port, nextA(61) => 
                           sigMatrix_12_125_port, nextA(60) => 
                           sigMatrix_12_124_port, nextA(59) => 
                           sigMatrix_12_123_port, nextA(58) => 
                           sigMatrix_12_122_port, nextA(57) => 
                           sigMatrix_12_121_port, nextA(56) => 
                           sigMatrix_12_120_port, nextA(55) => 
                           sigMatrix_12_119_port, nextA(54) => 
                           sigMatrix_12_118_port, nextA(53) => 
                           sigMatrix_12_117_port, nextA(52) => 
                           sigMatrix_12_116_port, nextA(51) => 
                           sigMatrix_12_115_port, nextA(50) => 
                           sigMatrix_12_114_port, nextA(49) => 
                           sigMatrix_12_113_port, nextA(48) => 
                           sigMatrix_12_112_port, nextA(47) => 
                           sigMatrix_12_111_port, nextA(46) => 
                           sigMatrix_12_110_port, nextA(45) => 
                           sigMatrix_12_109_port, nextA(44) => 
                           sigMatrix_12_108_port, nextA(43) => 
                           sigMatrix_12_107_port, nextA(42) => 
                           sigMatrix_12_106_port, nextA(41) => 
                           sigMatrix_12_105_port, nextA(40) => 
                           sigMatrix_12_104_port, nextA(39) => 
                           sigMatrix_12_103_port, nextA(38) => 
                           sigMatrix_12_102_port, nextA(37) => 
                           sigMatrix_12_101_port, nextA(36) => 
                           sigMatrix_12_100_port, nextA(35) => 
                           sigMatrix_12_99_port, nextA(34) => 
                           sigMatrix_12_98_port, nextA(33) => 
                           sigMatrix_12_97_port, nextA(32) => 
                           sigMatrix_12_96_port, nextA(31) => 
                           sigMatrix_12_95_port, nextA(30) => 
                           sigMatrix_12_94_port, nextA(29) => 
                           sigMatrix_12_93_port, nextA(28) => 
                           sigMatrix_12_92_port, nextA(27) => 
                           sigMatrix_12_91_port, nextA(26) => 
                           sigMatrix_12_90_port, nextA(25) => 
                           sigMatrix_12_89_port, nextA(24) => 
                           sigMatrix_12_88_port, nextA(23) => 
                           sigMatrix_12_87_port, nextA(22) => 
                           sigMatrix_12_86_port, nextA(21) => 
                           sigMatrix_12_85_port, nextA(20) => 
                           sigMatrix_12_84_port, nextA(19) => 
                           sigMatrix_12_83_port, nextA(18) => 
                           sigMatrix_12_82_port, nextA(17) => 
                           sigMatrix_12_81_port, nextA(16) => 
                           sigMatrix_12_80_port, nextA(15) => 
                           sigMatrix_12_79_port, nextA(14) => 
                           sigMatrix_12_78_port, nextA(13) => 
                           sigMatrix_12_77_port, nextA(12) => 
                           sigMatrix_12_76_port, nextA(11) => 
                           sigMatrix_12_75_port, nextA(10) => 
                           sigMatrix_12_74_port, nextA(9) => 
                           sigMatrix_12_73_port, nextA(8) => 
                           sigMatrix_12_72_port, nextA(7) => 
                           sigMatrix_12_71_port, nextA(6) => 
                           sigMatrix_12_70_port, nextA(5) => 
                           sigMatrix_12_69_port, nextA(4) => 
                           sigMatrix_12_68_port, nextA(3) => 
                           sigMatrix_12_67_port, nextA(2) => 
                           sigMatrix_12_66_port, nextA(1) => 
                           sigMatrix_12_65_port, nextA(0) => n_3233, 
                           nextSum(63) => sigMatrix_12_63_port, nextSum(62) => 
                           sigMatrix_12_62_port, nextSum(61) => 
                           sigMatrix_12_61_port, nextSum(60) => 
                           sigMatrix_12_60_port, nextSum(59) => 
                           sigMatrix_12_59_port, nextSum(58) => 
                           sigMatrix_12_58_port, nextSum(57) => 
                           sigMatrix_12_57_port, nextSum(56) => 
                           sigMatrix_12_56_port, nextSum(55) => 
                           sigMatrix_12_55_port, nextSum(54) => 
                           sigMatrix_12_54_port, nextSum(53) => 
                           sigMatrix_12_53_port, nextSum(52) => 
                           sigMatrix_12_52_port, nextSum(51) => 
                           sigMatrix_12_51_port, nextSum(50) => 
                           sigMatrix_12_50_port, nextSum(49) => 
                           sigMatrix_12_49_port, nextSum(48) => 
                           sigMatrix_12_48_port, nextSum(47) => 
                           sigMatrix_12_47_port, nextSum(46) => 
                           sigMatrix_12_46_port, nextSum(45) => 
                           sigMatrix_12_45_port, nextSum(44) => 
                           sigMatrix_12_44_port, nextSum(43) => 
                           sigMatrix_12_43_port, nextSum(42) => 
                           sigMatrix_12_42_port, nextSum(41) => 
                           sigMatrix_12_41_port, nextSum(40) => 
                           sigMatrix_12_40_port, nextSum(39) => 
                           sigMatrix_12_39_port, nextSum(38) => 
                           sigMatrix_12_38_port, nextSum(37) => 
                           sigMatrix_12_37_port, nextSum(36) => 
                           sigMatrix_12_36_port, nextSum(35) => 
                           sigMatrix_12_35_port, nextSum(34) => 
                           sigMatrix_12_34_port, nextSum(33) => 
                           sigMatrix_12_33_port, nextSum(32) => 
                           sigMatrix_12_32_port, nextSum(31) => 
                           sigMatrix_12_31_port, nextSum(30) => 
                           sigMatrix_12_30_port, nextSum(29) => 
                           sigMatrix_12_29_port, nextSum(28) => 
                           sigMatrix_12_28_port, nextSum(27) => 
                           sigMatrix_12_27_port, nextSum(26) => 
                           sigMatrix_12_26_port, nextSum(25) => 
                           sigMatrix_12_25_port, nextSum(24) => 
                           sigMatrix_12_24_port, nextSum(23) => 
                           sigMatrix_12_23_port, nextSum(22) => 
                           sigMatrix_12_22_port, nextSum(21) => 
                           sigMatrix_12_21_port, nextSum(20) => 
                           sigMatrix_12_20_port, nextSum(19) => 
                           sigMatrix_12_19_port, nextSum(18) => 
                           sigMatrix_12_18_port, nextSum(17) => 
                           sigMatrix_12_17_port, nextSum(16) => 
                           sigMatrix_12_16_port, nextSum(15) => 
                           sigMatrix_12_15_port, nextSum(14) => 
                           sigMatrix_12_14_port, nextSum(13) => 
                           sigMatrix_12_13_port, nextSum(12) => 
                           sigMatrix_12_12_port, nextSum(11) => 
                           sigMatrix_12_11_port, nextSum(10) => 
                           sigMatrix_12_10_port, nextSum(9) => 
                           sigMatrix_12_9_port, nextSum(8) => 
                           sigMatrix_12_8_port, nextSum(7) => 
                           sigMatrix_12_7_port, nextSum(6) => 
                           sigMatrix_12_6_port, nextSum(5) => 
                           sigMatrix_12_5_port, nextSum(4) => 
                           sigMatrix_12_4_port, nextSum(3) => 
                           sigMatrix_12_3_port, nextSum(2) => 
                           sigMatrix_12_2_port, nextSum(1) => 
                           sigMatrix_12_1_port, nextSum(0) => 
                           sigMatrix_12_0_port);
   booth_mul_row_1_13 : booth_mul_row_N64_RADIX3_3 port map( prevA(63) => 
                           sigMatrix_12_127_port, prevA(62) => 
                           sigMatrix_12_126_port, prevA(61) => 
                           sigMatrix_12_125_port, prevA(60) => 
                           sigMatrix_12_124_port, prevA(59) => 
                           sigMatrix_12_123_port, prevA(58) => 
                           sigMatrix_12_122_port, prevA(57) => 
                           sigMatrix_12_121_port, prevA(56) => 
                           sigMatrix_12_120_port, prevA(55) => 
                           sigMatrix_12_119_port, prevA(54) => 
                           sigMatrix_12_118_port, prevA(53) => 
                           sigMatrix_12_117_port, prevA(52) => 
                           sigMatrix_12_116_port, prevA(51) => 
                           sigMatrix_12_115_port, prevA(50) => 
                           sigMatrix_12_114_port, prevA(49) => 
                           sigMatrix_12_113_port, prevA(48) => 
                           sigMatrix_12_112_port, prevA(47) => 
                           sigMatrix_12_111_port, prevA(46) => 
                           sigMatrix_12_110_port, prevA(45) => 
                           sigMatrix_12_109_port, prevA(44) => 
                           sigMatrix_12_108_port, prevA(43) => 
                           sigMatrix_12_107_port, prevA(42) => 
                           sigMatrix_12_106_port, prevA(41) => 
                           sigMatrix_12_105_port, prevA(40) => 
                           sigMatrix_12_104_port, prevA(39) => 
                           sigMatrix_12_103_port, prevA(38) => 
                           sigMatrix_12_102_port, prevA(37) => 
                           sigMatrix_12_101_port, prevA(36) => 
                           sigMatrix_12_100_port, prevA(35) => 
                           sigMatrix_12_99_port, prevA(34) => 
                           sigMatrix_12_98_port, prevA(33) => 
                           sigMatrix_12_97_port, prevA(32) => 
                           sigMatrix_12_96_port, prevA(31) => 
                           sigMatrix_12_95_port, prevA(30) => 
                           sigMatrix_12_94_port, prevA(29) => 
                           sigMatrix_12_93_port, prevA(28) => 
                           sigMatrix_12_92_port, prevA(27) => 
                           sigMatrix_12_91_port, prevA(26) => 
                           sigMatrix_12_90_port, prevA(25) => 
                           sigMatrix_12_89_port, prevA(24) => 
                           sigMatrix_12_88_port, prevA(23) => 
                           sigMatrix_12_87_port, prevA(22) => 
                           sigMatrix_12_86_port, prevA(21) => 
                           sigMatrix_12_85_port, prevA(20) => 
                           sigMatrix_12_84_port, prevA(19) => 
                           sigMatrix_12_83_port, prevA(18) => 
                           sigMatrix_12_82_port, prevA(17) => 
                           sigMatrix_12_81_port, prevA(16) => 
                           sigMatrix_12_80_port, prevA(15) => 
                           sigMatrix_12_79_port, prevA(14) => 
                           sigMatrix_12_78_port, prevA(13) => 
                           sigMatrix_12_77_port, prevA(12) => 
                           sigMatrix_12_76_port, prevA(11) => 
                           sigMatrix_12_75_port, prevA(10) => 
                           sigMatrix_12_74_port, prevA(9) => 
                           sigMatrix_12_73_port, prevA(8) => 
                           sigMatrix_12_72_port, prevA(7) => 
                           sigMatrix_12_71_port, prevA(6) => 
                           sigMatrix_12_70_port, prevA(5) => 
                           sigMatrix_12_69_port, prevA(4) => 
                           sigMatrix_12_68_port, prevA(3) => 
                           sigMatrix_12_67_port, prevA(2) => 
                           sigMatrix_12_66_port, prevA(1) => 
                           sigMatrix_12_65_port, prevA(0) => n1, prevSum(63) =>
                           sigMatrix_12_63_port, prevSum(62) => 
                           sigMatrix_12_62_port, prevSum(61) => 
                           sigMatrix_12_61_port, prevSum(60) => 
                           sigMatrix_12_60_port, prevSum(59) => 
                           sigMatrix_12_59_port, prevSum(58) => 
                           sigMatrix_12_58_port, prevSum(57) => 
                           sigMatrix_12_57_port, prevSum(56) => 
                           sigMatrix_12_56_port, prevSum(55) => 
                           sigMatrix_12_55_port, prevSum(54) => 
                           sigMatrix_12_54_port, prevSum(53) => 
                           sigMatrix_12_53_port, prevSum(52) => 
                           sigMatrix_12_52_port, prevSum(51) => 
                           sigMatrix_12_51_port, prevSum(50) => 
                           sigMatrix_12_50_port, prevSum(49) => 
                           sigMatrix_12_49_port, prevSum(48) => 
                           sigMatrix_12_48_port, prevSum(47) => 
                           sigMatrix_12_47_port, prevSum(46) => 
                           sigMatrix_12_46_port, prevSum(45) => 
                           sigMatrix_12_45_port, prevSum(44) => 
                           sigMatrix_12_44_port, prevSum(43) => 
                           sigMatrix_12_43_port, prevSum(42) => 
                           sigMatrix_12_42_port, prevSum(41) => 
                           sigMatrix_12_41_port, prevSum(40) => 
                           sigMatrix_12_40_port, prevSum(39) => 
                           sigMatrix_12_39_port, prevSum(38) => 
                           sigMatrix_12_38_port, prevSum(37) => 
                           sigMatrix_12_37_port, prevSum(36) => 
                           sigMatrix_12_36_port, prevSum(35) => 
                           sigMatrix_12_35_port, prevSum(34) => 
                           sigMatrix_12_34_port, prevSum(33) => 
                           sigMatrix_12_33_port, prevSum(32) => 
                           sigMatrix_12_32_port, prevSum(31) => 
                           sigMatrix_12_31_port, prevSum(30) => 
                           sigMatrix_12_30_port, prevSum(29) => 
                           sigMatrix_12_29_port, prevSum(28) => 
                           sigMatrix_12_28_port, prevSum(27) => 
                           sigMatrix_12_27_port, prevSum(26) => 
                           sigMatrix_12_26_port, prevSum(25) => 
                           sigMatrix_12_25_port, prevSum(24) => 
                           sigMatrix_12_24_port, prevSum(23) => 
                           sigMatrix_12_23_port, prevSum(22) => 
                           sigMatrix_12_22_port, prevSum(21) => 
                           sigMatrix_12_21_port, prevSum(20) => 
                           sigMatrix_12_20_port, prevSum(19) => 
                           sigMatrix_12_19_port, prevSum(18) => 
                           sigMatrix_12_18_port, prevSum(17) => 
                           sigMatrix_12_17_port, prevSum(16) => 
                           sigMatrix_12_16_port, prevSum(15) => 
                           sigMatrix_12_15_port, prevSum(14) => 
                           sigMatrix_12_14_port, prevSum(13) => 
                           sigMatrix_12_13_port, prevSum(12) => 
                           sigMatrix_12_12_port, prevSum(11) => 
                           sigMatrix_12_11_port, prevSum(10) => 
                           sigMatrix_12_10_port, prevSum(9) => 
                           sigMatrix_12_9_port, prevSum(8) => 
                           sigMatrix_12_8_port, prevSum(7) => 
                           sigMatrix_12_7_port, prevSum(6) => 
                           sigMatrix_12_6_port, prevSum(5) => 
                           sigMatrix_12_5_port, prevSum(4) => 
                           sigMatrix_12_4_port, prevSum(3) => 
                           sigMatrix_12_3_port, prevSum(2) => 
                           sigMatrix_12_2_port, prevSum(1) => 
                           sigMatrix_12_1_port, prevSum(0) => 
                           sigMatrix_12_0_port, encoderIn(2) => B(27), 
                           encoderIn(1) => B(26), encoderIn(0) => B(25), 
                           nextA(63) => sigMatrix_13_127_port, nextA(62) => 
                           sigMatrix_13_126_port, nextA(61) => 
                           sigMatrix_13_125_port, nextA(60) => 
                           sigMatrix_13_124_port, nextA(59) => 
                           sigMatrix_13_123_port, nextA(58) => 
                           sigMatrix_13_122_port, nextA(57) => 
                           sigMatrix_13_121_port, nextA(56) => 
                           sigMatrix_13_120_port, nextA(55) => 
                           sigMatrix_13_119_port, nextA(54) => 
                           sigMatrix_13_118_port, nextA(53) => 
                           sigMatrix_13_117_port, nextA(52) => 
                           sigMatrix_13_116_port, nextA(51) => 
                           sigMatrix_13_115_port, nextA(50) => 
                           sigMatrix_13_114_port, nextA(49) => 
                           sigMatrix_13_113_port, nextA(48) => 
                           sigMatrix_13_112_port, nextA(47) => 
                           sigMatrix_13_111_port, nextA(46) => 
                           sigMatrix_13_110_port, nextA(45) => 
                           sigMatrix_13_109_port, nextA(44) => 
                           sigMatrix_13_108_port, nextA(43) => 
                           sigMatrix_13_107_port, nextA(42) => 
                           sigMatrix_13_106_port, nextA(41) => 
                           sigMatrix_13_105_port, nextA(40) => 
                           sigMatrix_13_104_port, nextA(39) => 
                           sigMatrix_13_103_port, nextA(38) => 
                           sigMatrix_13_102_port, nextA(37) => 
                           sigMatrix_13_101_port, nextA(36) => 
                           sigMatrix_13_100_port, nextA(35) => 
                           sigMatrix_13_99_port, nextA(34) => 
                           sigMatrix_13_98_port, nextA(33) => 
                           sigMatrix_13_97_port, nextA(32) => 
                           sigMatrix_13_96_port, nextA(31) => 
                           sigMatrix_13_95_port, nextA(30) => 
                           sigMatrix_13_94_port, nextA(29) => 
                           sigMatrix_13_93_port, nextA(28) => 
                           sigMatrix_13_92_port, nextA(27) => 
                           sigMatrix_13_91_port, nextA(26) => 
                           sigMatrix_13_90_port, nextA(25) => 
                           sigMatrix_13_89_port, nextA(24) => 
                           sigMatrix_13_88_port, nextA(23) => 
                           sigMatrix_13_87_port, nextA(22) => 
                           sigMatrix_13_86_port, nextA(21) => 
                           sigMatrix_13_85_port, nextA(20) => 
                           sigMatrix_13_84_port, nextA(19) => 
                           sigMatrix_13_83_port, nextA(18) => 
                           sigMatrix_13_82_port, nextA(17) => 
                           sigMatrix_13_81_port, nextA(16) => 
                           sigMatrix_13_80_port, nextA(15) => 
                           sigMatrix_13_79_port, nextA(14) => 
                           sigMatrix_13_78_port, nextA(13) => 
                           sigMatrix_13_77_port, nextA(12) => 
                           sigMatrix_13_76_port, nextA(11) => 
                           sigMatrix_13_75_port, nextA(10) => 
                           sigMatrix_13_74_port, nextA(9) => 
                           sigMatrix_13_73_port, nextA(8) => 
                           sigMatrix_13_72_port, nextA(7) => 
                           sigMatrix_13_71_port, nextA(6) => 
                           sigMatrix_13_70_port, nextA(5) => 
                           sigMatrix_13_69_port, nextA(4) => 
                           sigMatrix_13_68_port, nextA(3) => 
                           sigMatrix_13_67_port, nextA(2) => 
                           sigMatrix_13_66_port, nextA(1) => 
                           sigMatrix_13_65_port, nextA(0) => n_3234, 
                           nextSum(63) => sigMatrix_13_63_port, nextSum(62) => 
                           sigMatrix_13_62_port, nextSum(61) => 
                           sigMatrix_13_61_port, nextSum(60) => 
                           sigMatrix_13_60_port, nextSum(59) => 
                           sigMatrix_13_59_port, nextSum(58) => 
                           sigMatrix_13_58_port, nextSum(57) => 
                           sigMatrix_13_57_port, nextSum(56) => 
                           sigMatrix_13_56_port, nextSum(55) => 
                           sigMatrix_13_55_port, nextSum(54) => 
                           sigMatrix_13_54_port, nextSum(53) => 
                           sigMatrix_13_53_port, nextSum(52) => 
                           sigMatrix_13_52_port, nextSum(51) => 
                           sigMatrix_13_51_port, nextSum(50) => 
                           sigMatrix_13_50_port, nextSum(49) => 
                           sigMatrix_13_49_port, nextSum(48) => 
                           sigMatrix_13_48_port, nextSum(47) => 
                           sigMatrix_13_47_port, nextSum(46) => 
                           sigMatrix_13_46_port, nextSum(45) => 
                           sigMatrix_13_45_port, nextSum(44) => 
                           sigMatrix_13_44_port, nextSum(43) => 
                           sigMatrix_13_43_port, nextSum(42) => 
                           sigMatrix_13_42_port, nextSum(41) => 
                           sigMatrix_13_41_port, nextSum(40) => 
                           sigMatrix_13_40_port, nextSum(39) => 
                           sigMatrix_13_39_port, nextSum(38) => 
                           sigMatrix_13_38_port, nextSum(37) => 
                           sigMatrix_13_37_port, nextSum(36) => 
                           sigMatrix_13_36_port, nextSum(35) => 
                           sigMatrix_13_35_port, nextSum(34) => 
                           sigMatrix_13_34_port, nextSum(33) => 
                           sigMatrix_13_33_port, nextSum(32) => 
                           sigMatrix_13_32_port, nextSum(31) => 
                           sigMatrix_13_31_port, nextSum(30) => 
                           sigMatrix_13_30_port, nextSum(29) => 
                           sigMatrix_13_29_port, nextSum(28) => 
                           sigMatrix_13_28_port, nextSum(27) => 
                           sigMatrix_13_27_port, nextSum(26) => 
                           sigMatrix_13_26_port, nextSum(25) => 
                           sigMatrix_13_25_port, nextSum(24) => 
                           sigMatrix_13_24_port, nextSum(23) => 
                           sigMatrix_13_23_port, nextSum(22) => 
                           sigMatrix_13_22_port, nextSum(21) => 
                           sigMatrix_13_21_port, nextSum(20) => 
                           sigMatrix_13_20_port, nextSum(19) => 
                           sigMatrix_13_19_port, nextSum(18) => 
                           sigMatrix_13_18_port, nextSum(17) => 
                           sigMatrix_13_17_port, nextSum(16) => 
                           sigMatrix_13_16_port, nextSum(15) => 
                           sigMatrix_13_15_port, nextSum(14) => 
                           sigMatrix_13_14_port, nextSum(13) => 
                           sigMatrix_13_13_port, nextSum(12) => 
                           sigMatrix_13_12_port, nextSum(11) => 
                           sigMatrix_13_11_port, nextSum(10) => 
                           sigMatrix_13_10_port, nextSum(9) => 
                           sigMatrix_13_9_port, nextSum(8) => 
                           sigMatrix_13_8_port, nextSum(7) => 
                           sigMatrix_13_7_port, nextSum(6) => 
                           sigMatrix_13_6_port, nextSum(5) => 
                           sigMatrix_13_5_port, nextSum(4) => 
                           sigMatrix_13_4_port, nextSum(3) => 
                           sigMatrix_13_3_port, nextSum(2) => 
                           sigMatrix_13_2_port, nextSum(1) => 
                           sigMatrix_13_1_port, nextSum(0) => 
                           sigMatrix_13_0_port);
   booth_mul_row_1_14 : booth_mul_row_N64_RADIX3_2 port map( prevA(63) => 
                           sigMatrix_13_127_port, prevA(62) => 
                           sigMatrix_13_126_port, prevA(61) => 
                           sigMatrix_13_125_port, prevA(60) => 
                           sigMatrix_13_124_port, prevA(59) => 
                           sigMatrix_13_123_port, prevA(58) => 
                           sigMatrix_13_122_port, prevA(57) => 
                           sigMatrix_13_121_port, prevA(56) => 
                           sigMatrix_13_120_port, prevA(55) => 
                           sigMatrix_13_119_port, prevA(54) => 
                           sigMatrix_13_118_port, prevA(53) => 
                           sigMatrix_13_117_port, prevA(52) => 
                           sigMatrix_13_116_port, prevA(51) => 
                           sigMatrix_13_115_port, prevA(50) => 
                           sigMatrix_13_114_port, prevA(49) => 
                           sigMatrix_13_113_port, prevA(48) => 
                           sigMatrix_13_112_port, prevA(47) => 
                           sigMatrix_13_111_port, prevA(46) => 
                           sigMatrix_13_110_port, prevA(45) => 
                           sigMatrix_13_109_port, prevA(44) => 
                           sigMatrix_13_108_port, prevA(43) => 
                           sigMatrix_13_107_port, prevA(42) => 
                           sigMatrix_13_106_port, prevA(41) => 
                           sigMatrix_13_105_port, prevA(40) => 
                           sigMatrix_13_104_port, prevA(39) => 
                           sigMatrix_13_103_port, prevA(38) => 
                           sigMatrix_13_102_port, prevA(37) => 
                           sigMatrix_13_101_port, prevA(36) => 
                           sigMatrix_13_100_port, prevA(35) => 
                           sigMatrix_13_99_port, prevA(34) => 
                           sigMatrix_13_98_port, prevA(33) => 
                           sigMatrix_13_97_port, prevA(32) => 
                           sigMatrix_13_96_port, prevA(31) => 
                           sigMatrix_13_95_port, prevA(30) => 
                           sigMatrix_13_94_port, prevA(29) => 
                           sigMatrix_13_93_port, prevA(28) => 
                           sigMatrix_13_92_port, prevA(27) => 
                           sigMatrix_13_91_port, prevA(26) => 
                           sigMatrix_13_90_port, prevA(25) => 
                           sigMatrix_13_89_port, prevA(24) => 
                           sigMatrix_13_88_port, prevA(23) => 
                           sigMatrix_13_87_port, prevA(22) => 
                           sigMatrix_13_86_port, prevA(21) => 
                           sigMatrix_13_85_port, prevA(20) => 
                           sigMatrix_13_84_port, prevA(19) => 
                           sigMatrix_13_83_port, prevA(18) => 
                           sigMatrix_13_82_port, prevA(17) => 
                           sigMatrix_13_81_port, prevA(16) => 
                           sigMatrix_13_80_port, prevA(15) => 
                           sigMatrix_13_79_port, prevA(14) => 
                           sigMatrix_13_78_port, prevA(13) => 
                           sigMatrix_13_77_port, prevA(12) => 
                           sigMatrix_13_76_port, prevA(11) => 
                           sigMatrix_13_75_port, prevA(10) => 
                           sigMatrix_13_74_port, prevA(9) => 
                           sigMatrix_13_73_port, prevA(8) => 
                           sigMatrix_13_72_port, prevA(7) => 
                           sigMatrix_13_71_port, prevA(6) => 
                           sigMatrix_13_70_port, prevA(5) => 
                           sigMatrix_13_69_port, prevA(4) => 
                           sigMatrix_13_68_port, prevA(3) => 
                           sigMatrix_13_67_port, prevA(2) => 
                           sigMatrix_13_66_port, prevA(1) => 
                           sigMatrix_13_65_port, prevA(0) => n1, prevSum(63) =>
                           sigMatrix_13_63_port, prevSum(62) => 
                           sigMatrix_13_62_port, prevSum(61) => 
                           sigMatrix_13_61_port, prevSum(60) => 
                           sigMatrix_13_60_port, prevSum(59) => 
                           sigMatrix_13_59_port, prevSum(58) => 
                           sigMatrix_13_58_port, prevSum(57) => 
                           sigMatrix_13_57_port, prevSum(56) => 
                           sigMatrix_13_56_port, prevSum(55) => 
                           sigMatrix_13_55_port, prevSum(54) => 
                           sigMatrix_13_54_port, prevSum(53) => 
                           sigMatrix_13_53_port, prevSum(52) => 
                           sigMatrix_13_52_port, prevSum(51) => 
                           sigMatrix_13_51_port, prevSum(50) => 
                           sigMatrix_13_50_port, prevSum(49) => 
                           sigMatrix_13_49_port, prevSum(48) => 
                           sigMatrix_13_48_port, prevSum(47) => 
                           sigMatrix_13_47_port, prevSum(46) => 
                           sigMatrix_13_46_port, prevSum(45) => 
                           sigMatrix_13_45_port, prevSum(44) => 
                           sigMatrix_13_44_port, prevSum(43) => 
                           sigMatrix_13_43_port, prevSum(42) => 
                           sigMatrix_13_42_port, prevSum(41) => 
                           sigMatrix_13_41_port, prevSum(40) => 
                           sigMatrix_13_40_port, prevSum(39) => 
                           sigMatrix_13_39_port, prevSum(38) => 
                           sigMatrix_13_38_port, prevSum(37) => 
                           sigMatrix_13_37_port, prevSum(36) => 
                           sigMatrix_13_36_port, prevSum(35) => 
                           sigMatrix_13_35_port, prevSum(34) => 
                           sigMatrix_13_34_port, prevSum(33) => 
                           sigMatrix_13_33_port, prevSum(32) => 
                           sigMatrix_13_32_port, prevSum(31) => 
                           sigMatrix_13_31_port, prevSum(30) => 
                           sigMatrix_13_30_port, prevSum(29) => 
                           sigMatrix_13_29_port, prevSum(28) => 
                           sigMatrix_13_28_port, prevSum(27) => 
                           sigMatrix_13_27_port, prevSum(26) => 
                           sigMatrix_13_26_port, prevSum(25) => 
                           sigMatrix_13_25_port, prevSum(24) => 
                           sigMatrix_13_24_port, prevSum(23) => 
                           sigMatrix_13_23_port, prevSum(22) => 
                           sigMatrix_13_22_port, prevSum(21) => 
                           sigMatrix_13_21_port, prevSum(20) => 
                           sigMatrix_13_20_port, prevSum(19) => 
                           sigMatrix_13_19_port, prevSum(18) => 
                           sigMatrix_13_18_port, prevSum(17) => 
                           sigMatrix_13_17_port, prevSum(16) => 
                           sigMatrix_13_16_port, prevSum(15) => 
                           sigMatrix_13_15_port, prevSum(14) => 
                           sigMatrix_13_14_port, prevSum(13) => 
                           sigMatrix_13_13_port, prevSum(12) => 
                           sigMatrix_13_12_port, prevSum(11) => 
                           sigMatrix_13_11_port, prevSum(10) => 
                           sigMatrix_13_10_port, prevSum(9) => 
                           sigMatrix_13_9_port, prevSum(8) => 
                           sigMatrix_13_8_port, prevSum(7) => 
                           sigMatrix_13_7_port, prevSum(6) => 
                           sigMatrix_13_6_port, prevSum(5) => 
                           sigMatrix_13_5_port, prevSum(4) => 
                           sigMatrix_13_4_port, prevSum(3) => 
                           sigMatrix_13_3_port, prevSum(2) => 
                           sigMatrix_13_2_port, prevSum(1) => 
                           sigMatrix_13_1_port, prevSum(0) => 
                           sigMatrix_13_0_port, encoderIn(2) => B(29), 
                           encoderIn(1) => B(28), encoderIn(0) => B(27), 
                           nextA(63) => sigMatrix_14_127_port, nextA(62) => 
                           sigMatrix_14_126_port, nextA(61) => 
                           sigMatrix_14_125_port, nextA(60) => 
                           sigMatrix_14_124_port, nextA(59) => 
                           sigMatrix_14_123_port, nextA(58) => 
                           sigMatrix_14_122_port, nextA(57) => 
                           sigMatrix_14_121_port, nextA(56) => 
                           sigMatrix_14_120_port, nextA(55) => 
                           sigMatrix_14_119_port, nextA(54) => 
                           sigMatrix_14_118_port, nextA(53) => 
                           sigMatrix_14_117_port, nextA(52) => 
                           sigMatrix_14_116_port, nextA(51) => 
                           sigMatrix_14_115_port, nextA(50) => 
                           sigMatrix_14_114_port, nextA(49) => 
                           sigMatrix_14_113_port, nextA(48) => 
                           sigMatrix_14_112_port, nextA(47) => 
                           sigMatrix_14_111_port, nextA(46) => 
                           sigMatrix_14_110_port, nextA(45) => 
                           sigMatrix_14_109_port, nextA(44) => 
                           sigMatrix_14_108_port, nextA(43) => 
                           sigMatrix_14_107_port, nextA(42) => 
                           sigMatrix_14_106_port, nextA(41) => 
                           sigMatrix_14_105_port, nextA(40) => 
                           sigMatrix_14_104_port, nextA(39) => 
                           sigMatrix_14_103_port, nextA(38) => 
                           sigMatrix_14_102_port, nextA(37) => 
                           sigMatrix_14_101_port, nextA(36) => 
                           sigMatrix_14_100_port, nextA(35) => 
                           sigMatrix_14_99_port, nextA(34) => 
                           sigMatrix_14_98_port, nextA(33) => 
                           sigMatrix_14_97_port, nextA(32) => 
                           sigMatrix_14_96_port, nextA(31) => 
                           sigMatrix_14_95_port, nextA(30) => 
                           sigMatrix_14_94_port, nextA(29) => 
                           sigMatrix_14_93_port, nextA(28) => 
                           sigMatrix_14_92_port, nextA(27) => 
                           sigMatrix_14_91_port, nextA(26) => 
                           sigMatrix_14_90_port, nextA(25) => 
                           sigMatrix_14_89_port, nextA(24) => 
                           sigMatrix_14_88_port, nextA(23) => 
                           sigMatrix_14_87_port, nextA(22) => 
                           sigMatrix_14_86_port, nextA(21) => 
                           sigMatrix_14_85_port, nextA(20) => 
                           sigMatrix_14_84_port, nextA(19) => 
                           sigMatrix_14_83_port, nextA(18) => 
                           sigMatrix_14_82_port, nextA(17) => 
                           sigMatrix_14_81_port, nextA(16) => 
                           sigMatrix_14_80_port, nextA(15) => 
                           sigMatrix_14_79_port, nextA(14) => 
                           sigMatrix_14_78_port, nextA(13) => 
                           sigMatrix_14_77_port, nextA(12) => 
                           sigMatrix_14_76_port, nextA(11) => 
                           sigMatrix_14_75_port, nextA(10) => 
                           sigMatrix_14_74_port, nextA(9) => 
                           sigMatrix_14_73_port, nextA(8) => 
                           sigMatrix_14_72_port, nextA(7) => 
                           sigMatrix_14_71_port, nextA(6) => 
                           sigMatrix_14_70_port, nextA(5) => 
                           sigMatrix_14_69_port, nextA(4) => 
                           sigMatrix_14_68_port, nextA(3) => 
                           sigMatrix_14_67_port, nextA(2) => 
                           sigMatrix_14_66_port, nextA(1) => 
                           sigMatrix_14_65_port, nextA(0) => n_3235, 
                           nextSum(63) => sigMatrix_14_63_port, nextSum(62) => 
                           sigMatrix_14_62_port, nextSum(61) => 
                           sigMatrix_14_61_port, nextSum(60) => 
                           sigMatrix_14_60_port, nextSum(59) => 
                           sigMatrix_14_59_port, nextSum(58) => 
                           sigMatrix_14_58_port, nextSum(57) => 
                           sigMatrix_14_57_port, nextSum(56) => 
                           sigMatrix_14_56_port, nextSum(55) => 
                           sigMatrix_14_55_port, nextSum(54) => 
                           sigMatrix_14_54_port, nextSum(53) => 
                           sigMatrix_14_53_port, nextSum(52) => 
                           sigMatrix_14_52_port, nextSum(51) => 
                           sigMatrix_14_51_port, nextSum(50) => 
                           sigMatrix_14_50_port, nextSum(49) => 
                           sigMatrix_14_49_port, nextSum(48) => 
                           sigMatrix_14_48_port, nextSum(47) => 
                           sigMatrix_14_47_port, nextSum(46) => 
                           sigMatrix_14_46_port, nextSum(45) => 
                           sigMatrix_14_45_port, nextSum(44) => 
                           sigMatrix_14_44_port, nextSum(43) => 
                           sigMatrix_14_43_port, nextSum(42) => 
                           sigMatrix_14_42_port, nextSum(41) => 
                           sigMatrix_14_41_port, nextSum(40) => 
                           sigMatrix_14_40_port, nextSum(39) => 
                           sigMatrix_14_39_port, nextSum(38) => 
                           sigMatrix_14_38_port, nextSum(37) => 
                           sigMatrix_14_37_port, nextSum(36) => 
                           sigMatrix_14_36_port, nextSum(35) => 
                           sigMatrix_14_35_port, nextSum(34) => 
                           sigMatrix_14_34_port, nextSum(33) => 
                           sigMatrix_14_33_port, nextSum(32) => 
                           sigMatrix_14_32_port, nextSum(31) => 
                           sigMatrix_14_31_port, nextSum(30) => 
                           sigMatrix_14_30_port, nextSum(29) => 
                           sigMatrix_14_29_port, nextSum(28) => 
                           sigMatrix_14_28_port, nextSum(27) => 
                           sigMatrix_14_27_port, nextSum(26) => 
                           sigMatrix_14_26_port, nextSum(25) => 
                           sigMatrix_14_25_port, nextSum(24) => 
                           sigMatrix_14_24_port, nextSum(23) => 
                           sigMatrix_14_23_port, nextSum(22) => 
                           sigMatrix_14_22_port, nextSum(21) => 
                           sigMatrix_14_21_port, nextSum(20) => 
                           sigMatrix_14_20_port, nextSum(19) => 
                           sigMatrix_14_19_port, nextSum(18) => 
                           sigMatrix_14_18_port, nextSum(17) => 
                           sigMatrix_14_17_port, nextSum(16) => 
                           sigMatrix_14_16_port, nextSum(15) => 
                           sigMatrix_14_15_port, nextSum(14) => 
                           sigMatrix_14_14_port, nextSum(13) => 
                           sigMatrix_14_13_port, nextSum(12) => 
                           sigMatrix_14_12_port, nextSum(11) => 
                           sigMatrix_14_11_port, nextSum(10) => 
                           sigMatrix_14_10_port, nextSum(9) => 
                           sigMatrix_14_9_port, nextSum(8) => 
                           sigMatrix_14_8_port, nextSum(7) => 
                           sigMatrix_14_7_port, nextSum(6) => 
                           sigMatrix_14_6_port, nextSum(5) => 
                           sigMatrix_14_5_port, nextSum(4) => 
                           sigMatrix_14_4_port, nextSum(3) => 
                           sigMatrix_14_3_port, nextSum(2) => 
                           sigMatrix_14_2_port, nextSum(1) => 
                           sigMatrix_14_1_port, nextSum(0) => 
                           sigMatrix_14_0_port);
   booth_mul_row_1_15 : booth_mul_row_N64_RADIX3_1 port map( prevA(63) => 
                           sigMatrix_14_127_port, prevA(62) => 
                           sigMatrix_14_126_port, prevA(61) => 
                           sigMatrix_14_125_port, prevA(60) => 
                           sigMatrix_14_124_port, prevA(59) => 
                           sigMatrix_14_123_port, prevA(58) => 
                           sigMatrix_14_122_port, prevA(57) => 
                           sigMatrix_14_121_port, prevA(56) => 
                           sigMatrix_14_120_port, prevA(55) => 
                           sigMatrix_14_119_port, prevA(54) => 
                           sigMatrix_14_118_port, prevA(53) => 
                           sigMatrix_14_117_port, prevA(52) => 
                           sigMatrix_14_116_port, prevA(51) => 
                           sigMatrix_14_115_port, prevA(50) => 
                           sigMatrix_14_114_port, prevA(49) => 
                           sigMatrix_14_113_port, prevA(48) => 
                           sigMatrix_14_112_port, prevA(47) => 
                           sigMatrix_14_111_port, prevA(46) => 
                           sigMatrix_14_110_port, prevA(45) => 
                           sigMatrix_14_109_port, prevA(44) => 
                           sigMatrix_14_108_port, prevA(43) => 
                           sigMatrix_14_107_port, prevA(42) => 
                           sigMatrix_14_106_port, prevA(41) => 
                           sigMatrix_14_105_port, prevA(40) => 
                           sigMatrix_14_104_port, prevA(39) => 
                           sigMatrix_14_103_port, prevA(38) => 
                           sigMatrix_14_102_port, prevA(37) => 
                           sigMatrix_14_101_port, prevA(36) => 
                           sigMatrix_14_100_port, prevA(35) => 
                           sigMatrix_14_99_port, prevA(34) => 
                           sigMatrix_14_98_port, prevA(33) => 
                           sigMatrix_14_97_port, prevA(32) => 
                           sigMatrix_14_96_port, prevA(31) => 
                           sigMatrix_14_95_port, prevA(30) => 
                           sigMatrix_14_94_port, prevA(29) => 
                           sigMatrix_14_93_port, prevA(28) => 
                           sigMatrix_14_92_port, prevA(27) => 
                           sigMatrix_14_91_port, prevA(26) => 
                           sigMatrix_14_90_port, prevA(25) => 
                           sigMatrix_14_89_port, prevA(24) => 
                           sigMatrix_14_88_port, prevA(23) => 
                           sigMatrix_14_87_port, prevA(22) => 
                           sigMatrix_14_86_port, prevA(21) => 
                           sigMatrix_14_85_port, prevA(20) => 
                           sigMatrix_14_84_port, prevA(19) => 
                           sigMatrix_14_83_port, prevA(18) => 
                           sigMatrix_14_82_port, prevA(17) => 
                           sigMatrix_14_81_port, prevA(16) => 
                           sigMatrix_14_80_port, prevA(15) => 
                           sigMatrix_14_79_port, prevA(14) => 
                           sigMatrix_14_78_port, prevA(13) => 
                           sigMatrix_14_77_port, prevA(12) => 
                           sigMatrix_14_76_port, prevA(11) => 
                           sigMatrix_14_75_port, prevA(10) => 
                           sigMatrix_14_74_port, prevA(9) => 
                           sigMatrix_14_73_port, prevA(8) => 
                           sigMatrix_14_72_port, prevA(7) => 
                           sigMatrix_14_71_port, prevA(6) => 
                           sigMatrix_14_70_port, prevA(5) => 
                           sigMatrix_14_69_port, prevA(4) => 
                           sigMatrix_14_68_port, prevA(3) => 
                           sigMatrix_14_67_port, prevA(2) => 
                           sigMatrix_14_66_port, prevA(1) => 
                           sigMatrix_14_65_port, prevA(0) => n1, prevSum(63) =>
                           sigMatrix_14_63_port, prevSum(62) => 
                           sigMatrix_14_62_port, prevSum(61) => 
                           sigMatrix_14_61_port, prevSum(60) => 
                           sigMatrix_14_60_port, prevSum(59) => 
                           sigMatrix_14_59_port, prevSum(58) => 
                           sigMatrix_14_58_port, prevSum(57) => 
                           sigMatrix_14_57_port, prevSum(56) => 
                           sigMatrix_14_56_port, prevSum(55) => 
                           sigMatrix_14_55_port, prevSum(54) => 
                           sigMatrix_14_54_port, prevSum(53) => 
                           sigMatrix_14_53_port, prevSum(52) => 
                           sigMatrix_14_52_port, prevSum(51) => 
                           sigMatrix_14_51_port, prevSum(50) => 
                           sigMatrix_14_50_port, prevSum(49) => 
                           sigMatrix_14_49_port, prevSum(48) => 
                           sigMatrix_14_48_port, prevSum(47) => 
                           sigMatrix_14_47_port, prevSum(46) => 
                           sigMatrix_14_46_port, prevSum(45) => 
                           sigMatrix_14_45_port, prevSum(44) => 
                           sigMatrix_14_44_port, prevSum(43) => 
                           sigMatrix_14_43_port, prevSum(42) => 
                           sigMatrix_14_42_port, prevSum(41) => 
                           sigMatrix_14_41_port, prevSum(40) => 
                           sigMatrix_14_40_port, prevSum(39) => 
                           sigMatrix_14_39_port, prevSum(38) => 
                           sigMatrix_14_38_port, prevSum(37) => 
                           sigMatrix_14_37_port, prevSum(36) => 
                           sigMatrix_14_36_port, prevSum(35) => 
                           sigMatrix_14_35_port, prevSum(34) => 
                           sigMatrix_14_34_port, prevSum(33) => 
                           sigMatrix_14_33_port, prevSum(32) => 
                           sigMatrix_14_32_port, prevSum(31) => 
                           sigMatrix_14_31_port, prevSum(30) => 
                           sigMatrix_14_30_port, prevSum(29) => 
                           sigMatrix_14_29_port, prevSum(28) => 
                           sigMatrix_14_28_port, prevSum(27) => 
                           sigMatrix_14_27_port, prevSum(26) => 
                           sigMatrix_14_26_port, prevSum(25) => 
                           sigMatrix_14_25_port, prevSum(24) => 
                           sigMatrix_14_24_port, prevSum(23) => 
                           sigMatrix_14_23_port, prevSum(22) => 
                           sigMatrix_14_22_port, prevSum(21) => 
                           sigMatrix_14_21_port, prevSum(20) => 
                           sigMatrix_14_20_port, prevSum(19) => 
                           sigMatrix_14_19_port, prevSum(18) => 
                           sigMatrix_14_18_port, prevSum(17) => 
                           sigMatrix_14_17_port, prevSum(16) => 
                           sigMatrix_14_16_port, prevSum(15) => 
                           sigMatrix_14_15_port, prevSum(14) => 
                           sigMatrix_14_14_port, prevSum(13) => 
                           sigMatrix_14_13_port, prevSum(12) => 
                           sigMatrix_14_12_port, prevSum(11) => 
                           sigMatrix_14_11_port, prevSum(10) => 
                           sigMatrix_14_10_port, prevSum(9) => 
                           sigMatrix_14_9_port, prevSum(8) => 
                           sigMatrix_14_8_port, prevSum(7) => 
                           sigMatrix_14_7_port, prevSum(6) => 
                           sigMatrix_14_6_port, prevSum(5) => 
                           sigMatrix_14_5_port, prevSum(4) => 
                           sigMatrix_14_4_port, prevSum(3) => 
                           sigMatrix_14_3_port, prevSum(2) => 
                           sigMatrix_14_2_port, prevSum(1) => 
                           sigMatrix_14_1_port, prevSum(0) => 
                           sigMatrix_14_0_port, encoderIn(2) => B(31), 
                           encoderIn(1) => B(30), encoderIn(0) => B(29), 
                           nextA(63) => n_3236, nextA(62) => n_3237, nextA(61) 
                           => n_3238, nextA(60) => n_3239, nextA(59) => n_3240,
                           nextA(58) => n_3241, nextA(57) => n_3242, nextA(56) 
                           => n_3243, nextA(55) => n_3244, nextA(54) => n_3245,
                           nextA(53) => n_3246, nextA(52) => n_3247, nextA(51) 
                           => n_3248, nextA(50) => n_3249, nextA(49) => n_3250,
                           nextA(48) => n_3251, nextA(47) => n_3252, nextA(46) 
                           => n_3253, nextA(45) => n_3254, nextA(44) => n_3255,
                           nextA(43) => n_3256, nextA(42) => n_3257, nextA(41) 
                           => n_3258, nextA(40) => n_3259, nextA(39) => n_3260,
                           nextA(38) => n_3261, nextA(37) => n_3262, nextA(36) 
                           => n_3263, nextA(35) => n_3264, nextA(34) => n_3265,
                           nextA(33) => n_3266, nextA(32) => n_3267, nextA(31) 
                           => n_3268, nextA(30) => n_3269, nextA(29) => n_3270,
                           nextA(28) => n_3271, nextA(27) => n_3272, nextA(26) 
                           => n_3273, nextA(25) => n_3274, nextA(24) => n_3275,
                           nextA(23) => n_3276, nextA(22) => n_3277, nextA(21) 
                           => n_3278, nextA(20) => n_3279, nextA(19) => n_3280,
                           nextA(18) => n_3281, nextA(17) => n_3282, nextA(16) 
                           => n_3283, nextA(15) => n_3284, nextA(14) => n_3285,
                           nextA(13) => n_3286, nextA(12) => n_3287, nextA(11) 
                           => n_3288, nextA(10) => n_3289, nextA(9) => n_3290, 
                           nextA(8) => n_3291, nextA(7) => n_3292, nextA(6) => 
                           n_3293, nextA(5) => n_3294, nextA(4) => n_3295, 
                           nextA(3) => n_3296, nextA(2) => n_3297, nextA(1) => 
                           n_3298, nextA(0) => n_3299, nextSum(63) => P(63), 
                           nextSum(62) => P(62), nextSum(61) => P(61), 
                           nextSum(60) => P(60), nextSum(59) => P(59), 
                           nextSum(58) => P(58), nextSum(57) => P(57), 
                           nextSum(56) => P(56), nextSum(55) => P(55), 
                           nextSum(54) => P(54), nextSum(53) => P(53), 
                           nextSum(52) => P(52), nextSum(51) => P(51), 
                           nextSum(50) => P(50), nextSum(49) => P(49), 
                           nextSum(48) => P(48), nextSum(47) => P(47), 
                           nextSum(46) => P(46), nextSum(45) => P(45), 
                           nextSum(44) => P(44), nextSum(43) => P(43), 
                           nextSum(42) => P(42), nextSum(41) => P(41), 
                           nextSum(40) => P(40), nextSum(39) => P(39), 
                           nextSum(38) => P(38), nextSum(37) => P(37), 
                           nextSum(36) => P(36), nextSum(35) => P(35), 
                           nextSum(34) => P(34), nextSum(33) => P(33), 
                           nextSum(32) => P(32), nextSum(31) => P(31), 
                           nextSum(30) => P(30), nextSum(29) => P(29), 
                           nextSum(28) => P(28), nextSum(27) => P(27), 
                           nextSum(26) => P(26), nextSum(25) => P(25), 
                           nextSum(24) => P(24), nextSum(23) => P(23), 
                           nextSum(22) => P(22), nextSum(21) => P(21), 
                           nextSum(20) => P(20), nextSum(19) => P(19), 
                           nextSum(18) => P(18), nextSum(17) => P(17), 
                           nextSum(16) => P(16), nextSum(15) => P(15), 
                           nextSum(14) => P(14), nextSum(13) => P(13), 
                           nextSum(12) => P(12), nextSum(11) => P(11), 
                           nextSum(10) => P(10), nextSum(9) => P(9), nextSum(8)
                           => P(8), nextSum(7) => P(7), nextSum(6) => P(6), 
                           nextSum(5) => P(5), nextSum(4) => P(4), nextSum(3) 
                           => P(3), nextSum(2) => P(2), nextSum(1) => P(1), 
                           nextSum(0) => P(0));

end SYN_booth_struct;
